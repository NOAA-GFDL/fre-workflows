netcdf \00010101.atmos_daily.tile3.ps {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float ps(time, grid_yt, grid_xt) ;
		ps:_FillValue = 1.e+20f ;
		ps:missing_value = 1.e+20f ;
		ps:units = "Pa" ;
		ps:long_name = "Surface Air Pressure" ;
		ps:cell_methods = "time: mean" ;
		ps:cell_measures = "area: area" ;
		ps:time_avg_info = "average_T1,average_T2,average_DT" ;
		ps:standard_name = "surface_air_pressure" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile3.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.0008770345, 0.4596241, 0.9892928, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.01035247, 0.004304647, 0.6546783, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.8534847, 0.8118016, 0.9951549, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9894952, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4452189, 0.3028796, 0.7140614, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9903189, 0.3150955, 0.0007410151, 0, 0.02645395, 
    0.9012984, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.681631, 0, 0, 0, 0.004980796, 0.7708192, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5536854, 0, 0, 0, 0.004666397, 0.9395298, 1,
  1, 1, 1, 1, 1, 1, 1, 0.9995009, 0.3626226, 0, 0, 0, 0, 0.8367797, 1,
  1, 1, 1, 1, 1, 0.8451425, 0.7016711, 0.3953246, 0, 0, 0, 0, 0.006316811, 
    0.8673657, 1 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 ps =
  102725.9, 102528.7, 98586.38, 96061.5, 96037.18, 94948.3, 92511.11, 
    93080.79, 86992.27, 82241.31, 79864.66, 80168.27, 83153.2, 81662.26, 
    92132.42,
  102801.9, 102847.9, 100454, 95164.36, 92360.48, 90441.01, 89173.73, 
    89488.77, 84384.66, 81596.21, 80756.05, 81452.87, 83664.66, 82508.3, 
    93602.62,
  93437.3, 89954.59, 95113.65, 93655.62, 86971.98, 85888.8, 88243.92, 
    87513.95, 82461.68, 80152.55, 79148.66, 79875.7, 81247.3, 82858.38, 
    95664.15,
  87229.85, 87364.13, 86455, 84795.25, 84514.4, 83015.91, 83914.03, 84264.99, 
    81871.01, 80545.11, 80241.02, 81801.64, 81307.41, 83403.87, 89431.2,
  88907.26, 87861.05, 88932.03, 88126.96, 87969.02, 86351.78, 85288.23, 
    84792.91, 83788.52, 85900.05, 101105.9, 101759.9, 91776.24, 92144.66, 
    84449.05,
  89198.58, 87365.05, 89850.87, 90759.34, 89860.98, 89429.14, 88675.27, 
    89076.17, 90665.34, 101759.6, 102652.5, 102695.1, 102467.9, 94264.06, 
    78802.7,
  88269.84, 87543.18, 89685.59, 91022.54, 90807.66, 90856.37, 90767.55, 
    92769.34, 96723.77, 102513.7, 102480.4, 102588, 102495.9, 88072.9, 
    78526.11,
  92049.99, 88810.77, 89255.62, 91129.02, 90816.2, 89804.95, 90397.95, 
    92232.53, 96464.91, 102372.4, 102351, 102514.5, 102400, 86771.23, 88512.46,
  95021.39, 90713, 89749.78, 90890.13, 90083.88, 87707.2, 88968.84, 91579.81, 
    101789.7, 102306.5, 102264.1, 102337.9, 102284.3, 94379.68, 96809.1,
  98213.41, 93543.38, 91879, 94293.34, 94557.85, 94708.63, 95624.86, 
    101621.4, 102193.4, 102168.8, 102151.9, 102170.5, 102178.4, 99864.89, 
    100940.6,
  102913, 102709.8, 98750.66, 96222.44, 96208.45, 95113.62, 92664.87, 
    93233.06, 87153.84, 82419.27, 80047.42, 80345.43, 83325.56, 81828.58, 
    92303.23,
  102847.4, 102941.8, 100600.8, 95315.88, 92495.01, 90587.91, 89330.8, 
    89636.45, 84562.96, 81768.54, 80929.61, 81622.12, 83836.64, 82658.89, 
    93760.24,
  93627.52, 90104.57, 95227.48, 93805.87, 87146.97, 86033, 88379.26, 
    87660.85, 82635.66, 80329.47, 79323.84, 80040.05, 81405.98, 83002.95, 
    95848.38,
  87393.75, 87407.99, 86596.42, 84931, 84641.26, 83147.23, 84042.85, 
    84396.09, 82033.97, 80706.84, 80404.96, 81973, 81463.43, 83578.58, 
    89581.94,
  89068.97, 87887.55, 89018.02, 88202.85, 88062.31, 86439.68, 85393.3, 
    84903.19, 83920.84, 85996.55, 101170, 101830.9, 91884.35, 92273.03, 
    84585.12,
  89283.08, 87398.5, 89902.91, 90815.76, 89935.55, 89494.55, 88751.24, 
    89153.43, 90745.38, 101797, 102767.2, 102798.5, 102568.9, 94381.1, 
    78980.23,
  88264.84, 87569.35, 89706.79, 91061.79, 90859.95, 90918.9, 90831.22, 
    92842.95, 96800.16, 102605.8, 102570.8, 102698.1, 102592.4, 88194.24, 
    78716.21,
  91974.26, 88778.63, 89243.98, 91121.76, 90832.38, 89836.19, 90429.56, 
    92314.63, 96533.95, 102482.9, 102448.6, 102665.5, 102514.6, 86922.94, 
    88665.01,
  94918.41, 90660.12, 89718.55, 90867.02, 90108.16, 87764.52, 89032.36, 
    91628.83, 101833.2, 102412.7, 102361.1, 102482.2, 102428.2, 94529.58, 
    96973.84,
  98090.34, 93461.03, 91796.64, 94212.03, 94519.91, 94690.29, 95641.7, 
    101679.7, 102323.1, 102296.4, 102282.9, 102325.2, 102349.8, 100037.2, 
    101079.4,
  102771.8, 102546.2, 98624.88, 96085.4, 96071.85, 95010.2, 92590.36, 
    93104.56, 87090.88, 82355.2, 79985.2, 80276.9, 83200.39, 81739.34, 92044.7,
  102640.8, 102737.6, 100430.6, 95182.19, 92382.81, 90464.73, 89217.42, 
    89523.56, 84488.28, 81665.7, 80828.47, 81509.17, 83698.01, 82568.52, 
    93523.82,
  93481.22, 89953.37, 95035.09, 93642.77, 87024.03, 85887.12, 88247.98, 
    87551.12, 82534.88, 80217.3, 79249.54, 79927.93, 81283.54, 82857.32, 
    95601.01,
  87270.01, 87123.18, 86399.75, 84779.54, 84492.71, 82989.17, 83895.71, 
    84249.41, 81912.48, 80605.52, 80257.64, 81788.11, 81344.56, 83349.13, 
    89391,
  88869.38, 87559.92, 88758.66, 87930.27, 87838.91, 86224.3, 85200.14, 
    84729.2, 83763.51, 85773.62, 100835.2, 101564.1, 91669.64, 92000.16, 
    84482.6,
  88984.41, 87056.33, 89596.9, 90521.12, 89682.98, 89228.73, 88500.98, 
    88895.64, 90477.16, 101455.7, 102447.2, 102480.3, 102241.2, 94132.74, 
    78816.07,
  87855.49, 87153.72, 89369.8, 90739.51, 90587.67, 90646.22, 90557.22, 
    92548.16, 96483.4, 102221, 102198.9, 102389.6, 102268.6, 87984.88, 
    78501.71,
  91484.62, 88298.62, 88837.44, 90736.17, 90517.58, 89529.61, 90121.29, 
    91998.96, 96187.06, 102069.9, 102052.7, 102311.2, 102156.5, 86727.32, 
    88339.76,
  94398.47, 90160.9, 89286.77, 90438.91, 89765.1, 87447.17, 88733.16, 
    91285.51, 101405.1, 101995.4, 101927.1, 102074.1, 102041.5, 94199.39, 
    96644.72,
  97518.66, 92930.19, 91312.92, 93714.59, 94105.16, 94264.98, 95225.12, 
    101223.3, 101879.9, 101859.1, 101851, 101899.6, 101952.4, 99675.77, 
    100739.4,
  102242.3, 102018, 98134.16, 95614.66, 95623.11, 94599.45, 92233.59, 
    92730.15, 86760.82, 82012.91, 79638.91, 79925.24, 82808.14, 81372.05, 
    91570.95,
  102071.9, 102238.2, 99949.75, 94708.59, 91963.96, 90085.52, 88839.5, 
    89166.88, 84157.74, 81327.8, 80477, 81137.84, 83310.3, 82207.35, 93046.82,
  93026.77, 89437.83, 94554.13, 93183.65, 86601.1, 85462.68, 87850.71, 
    87190.02, 82152.51, 79847.84, 78879.38, 79552.82, 80877.54, 82438.95, 
    95095.23,
  86761.28, 86596.86, 85968.94, 84304.17, 84051.69, 82591.38, 83514.47, 
    83864.16, 81518.24, 80260.82, 79905.92, 81404.68, 80969.8, 82960.61, 
    88937.89,
  88323.19, 87023.09, 88278.19, 87429.59, 87391.21, 85783.85, 84765.34, 
    84316.01, 83353.09, 85354.36, 100386.5, 101242.5, 91263.98, 91531.2, 
    84086.13,
  88385.76, 86575.14, 89074.27, 90021.68, 89201.11, 88777.8, 88061.3, 
    88463.82, 90022.24, 101091.5, 102113, 102146, 101933.4, 93763.39, 78397.71,
  87456.04, 86701.06, 88858.12, 90231.54, 90041.69, 90150.3, 90082.38, 
    92097.22, 96085.1, 101856.6, 101830.3, 102002.4, 101906.6, 87605.29, 
    77999.56,
  91221.91, 87950.54, 88424.44, 90295.98, 90007.67, 89015.8, 89650.51, 
    91555.46, 95783.69, 101709.3, 101691.9, 101887.8, 101754.4, 86360.69, 
    87700.86,
  94242.91, 89867.89, 88962.66, 90074.8, 89312.1, 86926.8, 88243.75, 
    90816.59, 101075.4, 101643.4, 101566.2, 101659.5, 101614.1, 93768.12, 
    96185.42,
  97461.22, 92750.79, 91094.76, 93536.92, 93826.66, 93966.7, 94909.93, 
    100965.1, 101567, 101507.7, 101486.7, 101499, 101496.9, 99213.27, 100290.9,
  102019.7, 101705.7, 97816.3, 95355.1, 95390.13, 94411.27, 92043.67, 
    92571.69, 86541.18, 81721.86, 79301.35, 79605.14, 82512.49, 81104.91, 
    91333.54,
  101959.2, 101986.6, 99741.37, 94491.32, 91725.24, 89850.69, 88604.95, 
    88954.66, 83893.2, 81047.66, 80176.41, 80851.45, 83044.8, 81943.48, 
    92870.12,
  92816.25, 89234.46, 94264.1, 92962.81, 86344.89, 85237.98, 87611.85, 
    86950.91, 81874.99, 79554.32, 78560.04, 79247.01, 80598.61, 82175.85, 
    94903.92,
  86584.61, 86590.26, 85790.66, 84094.92, 83826.23, 82331.38, 83232.08, 
    83602.82, 81237.1, 79959.83, 79578, 81102.11, 80687.95, 82708.84, 88737.02,
  88161.89, 87045.41, 88170.68, 87339.38, 87203.74, 85579.8, 84528.28, 
    84063.47, 83091.28, 85103.45, 100300, 101067.3, 91065.42, 91348.08, 
    83835.26,
  88388.16, 86548.04, 89017.12, 89921.86, 89015.29, 88566.53, 87826.29, 
    88235.12, 89835, 100985.3, 101989.9, 102026.3, 101740.8, 93560.23, 
    78134.27,
  87495.68, 86741.83, 88836.88, 90161.31, 89923.4, 89962.12, 89871.48, 
    91879.37, 95882.34, 101707.2, 101684.6, 101870.8, 101781, 87371.28, 
    77808.05,
  91232.83, 87957.15, 88359.91, 90226.45, 89894.79, 88866.51, 89474.29, 
    91356.74, 95606.46, 101593.2, 101581, 101767.4, 101680.3, 86053.66, 
    87792.38,
  94203.25, 89823.99, 88862.76, 90002.48, 89191.14, 86790.43, 88067.96, 
    90686.36, 100945, 101538.8, 101496.3, 101601.3, 101615.6, 93684.28, 
    96335.27,
  97359.37, 92637.62, 90967, 93392.87, 93675.07, 93817.83, 94740.23, 
    100794.5, 101424.6, 101441.1, 101469.8, 101513.5, 101570.2, 99276.15, 
    100465.9,
  102711.2, 102348.8, 98352.92, 95776.52, 95769.38, 94702.88, 92230.26, 
    92790.06, 86658.16, 81843.12, 79385.63, 79649.56, 82544.15, 81066.14, 
    91404.8,
  102685.5, 102636.2, 100399.6, 95077.95, 92128.88, 90156.49, 88906.48, 
    89183.26, 84033.72, 81212.76, 80334.89, 80986.95, 83130.52, 81909.53, 
    92907.33,
  93327.73, 89780.59, 94774.63, 93389.5, 86709.93, 85571.25, 87887.54, 
    87141.9, 82073.2, 79712.58, 78588.05, 79256.46, 80614.27, 82190.21, 
    94990.01,
  87157.9, 87265.09, 86338.01, 84592.62, 84284.69, 82747.37, 83562.25, 
    83865.97, 81458.76, 80069.98, 79808.99, 81376.67, 80723.38, 82801.62, 
    88795.35,
  88771.16, 87686.89, 88732.3, 87894.55, 87682.9, 86034.1, 84909.83, 
    84386.35, 83320.71, 85452.38, 100656.6, 101297.9, 91296.04, 91576.08, 
    83800.85,
  89029.44, 87171.72, 89618.3, 90458.69, 89506.72, 89031.16, 88240.55, 
    88628.73, 90206.22, 101362.4, 102286.1, 102307.7, 102047.2, 93733.66, 
    78109.37,
  88112.02, 87340.45, 89422.91, 90691.7, 90435.2, 90412.27, 90294.9, 
    92257.17, 96257.01, 102106.9, 102089.4, 102121.1, 102077, 87444.38, 
    77847.65,
  91875.02, 88565.68, 88964.09, 90781.21, 90422.89, 89343.53, 89929.81, 
    91728.62, 96078.01, 102051.8, 102039.9, 102096.4, 101996.9, 86135.28, 
    88002.48,
  94838.6, 90446.73, 89476.27, 90579.31, 89724, 87288.58, 88526.44, 91181.53, 
    101496.3, 102019.6, 101975.3, 102004.4, 101941.1, 93949.52, 96499.84,
  98004.79, 93297.55, 91624.09, 94018.43, 94261.77, 94435.49, 95353.2, 
    101387, 101957.3, 101950.1, 101936.7, 101951.2, 101927.3, 99569.59, 
    100680.5,
  102566.2, 102216.1, 98192.67, 95614.02, 95593.33, 94531.5, 92081.19, 
    92626.5, 86579.88, 81754.35, 79314.48, 79560.75, 82484.68, 81040.32, 
    91374.25,
  102435.8, 102378.5, 100136.6, 94856.54, 91964.55, 90003.33, 88721.27, 
    88994.26, 83914.16, 81080.91, 80205.45, 80844.11, 83022.2, 81842.84, 
    92816.99,
  93259.28, 89571.27, 94524.21, 93213.5, 86548.98, 85419.85, 87697.46, 
    86963.45, 81942.62, 79592.05, 78503.13, 79144.94, 80495.54, 82068.85, 
    94845.07,
  87056.52, 87014.67, 86147.59, 84432.25, 84112.04, 82581.66, 83403.07, 
    83706.51, 81313.77, 79939.75, 79642.3, 81193.42, 80581.43, 82614.09, 
    88617.84,
  88649.2, 87462.35, 88515.58, 87680.69, 87493.83, 85857.83, 84750.12, 
    84217.91, 83168.61, 85249.67, 100230.9, 100856.8, 90985.01, 91278.41, 
    83610.7,
  88799.27, 86931.73, 89370.05, 90248.19, 89304.55, 88821.55, 88033.4, 
    88402.15, 89938.37, 100875.1, 101735.3, 101786.8, 101576.9, 93399.62, 
    77957.82,
  87885.73, 87112.58, 89183.2, 90458.12, 90200.92, 90183.48, 90051.12, 
    91986.07, 95888.08, 101580.8, 101532.1, 101598.1, 101601.3, 87156.94, 
    77649.44,
  91608.98, 88323.78, 88697.76, 90526.94, 90177.51, 89091.2, 89644.63, 
    91411.52, 95619.82, 101454.6, 101427.8, 101506.2, 101453.6, 85809.84, 
    87657.48,
  94584.26, 90214.01, 89175.16, 90277.18, 89441.7, 86999.88, 88213.2, 
    90770.29, 100886.9, 101363.3, 101324.8, 101358.6, 101314.5, 93452.11, 
    95934.73,
  97725.96, 93010.81, 91282.64, 93641.55, 93876.98, 94009.52, 94864.17, 
    100754.9, 101295.3, 101267.8, 101232.8, 101211.4, 101190.7, 98897.28, 
    100025.5,
  101683, 101333.2, 97352.77, 94728.16, 94681.43, 93641.9, 91253.42, 
    91773.16, 85860.14, 81024.42, 78600.12, 78844.32, 81663.99, 80254.95, 
    90281.84,
  101582.3, 101453.2, 99199.74, 93961.31, 91098.68, 89144.12, 87864, 
    88152.28, 83151.71, 80296.71, 79434.52, 80039.93, 82178.73, 81054.68, 
    91705.01,
  92435.84, 88781.62, 93676.38, 92353.05, 85759.09, 84595.24, 86873.4, 
    86154.54, 81147.8, 78818.15, 77798.48, 78409.39, 79725.19, 81234.9, 
    93714.93,
  86310.85, 86352.06, 85432.54, 83676.41, 83365.43, 81832.1, 82610.97, 
    82894.48, 80522.88, 79192.05, 78808.89, 80320.19, 79802.2, 81746.25, 
    87677.1,
  87878.01, 86817.38, 87819.53, 86977.25, 86769.56, 85101.68, 83979.96, 
    83443.75, 82386.67, 84394.64, 99457.6, 100139.3, 90152.99, 90353.55, 
    82796.88,
  88197.59, 86347.6, 88740.29, 89576.12, 88596.34, 88110.99, 87300.34, 
    87644.02, 89158.96, 100183.1, 101022.6, 100982.9, 100701.6, 92459.06, 
    77144.21,
  87365.59, 86568.27, 88606.19, 89847.14, 89555.3, 89517.27, 89359.92, 
    91287.87, 95203.48, 100930.6, 100802.8, 100806.7, 100676.8, 86291.16, 
    76794.79,
  91171.84, 87827.7, 88187.07, 89985.05, 89585.9, 88481.85, 89026.26, 
    90769.12, 95039.46, 100855.9, 100734.1, 100725.1, 100538.2, 84964.64, 
    86674.4,
  94197.95, 89770.71, 88774.88, 89839.68, 88931.14, 86468.8, 87665.9, 
    90263.83, 100452.1, 100832.3, 100663.6, 100598.2, 100447.9, 92508.66, 
    95025.81,
  97419.21, 92701.72, 91005.48, 93355.08, 93570.12, 93705.05, 94536.03, 
    100505.3, 100907.7, 100769.5, 100627, 100532.1, 100412.2, 98053.6, 99136.7,
  101370.9, 101028.8, 97059.93, 94512.15, 94520.78, 93498.12, 91108.25, 
    91621.95, 85678.68, 80888.47, 78461.23, 78752.13, 81622.02, 80234.4, 
    90490.84,
  101319.1, 101233.4, 98981.48, 93771.1, 90956.09, 89020.27, 87768.22, 
    88078.26, 83027.61, 80207, 79372.13, 80029.37, 82206.11, 81044.95, 
    91981.56,
  92170.92, 88591.45, 93561.98, 92220, 85629.79, 84528.5, 86845.3, 86116.2, 
    81083.38, 78775.41, 77731.18, 78384.77, 79761.82, 81314.9, 94120.44,
  86018.4, 86106.97, 85198.07, 83480.01, 83209.61, 81716.83, 82560.16, 
    82867.41, 80498.93, 79141.73, 78803.61, 80424.56, 79869.75, 81957.7, 
    87940.09,
  87602.48, 86578.51, 87651.55, 86830.18, 86663.14, 85040.27, 83960.52, 
    83447.65, 82404, 84511.48, 99977.1, 100602.5, 90484.39, 90751.85, 82971.72,
  87932.59, 86112.4, 88600.8, 89477.22, 88545.01, 88094.2, 87327.97, 
    87727.79, 89342.55, 100745, 101646.6, 101626.2, 101329, 92946.49, 77253.31,
  87071.8, 86311.42, 88456.92, 89755.09, 89503.95, 89531.63, 89456.92, 
    91490.66, 95596.8, 101560.5, 101471.7, 101516.9, 101388, 86646.66, 
    76956.62,
  90835.83, 87552.35, 88008.45, 89870.43, 89540.38, 88530.41, 89153.81, 
    91005.32, 95435.04, 101517.8, 101459.5, 101541.9, 101359.1, 85353.26, 
    87170.08,
  93807.46, 89471.77, 88550.09, 89672.75, 88857.04, 86468.88, 87751.08, 
    90469.23, 100971.2, 101522.8, 101441.2, 101486.2, 101366.4, 93198.03, 
    95847.66,
  96963.26, 92319.72, 90705.34, 93159.12, 93452.86, 93675.52, 94635.06, 
    100825, 101448.5, 101474.6, 101435.3, 101472.7, 101455.5, 99106.46, 
    100301.5,
  101111.8, 100806.9, 96934.14, 94446.65, 94467.26, 93487.09, 91151.97, 
    91688.83, 85810.83, 81030.62, 78660.09, 78947.8, 81904.44, 80535.66, 
    90847.04,
  100815.4, 100895.6, 98682.76, 93531.64, 90797.12, 88945.4, 87693.9, 
    88065.84, 83127.71, 80304.51, 79491.2, 80157.83, 82397.2, 81318.6, 92255.7,
  91858.09, 88229.02, 93178.29, 91954.3, 85399.1, 84314.23, 86653.92, 
    86042.01, 81076.87, 78784.84, 77836.74, 78520.24, 79927.15, 81508.61, 
    94285.25,
  85594.88, 85454.59, 84733.65, 83109.78, 82828.88, 81398.72, 82303.53, 
    82688.46, 80366.7, 79127.95, 78783.95, 80331.73, 79925.6, 81964.08, 
    88103.29,
  87081.4, 85878.9, 87024.23, 86211.61, 86115.35, 84537.53, 83522.75, 
    83097.74, 82143.16, 84116.42, 99108.14, 99987.87, 90169.95, 90564.78, 
    83097.8,
  87101.73, 85329.98, 87775.38, 88718.61, 87868.66, 87445.88, 86736.31, 
    87158.09, 88719.57, 99742.08, 100844.2, 100902.8, 100758.5, 92714.05, 
    77428.8,
  86135.67, 85419.44, 87532.28, 88889.02, 88698.39, 88778.72, 88712.22, 
    90719.92, 94723.75, 100512.6, 100613.1, 100775.9, 100808.4, 86529.03, 
    77059.92,
  89749.77, 86583.17, 87020.99, 88888.5, 88623.24, 87654.87, 88273.3, 
    90168.49, 94413.34, 100388.1, 100513, 100716, 100697.3, 85189.18, 86992.78,
  92615, 88367.37, 87447.12, 88579.07, 87862.36, 85545.58, 86833.6, 89402.34, 
    99551.09, 100281.9, 100335.7, 100525.5, 100590.5, 92742.53, 95404.46,
  95675.99, 91072.53, 89460.87, 91848.1, 92172.95, 92317.54, 93269.54, 
    99284.98, 100003.5, 100086.6, 100207.7, 100374.6, 100531.3, 98339.62, 
    99690.76,
  100626.6, 100288.4, 96512.05, 94055.66, 94074.85, 93149.83, 90905.5, 
    91415.37, 85682.12, 80877, 78557.49, 78825.28, 81744.61, 80433.92, 
    90451.12,
  100234.9, 100326.1, 98163.27, 93056.3, 90394.29, 88584.04, 87356.43, 
    87788.04, 82954.91, 80131.03, 79362.91, 79989.77, 82203.62, 81156.14, 
    91804.48,
  91408.4, 87693.46, 92647.18, 91440.76, 84948.39, 83882.28, 86252.21, 
    85712.55, 80788.52, 78548.52, 77674.45, 78359.26, 79750.24, 81263.62, 
    93753.62,
  85040.95, 84933.6, 84195.18, 82570.83, 82288.36, 80920.36, 81866.59, 
    82273.12, 80010.53, 78878.26, 78534.47, 80025.43, 79697.36, 81693.23, 
    87730.69,
  86488.02, 85394.58, 86495.72, 85647.42, 85537.98, 83965.71, 82994.27, 
    82611.55, 81736.98, 83584.84, 98177.09, 99282.89, 89720.91, 90132.3, 
    82848.52,
  86648.13, 84845.05, 87297.36, 88207.63, 87314.76, 86863.07, 86153.96, 
    86570.88, 88112.77, 98963.75, 100227.8, 100207.1, 100195.1, 92273.32, 
    77220.04,
  85852.99, 85062.76, 87151.26, 88455.38, 88179.34, 88227.13, 88132.48, 
    90184.77, 94248.66, 99980.12, 99912.12, 100030, 100168.7, 86190.41, 
    76753.8,
  89667.01, 86317.12, 86746.92, 88578.63, 88196.46, 87174.81, 87771.53, 
    89738.67, 94054.34, 99936.98, 99892.34, 100017.8, 99934.88, 84792.23, 
    86288.67,
  92779.22, 88305.36, 87378.27, 88499.08, 87640.11, 85248.01, 86542.52, 
    89212.23, 99481.62, 100038.6, 99894.02, 99895.11, 99816.81, 92031.8, 
    94547.07,
  96128.74, 91347.09, 89731.83, 92190.27, 92455.21, 92551.57, 93478.89, 
    99622.35, 100151.6, 99998.87, 99892.09, 99869.19, 99849.27, 97521.44, 
    98649.88,
  101395.5, 100976.8, 96942.62, 94271.46, 94165.33, 93064.95, 90633.69, 
    91104.27, 85171.29, 80329.97, 77979.66, 78300.82, 81183.39, 79833.21, 
    89840.16,
  101456.8, 101221.9, 98939.95, 93563.97, 90573.96, 88568.9, 87242.55, 
    87515.63, 82453.5, 79580.39, 78780.77, 79473.84, 81669.88, 80629.91, 
    91226.14,
  91961.91, 88435.41, 93366.32, 91911.07, 85149.59, 83974.29, 86290.46, 
    85552.95, 80444.92, 78121.47, 77208.31, 77894.52, 79275.37, 80799.12, 
    93283.72,
  85869.93, 86004.2, 84985.57, 83186.01, 82830.75, 81211.95, 82011.78, 
    82275.41, 79835.97, 78538.95, 78249.25, 79746.37, 79353.6, 81343.62, 
    87332.2,
  87558.37, 86470.95, 87525.77, 86673.78, 86410.66, 84678.2, 83495.89, 
    82918.29, 81871.06, 84060.27, 99554.03, 100168.8, 89914.63, 90038.03, 
    82552.91,
  87954.34, 86018.47, 88541.21, 89402.43, 88390.84, 87862.99, 87004.77, 
    87358.47, 89005.23, 100493.3, 101352.5, 101229.2, 100847.8, 92385.45, 
    76911.19,
  87093.13, 86243.09, 88381.48, 89693.61, 89403.86, 89356.31, 89210.38, 
    91257.78, 95368.42, 101292, 101088.9, 101098.2, 100756.5, 86137.54, 
    76418.44,
  90999.15, 87568.95, 87963.71, 89852.27, 89453.52, 88300.71, 88867.39, 
    90716.93, 95143.62, 101236.3, 101116.7, 101186.6, 100842.6, 84943.28, 
    86330.94,
  94062.66, 89555.02, 88530.95, 89667.13, 88747.77, 86229.42, 87458.8, 
    90185.31, 100737.6, 101221, 101059.8, 101055.5, 100878.9, 92674.48, 
    95247.23,
  97319.53, 92534.18, 90826.02, 93272.92, 93509.52, 93668.43, 94534.47, 
    100726.3, 101215.4, 101104, 100994.1, 100950.8, 100904.5, 98495.38, 
    99588.64,
  102056.2, 101743.1, 97740.05, 95175.7, 95162.77, 94145.69, 91724.32, 
    92276.27, 86122, 81211.3, 78681.38, 78902.37, 81778.2, 80319.09, 90663.12,
  101838.8, 101784.5, 99614.72, 94359.1, 91456.3, 89505.52, 88252.77, 
    88584.76, 83403.56, 80492.03, 79571.47, 80193.34, 82348.44, 81156.64, 
    92150.4,
  92694.55, 88970.49, 93866.41, 92622.1, 85957.7, 84749.3, 87102.26, 
    86461.55, 81347.13, 78931.98, 77783.56, 78408.66, 79778.62, 81350.23, 
    94226.69,
  86396.05, 86222.11, 85390.28, 83682.06, 83342.29, 81803.6, 82636.13, 
    83013.88, 80580.18, 79201.77, 78879.24, 80400.92, 79764.59, 81831.23, 
    87950.45,
  87892.31, 86601.7, 87618.48, 86780.53, 86584.98, 84959.23, 83846.84, 
    83355.66, 82321.04, 84365.08, 99352.32, 100240.9, 90248.58, 90539.88, 
    82884.2,
  87889.13, 86009.23, 88364.91, 89261.52, 88313.09, 87842.16, 87042.17, 
    87433.13, 88947.23, 100015.9, 101073.8, 101151.7, 100961.2, 92658.45, 
    77108.38,
  86909.49, 86102.59, 88120.57, 89387.3, 89123.62, 89111.94, 88981.68, 
    90923.75, 94909.15, 100764.8, 100796.5, 100883.6, 100882.7, 86344.24, 
    76667.26,
  90530.38, 87252.05, 87593.33, 89367.71, 89038.79, 87960.66, 88525.63, 
    90317.45, 94611.15, 100574.1, 100623.1, 100767.2, 100682.9, 84953.84, 
    86537.16,
  93400.16, 89049.84, 88028.15, 89112.28, 88296.6, 85841.27, 87036.02, 
    89601.38, 99915.16, 100509.7, 100457.1, 100537.3, 100509.2, 92481.4, 
    94924.46,
  96504.27, 91790.95, 90067.7, 92411.53, 92677.4, 92841.5, 93703.34, 
    99808.31, 100384.6, 100360.8, 100342.3, 100374, 100380.1, 98023.53, 
    99161.98,
  101980.2, 101647.8, 97726.67, 95205.63, 95227.43, 94280.2, 91984.85, 
    92531.95, 86559.26, 81635.45, 79152.15, 79394.16, 82190.45, 80810.04, 
    90731.63,
  101635.4, 101725.3, 99538.05, 94339.57, 91580.21, 89691.42, 88452.13, 
    88845.65, 83788.01, 80841.88, 79959.02, 80536.34, 82670.91, 81574.12, 
    92174.7,
  92700.66, 88996.45, 93944.95, 92673.42, 86126.88, 84946.47, 87334.33, 
    86724.88, 81645.31, 79263.45, 78235.34, 78854.7, 80180.12, 81683.64, 
    94226.31,
  86415.77, 86192.04, 85510.97, 83773.4, 83497.65, 82014.02, 82869.84, 
    83225.28, 80850.43, 79532.9, 79084.93, 80584.2, 80101.51, 82072.87, 
    88155.59,
  87893.84, 86615.33, 87737.65, 86857.23, 86754.62, 85142.74, 84085.96, 
    83608.12, 82568.85, 84452, 99449.61, 100476.8, 90475.24, 90707.98, 
    83227.92,
  87902.14, 86079.79, 88462.07, 89371.87, 88457.77, 88016.8, 87259.82, 
    87645.36, 89177.01, 100323.5, 101501.6, 101376.5, 101098.3, 92889.37, 
    77457.12,
  86908.06, 86134.05, 88238.73, 89540, 89281.62, 89322.22, 89224.13, 
    91210.55, 95337.59, 101362.7, 101295.1, 101410.8, 101256.1, 86649.56, 
    77064.63,
  90536.88, 87283.43, 87735.57, 89528.55, 89222.88, 88202.5, 88825.42, 
    90726.38, 95195.64, 101369.1, 101318.5, 101473.1, 101212.2, 85360.33, 
    87024.43,
  93389.19, 89127.49, 88214.39, 89310.55, 88555.34, 86166.23, 87500.79, 
    90162.09, 100716.3, 101361.1, 101295.4, 101422.1, 101276.7, 93125.42, 
    95671.54,
  96498.73, 91893.43, 90258.91, 92760.82, 93103.8, 93330.13, 94329.9, 
    100630.3, 101254.9, 101294.4, 101332, 101409.1, 101388.2, 98986.34, 
    100199.9,
  101972.8, 101633.4, 97722.78, 95259.41, 95287.3, 94284.74, 91943.3, 
    92484.3, 86557.62, 81693.31, 79265.96, 79517.41, 82364.4, 80995.46, 
    91046.73,
  101839.7, 101856.4, 99680.84, 94461.25, 91665.81, 89790.38, 88558.73, 
    88917.64, 83884.84, 81011.14, 80157.1, 80770.12, 82920.18, 81800.85, 
    92531.26,
  92712.32, 89173.59, 94156.16, 92860.23, 86264.02, 85163.08, 87548.87, 
    86888.87, 81841.49, 79498.62, 78468.71, 79110.68, 80432.66, 81957.73, 
    94562.98,
  86509.6, 86593.31, 85721.95, 84052.13, 83764.16, 82291.2, 83173.3, 
    83543.59, 81144.56, 79838.52, 79479.59, 80967.21, 80445.75, 82458.05, 
    88469.41,
  88066.05, 87022.03, 88069.88, 87240.42, 87084.84, 85478.02, 84413.17, 
    83952.17, 82952.35, 84966.34, 99932.72, 100723.9, 90807.45, 91128.34, 
    83527.41,
  88303.33, 86486.66, 88930.29, 89813.84, 88897.95, 88442.95, 87686.23, 
    88081.91, 89592.43, 100633.7, 101563.7, 101578.6, 101400.4, 93265.8, 
    77801.2,
  87441.3, 86680.75, 88752.03, 90034.7, 89787.56, 89794.53, 89694.2, 
    91660.56, 95613.51, 101421.4, 101422.5, 101470.4, 101418.8, 87021.3, 
    77442.63,
  91201.25, 87913.6, 88319.04, 90134.7, 89799.34, 88750.26, 89328.75, 
    91127.41, 95432.25, 101432.4, 101398.5, 101469.1, 101318, 85605.79, 
    87422.68,
  94218.09, 89821.02, 88836.3, 89927.63, 89103.66, 86703.97, 87943.86, 
    90564.75, 100860.5, 101465.3, 101387.9, 101450.4, 101292.6, 93325.33, 
    96005.25,
  97437.12, 92698.01, 91015.45, 93392.45, 93637.59, 93784.02, 94686.27, 
    100779.6, 101404.9, 101440.2, 101430.7, 101483.5, 101458.9, 99130.59, 
    100363.6,
  102588, 102282.7, 98422.82, 95919.98, 95926.59, 94863.75, 92438.74, 
    92978.23, 86930.51, 82151.58, 79771.55, 80054.95, 82986.43, 81536.77, 
    91861.27,
  102443.2, 102511.2, 100253.1, 95020.5, 92235.77, 90317.88, 89097, 89414.15, 
    84320.81, 81483.87, 80636.48, 81300.35, 83501.95, 82350.81, 93320.51,
  93344.37, 89777.49, 94819.61, 93471.3, 86850.28, 85696.37, 88061.88, 
    87372.98, 82346.53, 80007.4, 78978.14, 79644.11, 81018.02, 82593.55, 
    95376.78,
  87073.05, 86951.34, 86203.08, 84556.11, 84272.44, 82790.08, 83691.77, 
    84044.59, 81687.12, 80352.88, 80032.7, 81579.9, 81061.58, 83099.54, 
    89147.77,
  88743.38, 87392.7, 88539.34, 87688.21, 87571.44, 85961.02, 84931.95, 
    84475.39, 83484.62, 85511.55, 100449.4, 101202.2, 91369.9, 91726.22, 
    84166.51,
  88792.88, 86898.06, 89373.41, 90261.99, 89384.67, 88923.99, 88183.16, 
    88568.88, 90123.96, 101069, 102050.5, 102139.2, 101916.3, 93826.18, 
    78514.44,
  87720.41, 86992.76, 89131.48, 90463.8, 90264.54, 90296.39, 90182.09, 
    92125.66, 96054.49, 101782.1, 101786.4, 101975.9, 101932.3, 87662.2, 
    78169.44,
  91396.53, 88172.3, 88617.27, 90473.59, 90194.8, 89176.98, 89733.09, 
    91572.5, 95743.84, 101598.3, 101628, 101852.7, 101755.3, 86357.06, 
    87922.26,
  94317.59, 90033.54, 89066.51, 90167.52, 89421.83, 87062.65, 88288.49, 
    90819.95, 100841.5, 101528.5, 101472.8, 101605.1, 101597.3, 93751.36, 
    96080.11,
  97426.27, 92760.71, 91063.9, 93432.46, 93710.76, 93820.8, 94705.55, 
    100645.1, 101339.1, 101352.5, 101361, 101410.1, 101454.2, 99155.74, 
    100189.8,
  102021.6, 101670.1, 97822.08, 95413.16, 95449.81, 94441.74, 92102.55, 
    92574.04, 86644.12, 81879.77, 79503.08, 79802.65, 82665.76, 81310.3, 
    91379.5,
  101923.9, 101994.8, 99683.45, 94481.7, 91781.73, 89907.55, 88688.28, 
    89033.61, 84038.66, 81193.91, 80344.01, 81001.27, 83157.93, 82096.91, 
    92830.13,
  92824.48, 89278.18, 94349.78, 92994.26, 86444.82, 85300.17, 87701.9, 
    87044.16, 82028.42, 79710.57, 78760.83, 79420.73, 80761.2, 82307.59, 
    94883.28,
  86645.08, 86513.86, 85814.2, 84139.28, 83871.66, 82399.77, 83336.04, 
    83694.86, 81381.46, 80090.24, 79717.56, 81178.91, 80798.48, 82766.37, 
    88761.52,
  88286, 86965.95, 88184.86, 87306.1, 87211.06, 85579.27, 84569.13, 84144.05, 
    83185.12, 85188.84, 100165.2, 101017.9, 91062.59, 91328.24, 83924.16,
  88329.01, 86493.72, 89042.97, 89914.77, 89054.2, 88587.06, 87869.56, 
    88266.81, 89867.12, 100914, 101883.8, 101888.8, 101665.8, 93499.62, 
    78273.68,
  87339.33, 86604.12, 88782.11, 90119.31, 89911.49, 89960.86, 89867.91, 
    91858.38, 95889.95, 101610.9, 101580.1, 101740.8, 101650.2, 87417.06, 
    77831.13,
  91079.37, 87827.48, 88311.47, 90183.86, 89870.06, 88874.12, 89464.81, 
    91363.2, 95588.42, 101512, 101504.7, 101684.1, 101525, 86138.51, 87515.36,
  93993.14, 89677.4, 88783.32, 89902.68, 89155.43, 86786.58, 88071.05, 
    90669.35, 100894.7, 101523.9, 101428.1, 101520.8, 101460.1, 93563.18, 
    96006.23,
  97157.3, 92505.57, 90866.55, 93298.18, 93593.27, 93723.07, 94669.67, 
    100757.8, 101406.8, 101356.7, 101340, 101343.5, 101353.1, 99026.38, 
    100100.6,
  101320.4, 100956, 97123.36, 94670.62, 94715.55, 93775.21, 91547.99, 
    92037.13, 86222.05, 81455.88, 79113.11, 79422.81, 82327.62, 80989.62, 
    91122.73,
  100999, 101142, 98926.9, 93727.5, 91070.55, 89257.84, 88047.26, 88457.17, 
    83570.11, 80758.02, 79951.42, 80646.17, 82846.34, 81805.19, 92585.95,
  92066.61, 88472.11, 93471.94, 92182.48, 85656.74, 84607.57, 86987.84, 
    86425.47, 81461.09, 79213.75, 78299.53, 79019.52, 80413.34, 81976, 
    94596.47,
  85722.34, 85539.58, 84917.16, 83311.18, 83037.34, 81651.1, 82622.36, 
    83006.48, 80727.14, 79546.27, 79205.31, 80740.16, 80431.49, 82426.38, 
    88501.89,
  87172.7, 85963.1, 87148.12, 86266.24, 86230.68, 84671.88, 83717.19, 
    83355.95, 82487.54, 84420.7, 99267.12, 100303.7, 90497.06, 90895.88, 
    83594.7,
  87205.46, 85386.97, 87892.59, 88851.49, 88004.05, 87568.98, 86899.05, 
    87342.53, 88938.34, 99890.1, 101079.2, 101176.1, 101049.6, 93075.82, 
    77921.48,
  86175.23, 85441.51, 87613.76, 88993.85, 88796.73, 88904.35, 88866.95, 
    90871.86, 94942.54, 100687.5, 100780.1, 101047.9, 101056, 86941.73, 
    77529.05,
  89869.85, 86610.16, 87073.07, 88989.08, 88709.88, 87758.86, 88401.63, 
    90343.73, 94589.24, 100528, 100703.1, 100945.1, 100914.9, 85670.66, 
    87248.86,
  92774.36, 88439.4, 87539.48, 88697.66, 87979.08, 85660.68, 87000.94, 
    89561.78, 99738.3, 100492.3, 100523.2, 100723.2, 100793.1, 93023.12, 
    95653.61,
  95900.2, 91200.29, 89559.56, 92022.94, 92330.47, 92462.4, 93463.53, 
    99511.59, 100288.5, 100326.4, 100455.3, 100607.9, 100727.4, 98526.12, 
    99789.72,
  101820.4, 101429.5, 97442.3, 94843.42, 94810.71, 93797.98, 91469.19, 
    91947.6, 86094.17, 81182.48, 78831.37, 79080.12, 82003.6, 80678.27, 
    90760.85,
  101601.5, 101609.1, 99305.25, 93980.19, 91151.38, 89232.51, 87953.69, 
    88299.25, 83335.51, 80409.59, 79634.05, 80276.99, 82496.14, 81446.91, 
    92203.13,
  92383.81, 88654.72, 93661.69, 92344.93, 85671.91, 84523.07, 86876.09, 
    86242.58, 81196.35, 78872.81, 77975.1, 78616.18, 80039.85, 81573.97, 
    94223.9,
  86063.64, 85971.33, 85216.7, 83416.38, 83101.15, 81607.52, 82471.23, 
    82804.91, 80463.32, 79213.42, 78847.8, 80377.95, 80032.77, 82011.68, 
    88093.52,
  87664.51, 86392.53, 87576.38, 86672.34, 86545.09, 84868.74, 83783.59, 
    83305.55, 82341.19, 84276.74, 99539.66, 100371.4, 90358.19, 90609.88, 
    83183.8,
  87796.84, 85915.24, 88413.28, 89301.23, 88360.16, 87863.81, 87090.42, 
    87498.45, 89066.61, 100409.3, 101442.4, 101294.5, 101067.6, 92833.45, 
    77494.77,
  86798.82, 86004.37, 88173.19, 89523.15, 89260.54, 89285.71, 89160.51, 
    91189.47, 95300.06, 101202.8, 101117.4, 101216.6, 101093.5, 86611.07, 
    77024.42,
  90562.28, 87254.17, 87675.59, 89577.45, 89230.33, 88168.26, 88754.05, 
    90663.31, 95026.52, 101181.1, 101146.9, 101245.9, 101018.1, 85262.14, 
    86830.83,
  93528.73, 89116.24, 88135.89, 89307.65, 88476.28, 86028.21, 87330.09, 
    90028.88, 100596.4, 101202.1, 101056.3, 101086.7, 101000.1, 92919.8, 
    95445.73,
  96766.61, 92000.5, 90307.09, 92810.42, 93123.9, 93310.94, 94280.77, 
    100563.4, 101174.5, 101073.8, 100998.6, 100958.1, 100897.4, 98485.87, 
    99560.41,
  101733.1, 101375.1, 97530.58, 95129.59, 95175.38, 94198.26, 91921.88, 
    92400.09, 86553.82, 81714.84, 79355.87, 79640.88, 82570.41, 81277.06, 
    91475.8,
  101496.5, 101642.9, 99372.35, 94174.94, 91510.19, 89678.95, 88443.23, 
    88826.75, 83870.77, 81022.08, 80193.93, 80871.16, 83105.72, 82073.62, 
    92920.94,
  92476.21, 88937.41, 93965.83, 92638.29, 86095.96, 84971.71, 87387.1, 
    86788.03, 81733, 79449.7, 78518.92, 79248.27, 80644.84, 82192.38, 94957.71,
  86107.05, 86022.02, 85372.16, 83723.54, 83443.5, 82029.19, 82976.78, 
    83353.79, 81007.19, 79837.19, 79441.46, 80947.54, 80600.32, 82619.37, 
    88770.74,
  87666.1, 86438.19, 87630.18, 86744.59, 86700.34, 85113.33, 84116.77, 
    83730.17, 82781.77, 84675.81, 99718.95, 100783.5, 90897.94, 91199.95, 
    83805.65,
  87743.55, 85957.82, 88416.64, 89396.23, 88548.66, 88109.59, 87396.96, 
    87823.02, 89411.31, 100595.1, 101756.8, 101720.5, 101609.1, 93387.55, 
    78154.58,
  86770.37, 86023.52, 88199.26, 89586.6, 89360.87, 89470.08, 89410.37, 
    91462.42, 95621.19, 101435.8, 101440.4, 101585.3, 101519.1, 87206.28, 
    77616.72,
  90574.48, 87258.59, 87789.61, 89717.34, 89381.22, 88393.62, 88978.45, 
    90973.13, 95333.96, 101399.5, 101438.2, 101622.9, 101445.1, 85797.41, 
    87322.78,
  93693.05, 89222.45, 88342.59, 89499.23, 88704.48, 86290.73, 87586.19, 
    90260.18, 100674.5, 101362.7, 101307, 101463.6, 101447.7, 93355.97, 
    95918.59,
  96973.98, 92202.01, 90592.7, 93105.19, 93419.34, 93475.54, 94445.27, 
    100628.5, 101370.8, 101303, 101307.5, 101342.7, 101359.5, 99008.11, 
    100185.4,
  101146.7, 100753.9, 96910.13, 94415.91, 94433.33, 93453.86, 91221.86, 
    91673.86, 85966.33, 81129.3, 78868.46, 79123.21, 82088.97, 80792.62, 
    90916.7,
  100780.6, 100881.2, 98696.34, 93502.18, 90812.42, 88971.05, 87735.24, 
    88127.38, 83296.01, 80440.67, 79681.8, 80318.45, 82598.02, 81590.31, 
    92340.02,
  91866.67, 88198.26, 93194.13, 91914.27, 85368.62, 84276.26, 86690.47, 
    86097.7, 81154.13, 78895.23, 78042.24, 78724.12, 80166.91, 81702.6, 
    94301.34,
  85432.88, 85293.95, 84653.79, 83041.49, 82728.17, 81356.2, 82300.39, 
    82683.57, 80392.8, 79251.22, 78887.06, 80352.98, 80110.09, 82167.34, 
    88298.35,
  86889.52, 85754.4, 86929.59, 86027.8, 85976.83, 84409.39, 83410.78, 
    83067.96, 82163.54, 84037.74, 98875.1, 99940.12, 90232.43, 90624.89, 
    83349.16,
  86952.65, 85232.19, 87696.61, 88659.45, 87805.13, 87361.84, 86652.53, 
    87099.1, 88682.65, 99809.55, 100951.2, 100921.4, 100830.2, 92810.91, 
    77773.3,
  86067.41, 85337.84, 87497.44, 88858.02, 88617.5, 88741.7, 88696.41, 
    90761.7, 94890.4, 100717, 100646.7, 100803.9, 100748.3, 86674.47, 77238.73,
  89913.11, 86575.24, 87080.3, 88955.25, 88610.25, 87620.51, 88245.73, 
    90244.62, 94581.72, 100655, 100646.9, 100854.6, 100615.1, 85372.62, 
    86948.69,
  93021.43, 88562.59, 87666.31, 88792.43, 88003.79, 85635.93, 86956.66, 
    89633.73, 100024.9, 100665.9, 100587.4, 100729.6, 100651, 92824.73, 
    95497.01,
  96382.83, 91533.39, 89940.45, 92414.94, 92658.2, 92735.02, 93736.52, 
    99933.15, 100679.4, 100684.7, 100709.7, 100770, 100783.7, 98539.5, 
    99862.41,
  100858.1, 100470.5, 96517.47, 93951.55, 93922.2, 92913.04, 90580.21, 
    91063.41, 85175.28, 80333.02, 77993.55, 78288.62, 81187.36, 79818.34, 
    89907.59,
  100614, 100634.5, 98332.45, 93053.89, 90266.23, 88386.95, 87101.83, 
    87451.11, 82489.77, 79611.1, 78840.7, 79508.23, 81699.83, 80637.94, 
    91369.86,
  91519.63, 87753.46, 92786.09, 91475.28, 84822.77, 83706.11, 86076.89, 
    85420.34, 80397.58, 78105.5, 77246.42, 77925.23, 79295.45, 80857.05, 
    93374.97,
  85174.88, 85132.83, 84372.63, 82610.86, 82329.48, 80867.84, 81755.63, 
    82101.55, 79744.46, 78533.04, 78198.67, 79699.93, 79339.73, 81357.74, 
    87322.04,
  86795.83, 85660.6, 86817.05, 85926.6, 85825.76, 84158.3, 83097.23, 
    82625.55, 81660.61, 83709.34, 99083.35, 99777.26, 89724.55, 89981.09, 
    82509.35,
  87124.09, 85247.43, 87790.39, 88649.79, 87704.03, 87235.77, 86476.91, 
    86905.46, 88605.99, 100010, 100878.4, 100703.8, 100465, 92203.11, 76867.2,
  86304.01, 85504.65, 87709.64, 89029.64, 88722.91, 88730.59, 88640.36, 
    90816.12, 95012.86, 100883.5, 100674.2, 100631.3, 100430.9, 85980.12, 
    76465.26,
  90238.3, 86846.61, 87343.1, 89239.15, 88854.92, 87781.88, 88419.49, 
    90409.23, 94893.62, 100913.8, 100753.3, 100738.3, 100393.1, 84704.34, 
    86324.53,
  93407.34, 88888.9, 87973.23, 89108.45, 88226.17, 85769.57, 87139.1, 
    89972.03, 100614.4, 101018.5, 100810.1, 100722, 100507.5, 92337.62, 
    94997.09,
  96785.35, 91947.87, 90329, 92899.79, 93157.12, 93249.11, 94314.84, 
    100646.1, 101167.4, 101081.7, 100968.5, 100850.4, 100703.5, 98234.85, 
    99357.71,
  101049.8, 100666.2, 96699.11, 94107.07, 94095.43, 93094.45, 90759.09, 
    91275.42, 85373.83, 80474.13, 78106.76, 78461.23, 81421.29, 80062.58, 
    90328.65,
  100909.5, 100916.8, 98595.48, 93212.96, 90384.62, 88499.91, 87223.62, 
    87588.64, 82602.01, 79727.55, 78955.16, 79661.73, 81911.16, 80854.47, 
    91776.1,
  91736.04, 87955.65, 93070.15, 91681.52, 84982.01, 83823.77, 86177.47, 
    85529.33, 80481.85, 78193.02, 77308.05, 78027.13, 79450.86, 81049.62, 
    93900.12,
  85425.84, 85366.97, 84592.86, 82768.03, 82467.56, 80970.53, 81858.63, 
    82210.52, 79848.4, 78638.73, 78315.65, 79884.27, 79541.93, 81590.11, 
    87745.64,
  87070.47, 85897.38, 87088.34, 86160.11, 86032.3, 84336.02, 83262.87, 
    82801.91, 81836.66, 83998.76, 99648.8, 100418.2, 90096.68, 90385.34, 
    82772.98,
  87391.37, 85520.8, 88125.77, 88952.97, 87988.09, 87502.16, 86767.52, 
    87217.62, 89005.69, 100642.6, 101559.9, 101415.3, 101081.9, 92661.8, 
    76976.2,
  86556.34, 85767.37, 88050.35, 89401.97, 89130.09, 89204.21, 89135.47, 
    91313.41, 95554.84, 101530.9, 101381.1, 101433, 101185.9, 86334.51, 
    76648.8,
  90552.26, 87131.08, 87668.87, 89582.09, 89223.92, 88165.36, 88841, 
    90867.53, 95395.98, 101626.4, 101533.3, 101602.5, 101300.4, 85104.62, 
    86906.9,
  93744.98, 89233.39, 88329.52, 89527.07, 88658.3, 86160.75, 87559.77, 
    90387.42, 101203.1, 101715, 101611.1, 101634.2, 101466.7, 93178.73, 
    95952.36,
  97189.91, 92347.3, 90707.19, 93288.3, 93521.37, 93623.45, 94700.23, 
    101132.6, 101765.1, 101769.6, 101733.9, 101722.1, 101669.4, 99238.49, 
    100374.2,
  101098.1, 100821.2, 96761.67, 94205.1, 94168.09, 93118.45, 90706.74, 
    91244.92, 85258.07, 80368.41, 77972.82, 78301.34, 81267.44, 79893.45, 
    90282.13,
  101093.5, 101190.9, 98773.3, 93389.59, 90495.27, 88549.51, 87237.22, 
    87571.09, 82490.51, 79599.25, 78790.99, 79491.78, 81750.97, 80679.32, 
    91764.86,
  91800.64, 88152.23, 93318.03, 91830.09, 85094.94, 83925.96, 86296.16, 
    85570.37, 80463.66, 78137.1, 77205.38, 77903.23, 79338.49, 80963.32, 
    93948.89,
  85473.48, 85585.52, 84760.96, 82934.12, 82659.58, 81104.7, 82006.84, 
    82313.84, 79876.01, 78608.23, 78306.27, 79896.16, 79460.94, 81530.44, 
    87729.76,
  87241.93, 86184.74, 87376.98, 86465.59, 86323.59, 84606.41, 83541.66, 
    83062.48, 82027.11, 84287.43, 100147.7, 100728.9, 90270.49, 90513.51, 
    82719.51,
  87638.12, 85758.22, 88400.84, 89272.56, 88305.78, 87851.31, 87107.45, 
    87547.29, 89345.98, 101020.3, 101872, 101784.8, 101449.6, 92805.36, 
    76955.85,
  86811.78, 86034.1, 88324.1, 89664.12, 89416.21, 89500.56, 89437.1, 
    91607.29, 95831.51, 101851.7, 101721.4, 101753.8, 101500.6, 86443.32, 
    76632.98,
  90844.71, 87430.34, 87991.83, 89894.83, 89537.02, 88502.16, 89213.41, 
    91164.91, 95713.13, 101929.3, 101819.4, 101863.2, 101601.2, 85232.99, 
    87030.45,
  94091.39, 89543.5, 88656.31, 89832.55, 88935.34, 86459.66, 87859.34, 
    90680.45, 101522.2, 101943.2, 101824, 101817.7, 101642.8, 93278.85, 
    95973.33,
  97601.31, 92679.38, 91096.13, 93699.01, 93920.14, 94063.23, 95145.91, 
    101529.3, 102021.5, 101989.4, 101906.3, 101868.7, 101771.6, 99323.9, 
    100491.1,
  101161.3, 100784.5, 96656.86, 93958.57, 93862.21, 92691, 90171.18, 
    90668.45, 84646.84, 79900.42, 77572.14, 77988, 81043.65, 79680.55, 
    90453.61,
  101387, 101184.3, 98758.41, 93302.08, 90328.38, 88291.2, 86970.87, 
    87234.69, 82078.34, 79335.55, 78547.38, 79323.73, 81622.42, 80505.05, 
    92011.68,
  91848.48, 88225.59, 93354.48, 91767.35, 84951.7, 83857.37, 86189.42, 
    85361.19, 80257.62, 78011.66, 77054.27, 77839.95, 79276.98, 80977.53, 
    94169.7,
  85721.48, 85841.33, 84801.91, 83046.59, 82716.2, 81120.18, 82005.95, 
    82302.38, 79847.34, 78532.15, 78291.71, 79921.12, 79391.23, 81545.95, 
    87704.8,
  87461.86, 86478.56, 87559.23, 86652.83, 86465.73, 84711.6, 83598.38, 
    83044.18, 81980.72, 84339.35, 100205, 100726, 90313.12, 90643.3, 82618.18,
  87905.2, 86041.91, 88685.69, 89515.23, 88553.39, 88042.93, 87259.8, 
    87638.17, 89404.6, 100968.5, 101751.6, 101670.4, 101458.3, 92822.05, 
    76766.4,
  87205.24, 86379.16, 88632.24, 89939.71, 89707.91, 89670.66, 89613.77, 
    91660.8, 95834, 101746.5, 101705.1, 101629.5, 101598.1, 86328.86, 76572.66,
  91284.69, 87800.73, 88286.41, 90205.29, 89812.71, 88669.95, 89284.62, 
    91111.28, 95711.57, 101781.7, 101685.9, 101652.6, 101507.5, 85073.02, 
    87046.54,
  94611.73, 89935.28, 88965.7, 90132.43, 89173.48, 86626.54, 87893.99, 
    90744.48, 101353.4, 101764.8, 101633.8, 101634.4, 101499.8, 93147.13, 
    95810.78,
  98125.12, 93099.08, 91423.82, 93916.67, 94139.67, 94260.77, 95168.13, 
    101352.3, 101827.6, 101753.7, 101618.6, 101580.1, 101496.5, 99093.38, 
    100225.3,
  101916.3, 101568.9, 97390.68, 94663.97, 94569.32, 93411.63, 90869.69, 
    91394.28, 85199.81, 80315.66, 77806.2, 78055.64, 81024.47, 79534.84, 
    90081.24,
  101936.2, 101713.2, 99485.7, 94014.9, 90921.84, 88839.1, 87540.56, 87779.3, 
    82539.38, 79635.92, 78725.46, 79376.38, 81579.8, 80382.2, 91608.89,
  92325.18, 88733.76, 93630.35, 92172.42, 85358.96, 84140.92, 86441.87, 
    85682.3, 80526.7, 78096.57, 76963.52, 77638.5, 79034.45, 80655.23, 93682.2,
  86178.35, 86221.12, 85162.7, 83368.71, 82944.52, 81297.02, 82072.61, 
    82380.19, 79888.32, 78428.89, 78146.73, 79689.88, 79075.3, 81212.05, 
    87333.45,
  87784.28, 86619.31, 87596.02, 86715.04, 86395.84, 84669.98, 83459.73, 
    82876.48, 81738.85, 83910.7, 99202.44, 99921.66, 89724.74, 90070.35, 
    82218.77,
  88079.14, 86118.6, 88545.11, 89356.4, 88302.02, 87732.44, 86857.77, 
    87197.51, 88729.64, 99918.46, 100907.4, 100961.7, 100682.2, 92258.55, 
    76457.12,
  87204.52, 86312.46, 88326.23, 89570.66, 89234.91, 89130.39, 88975, 
    90875.42, 94822.09, 100714.3, 100665.1, 100688.6, 100655.8, 85879.41, 
    76118.01,
  91077.82, 87609.16, 87904.22, 89694.87, 89212.91, 88005.4, 88492.63, 
    90207.55, 94588.7, 100538.9, 100489.8, 100564.9, 100481.1, 84552.97, 
    86184.62,
  94165.98, 89587.81, 88484.99, 89506.53, 88499.7, 85932.08, 87042.34, 
    89698.13, 99985.97, 100445.2, 100315.7, 100299.8, 100258.2, 92193.96, 
    94644.76,
  97434.81, 92581.53, 90777.06, 93063.19, 93185.35, 93268.44, 94009.13, 
    99907.52, 100375.5, 100253, 100112.3, 100063.7, 100030.6, 97718.86, 
    98841.8,
  101442.4, 101088.7, 97036.82, 94336.79, 94260.79, 93200.55, 90765.77, 
    91303.93, 85273.95, 80386.24, 77897.95, 78188.28, 81047.43, 79663.3, 
    89914.02,
  101509.1, 101285.7, 98982.48, 93673.55, 90735.2, 88724.6, 87419.34, 
    87693.34, 82551.86, 79681.84, 78827.85, 79487.98, 81656.84, 80529.43, 
    91433.66,
  92100, 88558.07, 93449.78, 92018.32, 85318.83, 84151.15, 86461.81, 
    85710.42, 80603.02, 78245.7, 77167.2, 77796.33, 79176.34, 80736.94, 
    93530.65,
  86052.93, 86160.88, 85142.12, 83336.46, 83004.9, 81406.34, 82185.91, 
    82454.7, 80013.56, 78616.86, 78313.92, 79872.84, 79269.25, 81263.57, 
    87328.66,
  87700.02, 86628.14, 87628.37, 86754.49, 86505.91, 84802.79, 83640.95, 
    83083.86, 81965.88, 84120.55, 99473.05, 100056.2, 89810.94, 90014.49, 
    82291.73,
  88057.1, 86168.96, 88651.51, 89461.27, 88461.08, 87940.59, 87090.36, 
    87432.73, 88998.84, 100234.6, 101003.3, 100921.7, 100599.2, 92203.59, 
    76546.45,
  87268.62, 86417.16, 88524.06, 89789.7, 89512.98, 89438.16, 89292.64, 
    91225.16, 95192.22, 101002.2, 100852.1, 100783.8, 100596.3, 85899.95, 
    76231.65,
  91175.56, 87746.23, 88169.46, 90013.41, 89574.12, 88395.19, 88925.88, 
    90655.47, 95072.3, 100976.1, 100805.8, 100744.9, 100520.8, 84555.51, 
    86419.23,
  94295.02, 89790.64, 88789.86, 89894.87, 88942.42, 86414.05, 87590.48, 
    90282.49, 100593.8, 100945.9, 100745.7, 100663.4, 100478.5, 92381.99, 
    94964.24,
  97625.62, 92819.36, 91143.58, 93542.12, 93723.72, 93823.94, 94626.95, 
    100639.6, 101036.5, 100917.3, 100729, 100626.5, 100489.8, 98112.73, 
    99187.05,
  102317.5, 102122.3, 97967.33, 95332.03, 95299.83, 94164.5, 91631.41, 
    92200.73, 85920.08, 81094.45, 78608.36, 78887.94, 81872.86, 80408.73, 
    90999.35,
  102485.7, 102331.6, 100068, 94640.62, 91596.51, 89602.59, 88342.73, 
    88599.11, 83328.2, 80530.36, 79637.66, 80327.98, 82533.89, 81283.1, 
    92504.98,
  92928.81, 89305.12, 94349.22, 92873.05, 86155.21, 85015.42, 87340.6, 
    86544.12, 81409.06, 79014.74, 77820.43, 78541.18, 79954.9, 81567.92, 
    94645.83,
  86725.88, 86845.07, 85869.36, 84107.41, 83793.62, 82199.59, 83035.69, 
    83347.82, 80854.1, 79422.3, 79275.88, 80857.3, 80080.26, 82223.19, 
    88293.75,
  88304.63, 87294.81, 88372.55, 87555.16, 87349.34, 85670.75, 84504.38, 
    83954.18, 82825.07, 85149.25, 100593.4, 101187.5, 90914.5, 91189.16, 
    83179.69,
  88700.4, 86834.1, 89398.85, 90289.93, 89341.62, 88844.05, 88038.18, 
    88413.23, 90064.58, 101399, 102308.3, 102289.4, 101992.1, 93365.11, 
    77428.89,
  87824.6, 87044.71, 89239.05, 90587.1, 90337.45, 90330.09, 90249.81, 
    92236.13, 96313.64, 102215.9, 102143.2, 102069.6, 102030.4, 86923.45, 
    77207.08,
  91733.11, 88371.56, 88834.28, 90734.79, 90373.73, 89283.44, 89860.55, 
    91649.41, 96138.35, 102144.8, 102094, 102118.2, 101978.3, 85649.05, 
    87659.98,
  94781.27, 90337.86, 89385.25, 90547.52, 89653.03, 87167.33, 88404.47, 
    91216.73, 101627, 102139.6, 102026.4, 102065, 101925.1, 93723.37, 96319.26,
  98043.22, 93298.92, 91659.7, 94124.84, 94364.82, 94553.76, 95454.6, 
    101541.4, 102103.3, 102079.5, 102002.8, 102046.8, 101980.7, 99593.91, 
    100743.4,
  102351.5, 102079.1, 98069.93, 95549.95, 95549.73, 94476.48, 92009.73, 
    92578.53, 86409.12, 81511.88, 79086.23, 79377.03, 82375.03, 80911.9, 
    91496.9,
  102290.1, 102381, 100058.2, 94698.3, 91826.73, 89868.97, 88613.44, 
    88920.41, 83742.42, 80872.09, 80021.42, 80705.96, 82954.43, 81749.7, 
    92984.31,
  93020.62, 89346.74, 94510.26, 93126.08, 86391.15, 85233.4, 87613.62, 
    86870.66, 81750.65, 79382.84, 78290.75, 78981.05, 80397.4, 82018.7, 
    95142.8,
  86662.07, 86681.1, 85872.8, 84134.56, 83850.99, 82333.73, 83221.23, 
    83557.55, 81142.84, 79750.8, 79505.8, 81142.98, 80479.06, 82643.97, 
    88769.28,
  88307.59, 87155.06, 88313.18, 87475.29, 87344.69, 85703.09, 84612.45, 
    84079.66, 83056.57, 85198.93, 100664.6, 101273.6, 91172.95, 91549.39, 
    83595.49,
  88450.83, 86656.66, 89182.85, 90100.31, 89191.81, 88759.66, 88014.12, 
    88435.89, 90053.01, 101336.7, 102345.2, 102357.1, 102157.9, 93707.09, 
    77898.31,
  87525.2, 86796.13, 88984.7, 90351.05, 90140.38, 90213.98, 90147.84, 
    92178.77, 96229.34, 102130.3, 102132.4, 102166.9, 102208.1, 87293.5, 
    77719.61,
  91315.9, 88030.64, 88521.99, 90424.2, 90123.78, 89112.92, 89748.22, 
    91654.1, 95985.23, 102006.6, 102056.8, 102179.7, 102130.1, 86036.65, 
    88098.51,
  94297.95, 89939.57, 89025.92, 90183.06, 89409.02, 86998.41, 88299.2, 
    90950.27, 101367.2, 101936.2, 101952.9, 102052.2, 102068.4, 93991.77, 
    96696.35,
  97473.55, 92784.53, 91150.91, 93620.06, 93918.12, 94077.06, 95048.98, 
    101177.6, 101811.3, 101828.4, 101874.7, 101961.9, 102042.4, 99744.01, 
    101019.4,
  101522.4, 101252.7, 97422.89, 94976, 95029.34, 94023.2, 91679.02, 92182.34, 
    86181.48, 81339.16, 78953.7, 79285.9, 82228.97, 80839.41, 91352.28,
  101468.7, 101598.4, 99294.55, 94036.52, 91334.94, 89453.34, 88214.59, 
    88571.08, 83507.51, 80642.16, 79827.38, 80523.61, 82768.41, 81670.04, 
    92828.37,
  92328.09, 88748.3, 93916.59, 92534.67, 85913.53, 84806.37, 87227.14, 
    86554.6, 81462.16, 79150.78, 78199.9, 78911.4, 80314.45, 81909.91, 
    94995.37,
  85956.48, 86005.69, 85264.23, 83571.42, 83318.99, 81852.14, 82812.25, 
    83185.01, 80824.41, 79532.84, 79176.64, 80744.18, 80377.96, 82405.39, 
    88715.24,
  87548.21, 86503.29, 87666.92, 86811.42, 86715.98, 85095.85, 84081.38, 
    83654.08, 82684.12, 84663.73, 100033.7, 100791.5, 90739.11, 91138.08, 
    83608.88,
  87754.27, 85974.91, 88505.02, 89446.38, 88579.05, 88154.95, 87459.23, 
    87896.92, 89490.95, 100698.9, 101705.2, 101700.3, 101496.8, 93313.83, 
    77865.59,
  86888.67, 86167.74, 88334.05, 89696.96, 89504.49, 89599.3, 89553.44, 
    91622.12, 95659.87, 101464.6, 101471.2, 101607.4, 101552.5, 87060.12, 
    77571.48,
  90708.12, 87417.95, 87907.82, 89799.66, 89520.75, 88543.67, 89187.8, 
    91101.87, 95376.82, 101366.6, 101391.5, 101581.3, 101507.8, 85786.64, 
    87716.89,
  93785.84, 89376.74, 88493.38, 89632.95, 88842.23, 86480.8, 87790.17, 
    90431.04, 100762.9, 101323.9, 101297.2, 101432.1, 101474.1, 93481.54, 
    96223.6,
  97042.87, 92299.66, 90715.33, 93166.46, 93457.34, 93593.87, 94546.79, 
    100641, 101232.5, 101244.7, 101263.7, 101329, 101431.4, 99184.54, 100425.3,
  101167.3, 101027, 97037.93, 94512.98, 94481.09, 93470.78, 91137.35, 
    91680.51, 85693.6, 80922.91, 78603.28, 78910.12, 81963.76, 80499.23, 
    91097.85,
  101300.7, 101324.7, 98940.62, 93673.21, 90868.21, 88987.55, 87719.76, 
    88113.24, 83069.32, 80262.77, 79475.24, 80183.67, 82452.77, 81357.95, 
    92555.73,
  91988.09, 88499.5, 93572.35, 92182.34, 85514.05, 84451.55, 86832.52, 
    86121.68, 81074.26, 78813.47, 77902.92, 78631.73, 80040.12, 81670.39, 
    94644.6,
  85826.38, 86026.99, 85046.6, 83343.72, 83074.09, 81568.65, 82503.35, 
    82871.75, 80527.75, 79255.38, 78889.02, 80465.84, 80120.11, 82185.72, 
    88438.81,
  87492.09, 86546.05, 87645.53, 86779.36, 86613.95, 84948.8, 83897.31, 
    83425.53, 82449.66, 84545.66, 100044.6, 100680.4, 90544.86, 90919.06, 
    83375.38,
  87919.3, 86071.55, 88625.08, 89477.86, 88558.17, 88105.3, 87386.43, 
    87800.69, 89483.85, 100854.8, 101639.4, 101612.7, 101454.4, 93149.16, 
    77680.77,
  87164.98, 86395.87, 88592.58, 89829.72, 89594.16, 89628.47, 89592.8, 
    91681.16, 95791.65, 101591.7, 101479.7, 101522.4, 101499.6, 86849.67, 
    77434.88,
  91094.71, 87745.98, 88267.66, 90117.78, 89731.54, 88694.81, 89363.16, 
    91234.25, 95649.63, 101608.9, 101503.3, 101545.5, 101491.1, 85658.3, 
    87676.84,
  94260.86, 89803.95, 88904.4, 90051.54, 89175.29, 86714.2, 88027.3, 
    90753.55, 101234.1, 101627.4, 101483.8, 101484.2, 101485.7, 93449.01, 
    96261.55,
  97623.27, 92830.57, 91279.38, 93762.82, 94026.02, 94186.32, 95126.21, 
    101283.5, 101736.4, 101613.7, 101508.2, 101473.9, 101504.5, 99199.54, 
    100428.4,
  101470.4, 101212.5, 97210.38, 94676.77, 94671.52, 93608.26, 91201.2, 
    91728.84, 85707.78, 80927.23, 78600.23, 78895.27, 81934.87, 80465.98, 
    91105.48,
  101477.3, 101518.2, 99164.91, 93896.51, 91031.04, 89110.68, 87842.9, 
    88157.09, 83081.83, 80281.23, 79480.66, 80170.37, 82444.56, 81297.41, 
    92535.46,
  92239.72, 88645.94, 93730.81, 92321.82, 85658.45, 84555.2, 86927.32, 
    86187.72, 81119.29, 78841.09, 77910.77, 78646.45, 80053.22, 81696.79, 
    94711.39,
  86016.91, 86126.66, 85222.27, 83513.67, 83233.54, 81695.55, 82568.55, 
    82923.48, 80576.18, 79280.07, 78931.52, 80545.89, 80148.27, 82269.05, 
    88480.75,
  87640.16, 86626.02, 87750.78, 86936.61, 86783.91, 85105.22, 84024.89, 
    83496.4, 82517.75, 84665.52, 100436.5, 100975.7, 90685.3, 91088.17, 
    83408.19,
  87952.34, 86133.02, 88741.61, 89646.05, 88725.38, 88268.7, 87547.01, 
    87967.14, 89650.06, 101191.4, 102016, 101902.3, 101693.8, 93333.16, 
    77700.12,
  87098.37, 86367.64, 88617.85, 89981.9, 89770.59, 89804.01, 89772.45, 
    91880.97, 96064.54, 101999.9, 101873.5, 101791.5, 101721.1, 86991.72, 
    77503.45,
  90922.41, 87641.36, 88195.04, 90148.17, 89868.12, 88834.05, 89502.71, 
    91406.2, 95872.2, 101944.9, 101900.5, 101844, 101769, 85734.05, 87838.29,
  94004.02, 89638.24, 88775.95, 89987.84, 89187.01, 86744.8, 88104.85, 
    90851.04, 101514.5, 101955.6, 101876.6, 101793.4, 101773.5, 93545.09, 
    96486.96,
  97295.45, 92554.15, 91030.76, 93614.76, 93947.02, 94174.81, 95163.55, 
    101442.5, 101984.8, 101931, 101877.3, 101810, 101760.4, 99417.17, 100695.9,
  101007, 100702.9, 96838.95, 94399.64, 94431.11, 93378.48, 91027.98, 
    91574.51, 85607.16, 80845.37, 78494.52, 78829.82, 81897.43, 80498.71, 
    91066.36,
  100850.4, 100938.8, 98688.27, 93491.77, 90781.21, 88902.25, 87652.69, 
    88010.9, 82974.57, 80177.8, 79402.75, 80118.43, 82406.08, 81314.81, 
    92479.89,
  91770.42, 88207.64, 93416.29, 92034.28, 85401.03, 84344.77, 86742.66, 
    86030.99, 80995.91, 78712.04, 77812.93, 78562.13, 80002.95, 81645.51, 
    94677.7,
  85487.55, 85636.3, 84770.81, 83163.89, 82935.41, 81477.3, 82413.25, 
    82758.1, 80416.67, 79151, 78825.71, 80406.91, 80095.27, 82153.62, 88469.93,
  87132.66, 86232.02, 87317.79, 86482.91, 86385.84, 84787.87, 83778.34, 
    83315.77, 82373.48, 84451.02, 99959.41, 100605.7, 90449.76, 90890.95, 
    83392.73,
  87453.02, 85668.34, 88244.41, 89168.32, 88304.26, 87885.32, 87176.77, 
    87622.07, 89286.1, 100698.1, 101690.9, 101623.6, 101408.8, 93121.25, 
    77654.25,
  86670.41, 85939.07, 88162.01, 89493.28, 89305.99, 89395.09, 89345.55, 
    91432.84, 95598.45, 101587.3, 101501, 101569.7, 101459.6, 86887.34, 
    77398.9,
  90484.88, 87222.2, 87751.38, 89667.59, 89417.76, 88409.64, 89067, 91013.05, 
    95425.61, 101577.4, 101555.7, 101666, 101518.2, 85640.89, 87600.05,
  93584.3, 89239.95, 88364.58, 89526.1, 88751.56, 86356.04, 87686, 90418.86, 
    101006.4, 101585.7, 101576, 101620.4, 101627.8, 93444.65, 96297.73,
  96864.16, 92146.28, 90586.56, 93082.59, 93382.04, 93594.35, 94639.63, 
    100899.3, 101549.2, 101574.4, 101615.2, 101611.1, 101645.4, 99265.62, 
    100584,
  101247.6, 100937.5, 97053.03, 94560.3, 94566.8, 93536.13, 91126.03, 
    91681.83, 85657.26, 80927.74, 78568.76, 78881.52, 82015.03, 80540.49, 
    91250.09,
  101176.4, 101202.4, 98919.75, 93660.74, 90909.18, 89025.45, 87772.35, 
    88149.36, 83062.17, 80299.68, 79481.49, 80200.62, 82511.88, 81384.01, 
    92714.4,
  92042.54, 88413.04, 93594.34, 92208.43, 85561.75, 84507.34, 86874.02, 
    86164.58, 81124.51, 78864.02, 77937, 78678.12, 80114.89, 81796.53, 
    94850.11,
  85752.73, 85884.52, 85006.05, 83333.81, 83102.9, 81627.62, 82556.45, 
    82911.02, 80572.47, 79289.06, 78960.16, 80548.38, 80219.95, 82333.43, 
    88645.1,
  87375.8, 86433.31, 87515.18, 86685.59, 86578.82, 84965.2, 83938.02, 
    83479.38, 82516.72, 84613.66, 100102.3, 100686.8, 90576.53, 91068.9, 
    83526.12,
  87680.92, 85887.89, 88417.3, 89334.17, 88464.05, 88037.68, 87330.59, 
    87765.66, 89421.91, 100715.7, 101664.7, 101604.5, 101486.1, 93241.29, 
    77821.96,
  86850.55, 86106.95, 88317.5, 89652.85, 89474.72, 89557.35, 89494.45, 
    91553.16, 95703.51, 101619.6, 101565.4, 101592.7, 101523.2, 86991.86, 
    77566.66,
  90634.79, 87348.55, 87900.83, 89831.4, 89541.89, 88548.02, 89216.14, 
    91171.41, 95556.07, 101621.4, 101594.9, 101688.5, 101560.3, 85811.73, 
    87807.93,
  93670.45, 89335.62, 88478.84, 89672.57, 88912.8, 86543.09, 87873.92, 
    90558.58, 101087.1, 101643.7, 101636.9, 101676.9, 101634.9, 93567.95, 
    96382.16,
  96893.52, 92223.14, 90695.82, 93230.99, 93526.84, 93687.68, 94744.97, 
    100981.7, 101620.4, 101634.7, 101692.6, 101713.4, 101753.3, 99427.95, 
    100681,
  101688.5, 101427.6, 97501.8, 95023.83, 95074.24, 94076.18, 91683.68, 
    92241.55, 86224.88, 81461.76, 79091.45, 79452.05, 82632.07, 81171.64, 
    92091.27,
  101574, 101639.5, 99340.66, 94126.91, 91405.76, 89539.4, 88289.32, 88676.9, 
    83599.96, 80827.63, 80005.28, 80737.62, 83106.63, 81974.06, 93417.41,
  92481.58, 88829.85, 94045.33, 92653.98, 86007.84, 84966.24, 87356.32, 
    86670.76, 81618.3, 79352.23, 78422.34, 79179.68, 80645.91, 82342.39, 
    95544.82,
  86138.29, 86247.77, 85424.7, 83772.24, 83527.88, 82078.77, 83035.84, 
    83393.62, 81047.38, 79769.34, 79444.62, 81043.18, 80724.27, 82856.71, 
    89270.62,
  87726.33, 86794.91, 87906.07, 87099.23, 87012.88, 85402.41, 84403.43, 
    83951.12, 82983.24, 85071.08, 100570.6, 101178.7, 91103.93, 91593.01, 
    84087.62,
  88005.17, 86242.28, 88809.63, 89743.98, 88902.2, 88486.23, 87798.61, 88243, 
    89906.09, 101192.3, 102117.6, 102080.6, 101968.3, 93759.77, 78325.46,
  87172.07, 86466.85, 88688.34, 90046.45, 89885.8, 89985.8, 89948.16, 
    92016.45, 96137.55, 102038.2, 102001.8, 102038.1, 101997.7, 87502.91, 
    78029.53,
  90933.05, 87714.27, 88275.26, 90195.62, 89929.36, 88968.08, 89649.44, 
    91550.29, 95970.79, 102044.2, 102029.9, 102107.7, 102013.7, 86262.62, 
    88268.14,
  93969.91, 89682.84, 88855.24, 90035.19, 89290.11, 86959.11, 88322.84, 
    90994.83, 101459.9, 102060.5, 102051.2, 102096, 102074.1, 94024.48, 
    96870.26,
  97180.55, 92567.76, 91051.96, 93572.97, 93870.87, 94042.03, 95081.02, 
    101272.2, 102010.1, 102074.7, 102133, 102153.5, 102141, 99797.91, 101068.6,
  101854.6, 101575.3, 97686.3, 95230.16, 95266.2, 94245.54, 91864.55, 
    92425.81, 86405.32, 81616.16, 79247.11, 79534.64, 82651.38, 81200.03, 
    92058.01,
  101638.2, 101729.9, 99464.73, 94284.52, 91575.45, 89708.16, 88455.66, 
    88829.69, 83770.77, 80953.76, 80138.78, 80830.91, 83138.71, 82009.28, 
    93432.55,
  92558.39, 88992.03, 94158.56, 92782.63, 86174.6, 85126.11, 87515.62, 
    86829.59, 81781.29, 79475.52, 78522.88, 79244.12, 80687.05, 82343.08, 
    95589.24,
  86170.04, 86302.78, 85517.12, 83891.48, 83669.44, 82222.77, 83174.65, 
    83540.52, 81180.01, 79876.83, 79531.18, 81125.23, 80712.97, 82824.03, 
    89244.02,
  87765.45, 86847.68, 87993.75, 87178.96, 87122.52, 85545, 84546.25, 
    84083.95, 83105.42, 85188.45, 100672, 101327, 91214.99, 91638.42, 84029.89,
  88027.02, 86287.16, 88907.27, 89856.82, 89039.05, 88643.23, 87961.59, 
    88406.04, 90054.79, 101444.8, 102318, 102237.8, 102038.8, 93793.31, 
    78271.17,
  87200.76, 86524.7, 88809.3, 90166.59, 90039.12, 90150.82, 90134.63, 
    92224.33, 96386.78, 102292.1, 102143.2, 102186.8, 102104.4, 87517.84, 
    78000.46,
  91052.85, 87786.41, 88405.6, 90360.65, 90126.85, 89161.45, 89862.84, 
    91793.44, 96239.74, 102311, 102242.1, 102287.9, 102140.1, 86258.23, 
    88279.03,
  94181.19, 89838.6, 89051.78, 90273.44, 89512.53, 87164.3, 88538.44, 
    91272.83, 101896.5, 102386.6, 102310.8, 102311.9, 102187.8, 94072.69, 
    96857.75,
  97509.63, 92863.11, 91380.14, 93949.52, 94242.3, 94446.61, 95529.41, 
    101863.6, 102454.2, 102461, 102438.2, 102426.1, 102338.3, 99972.2, 
    101184.4,
  101560.7, 101264.6, 97313.79, 94767.93, 94758.15, 93755.75, 91415.59, 
    91957.24, 85972.72, 81192.01, 78830.57, 79118.46, 82111.72, 80679.5, 
    91220.48,
  101474.6, 101454.1, 99135.97, 93873.54, 91090.09, 89200.81, 87934.09, 
    88333.9, 83304.5, 80489.67, 79667.68, 80362.89, 82618.94, 81492.21, 
    92675.47,
  92252.39, 88652.13, 93741.78, 92380.66, 85695.71, 84625.34, 86988.39, 
    86314.75, 81292.09, 79017.68, 78068.67, 78785.73, 80202.74, 81801.78, 
    94879.8,
  86003.8, 86159.35, 85214.77, 83533.82, 83251.66, 81746.74, 82631.77, 
    82995.41, 80670.52, 79414.65, 79057.61, 80635.98, 80236.26, 82285.59, 
    88571.66,
  87630.52, 86716.2, 87783.3, 86929.77, 86774.8, 85115.15, 84039.78, 
    83550.31, 82587.78, 84684.05, 100327.2, 100990.6, 90763.89, 91087.75, 
    83464,
  88045.35, 86217.85, 88763.52, 89611.39, 88683.68, 88231.41, 87497.57, 
    87941.36, 89674.77, 101237.1, 102045.2, 101951.9, 101662.7, 93325.09, 
    77729.98,
  87286.03, 86505.44, 88723.16, 89972.33, 89761.31, 89813.55, 89778.63, 
    91928.41, 96127.84, 102067.8, 101900, 101918.4, 101750.6, 87017.91, 
    77469.43,
  91179.27, 87810.41, 88369.16, 90241.88, 89905.32, 88885.04, 89557.27, 
    91458.34, 95950.82, 102100.7, 102000.8, 102013, 101803.3, 85745.02, 
    87724.96,
  94342.84, 89928.66, 89056.67, 90196.34, 89327.79, 86894.48, 88242.44, 
    90998.32, 101690.3, 102154.3, 102050.7, 102028, 101819, 93633.62, 96406.96,
  97743.16, 92957.06, 91392.39, 93935.91, 94211, 94386.65, 95374.16, 
    101666.2, 102193, 102205, 102153.1, 102133.1, 102050.4, 99643.52, 100862.2,
  101149.3, 100812.3, 96822.41, 94219.33, 94201.62, 93114.45, 90692.38, 
    91214.99, 85233.73, 80434.55, 78081.58, 78384.44, 81385.98, 79970.16, 
    90356.09,
  101274.2, 101111.8, 98822.4, 93503.76, 90611.23, 88646.88, 87346.91, 
    87634.91, 82581.29, 79745.3, 78927.91, 79624.92, 81883.22, 80801.83, 
    91793.98,
  91901.45, 88434.73, 93396.67, 91951.17, 85289.16, 84148.63, 86446.05, 
    85679.1, 80609.37, 78303.57, 77362.62, 78082.94, 79479.89, 81096.95, 
    93955.2,
  85869.55, 86055.7, 85023.31, 83281.59, 82961.26, 81383.67, 82226.16, 
    82499.21, 80084.19, 78757.14, 78450.7, 80014.18, 79596.39, 81638.3, 
    87757.32,
  87529.98, 86555.54, 87621.56, 86759.82, 86542.67, 84848.13, 83711.96, 
    83159.47, 82094.88, 84310.84, 100001.6, 100611, 90264.84, 90505.3, 
    82835.45,
  87970.73, 86100.05, 88683.87, 89515.39, 88529.91, 88025, 87210.68, 
    87610.32, 89283.66, 100829.8, 101666.3, 101608.6, 101305.7, 92792.99, 
    77118.73,
  87216, 86393.41, 88593.39, 89873.76, 89602.41, 89552.05, 89452.23, 
    91486.48, 95603.15, 101592.1, 101470.5, 101513.4, 101296.2, 86493.79, 
    76756.62,
  91173.88, 87758.16, 88203.85, 90082.39, 89682.48, 88542.04, 89146.81, 
    90976.98, 95435.79, 101548.2, 101461.6, 101527.9, 101309.8, 85254.92, 
    86991.35,
  94350.71, 89799.71, 88812.79, 89950.66, 89010.31, 86509.54, 87742.92, 
    90513.62, 101010.5, 101491.9, 101374.9, 101401.9, 101304.5, 93103.67, 
    95812.15,
  97730.41, 92871.11, 91191.88, 93609.23, 93814.98, 93971.42, 94819.62, 
    100941.2, 101454.7, 101401.6, 101322.4, 101322.2, 101329.6, 98971.1, 
    100167.5,
  101455.8, 101161.7, 97161.09, 94499.55, 94414.34, 93297.15, 90829.4, 
    91329.41, 85302.27, 80463.2, 78042.41, 78335.23, 81271.16, 79873.3, 
    90323.82,
  101598.6, 101462.1, 99192.62, 93815.43, 90823.08, 88807.01, 87525.3, 
    87785.47, 82629.77, 79748.26, 78913.46, 79596.14, 81814.98, 80718.73, 
    91800.55,
  92109.77, 88595.99, 93569.49, 92124.2, 85400.7, 84234.46, 86553.93, 
    85787.78, 80670.03, 78336.21, 77327.98, 78022.18, 79423.06, 81057.46, 
    93932.11,
  86028.5, 86190.97, 85167.84, 83369.59, 83041.2, 81435.23, 82254.41, 
    82536.38, 80085.2, 78728.92, 78389.6, 79971.09, 79484.09, 81578.38, 
    87684.89,
  87707.66, 86673.95, 87701.86, 86832.5, 86581.67, 84878.16, 83725.13, 
    83150.99, 82065.31, 84179.53, 99691.66, 100349.8, 90118.05, 90428.19, 
    82720.2,
  88119.18, 86220.23, 88749.04, 89550.77, 88543.11, 88008.4, 87156.11, 
    87506.94, 89102.03, 100381.3, 101235.7, 101249.6, 101023.6, 92655.02, 
    76944.92,
  87338.54, 86495.75, 88640.91, 89876.03, 89586.68, 89505.49, 89369.86, 
    91313.23, 95284.03, 101103.6, 101021, 101067.4, 101015.4, 86304.6, 
    76628.16,
  91273.57, 87840.32, 88268.45, 90082.07, 89630.32, 88445.97, 88974.05, 
    90697.89, 95091.14, 100997.1, 100886.1, 100921.9, 100864.4, 84939.21, 
    86872.24,
  94411.23, 89881.42, 88897.43, 89993.12, 89015.67, 86475.73, 87641.08, 
    90328.01, 100598.3, 100923.8, 100748.7, 100721, 100729.4, 92684.67, 
    95414.65,
  97740.62, 92931.23, 91263.14, 93652.08, 93815.88, 93931.51, 94733.05, 
    100693.9, 101011.1, 100826.2, 100650.7, 100587, 100589.8, 98333.41, 
    99607.85,
  102180.1, 101898, 97726.14, 95026.5, 94933.74, 93760.59, 91232.38, 
    91753.64, 85547.03, 80757.41, 78335.77, 78667.06, 81687.73, 80243.78, 
    90823.72,
  102291.8, 102094.1, 99803.8, 94364.34, 91363.39, 89314.39, 88036.48, 
    88251.18, 83006.41, 80225.14, 79350.66, 80074.67, 82290.03, 81108.38, 
    92330.8,
  92677.41, 89214.29, 94219.98, 92678.48, 85882.49, 84784.11, 87091.4, 
    86273.74, 81146.45, 78788.52, 77694.94, 78464.11, 79861.02, 81494.46, 
    94468.15,
  86604.13, 86773.68, 85705.74, 83959.5, 83638.48, 81999.79, 82832.53, 
    83141.38, 80639.08, 79214.77, 79022.44, 80590.58, 79939.23, 82108.52, 
    88180.74,
  88217.71, 87216.36, 88272.86, 87403.23, 87170.14, 85476.91, 84325.75, 
    83744.45, 82619.55, 84982.88, 100484.2, 101089.6, 90754.87, 91074.52, 
    83081.86,
  88630.5, 86768.58, 89351.99, 90167.53, 89217.95, 88691.3, 87870.84, 
    88216.45, 89909.22, 101183.7, 102072.3, 102045.6, 101778.8, 93222.23, 
    77363.09,
  87812.2, 87007.32, 89189.81, 90471.88, 90227.07, 90166.85, 90108, 92063.77, 
    96116.34, 101990.5, 101964.4, 101840.5, 101768.7, 86757.8, 77154.3,
  91710.12, 88339.42, 88808.43, 90661.93, 90265.1, 89136.43, 89682.05, 91456, 
    95975.68, 101920.4, 101869.6, 101854.9, 101710.2, 85486.36, 87545.15,
  94810.66, 90341.8, 89361.09, 90495.45, 89571.08, 87090.05, 88306.11, 
    91117.14, 101383.9, 101890.9, 101790.5, 101775.1, 101652.5, 93473.45, 
    96146.16,
  98109.02, 93309.04, 91650.96, 94067.05, 94277.79, 94442.8, 95299.48, 
    101285.4, 101812.7, 101812.1, 101700.3, 101684.4, 101624.9, 99247.76, 
    100390.7,
  102480, 102116.7, 98072.41, 95461.39, 95433.52, 94324.91, 91845.7, 
    92440.77, 86206.36, 81395.95, 78959.53, 79269.79, 82290.3, 80777.82, 
    91463.38,
  102403, 102395.5, 100103.2, 94717.48, 91755.93, 89777.86, 88545.66, 
    88835.97, 83614.34, 80839.55, 79932.28, 80634.41, 82845.36, 81634.68, 
    92982.36,
  93086.8, 89426.87, 94481.98, 93054.45, 86353.28, 85212.45, 87520.85, 
    86760.77, 81684.17, 79306.68, 78163.88, 78939.97, 80335.77, 82036.2, 
    95109.3,
  86810.91, 86832.48, 85941.52, 84233.91, 83926.62, 82384.65, 83224.48, 
    83529.57, 81090.73, 79691.41, 79530.88, 81085.12, 80379.35, 82647.96, 
    88744,
  88502.67, 87309.49, 88395.34, 87556.34, 87386.73, 85729.92, 84614.37, 
    84080.41, 83011.8, 85262.55, 100498.7, 101148.8, 91131.1, 91594.09, 
    83542.06,
  88651.52, 86815.57, 89309.46, 90201.73, 89277.77, 88804.82, 88039.23, 
    88405.81, 90039.76, 101174.1, 102177.9, 102273.3, 102092.1, 93669.99, 
    77902.91,
  87739.35, 86993.79, 89125.95, 90450.12, 90223.1, 90232.07, 90145.09, 
    92102.08, 96130.31, 101963.2, 102001.3, 102038.1, 102157, 87285.03, 
    77745.18,
  91525.25, 88236.91, 88681.35, 90548.21, 90217.48, 89161.3, 89763.62, 
    91595.18, 95930.82, 101860.9, 101889.3, 102014.9, 101996.8, 86030.88, 
    88057.27,
  94540.52, 90163.64, 89190.89, 90323.65, 89495.43, 87077.32, 88337.46, 
    90983.37, 101273.8, 101808, 101773.8, 101844.7, 101851.6, 93836.96, 
    96395.67,
  97728.72, 92981.1, 91337.97, 93771.8, 94028.27, 94163.34, 95088.54, 
    101114.9, 101713.9, 101684.1, 101674.6, 101706.5, 101732.3, 99431.48, 
    100589.8,
  102053.1, 101658.6, 97733.66, 95215.16, 95249.74, 94219.32, 91808.59, 
    92311.36, 86275.52, 81451.27, 79064.86, 79337.9, 82284.14, 80810.8, 
    91270.76,
  101868.8, 101931.1, 99616.92, 94342.3, 91558.73, 89627.39, 88379.17, 
    88713.83, 83645.2, 80778.16, 79924.05, 80582.08, 82798.56, 81632.87, 
    92705.92,
  92706.58, 89087.24, 94204.7, 92846.09, 86190.43, 85033.27, 87407.05, 
    86705.55, 81647.32, 79303.72, 78319.36, 78991.2, 80365.94, 81953.2, 
    94859.05,
  86371.86, 86340.77, 85549.99, 83863.5, 83602.48, 82106.51, 83020.69, 
    83357.49, 80993.21, 79658.94, 79311.78, 80879.63, 80440.95, 82466.92, 
    88570.59,
  87952.8, 86834.73, 87980.09, 87138.38, 87006.33, 85376.25, 84328.1, 
    83859.34, 82864.07, 84885.78, 100110.1, 100813.8, 90821.83, 91172.02, 
    83581.29,
  88073.71, 86265.1, 88777.72, 89701.78, 88811.77, 88371.13, 87633.35, 
    88029.52, 89628.24, 100741.8, 101693.5, 101723.1, 101516.5, 93357.51, 
    77880.23,
  87179.12, 86437.97, 88584.77, 89929.6, 89708.66, 89766.16, 89680.83, 
    91688.74, 95670.81, 101473.6, 101434, 101591.2, 101501.6, 87163.2, 
    77579.41,
  90973.78, 87682.64, 88123.43, 89999.83, 89678.77, 88667.01, 89274.18, 
    91167.38, 95395.28, 101360.4, 101331.2, 101509.1, 101382.7, 85868.02, 
    87535.41,
  93994.32, 89594.83, 88637.8, 89762.42, 88959.65, 86546.98, 87828.26, 
    90439.06, 100720.3, 101321.1, 101250.3, 101352.2, 101310.3, 93394.16, 
    95950.66,
  97219.69, 92471.32, 90789.46, 93214.31, 93478.09, 93616.44, 94536.99, 
    100631.7, 101256.7, 101209.5, 101173.5, 101190.5, 101228.7, 98935.27, 
    100075.4,
  101642.4, 101314.5, 97403.12, 94929.55, 94979.18, 93987.53, 91628.41, 
    92149.1, 86147, 81366.07, 78972.73, 79270.05, 82231.45, 80745.88, 91248.3,
  101490.1, 101536.2, 99243.84, 94029.44, 91303.86, 89426, 88195.05, 
    88567.68, 83510.71, 80672.1, 79826.64, 80517.73, 82764.63, 81597.3, 
    92724.77,
  92364.23, 88786.18, 93880.77, 92519.48, 85939.32, 84857.09, 87223.78, 
    86555.54, 81514.31, 79193.28, 78230.2, 78939.8, 80325.9, 81912.66, 
    94826.84,
  86051.55, 86041.04, 85253.7, 83636.33, 83382.95, 81924.48, 82851.69, 
    83217.89, 80864.17, 79559.78, 79201.12, 80770.26, 80408.95, 82460.31, 
    88616.15,
  87644.34, 86507.55, 87642.48, 86810.25, 86712.81, 85125.77, 84114.13, 
    83678.84, 82713.69, 84742.01, 100013.5, 100719.2, 90731.8, 91132.67, 
    83602.62,
  87764.41, 85954.7, 88464.82, 89391.83, 88537.97, 88107.77, 87393.41, 
    87806.12, 89454.27, 100625.7, 101629.7, 101644.4, 101464.1, 93281.32, 
    77943.91,
  86819.95, 86115.02, 88261.23, 89600.77, 89408.27, 89474.02, 89426.01, 
    91429.58, 95467.01, 101276.1, 101376.9, 101528.8, 101476.3, 87084.55, 
    77670.55,
  90505.88, 87297.92, 87779.43, 89658.45, 89364.81, 88364.4, 88985.11, 
    90876.46, 95186.7, 101154.4, 101230.1, 101432, 101392.5, 85826.09, 87664.3,
  93425.23, 89134.28, 88228.81, 89394.68, 88635.97, 86286.36, 87579.15, 
    90192.8, 100398.5, 101063.6, 101074.8, 101231.8, 101287.6, 93395.85, 
    96052.16,
  96513.8, 91850.34, 90247.76, 92704.62, 93020.7, 93161.68, 94123.81, 
    100195.1, 100916, 100941, 101000.9, 101097, 101209.5, 98981.73, 100189.1,
  101514.5, 101200.1, 97329.45, 94877.62, 94926.02, 93947.44, 91630.58, 
    92149.01, 86207.75, 81440.59, 79097.41, 79404.88, 82393.66, 80966.87, 
    91492.53,
  101255.5, 101388.7, 99115, 93945.96, 91271.73, 89429.98, 88196.02, 
    88575.78, 83572.71, 80777.06, 79959.16, 80664.66, 82918.44, 81790.52, 
    92904.56,
  92183.56, 88618.48, 93778.33, 92447.91, 85868.62, 84823.06, 87211.88, 
    86565.98, 81556.79, 79267.53, 78334.74, 79062.02, 80471.09, 82074.3, 
    95019.26,
  85734.23, 85788.74, 85049.27, 83525.91, 83294.09, 81887.91, 82859.69, 
    83240.15, 80910.62, 79658.2, 79309.2, 80884.32, 80522.07, 82599.62, 
    88824.72,
  87270.38, 86299.93, 87400.5, 86600, 86568.95, 85033.49, 84081.34, 83678.84, 
    82745.66, 84755.56, 99971.52, 100709, 90815.95, 91236.87, 83747.9,
  87390.41, 85673.7, 88191.28, 89161.59, 88369.26, 88010.38, 87354.7, 
    87788.3, 89426.45, 100567.1, 101582.4, 101625.7, 101523.8, 93371.52, 
    78068.77,
  86464.66, 85820.95, 88009.84, 89389.81, 89259.61, 89398.29, 89384, 
    91420.98, 95448.61, 101257.4, 101343.8, 101524.2, 101547.7, 87131.74, 
    77791.02,
  90194.01, 86996.96, 87512, 89441.62, 89217.91, 88309.06, 88979.61, 
    90894.39, 95151.79, 101143.8, 101265.4, 101467.1, 101487, 85935.3, 
    87823.71,
  93222.31, 88890.5, 88039.62, 89204.7, 88501.66, 86219.91, 87578.98, 
    90161.6, 100328.5, 101010.8, 101079.1, 101258.7, 101386.7, 93519.79, 
    96205.95,
  96464.41, 91741.02, 90184.45, 92647.35, 92958.59, 93076.87, 94067.41, 
    100096.1, 100807.9, 100845.4, 100930.9, 101054.5, 101225.1, 99061.04, 
    100292.8,
  101479.9, 101182.7, 97276.08, 94839.38, 94873.9, 93836.35, 91477.2, 
    92000.5, 86021.23, 81284.52, 78958.39, 79280.45, 82389.77, 80984.1, 
    91676.25,
  101425.5, 101481.1, 99154.84, 93940.59, 91205.1, 89334.74, 88054.86, 
    88449.58, 83435.73, 80665.24, 79883.08, 80580.35, 82890.24, 81806.22, 
    93041.52,
  92248.84, 88756.92, 93846.87, 92464.73, 85831.96, 84780.31, 87137.39, 
    86458.47, 81442.61, 79172.23, 78283.34, 79020.69, 80461.44, 82107.27, 
    95149.66,
  85992.11, 86116.49, 85227.34, 83615.8, 83366.68, 81888.93, 82844.22, 
    83201.2, 80871.16, 79624.38, 79287.74, 80867.89, 80557.84, 82623.95, 
    88935.97,
  87606.12, 86616.88, 87693.47, 86863.73, 86770.15, 85162.1, 84147.18, 
    83704.76, 82767.05, 84789.56, 100068.8, 100755.7, 90821.99, 91252.72, 
    83832.82,
  87878.45, 86072.01, 88585.48, 89469.92, 88629.75, 88215.43, 87517.66, 
    87925.49, 89573.05, 100791, 101738.6, 101732.2, 101569.7, 93434.73, 
    78131.91,
  87031.68, 86290.18, 88439.08, 89751.66, 89570.41, 89671.35, 89635.82, 
    91679.59, 95703.47, 101515.3, 101538.4, 101663.3, 101600.3, 87191.96, 
    77851.52,
  90913.8, 87561.68, 88015.17, 89882.62, 89567.46, 88596.49, 89256.76, 
    91188.34, 95491.34, 101510.5, 101555, 101682.4, 101625.6, 85980.66, 
    87947.95,
  93979.34, 89562.77, 88622.58, 89745.82, 88914.77, 86555.22, 87889.42, 
    90540.59, 100894.2, 101472.2, 101461.3, 101554.9, 101614.4, 93637.48, 
    96431.41,
  97245.51, 92506.34, 90831.11, 93328.69, 93609.3, 93700.37, 94676.35, 
    100831.9, 101473.8, 101424.1, 101415.6, 101460, 101558.4, 99317.56, 
    100536.7,
  102214.1, 101872.2, 97838.65, 95279.16, 95282.62, 94111.56, 91689.6, 
    92183.6, 86115.95, 81375.42, 79034.11, 79399.29, 82566.41, 81095.03, 
    91903.69,
  102202.8, 102117.6, 99888.2, 94539.91, 91634.67, 89651.69, 88415.67, 
    88662.85, 83555.72, 80793.07, 79966.17, 80683, 83035.93, 81889.3, 93342.27,
  92841.05, 89289.07, 94355.41, 92979.33, 86276.34, 85154.02, 87482.88, 
    86736.05, 81656.59, 79360.38, 78438.54, 79177.46, 80634.97, 82303.53, 
    95453.76,
  86675.63, 86796.13, 85841.4, 84120.29, 83859.93, 82335.39, 83201.86, 
    83519.99, 81143.18, 79836.66, 79487.72, 81058.88, 80719.2, 82826.95, 
    89187.91,
  88279.55, 87252.32, 88312.46, 87489.4, 87334.24, 85704.05, 84615.34, 
    84095.88, 83084.35, 85191.46, 100624.4, 101242.2, 91108.3, 91544.9, 
    84019.86,
  88597.88, 86750.47, 89251.05, 90127.31, 89216.16, 88765.1, 88019.01, 
    88416.98, 90047.7, 101347.1, 102178.7, 102186.1, 101981.5, 93730.91, 
    78307.67,
  87693.55, 86947.98, 89090.81, 90406.96, 90183.27, 90213.1, 90153.95, 
    92166.05, 96235.21, 102102.5, 102025.8, 102061.2, 101988, 87489.52, 
    78031.55,
  91525.7, 88235.17, 88682.07, 90577.51, 90245.54, 89228.38, 89851.12, 
    91681.24, 96093.72, 102095.3, 102054.8, 102097.7, 102006.3, 86257.45, 
    88236.3,
  94515.98, 90162.43, 89237.07, 90380.49, 89554.59, 87160.18, 88459.4, 
    91151.85, 101651.3, 102120.2, 102052, 102057.1, 102048.5, 93969.51, 
    96794.58,
  97721.57, 93045.69, 91431.38, 93897.28, 94190.33, 94372.03, 95336, 
    101562.3, 102169.9, 102146.2, 102117.4, 102080.3, 102088.8, 99721.06, 
    100977.7,
  102424, 102157.3, 98115.62, 95532.86, 95503.79, 94380.44, 91918.59, 
    92465.18, 86357.06, 81647.4, 79286.5, 79614.06, 82825.19, 81305.6, 
    92233.65,
  102495.9, 102425.9, 100140.2, 94809.23, 91903.02, 89948.98, 88709.95, 
    88966.9, 83824.02, 81081, 80235.21, 80943.7, 83271.23, 82086.05, 93750.06,
  93154.95, 89576.19, 94639.3, 93179.38, 86587.05, 85457.02, 87794.28, 
    87013.84, 81959.79, 79656.05, 78637.64, 79422.81, 80884.89, 82553.08, 
    95883.73,
  86971.98, 87101.69, 86161.56, 84459.52, 84206.41, 82673.59, 83549.58, 
    83872.07, 81461.28, 80085.47, 79839.63, 81399.56, 80907.43, 83090.18, 
    89505.33,
  88595.94, 87558.2, 88620.71, 87805.7, 87654.67, 86043.01, 84950.64, 
    84466.34, 83421.02, 85637.59, 101148.1, 101771.1, 91542.59, 92006.28, 
    84250.02,
  88876, 87040.96, 89555.46, 90439.55, 89539.05, 89112.88, 88376.64, 88809.8, 
    90469.1, 101806.1, 102732, 102753.8, 102557.4, 94153.34, 78523.29,
  87933.31, 87212.41, 89380.76, 90710.53, 90516.83, 90568.71, 90539.25, 
    92557.3, 96642.64, 102649.3, 102651.5, 102638.5, 102618.5, 87834.55, 
    78291.03,
  91658.72, 88441.8, 88927.41, 90828.57, 90539.02, 89540.47, 90212.8, 
    92070.1, 96481.65, 102596.5, 102627.1, 102689.6, 102616, 86587.52, 
    88730.31,
  94589.2, 90312.1, 89433.16, 90600.85, 89842.87, 87488.73, 88816.32, 
    91496.77, 101890.7, 102583.8, 102599.4, 102646, 102637.9, 94449.41, 
    97309.62,
  97726.48, 93112.13, 91528.69, 94005.83, 94334.83, 94539.95, 95532.16, 
    101658.6, 102384.5, 102546.4, 102590.6, 102634.8, 102636, 100272, 101583.4,
  102402.3, 102109, 98142.3, 95637.77, 95651.79, 94570.09, 92104.85, 
    92705.14, 86612.88, 81850.34, 79456.17, 79765.38, 83020.27, 81560.73, 
    92553.29,
  102415.6, 102458.8, 100101.9, 94829.76, 91996.25, 90072.55, 88853.48, 
    89156.66, 84012.58, 81265.72, 80446.51, 81136.62, 83487.3, 82369.75, 
    94049.28,
  93212.88, 89615.06, 94702.94, 93322.34, 86670.12, 85567.56, 87872.23, 
    87135.15, 82102.22, 79778.48, 78712.61, 79490.52, 81023.57, 82797.46, 
    96154.12,
  87016.79, 87053.76, 86179.7, 84517.06, 84252.9, 82751.95, 83607.32, 
    83945.95, 81549.29, 80154.42, 79979.77, 81509.01, 81012.95, 83344.49, 
    89778.23,
  88704.26, 87542.91, 88628.09, 87829.85, 87675.18, 86059.2, 84987.92, 
    84489.62, 83459.69, 85685.53, 100903.6, 101565.9, 91539.16, 92156.49, 
    84502.29,
  88894.47, 87052.54, 89549.36, 90457.65, 89542.93, 89101.3, 88373.16, 
    88795.88, 90420.71, 101550.4, 102582.9, 102617.8, 102514.5, 94265.97, 
    78755.06,
  87930.39, 87224, 89365, 90688.97, 90499.89, 90541.45, 90478.1, 92483.71, 
    96493.41, 102391.2, 102488.9, 102508.4, 102638.7, 87906.27, 78459.83,
  91692.67, 88450.51, 88918.68, 90785.96, 90504.13, 89481.58, 90125.8, 
    91985.07, 96290.8, 102349.4, 102457.8, 102594.2, 102588.5, 86693.84, 
    88840.31,
  94678.24, 90370.95, 89449.17, 90594.32, 89835.95, 87476.84, 88777.31, 
    91393.53, 101674.4, 102319.9, 102402.2, 102546.2, 102616.5, 94570.11, 
    97386.73,
  97877.89, 93209.51, 91552.86, 94007.12, 94319.55, 94486.5, 95441.86, 
    101509.1, 102150.3, 102249.4, 102359.4, 102495.5, 102639.6, 100333.3, 
    101690.2,
  102239.9, 101968.6, 98164.61, 95707.27, 95738.56, 94699.51, 92243.02, 
    92832.06, 86727.91, 81956.73, 79588.9, 79880.41, 83080.7, 81602.41, 
    92604.58,
  102255.5, 102309, 100029.9, 94837.49, 92078.77, 90171.85, 88921.73, 
    89268.89, 84139.27, 81340.2, 80481.88, 81191.34, 83551.54, 82416.99, 
    94051.23,
  93159.52, 89647.23, 94741.25, 93364.23, 86743.57, 85646.67, 87978.71, 
    87232.68, 82200.45, 79876.84, 78804.73, 79571.96, 81078.04, 82829.73, 
    96162.26,
  86947.06, 87065.18, 86206.6, 84546.77, 84306.52, 82811.35, 83697.18, 
    84020.06, 81642.84, 80235.95, 79994.75, 81584.1, 81048.92, 83360.15, 
    89779.28,
  88578, 87576.47, 88675.98, 87871.5, 87763.93, 86151.29, 85094.76, 84590.7, 
    83555.84, 85697.96, 100992.6, 101508.6, 91587.61, 92110.38, 84559.56,
  88901.88, 87094.03, 89625.2, 90516.51, 89620.84, 89193.88, 88463.07, 
    88872.45, 90493.16, 101632.2, 102540.2, 102548.2, 102438, 94220.72, 
    78802.02,
  88053.92, 87321.84, 89488.81, 90804.55, 90592.98, 90653.22, 90583.66, 
    92604.65, 96624.57, 102451.5, 102475.4, 102517.8, 102573.8, 87921.71, 
    78484.81,
  91885.5, 88600.79, 89091.14, 90962.16, 90643.88, 89626.04, 90270.37, 
    92133.66, 96452.62, 102436.9, 102487.7, 102601.9, 102530.1, 86695.98, 
    88798.26,
  94878.17, 90537.16, 89628.94, 90773.13, 89969.46, 87609.81, 88930.26, 
    91578.7, 101917.8, 102428.5, 102462.3, 102585.5, 102584.5, 94579.3, 
    97348.78,
  98185.72, 93499.94, 91844.44, 94308.6, 94574.66, 94742.51, 95710.12, 
    101829.2, 102396.1, 102398.9, 102446.5, 102561.8, 102627.1, 100350.3, 
    101660.7,
  102028.3, 101846.9, 98015.3, 95547.03, 95535.73, 94475.93, 92037.85, 
    92606.69, 86545.42, 81773.52, 79411.95, 79695.52, 82753.15, 81353.41, 
    92120.57,
  102136.8, 102207.1, 99866.77, 94684.87, 91929.06, 90004.55, 88732.4, 
    89057.55, 83940.03, 81178.2, 80332.9, 80998, 83275.51, 82146.07, 93629.59,
  92961.96, 89528.3, 94651.62, 93238.68, 86570.3, 85493.83, 87849.24, 
    87057.55, 82047.53, 79750.82, 78702.56, 79427.92, 80864.81, 82548.55, 
    95860.99,
  86787.57, 86963.88, 86064.69, 84420.63, 84179.69, 82680.76, 83596.82, 
    83897.52, 81501.31, 80120.3, 79882.3, 81505.34, 80892.51, 83095.44, 
    89435.32,
  88432.65, 87495.66, 88608.89, 87791.94, 87694.31, 86048.4, 85006.59, 
    84500.12, 83447.93, 85632.77, 101110.9, 101553.9, 91562.26, 91931.99, 
    84216.99,
  88816.48, 86949.14, 89539.25, 90413.07, 89550.65, 89137.47, 88412.9, 
    88816.77, 90503.57, 101832.1, 102607.6, 102585.2, 102384.3, 94047.61, 
    78523.23,
  87981.22, 87224.02, 89454.18, 90746.64, 90558.41, 90629.35, 90600.27, 
    92641.13, 96792.43, 102611.7, 102538.2, 102527.9, 102530.6, 87753.02, 
    78303.39,
  91766.64, 88500.04, 89044.32, 90918.88, 90623.95, 89627.6, 90307.31, 
    92201.91, 96660.59, 102612.2, 102567.2, 102615.6, 102479.1, 86520.8, 
    88704.13,
  94808.05, 90483.87, 89637.15, 90774.42, 89973.17, 87634.7, 88955.41, 
    91698.65, 102227.5, 102647.9, 102573.2, 102613.8, 102538.6, 94529.49, 
    97315.51,
  98064.47, 93378.54, 91851.71, 94353.06, 94617.48, 94823.57, 95879.69, 
    102108.5, 102692.5, 102675.7, 102630.3, 102625, 102613.3, 100334.7, 
    101702.4,
  101857.1, 101651.1, 97793.67, 95320.94, 95305.35, 94264.52, 91851.69, 
    92416.67, 86391.04, 81638.8, 79260.1, 79551.73, 82526.86, 81109.8, 
    91741.37,
  102022.8, 102012, 99658.18, 94482.11, 91721.33, 89799.21, 88546.7, 
    88884.82, 83800.13, 81035.27, 80185.53, 80856.87, 83087.55, 81922.85, 
    93181.79,
  92773.83, 89362.13, 94449.17, 93025.45, 86382, 85304.41, 87643.75, 
    86874.24, 81884.01, 79574.26, 78516.73, 79225.46, 80656.7, 82253.16, 
    95383.02,
  86625.08, 86830.82, 85860.77, 84241.32, 83997.49, 82503.15, 83398.43, 
    83711.62, 81325.65, 79962.77, 79699.91, 81321.78, 80717.8, 82822.73, 
    89001.41,
  88271.84, 87403.02, 88464.16, 87634.98, 87497.98, 85856.58, 84821.09, 
    84312.77, 83288.8, 85475.31, 100961.3, 101504.1, 91395.45, 91714.84, 
    83876.16,
  88658.45, 86799.17, 89442.19, 90289.31, 89415.48, 88951.01, 88221.94, 
    88640.25, 90326.09, 101769.2, 102576.7, 102548.2, 102281.6, 93890.58, 
    78154.3,
  87877.81, 87071.92, 89323.89, 90612.96, 90424.88, 90469.23, 90441.24, 
    92527.48, 96691.17, 102592.2, 102462, 102403.6, 102352.4, 87550.33, 
    77941.17,
  91621, 88348.45, 88919.58, 90774.82, 90495.49, 89483.86, 90179, 92026.3, 
    96551.36, 102623.6, 102528.8, 102478.2, 102310.6, 86228.59, 88367.75,
  94634.73, 90334.87, 89479.9, 90634.57, 89834.63, 87474.96, 88789.43, 
    91560.45, 102211.8, 102701.8, 102601.8, 102538.7, 102327.2, 94299.65, 
    97274.21,
  97839.7, 93197.45, 91671.18, 94209.05, 94492.07, 94675.34, 95719.25, 
    102041.7, 102754.9, 102803.7, 102788.1, 102790.1, 102666.6, 100392.5, 
    101814.8,
  101531.1, 101305, 97472.28, 95026.04, 95042.89, 94001.33, 91603.78, 
    92145.27, 86149.75, 81355.52, 78957.86, 79255.98, 82217.23, 80823.01, 
    91338.97,
  101545.5, 101623.6, 99325.05, 94167.79, 91423.6, 89514.15, 88258.84, 
    88561.71, 83504.35, 80684.56, 79854.74, 80538.89, 82765.3, 81643.36, 
    92744.98,
  92498.64, 89023.54, 94083.48, 92702.97, 86106.22, 85009.24, 87303.23, 
    86566.7, 81540.23, 79225.91, 78197.9, 78889.75, 80310.17, 81938.47, 
    94959.78,
  86295.26, 86436.51, 85577.13, 83944.95, 83699.38, 82196.66, 83042.04, 
    83351, 80970.26, 79614.99, 79303.95, 80885.6, 80383.29, 82471.36, 88694.07,
  87911.62, 86958.36, 88060.29, 87261.19, 87151.27, 85524.17, 84435.94, 
    83928.96, 82884.56, 85100.68, 100745.7, 101412.8, 91094.9, 91387.46, 
    83677.6,
  88256.45, 86418.2, 89005.5, 89906.5, 89044.56, 88597.8, 87895.62, 88361.8, 
    90079.93, 101708.2, 102531.9, 102473.9, 102108.5, 93667.3, 77827.43,
  87392.09, 86652.78, 88901.92, 90229.47, 90066.84, 90140.62, 90171.75, 
    92291.57, 96546.59, 102566.6, 102340.4, 102242.7, 102103, 87297.31, 
    77541.48,
  91098.3, 87900.06, 88484.38, 90397.72, 90126.69, 89138.34, 89880.91, 
    91784.81, 96476.26, 102591.5, 102440.6, 102337.8, 102048, 85930.41, 
    87858.23,
  94094.78, 89858.16, 89052.2, 90247.99, 89463.92, 87152.85, 88467.58, 
    91465.2, 102239.1, 102715.3, 102550.3, 102419.6, 102138.9, 93946.79, 
    96989.48,
  97285.32, 92711.5, 91232.24, 93807.18, 94106.55, 94374.5, 95568.74, 
    102060.2, 102765.2, 102846.5, 102772.1, 102742.2, 102605, 100224.4, 
    101583.2,
  100408.7, 100152.1, 96300.64, 93868.9, 93884.93, 92896.77, 90603.97, 
    91134.26, 85290.52, 80563.09, 78255.76, 78599.63, 81614.36, 80288.68, 
    90775.17,
  100538.9, 100530.7, 98235.04, 93095.04, 90372.08, 88518.52, 87258.2, 
    87620.48, 82666.8, 79870.62, 79103.15, 79815.4, 82095.52, 81080.97, 
    92128.88,
  91493.92, 88054.84, 93070.95, 91679.05, 85121.97, 84082.02, 86408.12, 
    85685.69, 80692.01, 78438.29, 77561.12, 78276.13, 79711.35, 81334.52, 
    94298.06,
  85510.69, 85683.09, 84738.98, 83081.65, 82832.18, 81357.71, 82252.12, 
    82568.77, 80195.64, 78966.6, 78670.31, 80260.92, 79837.02, 81917.11, 
    88155.75,
  87167.63, 86296.05, 87394.3, 86571.74, 86443.2, 84809.4, 83773.28, 
    83291.88, 82307.89, 84565.26, 100331.7, 100981.4, 90582.29, 90782.64, 
    83159.06,
  87578.53, 85833.72, 88444.36, 89318.99, 88463.5, 88072.59, 87366.59, 
    87839.34, 89596.62, 101241.8, 102105.2, 102044.3, 101748.2, 93214.6, 
    77476.66,
  86834.59, 86142.8, 88424.16, 89748.77, 89612.66, 89693.69, 89739.95, 
    91877.77, 96093.07, 102032.3, 101822.2, 101825.4, 101713.5, 86892.23, 
    77101.45,
  90641.75, 87443.3, 88034.45, 89950.91, 89699.38, 88739.48, 89471.64, 
    91354.83, 96035.65, 102081.6, 101925.9, 101912.1, 101798.9, 85541.44, 
    87514.93,
  93744.38, 89467.55, 88666.77, 89841.72, 89039.87, 86692.42, 88098.83, 
    91171.67, 101798.3, 102208.6, 102026.7, 101938.5, 101829.2, 93680.9, 
    96731.18,
  97072.7, 92434.21, 91043.2, 93584.63, 93907.29, 94177.88, 95393.03, 
    101736.3, 102360.6, 102414, 102297, 102266.6, 102171.4, 99859.51, 101200.5,
  100948.4, 100664.4, 96507.28, 93773.73, 93619.78, 92384.2, 89898.43, 
    90262.89, 84364.41, 79693.61, 77462.02, 77868.38, 81011.38, 79592.99, 
    90295.27,
  101175.9, 100957.8, 98589.35, 93183.84, 90157.56, 88140.98, 86826.34, 
    86987.25, 81936.09, 79200.91, 78398.2, 79144.38, 81483.17, 80435.06, 
    91665.16,
  91640.99, 88243.38, 93161.65, 91545.91, 84827.2, 83776.04, 86064.38, 
    85182.32, 80133.89, 77941.04, 77086.23, 77849.87, 79270.17, 80907.3, 
    93752.09,
  85742.58, 85919.09, 84851.23, 83129.23, 82765.52, 81155.66, 82011.8, 
    82249.16, 79842.9, 78612.15, 78372.17, 79893.85, 79490.2, 81569.88, 
    87624.73,
  87398.24, 86487.33, 87552.27, 86686.67, 86479.08, 84763.53, 83647.27, 
    83066.02, 82046.44, 84366.41, 100101.1, 100612, 90253.12, 90485.17, 
    82679.65,
  87840.32, 86112.62, 88729.76, 89535.84, 88610.21, 88116.47, 87341.26, 
    87712.53, 89521.21, 100940.7, 101641.6, 101559.8, 101415.9, 92723.56, 
    77155.05,
  87111.41, 86383.75, 88637.14, 89933.77, 89747.41, 89750.25, 89729.11, 
    91752.17, 95925.8, 101743.7, 101552.6, 101444.9, 101353, 86508.82, 76906.7,
  90997.35, 87716.09, 88290.16, 90187.44, 89841.16, 88788.24, 89458.08, 
    91300.27, 95977.98, 101930.5, 101688.3, 101592.6, 101336.6, 85311.32, 
    87318.93,
  94142.21, 89742.98, 88906.01, 90077.77, 89216.1, 86803.51, 88149.57, 
    91116.54, 101675.3, 102102.8, 101896.1, 101794.6, 101472.8, 93437.27, 
    96490.69,
  97488.3, 92713.29, 91240.14, 93774.02, 94083.75, 94259.7, 95360.67, 
    101642.8, 102233.4, 102264.5, 102118.4, 102100.5, 101964.9, 99649.58, 
    100948.9,
  101577.3, 101273.1, 97152.83, 94411.91, 94302.1, 93118.28, 90634, 91161.68, 
    85062.76, 80268, 77839, 78154.72, 81246.41, 79786.98, 90295.56,
  101610, 101440.9, 99149.14, 93743.2, 90761.51, 88736.18, 87428.62, 
    87647.45, 82501.71, 79738.29, 78861.45, 79570.47, 81802.7, 80651.28, 
    91874.44,
  92150.27, 88613.54, 93579.28, 92065.36, 85337.68, 84245.21, 86551.23, 
    85705.18, 80613.44, 78347.07, 77373.89, 78133.38, 79477.36, 81141.33, 
    93992.38,
  86052.84, 86218.03, 85195.95, 83447.75, 83119.45, 81520.68, 82366.95, 
    82644.33, 80214.16, 78867.99, 78581.65, 80184.49, 79647.62, 81815.09, 
    87777.59,
  87659.81, 86684.3, 87739.35, 86891.67, 86702.45, 85004.35, 83866.96, 
    83300.59, 82217.2, 84559.98, 100273.6, 100802.8, 90450.91, 90797.47, 
    82776.43,
  88063.61, 86204.79, 88756.24, 89619.73, 88700.12, 88216.7, 87451.18, 
    87828.09, 89570.64, 100958, 101784.3, 101730.1, 101596.3, 92966.08, 
    77224.98,
  87203.55, 86422.02, 88586.81, 89913.4, 89722.59, 89736.86, 89666.64, 
    91659.71, 95816.28, 101764.1, 101677.2, 101539.7, 101523.8, 86620.58, 
    77008.52,
  91073.15, 87733.51, 88206.95, 90069.81, 89746.13, 88703.94, 89355.73, 
    91178.64, 95740.75, 101791, 101668.7, 101596, 101514, 85435.45, 87416.59,
  94122.47, 89708.2, 88770.11, 89908.59, 89066.92, 86640.27, 87920.54, 
    90686.28, 101287.9, 101832, 101706.4, 101611.3, 101437.9, 93295.24, 
    96249.58,
  97404.05, 92664.73, 91016.12, 93492.04, 93765.7, 93930.83, 94908.98, 
    101140.4, 101828.8, 101862.5, 101815, 101781.4, 101694, 99343.3, 100632.4,
  101820.9, 101515.8, 97537.62, 94995.35, 95007.93, 93955.33, 91534.88, 
    92070.62, 86004.23, 81159.66, 78729.41, 78994.94, 81943.87, 80437.4, 
    90902.55,
  101742.6, 101743.8, 99441.83, 94174.91, 91343.19, 89412.97, 88165.84, 
    88467.62, 83328.72, 80475.95, 79607.2, 80275.12, 82483.03, 81289.24, 
    92432.93,
  92500.4, 88901.49, 93976.75, 92612.28, 85928.24, 84811.66, 87179.73, 
    86444.16, 81346.77, 79015.72, 77984.73, 78687.18, 80040, 81666.27, 
    94575.27,
  86197.44, 86329.95, 85423.11, 83728.33, 83450.75, 81935.11, 82804.86, 
    83141.27, 80765.62, 79407.8, 79092.02, 80676.76, 80143.55, 82269.16, 
    88319.93,
  87807.72, 86818.41, 87879.76, 87055.98, 86912.02, 85280.09, 84191.01, 
    83677.37, 82675.19, 84801.13, 100373.7, 101032.2, 90814.58, 91176.45, 
    83299.66,
  88115.98, 86296.03, 88828.54, 89722.92, 88807.33, 88364.47, 87613.45, 
    88029.79, 89683.42, 101154.7, 102074.2, 102075.3, 101824.9, 93393.18, 
    77583.62,
  87272.43, 86526.33, 88710.55, 90022.02, 89789.61, 89834.69, 89769.99, 
    91859.94, 96027.28, 102018.1, 101932.6, 101992.3, 101884.1, 87052.82, 
    77332.26,
  91104.39, 87820.2, 88344.44, 90245.39, 89917.88, 88879.03, 89538.81, 
    91451.68, 95890.09, 102033.8, 101983, 102063.3, 101888.9, 85788.79, 
    87667.26,
  94195.82, 89828.76, 88952.59, 90134.06, 89291.49, 86837.52, 88179.34, 
    90934.44, 101570.8, 102092.3, 102005.7, 102011.2, 101904.9, 93677.48, 
    96400.88,
  97498.8, 92811.63, 91257.23, 93831.88, 94131.52, 94326.54, 95321.92, 
    101579, 102128.9, 102111, 102094.4, 102072.8, 101999.2, 99575.21, 100789,
  101715, 101422.3, 97484.31, 94934.23, 94957.52, 94008.71, 91689.65, 
    92263.7, 86242, 81372.11, 78965.3, 79269.3, 82242.9, 80827.63, 91285.31,
  101709.3, 101652.8, 99392.64, 94159.88, 91357.91, 89476.02, 88233.25, 
    88610.47, 83538.12, 80663.16, 79847.93, 80543.27, 82793.17, 81679.93, 
    92833.2,
  92450.5, 88944.29, 93996.75, 92613.81, 85968.1, 84889.98, 87291.93, 
    86612.13, 81539.38, 79205.08, 78229.76, 78933.35, 80347.51, 81970.51, 
    95003.09,
  86326.19, 86526.68, 85556.02, 83854.15, 83562.11, 82035.78, 82914.23, 
    83288.34, 80904.09, 79608.57, 79314.29, 80905.21, 80443.67, 82496.46, 
    88685.55,
  87972.92, 87082.38, 88156.45, 87323.24, 87148.67, 85487.24, 84400.52, 
    83910.1, 82925.87, 85148.18, 100939.6, 101639.4, 91219.2, 91464.86, 
    83722.66,
  88415.36, 86606.4, 89209.59, 90081.17, 89135.77, 88688.05, 87943.44, 
    88405.88, 90146.34, 101875.6, 102785.9, 102685.4, 102321.8, 93746.13, 
    77859.11,
  87615.54, 86868.87, 89138.47, 90456.17, 90238, 90277.35, 90253.32, 
    92434.46, 96702.91, 102751.8, 102609.2, 102630, 102413.1, 87374.33, 
    77559.9,
  91499.14, 88185.02, 88741.03, 90653.48, 90339.55, 89293.55, 89997.84, 
    91895.7, 96495.16, 102771.4, 102708.6, 102740.3, 102458.3, 85998.39, 
    87970.74,
  94628.8, 90201.74, 89327.68, 90510.78, 89659.44, 87237.88, 88589.34, 
    91458.73, 102252.9, 102815, 102736.6, 102763.1, 102534.3, 94203.31, 
    97071.48,
  97997.15, 93186.12, 91647.99, 94233.1, 94528.58, 94717.15, 95747.09, 
    102090.7, 102741.5, 102844.4, 102824.8, 102860, 102771.7, 100326.1, 
    101543.5,
  102199.2, 101913.7, 97861.64, 95276.11, 95269.77, 94235.27, 91822.95, 
    92363.5, 86313.05, 81450.85, 79034.64, 79329.1, 82320.88, 80926.26, 
    91557.69,
  102180.8, 102149.6, 99868.4, 94527.84, 91653.38, 89710.04, 88458.71, 
    88764.4, 83645.77, 80792.66, 79953.88, 80630.5, 82872.87, 81731.17, 
    93038.04,
  92878.81, 89295.47, 94253.97, 92919.47, 86232.61, 85103.48, 87456.97, 
    86733.61, 81663.13, 79305.65, 78251.21, 78955, 80400.26, 82015.84, 
    95167.52,
  86679.02, 86761.4, 85794.89, 84083.06, 83754.83, 82224.54, 83069.98, 
    83421.95, 81009.21, 79653.41, 79363.86, 80950.55, 80407.56, 82547.1, 
    88807.3,
  88245.77, 87201.27, 88213.55, 87380.06, 87176.44, 85531.78, 84418.2, 
    83898.46, 82879.77, 85000.54, 100379, 101122.1, 91016.16, 91418.3, 
    83651.56,
  88564.84, 86707.34, 89157.63, 90034.24, 89078.49, 88591.6, 87786.92, 
    88175.62, 89763.24, 101080.1, 102207.6, 102242.8, 101978.3, 93619.84, 
    77871.77,
  87672.42, 86892.32, 88979.58, 90281.26, 90020.98, 90014.69, 89908.02, 
    91903.84, 95972.09, 101980.3, 102010.7, 102072.1, 102050.4, 87231.46, 
    77587.31,
  91518.92, 88174.55, 88554.8, 90383.57, 90026.2, 88934.16, 89511.36, 
    91351.3, 95718.19, 101858.8, 101922.9, 102102.9, 102006.7, 85915, 87857.86,
  94537.6, 90086.34, 89070.8, 90147.77, 89291.02, 86846.91, 88077.3, 90717, 
    101074.4, 101764.5, 101809.1, 101974.9, 101975.1, 93809.6, 96550.55,
  97780.79, 93006.01, 91272.15, 93620.4, 93839.84, 93974.84, 94850.73, 
    100945.1, 101589.2, 101655.7, 101736.1, 101872.2, 101988.7, 99641.41, 
    100937,
  102030.7, 101672.3, 97639.67, 94965.6, 94902.89, 93852.59, 91441.58, 
    91935.14, 85992.52, 81126.38, 78684.7, 78964.55, 81859.67, 80482.04, 
    90727.24,
  101951.5, 101773.2, 99544.91, 94245.91, 91320.45, 89337.8, 88050.98, 
    88316.6, 83269.92, 80380.11, 79539.12, 80180.27, 82362.74, 81268.02, 
    92173.19,
  92684.12, 89054.84, 93922.11, 92567.51, 85920.2, 84772.59, 87060.12, 
    86327.43, 81296.2, 78960.29, 77949.56, 78578.68, 79927.05, 81493.44, 
    94247.52,
  86581.7, 86592.86, 85667.67, 83907.12, 83577.3, 82015.3, 82797.45, 
    83094.42, 80690.4, 79368.85, 79067.01, 80610.48, 80033.29, 81992.59, 
    88074.41,
  88158.34, 87046.66, 88092.41, 87254.56, 87028.76, 85365.6, 84240.65, 83712, 
    82664.18, 84826.85, 100196.3, 100860.1, 90605.51, 90770.57, 83149.55,
  88435.05, 86595.42, 89088.12, 89931.37, 88951.98, 88462.23, 87658.35, 
    88059.13, 89700.8, 101046.9, 101830.1, 101703.2, 101352.9, 92954.95, 
    77312.58,
  87598.06, 86822.52, 88950.96, 90234.77, 89973.1, 89956.62, 89889.91, 
    91901.67, 95993.95, 101816.1, 101601.9, 101541.5, 101339.4, 86673.38, 
    76914.94,
  91447.99, 88108.47, 88593.25, 90457.99, 90074.11, 88982.55, 89591.37, 
    91379.16, 95877.44, 101803.8, 101610.9, 101559.8, 101292.9, 85276.2, 
    87093.51,
  94534.42, 90116.27, 89211.44, 90378.95, 89480.97, 87005.66, 88257.41, 
    91075, 101514, 101813.5, 101602.5, 101538.1, 101327.4, 93205.48, 95868.2,
  97887.13, 93154.36, 91598.85, 94118.84, 94396.41, 94581.13, 95497.21, 
    101638, 101989.5, 101812.5, 101670, 101586.4, 101457.9, 99066.55, 100207.7,
  102133.1, 101943.9, 97871.21, 95293.46, 95256.41, 94102.7, 91612.66, 
    92087.59, 85935.33, 81199.17, 78818.27, 79178.07, 82218.71, 80747.67, 
    91473.98,
  102312.1, 102197.3, 99923.07, 94616.41, 91702.93, 89720.12, 88476.92, 
    88660.65, 83452.93, 80716.39, 79883.91, 80639.44, 82856.82, 81658.13, 
    93010.6,
  92800.66, 89444.96, 94466.75, 92976.99, 86263.74, 85225.61, 87580.48, 
    86734.94, 81622.87, 79296.76, 78228.72, 79015.58, 80421.15, 82067.07, 
    95191.59,
  86768.14, 87005.66, 86005.71, 84320.38, 84043.78, 82463.22, 83351.24, 
    83659.62, 81169.62, 79768.23, 79639.52, 81243.73, 80575.99, 82765.71, 
    88835.59,
  88403.12, 87481.93, 88584.74, 87751.18, 87573.88, 85915.07, 84826.64, 
    84313.44, 83236.11, 85610.41, 101381.6, 101906.5, 91545.23, 91844.88, 
    83704.66,
  88805.29, 87013.2, 89672.69, 90549, 89632.08, 89151.9, 88414.12, 88820.23, 
    90605.11, 102103.7, 103029.8, 103015, 102770.7, 94013.31, 77979.34,
  87969.48, 87230.73, 89529.57, 90883.3, 90693.77, 90731.19, 90696.68, 
    92751.45, 96958.11, 102954.9, 102960.8, 102876.5, 102853.2, 87497.59, 
    77819.46,
  91776.52, 88514.79, 89106.28, 91062.65, 90748.66, 89696.12, 90361.77, 
    92254.95, 96833.95, 102948.1, 102929.7, 102963.1, 102804.2, 86272.57, 
    88375.27,
  94845.98, 90497.8, 89651.57, 90868.05, 90066.04, 87665.86, 88993.7, 
    91815.11, 102433.6, 102970.3, 102900.2, 102935.3, 102789.2, 94517.6, 
    97138.35,
  98130.28, 93425.96, 91924.82, 94478.68, 94798.37, 94972.46, 96011.6, 
    102328, 102934.9, 102967.6, 102889.4, 102886.7, 102799.8, 100373.2, 
    101482.1,
  102245.8, 102026.8, 98135.73, 95644.9, 95633.45, 94557.88, 92137.98, 
    92681.28, 86592.66, 81793.31, 79374.29, 79660.31, 82674.94, 81204.45, 
    91814.52,
  102251.2, 102375.1, 100028.6, 94756.48, 91954.89, 90032.47, 88797.95, 
    89106.08, 83980.7, 81158.41, 80309.48, 80981.75, 83229.39, 82046.64, 
    93309.24,
  92994.05, 89483.01, 94623.96, 93214.23, 86536.64, 85433.51, 87800.45, 
    87081.61, 82012.14, 79656.52, 78593.21, 79301.02, 80720.23, 82342.53, 
    95441.33,
  86790.47, 86774.08, 86005.32, 84331.88, 84040.23, 82539.8, 83423.23, 
    83797.47, 81387.23, 80020.73, 79745.94, 81321.93, 80753.14, 82880.8, 
    89069.21,
  88426.36, 87190.01, 88350.54, 87546.04, 87426.09, 85816.82, 84757.22, 
    84277.33, 83270.2, 85393.33, 100691.1, 101423.3, 91360.81, 91749.2, 
    83957.33,
  88623.24, 86729.27, 89237.88, 90149.39, 89282.41, 88856.62, 88123.15, 
    88550.32, 90162.63, 101413.4, 102528.1, 102574.3, 102271, 93920.4, 78237.8,
  87601.93, 86904.2, 89051.32, 90401.05, 90209.79, 90286.69, 90230.75, 
    92276.42, 96319.83, 102331.2, 102346.3, 102400.4, 102387, 87568.02, 
    77953.85,
  91261.38, 88113.91, 88612.34, 90487.91, 90225.82, 89248.41, 89895.08, 
    91781.27, 96121.87, 102250.6, 102295.5, 102465.8, 102367.4, 86256.04, 
    88235.26,
  94192.67, 89987.16, 89144.27, 90280.87, 89549.51, 87192.95, 88493.23, 
    91160.6, 101621.2, 102244.1, 102254.5, 102395.1, 102356.9, 94252.71, 
    96869.57,
  97358.59, 92803.28, 91279.65, 93735.07, 94079.83, 94277.64, 95286.28, 
    101533.2, 102166.3, 102200, 102251.1, 102350.2, 102391.6, 100037.1, 
    101214.5,
  101016.7, 100784.4, 97028.07, 94699.84, 94768.7, 93819.95, 91560.75, 
    92092.89, 86186.49, 81401.92, 79022.66, 79325.32, 82243.65, 80861.88, 
    91105.16,
  101173, 101222.3, 98913.23, 93808.96, 91179.47, 89373.09, 88164.8, 
    88531.25, 83548.37, 80707.59, 79894.84, 80576.59, 82789.96, 81687.98, 
    92632.8,
  92106.44, 88689.73, 93748.95, 92374.07, 85875.07, 84813.64, 87205.86, 
    86533.96, 81543.42, 79240.84, 78295.67, 78971.76, 80357.96, 81926.02, 
    94744.34,
  86018.18, 86110.62, 85272.52, 83646.49, 83407.2, 81961.38, 82911.16, 
    83260.34, 80923.96, 79632.5, 79295.41, 80847.16, 80428.62, 82431, 88552.77,
  87616.52, 86632.94, 87770.69, 86933.19, 86823.12, 85211.73, 84216.72, 
    83781.31, 82823.55, 84847.92, 100139.9, 100828.6, 90816.71, 91133.02, 
    83575.59,
  87975.71, 86169.74, 88730.89, 89622.65, 88739.53, 88294.49, 87572.23, 
    88005.32, 89641.93, 100909.8, 101965.2, 101877, 101612.5, 93365.66, 
    77897.38,
  87138.64, 86422.77, 88608.77, 89926.61, 89730.28, 89796.93, 89747.86, 
    91820.45, 95917.13, 101824.9, 101717.6, 101771.8, 101699.8, 87110.93, 
    77636.86,
  90947.63, 87699.17, 88220.73, 90085.81, 89794.56, 88787.5, 89433.23, 
    91325.45, 95721.24, 101797.7, 101769.2, 101901.1, 101755.3, 85837.51, 
    87854.51,
  93983.29, 89676.68, 88827.32, 89964.43, 89148.85, 86787.02, 88107.92, 
    90840.44, 101354.6, 101858.3, 101825.4, 101882, 101752.3, 93691.31, 
    96495.13,
  97216.7, 92573.89, 91071.28, 93558.13, 93818.02, 93977.73, 95045.68, 
    101269.2, 101871, 101918.5, 101932.3, 101970.8, 101937.1, 99600.74, 
    100835.5,
  101253.6, 101001, 96976.4, 94424.39, 94370.34, 93308.22, 90914.25, 
    91456.47, 85503.24, 80840.7, 78530.87, 78875.11, 81858.91, 80413.3, 
    90770.04,
  101382.1, 101283.3, 98938.42, 93674.55, 90842.91, 88934.23, 87695.51, 
    88010.65, 82969.67, 80251.47, 79429.78, 80152.38, 82382.71, 81237.08, 
    92324.23,
  92108.34, 88601.7, 93596.65, 92151.48, 85589.32, 84535.24, 86846.68, 
    86066.42, 81088.46, 78871.4, 77921.62, 78660.11, 79995.23, 81625.67, 
    94424.29,
  86028.63, 86246.23, 85271.76, 83567.46, 83278.47, 81769.46, 82675.03, 
    82989.86, 80633.33, 79285.84, 79002.09, 80626.05, 80115.67, 82258.52, 
    88225.99,
  87634.09, 86718.86, 87791.53, 86951.74, 86801.21, 85146.52, 84092, 
    83592.43, 82588.8, 84790.38, 100447.5, 100923.4, 90777.93, 91098.31, 
    83251.59,
  88024.7, 86208.44, 88799.59, 89636.53, 88732.77, 88290.84, 87574.73, 
    88013.03, 89746.88, 101158.2, 101985.5, 101947.9, 101746.3, 93256.4, 
    77642.88,
  87210.44, 86440.08, 88666.75, 89963.01, 89774.59, 89838.26, 89812.28, 
    91885.3, 96059.69, 101965.8, 101895.1, 101846.4, 101810.3, 86915.84, 
    77503.69,
  90988.52, 87717.2, 88262.83, 90139.23, 89831.02, 88818.57, 89526.84, 91406, 
    95933.36, 101998, 101940.9, 101947, 101770.1, 85709.27, 87809.46,
  94019.55, 89708.92, 88865.24, 90027.13, 89224.89, 86845.88, 88196.73, 
    90949.49, 101573, 102032.4, 101961.6, 101966.2, 101771.4, 93643.81, 
    96371.54,
  97300.58, 92627.74, 91136.7, 93676.59, 93956.96, 94120.04, 95188.84, 
    101456.9, 102046.7, 102077.2, 102022.8, 102031, 101962.4, 99582.45, 
    100742.8,
  101448.1, 101129.9, 97190.05, 94639.34, 94630.02, 93598.71, 91188.26, 
    91679.1, 85772.43, 81056.98, 78749.54, 79076.73, 82104.89, 80703.15, 
    91250.91,
  101386.1, 101375.2, 99086.29, 93843.91, 91064.47, 89153.02, 87895.59, 
    88194.41, 83186.43, 80422.48, 79642.87, 80357.84, 82621.95, 81527.26, 
    92750.85,
  92261.56, 88698.54, 93728.39, 92343.54, 85775.09, 84685.82, 87014.96, 
    86233.03, 81269.7, 79038.27, 78120.35, 78881.92, 80269.44, 81896.3, 
    94875.84,
  86017.31, 86203.88, 85324.67, 83614.68, 83376.47, 81874.96, 82785.38, 
    83101.38, 80746.77, 79459.44, 79110.2, 80748.95, 80343.24, 82501.71, 
    88639.28,
  87644.32, 86695.55, 87801.37, 86966.98, 86868.87, 85243.27, 84202.09, 
    83690.66, 82713.8, 84857.33, 100592.6, 101125.8, 90880.59, 91354.55, 
    83559.27,
  87955.98, 86159.38, 88742.92, 89649.1, 88767.1, 88326.7, 87615.79, 
    88040.72, 89792.09, 101323, 102234.1, 102234.7, 102025.8, 93525.3, 
    77919.34,
  87150.39, 86403.69, 88658.84, 89967.9, 89795.55, 89887.8, 89862.88, 
    91987.26, 96164.6, 102158.6, 102114.2, 102119, 102068.2, 87169.04, 
    77732.68,
  90959.12, 87683.71, 88247.34, 90125.35, 89864.34, 88879.86, 89560.69, 
    91512.2, 96004.34, 102169.1, 102162.1, 102246, 102096.2, 85967.94, 
    88030.38,
  93992.3, 89668.32, 88857.63, 90024.2, 89247.09, 86892.3, 88245.19, 
    90952.05, 101602.7, 102178.6, 102169.9, 102215.1, 102120.6, 93857.21, 
    96724.52,
  97327.76, 92635.7, 91131.68, 93668.84, 93942.16, 94081.86, 95154.95, 
    101427.7, 102136, 102197.6, 102226.7, 102263.2, 102226.2, 99841.64, 
    101149.2,
  101413.2, 101079.9, 97136.79, 94602.91, 94593.26, 93580.86, 91207.99, 
    91741.71, 85834.72, 81088.84, 78763.19, 79085.92, 82044.02, 80667.24, 
    91208.35,
  101350.7, 101313.3, 99017.92, 93795.82, 91013.23, 89126.32, 87855.55, 
    88214.71, 83207.94, 80428.55, 79655.38, 80344.88, 82587.34, 81479.97, 
    92627.86,
  92192.45, 88614.65, 93645.34, 92310.78, 85712.83, 84624.71, 86956.53, 
    86242.28, 81269.72, 79022.14, 78098.7, 78809.28, 80236.66, 81830.35, 
    94785.6,
  86013.95, 86205.21, 85243.06, 83561.84, 83296.91, 81808.83, 82697.96, 
    83046.78, 80725.73, 79449.55, 79114.27, 80682.26, 80287.61, 82319.7, 
    88561.26,
  87646.21, 86740.53, 87771.95, 86928.89, 86791.41, 85149.15, 84094.4, 
    83613.24, 82667.34, 84740.11, 100261.9, 100859.5, 90771.95, 91059.99, 
    83516.63,
  88053.06, 86227.23, 88719.88, 89559.84, 88657.32, 88233.62, 87495.09, 
    87910.48, 89579.97, 101030.9, 102022, 101988.3, 101649.2, 93304.52, 
    77847.15,
  87277.48, 86490.04, 88692.2, 89975.71, 89770.83, 89819.58, 89755.05, 
    91878.19, 95956.7, 101960.3, 101832.4, 101895.2, 101719.6, 87048.19, 
    77594.29,
  91055.19, 87764.39, 88277.18, 90108.41, 89803.98, 88792.34, 89426.25, 
    91320.08, 95771.54, 101912.8, 101888.1, 102024.3, 101767.8, 85793.4, 
    87760.14,
  94171.09, 89801.48, 88931.64, 90078.34, 89228.41, 86824.73, 88163.93, 
    90908.68, 101428.5, 101957.5, 101938.8, 101985.6, 101858.6, 93649.57, 
    96336.71,
  97472.95, 92720.14, 91199.99, 93702.8, 93970.88, 94137.12, 95143.96, 
    101351.1, 101949.5, 101982.4, 101978.5, 101982.6, 101918, 99502.64, 
    100703.5,
  101498, 101137.7, 97158.32, 94568.36, 94494.1, 93411.88, 91012.88, 
    91525.03, 85629.39, 80916.71, 78590.88, 78857.8, 81819.56, 80440.77, 
    90890.6,
  101450.1, 101399.6, 99084.2, 93833.78, 90965.77, 89002.22, 87741.23, 
    88030.81, 83045, 80261.85, 79414.75, 80122.2, 82384.08, 81259.28, 92407.69,
  92256.71, 88738.16, 93688.89, 92290.62, 85707.74, 84569.98, 86872.23, 
    86089.97, 81132.25, 78859.39, 77929.55, 78677.74, 80074.04, 81658.09, 
    94520.49,
  86110.09, 86309.56, 85364.41, 83685.41, 83402.87, 81841.23, 82712.91, 
    82974.72, 80617.72, 79307.52, 79007.77, 80561.8, 80130.47, 82225.04, 
    88277.42,
  87748.81, 86823.6, 87867.5, 87044.69, 86912.05, 85229.38, 84149.12, 
    83600.6, 82600.55, 84745.28, 100453.8, 101011.5, 90782.81, 91091.86, 
    83353.45,
  88116.44, 86301.49, 88812.33, 89684.37, 88799.02, 88360.52, 87585.31, 
    87989.74, 89688.02, 101181.8, 102044.8, 102093.9, 101783.2, 93325.81, 
    77673.75,
  87340.84, 86542.62, 88696.51, 89974.58, 89747.41, 89797.97, 89741.62, 
    91850.59, 95951.7, 101989.1, 101928.3, 102016.8, 101827.6, 87002.34, 
    77432.45,
  91125.02, 87809.95, 88316.55, 90187.25, 89867.59, 88816.12, 89438.84, 
    91396.01, 95823.66, 102014.8, 101973.2, 102066.4, 101864.5, 85723.58, 
    87665.94,
  94234.7, 89818.23, 88918.45, 90081.88, 89248.05, 86805.91, 88118.81, 
    90875.42, 101469.8, 102017.5, 101967, 102014.1, 101887.2, 93636.68, 
    96347.7,
  97489.25, 92723.55, 91189.05, 93660.66, 93934.09, 94130.02, 95136.77, 
    101398.1, 102005.2, 102009.8, 101980.3, 101995.7, 101947, 99584.77, 
    100802.8,
  101509.5, 101167.3, 97196.88, 94623.39, 94575.83, 93478.99, 91062.84, 
    91569.95, 85660.6, 80950.2, 78606.62, 78900.52, 81831.54, 80436.93, 
    90857.11,
  101350.2, 101333.9, 99055.2, 93834.45, 91005.82, 89047.35, 87784.43, 
    88052.66, 83064.96, 80279.72, 79472.27, 80150.46, 82370.66, 81252.34, 
    92314.48,
  92238.92, 88570.05, 93615.64, 92280.62, 85669.75, 84527.89, 86849.32, 
    86085.27, 81125.17, 78859, 77895.42, 78581.75, 80002.8, 81592.13, 94427.54,
  86008.91, 86064.95, 85221.24, 83495.75, 83238.83, 81725.73, 82601.88, 
    82919.02, 80572.76, 79261.93, 78941.53, 80514.41, 80044.39, 82097.52, 
    88223.71,
  87570.34, 86523.01, 87615.7, 86784.34, 86676.84, 85060.34, 83992.99, 
    83485.74, 82509.16, 84584.99, 100081.7, 100721, 90615.42, 90932.9, 
    83269.55,
  87859.3, 86043.71, 88534.31, 89424.36, 88532.38, 88108.16, 87361.99, 
    87765.56, 89389.56, 100858.3, 101857, 101837.5, 101515, 93163.05, 77538.73,
  87012.62, 86254.9, 88394.07, 89697.66, 89488.04, 89549.07, 89464.77, 
    91587.05, 95745.93, 101765.2, 101680, 101773.9, 101652.1, 86850.73, 
    77268.59,
  90849.09, 87523.13, 87997.66, 89861.21, 89579.28, 88579.74, 89205.98, 
    91177.55, 95573.62, 101754.1, 101725.2, 101846.2, 101675.6, 85557.75, 
    87558.97,
  93924.23, 89526.44, 88639.24, 89789.13, 88961.84, 86566.18, 87884.78, 
    90610.41, 101224.7, 101791.8, 101754.9, 101816.8, 101721.9, 93542.04, 
    96267.52,
  97205.8, 92476.05, 90886.91, 93397.49, 93693.26, 93884.09, 94913.95, 
    101204.7, 101805.7, 101805.5, 101790.4, 101804.3, 101759.3, 99393.79, 
    100638.8,
  101105.6, 100719.2, 96777.41, 94194.69, 94146.55, 93137.94, 90781.53, 
    91299.01, 85442.11, 80678.31, 78355.94, 78640.61, 81570.39, 80244.8, 
    90475.75,
  101051.6, 100928.6, 98641.17, 93375.84, 90577.41, 88663.3, 87370.18, 
    87711.28, 82746.19, 79957.42, 79157.61, 79848.32, 82081.69, 81025.67, 
    91905.62,
  91851.41, 88286.48, 93247.6, 91836.02, 85239.73, 84128.21, 86437.56, 
    85715.51, 80731.75, 78510.14, 77610.92, 78324.63, 79713.53, 81314.16, 
    94113.74,
  85753.28, 85932.06, 84943.7, 83194.69, 82902.33, 81373.75, 82223.41, 
    82530.98, 80209.05, 78961.4, 78633.02, 80200.39, 79786.06, 81828.29, 
    87941.25,
  87416.49, 86480.46, 87516.82, 86641.83, 86449.66, 84789.59, 83720.85, 
    83225.28, 82246.78, 84428.45, 100107.2, 100671.1, 90424.3, 90685.14, 
    83003.56,
  87859.91, 86023.41, 88561.52, 89355.8, 88405.51, 87944.94, 87195.55, 
    87661.12, 89423.68, 100988.6, 101777, 101676.6, 101307.3, 92882.55, 
    77325.76,
  87129.18, 86332.2, 88551.18, 89756.98, 89477.29, 89524.16, 89532.45, 
    91679.36, 95857.4, 101801.1, 101631.5, 101621.5, 101363.8, 86654.73, 
    77086.56,
  91072.62, 87695.82, 88238.88, 90083.98, 89683.07, 88627.3, 89282.7, 
    91176.87, 95730.17, 101867.7, 101760.1, 101775.7, 101410.5, 85301.95, 
    87350.28,
  94259.92, 89784.16, 88903.38, 90037.27, 89142.88, 86688.47, 88012.37, 
    90863.59, 101467.5, 101939.5, 101833.2, 101845.6, 101617.4, 93477.83, 
    96307.6,
  97627.14, 92814.21, 91280.05, 93788.67, 94060.02, 94230.84, 95217.7, 
    101442.5, 101976.9, 102006.6, 101945.5, 101940.7, 101845.3, 99477.59, 
    100656.2,
  101505.9, 101219.2, 97200.76, 94563.69, 94512.05, 93422.55, 91031.97, 
    91511.07, 85576.55, 80823.41, 78492.52, 78829.22, 81851.6, 80459.27, 
    91103.01,
  101646.6, 101506.3, 99152.73, 93830.54, 90979.2, 89033.25, 87756.31, 
    87996.72, 82944.48, 80149.2, 79392.15, 80149.22, 82428.36, 81335.93, 
    92576.97,
  92262.18, 88682.12, 93760.51, 92296.15, 85645.62, 84573.63, 86920.09, 
    86099.9, 81062.53, 78844.74, 77943.93, 78713.05, 80082.7, 81758.86, 
    94689.7,
  86115.08, 86324.34, 85335.5, 83609.23, 83330.16, 81822.31, 82718.55, 
    83009.38, 80617.78, 79335.23, 79020.05, 80682.98, 80200.08, 82409.33, 
    88458.67,
  87767.12, 86869.97, 87951.36, 87112.71, 86968.76, 85268.11, 84220.45, 
    83691.8, 82675.41, 84936, 100927.8, 101456.2, 91035.11, 91409.74, 83438.26,
  88227.06, 86387.67, 89034.13, 89880.71, 88984.12, 88538.66, 87815.2, 
    88236.59, 90014.63, 101683, 102494.7, 102444.3, 102239.4, 93667.89, 
    77727.16,
  87405.94, 86636.12, 88923.65, 90234.05, 90050.72, 90109.87, 90072.02, 
    92183.62, 96443.35, 102433, 102371.8, 102310.8, 102307.5, 87195.1, 
    77562.59,
  91309.49, 87985.78, 88559.05, 90464.75, 90148.8, 89079.23, 89778.96, 
    91690.85, 96324.16, 102493.1, 102430.9, 102403.1, 102236.5, 85900.64, 
    88104.59,
  94474.1, 90021.28, 89151.97, 90331.07, 89468.95, 87039.73, 88395.02, 
    91212.77, 101966.3, 102510.5, 102449.4, 102451.4, 102265.7, 94048.08, 
    96970.14,
  97845.88, 93025.38, 91482.62, 94023.12, 94321.6, 94481.27, 95522.98, 
    101812.6, 102463.9, 102532.8, 102500.9, 102527.9, 102468.9, 100070, 
    101272.5,
  101773.6, 101497.4, 97465.38, 94883.16, 94858.45, 93788.75, 91394.68, 
    91905.12, 85944.07, 81193.35, 78829.71, 79162.46, 82308.25, 80912.95, 
    91747.9,
  101885.3, 101769.3, 99439.16, 94137.57, 91264.29, 89326.52, 88058.52, 
    88392.68, 83320.69, 80518.58, 79726.24, 80438.52, 82812.51, 81732.87, 
    93161.58,
  92502.57, 88931.27, 94007.73, 92583.95, 85926.48, 84825.67, 87169.05, 
    86397.55, 81365.24, 79092.77, 78190.88, 78927.21, 80400.7, 82084.63, 
    95296.17,
  86359.11, 86513.31, 85498.83, 83771.91, 83501.51, 81973.28, 82860.59, 
    83187.84, 80839.52, 79530.27, 79199.88, 80800.95, 80493.13, 82621.06, 
    88995.59,
  87958.84, 86992.06, 88084.37, 87254.31, 87109.2, 85417.75, 84318.87, 
    83793.67, 82794.12, 84956.95, 100748.9, 101274.1, 90980.88, 91412.27, 
    83840.1,
  88400.25, 86509.34, 89119.91, 89974.37, 89057.3, 88584.89, 87837.91, 
    88251.02, 89924.41, 101457.1, 102444.2, 102440.1, 102191.8, 93710.74, 
    78074.2,
  87560, 86761.19, 88963.49, 90293.53, 90078.02, 90118.95, 90029.05, 
    92085.72, 96295.03, 102330.2, 102290.2, 102299.2, 102208.4, 87337.06, 
    77830.48,
  91459.7, 88085.3, 88592.12, 90461.32, 90151.62, 89100.8, 89727.37, 
    91580.62, 96084.96, 102295.5, 102318.9, 102407.4, 102286.6, 86123.43, 
    88213.45,
  94561.76, 90098.72, 89180.49, 90318.09, 89475.31, 87029.08, 88346.74, 
    91046.29, 101653.8, 102289.6, 102290.6, 102330.5, 102312.2, 94018.26, 
    96931.85,
  97859.7, 93091.13, 91467.8, 93924.88, 94187.14, 94347.88, 95334.25, 
    101562.4, 102181, 102272.9, 102320.6, 102355.9, 102375.9, 99955.42, 
    101227.5,
  101899.5, 101574, 97490.49, 94885.5, 94837.34, 93736.29, 91289.7, 91817.23, 
    85753.53, 81039.12, 78661.34, 79025.46, 82148.77, 80668.89, 91493.81,
  101954.2, 101757, 99509.68, 94188.11, 91291.41, 89318.46, 88056.84, 
    88356.3, 83235.14, 80463.34, 79640.75, 80358.53, 82668.84, 81581.31, 
    93003.38,
  92532.91, 89088.23, 94035.3, 92591.77, 85953.98, 84867.25, 87171.98, 
    86387.52, 81377.3, 79095.17, 78156.38, 78896.04, 80323.41, 82010.53, 
    95095.89,
  86524.93, 86699.05, 85674.8, 83978.27, 83675.84, 82098.77, 82957.59, 
    83266.27, 80869.8, 79523.91, 79252.95, 80801.54, 80435.72, 82562.98, 
    88793.01,
  88137.7, 87131.65, 88201.88, 87355.97, 87183.09, 85514.95, 84402.91, 
    83870.23, 82852.37, 85057.88, 100667.1, 101225.7, 90993.84, 91340.9, 
    83732.99,
  88513.3, 86645.8, 89200.19, 90038.43, 89113.91, 88646.02, 87859.87, 
    88253.86, 89905.06, 101290.8, 102193.6, 102241.2, 102022.3, 93591.2, 
    78026.26,
  87649.42, 86859.61, 89028.28, 90331.81, 90106.12, 90106.9, 90043.66, 
    92034.8, 96122.88, 102109, 102120.1, 102157.3, 102036, 87288.5, 77797.55,
  91406.57, 88131.73, 88613.09, 90488.45, 90163.1, 89098.06, 89701.88, 
    91506.14, 95985.8, 102075.8, 102098.2, 102213.2, 102068.3, 86095.42, 
    88085.88,
  94393.59, 90064.48, 89149.94, 90301.8, 89479.27, 87079.82, 88350.19, 
    91073.88, 101457.7, 102059.4, 102082.3, 102158.7, 102109.7, 93908.2, 
    96691.81,
  97589.93, 92922.68, 91316.68, 93765.38, 94034.79, 94220.12, 95149.05, 
    101267.8, 101917.1, 102023.1, 102054, 102122, 102136.1, 99738.87, 100947.2,
  101520.3, 101244.9, 97255.36, 94675.1, 94636.73, 93525.38, 91060.16, 
    91591.18, 85596.83, 80913.44, 78576.9, 78849.29, 81904.54, 80359.33, 
    91012.34,
  101433.8, 101418.6, 99219.7, 93952.96, 91063.87, 89111.91, 87842.62, 
    88115.91, 83064.66, 80320.73, 79495.13, 80175.48, 82411.95, 81231.77, 
    92476.02,
  92252.25, 88718.09, 93709.45, 92346.19, 85700.45, 84582.07, 86891.3, 
    86127.08, 81157.61, 78876.1, 77891.91, 78644.97, 80047.54, 81669.82, 
    94484.59,
  86100.19, 86140.98, 85241.12, 83578.92, 83300.16, 81786.02, 82628.92, 
    82969.02, 80620.31, 79283.95, 79023.67, 80546.78, 80133.38, 82254.66, 
    88278.52,
  87725.11, 86603.32, 87662.48, 86844.3, 86696.77, 85077.73, 84008.83, 
    83491.09, 82488.01, 84631.09, 99816.03, 100479.7, 90476.5, 90939.59, 
    83338.95,
  87965.05, 86096.82, 88569.54, 89452.55, 88573.21, 88130.16, 87393.84, 
    87760.57, 89363.39, 100437.4, 101427, 101474.2, 101313.9, 93061.97, 
    77756.18,
  87085.02, 86289.58, 88414.68, 89716.59, 89517.85, 89547.04, 89474.62, 
    91450.49, 95423.77, 101253.9, 101326.2, 101347.3, 101396.3, 86825.53, 
    77522.41,
  90819.78, 87536.57, 87992.73, 89834.03, 89532.91, 88506.17, 89122.61, 
    90952.39, 95230.94, 101181.1, 101272, 101387.3, 101371.9, 85676.1, 
    87687.48,
  93803.38, 89473.13, 88545.29, 89650.41, 88849.92, 86463.5, 87719.16, 
    90332.1, 100521.5, 101119.7, 101194.5, 101312.3, 101364.1, 93376.93, 
    96122.82,
  96984.1, 92341, 90719.77, 93104.71, 93383.48, 93567.85, 94467.01, 100440.7, 
    101047.9, 101058.2, 101126.5, 101228.4, 101352.5, 99072.78, 100324.8,
  101677, 101369.8, 97360.32, 94785.5, 94762.45, 93709.51, 91271.94, 
    91821.03, 85778.48, 81053.84, 78651.23, 78911.38, 81817.7, 80314.77, 
    90614.19,
  101735.3, 101568.6, 99300.84, 94039.66, 91178.27, 89230.09, 87994.62, 
    88280.36, 83201.45, 80431.62, 79555.02, 80223.65, 82376.33, 81183.73, 
    92135.75,
  92402.7, 88997.66, 93874.33, 92443.61, 85881.56, 84786.15, 87058.79, 
    86288.22, 81298.02, 78994.71, 77930.55, 78631.04, 79945.3, 81557.27, 
    94230.97,
  86447.61, 86644.02, 85625.85, 83935.21, 83616.98, 82051.13, 82874.1, 
    83160.42, 80751.84, 79385.06, 79163.27, 80720.7, 80074.5, 82185.47, 
    88078.01,
  88044.92, 87076.3, 88101.66, 87275.25, 87076.59, 85427.73, 84309.39, 
    83759.98, 82697.34, 84926.98, 100127, 100649.2, 90630.88, 90918.44, 
    83131.06,
  88450.31, 86608, 89100.43, 89904.38, 88982.05, 88513.99, 87734.55, 
    88106.98, 89720.99, 100845.5, 101647.9, 101611.4, 101371.3, 93054.33, 
    77586.52,
  87634.03, 86847.58, 88975.7, 90202.38, 89966.27, 89960.3, 89889.53, 
    91832.23, 95848.59, 101638.3, 101554.8, 101506.3, 101426.1, 86823.28, 
    77389.78,
  91397.5, 88118.27, 88579.84, 90384.83, 90029.48, 88991.64, 89575.62, 
    91318.41, 95742.91, 101611.4, 101521.8, 101520.7, 101378.3, 85583.48, 
    87556.32,
  94367.38, 90054.34, 89136, 90236.21, 89370.23, 87000.26, 88242.07, 
    90963.95, 101167.1, 101619.7, 101494.6, 101467.6, 101351.9, 93348.42, 
    95970.15,
  97539.25, 92908.79, 91312.61, 93691.04, 93946.22, 94139.95, 95093.53, 
    101104.8, 101652.6, 101607.4, 101491.3, 101432.2, 101364, 99020.45, 
    100138.9,
  102017.8, 101689, 97670.81, 95154.34, 95162.98, 94122.42, 91698.34, 
    92273.5, 86209.83, 81479.3, 79080.3, 79356.51, 82315.19, 80829.18, 
    91255.01,
  101846.7, 101849.9, 99642.97, 94414, 91570.93, 89661.16, 88432.55, 
    88734.33, 83662.13, 80888.65, 80012.16, 80688.3, 82858.09, 81689.45, 
    92732.52,
  92782.55, 89301.05, 94188.09, 92826.61, 86271.14, 85157.17, 87429.82, 
    86690.09, 81735.4, 79410.56, 78325.74, 79054.84, 80420.52, 82048.23, 
    94807.04,
  86631.82, 86590.78, 85752.31, 84136.05, 83847.7, 82341.49, 83175.66, 
    83508.41, 81156.1, 79809.54, 79581.73, 81141.42, 80518.86, 82653.2, 
    88599.65,
  88199.27, 86960.77, 88040.68, 87225.8, 87098.78, 85523.91, 84475.84, 
    83994.77, 82981.73, 85160.79, 100158.3, 100882.6, 90986.73, 91374.02, 
    83580.53,
  88292.62, 86431.97, 88846.15, 89755.69, 88902.05, 88483.34, 87749.29, 
    88155.77, 89746.63, 100766.7, 101861.4, 101942.3, 101769.2, 93489.33, 
    78013.98,
  87224.42, 86497.07, 88604.61, 89946.12, 89770.29, 89831.34, 89776.25, 
    91739.41, 95719.6, 101602.3, 101710.3, 101769.5, 101846.8, 87202.11, 
    77823.42,
  90710.16, 87599.71, 88096.2, 89974, 89718.86, 88757.92, 89388.02, 91206.38, 
    95491.21, 101506.6, 101616.7, 101790.9, 101764.5, 85972.7, 87942.32,
  93545.48, 89384.81, 88541.15, 89687.63, 88993.66, 86701.66, 87985.08, 
    90565.77, 100683.5, 101453.1, 101531.9, 101706.9, 101703, 93739.22, 
    96345.12,
  96572.11, 92072.66, 90526.24, 92927.21, 93267.62, 93443.38, 94423.42, 
    100396.3, 101180.6, 101355.3, 101464.6, 101635.9, 101722.9, 99417.95, 
    100658.2,
  101314, 100954.4, 97126.62, 94683.25, 94693.65, 93792.85, 91577.25, 
    92109.66, 86322.68, 81543.71, 79166.78, 79409.97, 82268.18, 80876.49, 
    90930.16,
  101050.8, 101166, 98952.83, 93819.3, 91126.75, 89322.63, 88139.59, 
    88526.84, 83665.99, 80826.89, 79983.46, 80589.68, 82743.83, 81644.95, 
    92327.95,
  92289.7, 88604.01, 93532.76, 92246.74, 85828.19, 84717, 87045.98, 86477.78, 
    81571.77, 79300.59, 78303.91, 78934.25, 80292.52, 81807.34, 94305.8,
  86167.63, 85944.62, 85272.83, 83537.83, 83267.95, 81834.33, 82705.54, 
    83099.76, 80819.85, 79602.75, 79247.27, 80721.1, 80236.95, 82225.14, 
    88214.8,
  87677.78, 86307.98, 87496.27, 86576, 86480.27, 84884.86, 83857.21, 
    83455.98, 82529.29, 84467.14, 99059.8, 99925.91, 90336.79, 90660.56, 
    83300.41,
  87726.75, 85902.98, 88283.66, 89117.55, 88228.6, 87767.01, 87040.24, 
    87427.24, 88949.21, 99792.51, 100769.8, 100752.3, 100658, 92694.01, 
    77725.6,
  86813.91, 86016.9, 88088.99, 89375.13, 89116.06, 89135.33, 89046.56, 
    90951.66, 94903.77, 100445.3, 100459.6, 100606.7, 100647.3, 86673.68, 
    77327.73,
  90520.24, 87235.45, 87669.65, 89455.88, 89108.8, 88094.27, 88663.15, 
    90455.24, 94633.85, 100343.6, 100411.4, 100552.1, 100463.3, 85367.88, 
    86971.27,
  93405.33, 89079.76, 88121.66, 89191.62, 88389.37, 86039.18, 87248.3, 
    89771.53, 99700.62, 100317.1, 100262.1, 100377.6, 100387.7, 92738.7, 
    95221.2,
  96507.62, 91850.27, 90159.52, 92493.74, 92726.7, 92839.53, 93702.99, 
    99593.88, 100185.3, 100155.9, 100151.5, 100210.3, 100267.1, 98082.02, 
    99226.8,
  101034.1, 100618.1, 96719.62, 94193.87, 94124.73, 93124.52, 90872.22, 
    91350.45, 85673.02, 80948.09, 78675.34, 79005.2, 81882.09, 80573.87, 
    90495.85,
  100773.1, 100807.5, 98558.39, 93353.55, 90593.2, 88761.38, 87525.24, 
    87884.61, 83057.97, 80263.04, 79509.93, 80180.83, 82361.88, 81353.12, 
    91897.75,
  91872.13, 88115.62, 93122.52, 91816.19, 85341.96, 84220.7, 86536.69, 
    85902.88, 80996.39, 78785.91, 77920.84, 78629.26, 79985.09, 81530.84, 
    93931.2,
  85676.8, 85542.26, 84799.63, 83067.15, 82829.91, 81401.82, 82283.33, 
    82625.87, 80366.58, 79181.52, 78829.86, 80339.12, 80015.37, 81991.77, 
    87982.26,
  87189.92, 86018.32, 87160.37, 86284.2, 86199.62, 84590.17, 83571.83, 
    83120.23, 82205.23, 84174.55, 99051.37, 99876.35, 90113.66, 90459.86, 
    83135.77,
  87368.59, 85548.97, 88015.85, 88874.27, 87998.62, 87571.81, 86851.63, 
    87234.15, 88798.8, 99718.24, 100643.8, 100623.6, 100512.4, 92603.17, 
    77519.01,
  86504.84, 85717.84, 87845.78, 89139.74, 88914.59, 88977.8, 88904.05, 
    90883.38, 94833.14, 100492.4, 100422.2, 100566.9, 100546, 86539.78, 
    77214.67,
  90265.07, 86966.53, 87401.86, 89240.65, 88925.02, 87944.48, 88556.31, 
    90402.67, 94618.16, 100480.2, 100453.5, 100579.5, 100467.2, 85275.46, 
    87083.91,
  93238.49, 88862.5, 87932.72, 89035.55, 88254.84, 85928.18, 87220.79, 
    89805.77, 99935.98, 100468.8, 100423.4, 100510.7, 100477.4, 92764.18, 
    95361.75,
  96384.82, 91696.11, 90071.21, 92470.69, 92729.74, 92852.58, 93811.98, 
    99818.68, 100421.3, 100415.5, 100430.1, 100474.1, 100492.1, 98251.46, 
    99369.61,
  101128.7, 100706.3, 96719.21, 94052.48, 93955.76, 92862.02, 90464.2, 
    90928.71, 85006.24, 80309.21, 77971.54, 78227.62, 81146.73, 79759.86, 
    89937.86,
  101139.1, 100868.3, 98567.74, 93304.14, 90446.43, 88485.3, 87200.83, 
    87448.48, 82416.19, 79660.7, 78818.04, 79494.21, 81646.71, 80583.8, 
    91357.23,
  91867.69, 88379.43, 93250.88, 91754.09, 85183.12, 84113.34, 86365.08, 
    85549.88, 80527.88, 78217.07, 77236.69, 77905.22, 79260.57, 80874.7, 
    93366.85,
  85908.18, 86063.51, 85006.1, 83278.77, 82944.38, 81415.44, 82246.23, 
    82506.15, 80080.44, 78748.37, 78521.91, 79973.77, 79454.09, 81432.6, 
    87451.28,
  87551.73, 86580.04, 87564.41, 86681.23, 86451.82, 84810.9, 83735.72, 
    83170.41, 82131.4, 84333.19, 99326.84, 99708.2, 89770.03, 90005.37, 
    82565.55,
  88012.4, 86132.04, 88600.07, 89361.6, 88382.8, 87938.09, 87192.09, 
    87562.59, 89222.28, 100169.4, 100779.7, 100614, 100373.5, 92111.32, 
    77073.7,
  87266.33, 86432.07, 88544.18, 89739.02, 89444.95, 89450.04, 89397.3, 
    91375.02, 95390.16, 100995.6, 100765.2, 100588.4, 100359.5, 85963.54, 
    76879.91,
  91134.67, 87755.83, 88210.54, 90000.22, 89614.7, 88561.52, 89175.65, 
    90967.47, 95378.06, 101118, 100899.9, 100788, 100391.7, 85025.19, 87065.77,
  94200.05, 89762.37, 88829.98, 89909.74, 89017.92, 86603.88, 87906.96, 
    90639.4, 100892.6, 101231.2, 101037.2, 100932.8, 100631.4, 92790.63, 
    95549.65,
  97433.79, 92714.1, 91114.66, 93561.51, 93784.85, 93935.14, 94913.6, 
    100981.2, 101430.6, 101335.5, 101181.5, 101097.3, 100945.5, 98587.82, 
    99771.45,
  101727.5, 101437.9, 97428.17, 94867.15, 94795.31, 93672.52, 91207.16, 
    91703.72, 85621.37, 80931.4, 78557.97, 78832.14, 81720.2, 80235.12, 
    90602.57,
  101889.6, 101711.1, 99414.12, 94162.69, 91298.88, 89341.94, 88077.07, 
    88298.35, 83146.82, 80392.53, 79504.2, 80198.59, 82293.72, 81083.03, 
    92195.55,
  92532.71, 89146.98, 94096.81, 92628.5, 86006, 84943.22, 87220.84, 86360.09, 
    81277.51, 78973.67, 77922.9, 78634.59, 79880.39, 81555.98, 94293.32,
  86614.32, 86793.47, 85739.12, 84078.64, 83794.42, 82241.82, 83094.16, 
    83384.06, 80938.04, 79639.62, 79420.7, 80973.02, 80221.19, 82260.26, 
    88087.77,
  88232.69, 87295.95, 88336.09, 87487.67, 87315.32, 85677.61, 84609.66, 
    84063.75, 82964.72, 85363.86, 100843.6, 101272.5, 91054.6, 91239.16, 
    83112.95,
  88667.02, 86850.45, 89401.48, 90202.37, 89288.3, 88867.08, 88134.86, 
    88584.8, 90341.09, 101671.1, 102461.9, 102299.8, 102004.2, 93322.51, 
    77651.59,
  87919.06, 87132.5, 89325.05, 90573.14, 90371.91, 90401.73, 90409.27, 
    92465.92, 96633.83, 102512.9, 102358.4, 102171.3, 101911.7, 86889.57, 
    77604.48,
  91741.7, 88456.06, 88982.72, 90822.52, 90485.15, 89452.39, 90136.79, 
    91967.75, 96583.93, 102566.4, 102407.9, 102352, 101829.1, 85926.3, 
    88143.98,
  94828.98, 90452.03, 89582.31, 90739.15, 89843.27, 87466.6, 88770.12, 
    91661.92, 102157.7, 102627.6, 102468.8, 102441.2, 102104.9, 94001.29, 
    96830.98,
  98112.16, 93390.95, 91847.26, 94335.59, 94609.85, 94830.6, 95836.65, 
    102086.1, 102650.6, 102690.8, 102564.6, 102534.5, 102372.3, 100001.3, 
    101219.6,
  101902.2, 101672.1, 97582.34, 94971.69, 94888.34, 93784.02, 91328.89, 
    91837.45, 85790.49, 81146.23, 78824.5, 79138.23, 82221.95, 80759.21, 
    91424.09,
  102041.7, 101863, 99565.42, 94253.16, 91377.16, 89424.06, 88183.02, 
    88441.24, 83317.12, 80601.2, 79771.72, 80528.93, 82778.34, 81582.33, 
    92907.37,
  92586.4, 89200.15, 94141.14, 92677.07, 86031.98, 84992.86, 87296.27, 
    86482.21, 81468.89, 79188.12, 78175.43, 78978.4, 80353.27, 82049.48, 
    95068.34,
  86697.62, 86861.36, 85828.07, 84147.59, 83839.9, 82282.87, 83148.95, 
    83452.94, 81006.23, 79641.64, 79459.91, 81036.48, 80452.36, 82697.68, 
    88703.64,
  88267.96, 87330.43, 88389.94, 87550.95, 87394.56, 85712.3, 84631.12, 
    84084.34, 83013.69, 85439.03, 100946.1, 101535.2, 91233.2, 91697.05, 
    83535.26,
  88682.44, 86869.53, 89465.44, 90256.04, 89376.02, 88905.8, 88176.75, 
    88544.1, 90339.64, 101636, 102611.3, 102543.1, 102484.5, 93707.16, 
    78056.11,
  87887.05, 87104.36, 89313.46, 90596.61, 90422.21, 90445.35, 90414.68, 
    92410.54, 96587.97, 102524.3, 102478.4, 102289, 102405.6, 87299.73, 
    77936.08,
  91637.48, 88401.34, 88942.96, 90779.27, 90481.96, 89449.13, 90096.68, 
    91904.09, 96533.93, 102550.4, 102418.9, 102413.3, 102169.8, 86289.59, 
    88457.95,
  94646.27, 90364.26, 89485.01, 90641.93, 89820.45, 87448.15, 88742.09, 
    91531.48, 102077.2, 102608, 102450.8, 102453.2, 102185.5, 94223.76, 
    97167.52,
  97863.54, 93205.55, 91689.48, 94147.67, 94401.7, 94580.01, 95570.6, 
    101802.3, 102565.3, 102669.5, 102589.1, 102594.4, 102493.9, 100211, 
    101571.8,
  101792.6, 101454.5, 97436.94, 94906.7, 94881.91, 93770.88, 91370.95, 
    91912.23, 85969.89, 81294.31, 78953.06, 79231.95, 82369.48, 80940.24, 
    91617.84,
  101814.9, 101737.9, 99451.91, 94197.18, 91313.88, 89388.95, 88156.9, 
    88435.52, 83404.27, 80668.77, 79855.44, 80558.91, 82824.46, 81715.6, 
    93065.41,
  92545.38, 89057.68, 94040.96, 92537.46, 85994.27, 84925.89, 87224.27, 
    86459.52, 81520.39, 79261.85, 78288.85, 79044.27, 80471.41, 82103.62, 
    95178.95,
  86514.73, 86662.39, 85692.98, 84046.05, 83760.7, 82218, 83049.52, 83379.3, 
    81008.51, 79637.05, 79359.5, 80920.06, 80514.81, 82648.23, 88875.38,
  88098.8, 87174.9, 88226.68, 87394.46, 87240.61, 85562.3, 84484.75, 
    83950.43, 82898.48, 85164.88, 100573.1, 101203.6, 90983.56, 91482.91, 
    83718.16,
  88479.46, 86652.99, 89238.89, 90048.98, 89159.51, 88678.09, 87920.28, 
    88322.66, 90012.7, 101256.1, 102283.1, 102272.6, 102117.2, 93639.41, 
    78093.32,
  87670.25, 86884.91, 89087.95, 90368.18, 90159.07, 90147.65, 90080.02, 
    92095.97, 96188.38, 102141.1, 102199.1, 102134.5, 102204.4, 87214.42, 
    77909.76,
  91362.45, 88147.29, 88676.01, 90530, 90236.28, 89176.46, 89788.73, 
    91589.13, 96115.43, 102109.2, 102143.3, 102230.2, 102142.1, 86144.92, 
    88281.52,
  94361.86, 90112.84, 89232.02, 90377.84, 89583.76, 87235.09, 88499.01, 
    91214.45, 101580.2, 102133, 102100.7, 102203.2, 102167.9, 94017.89, 
    96871.05,
  97583.39, 92935.73, 91413.45, 93849.45, 94104.29, 94282.6, 95266.66, 
    101395.8, 102082.7, 102183.1, 102143.2, 102199.2, 102213.4, 99907.25, 
    101253.4,
  101515.7, 101237.8, 97349.59, 94896.84, 94916.15, 93873.09, 91503.62, 
    92064.54, 86123.53, 81427.55, 79081.82, 79373.18, 82411.02, 80976.51, 
    91539.8,
  101470.2, 101497, 99190.27, 94064.97, 91330.5, 89434.59, 88220.99, 
    88539.88, 83554.62, 80815.27, 79990.53, 80668.93, 82902.55, 81771.96, 
    92963.09,
  92482.85, 88986.47, 94034.43, 92580.85, 86043.68, 84969.96, 87259.89, 
    86510.91, 81626.47, 79354.79, 78350.38, 79084.67, 80535.56, 82145.11, 
    95104.39,
  86268.58, 86423.72, 85539.61, 83938.03, 83682.06, 82185.14, 83036.38, 
    83359.52, 81052.69, 79720.74, 79464.55, 81000.29, 80539.12, 82678.96, 
    88885.62,
  87889.38, 87028.77, 88057.4, 87232.11, 87122.35, 85488.21, 84427.15, 
    83909.53, 82903.38, 85080.16, 100385.3, 101006.5, 91001.86, 91362.53, 
    83796.34,
  88239.64, 86440.95, 88999.52, 89866.24, 89009.49, 88548.75, 87804.45, 
    88232.33, 89904.53, 101145, 102155.6, 102062.7, 101876.2, 93508.73, 
    78177.84,
  87467.83, 86695.91, 88903.8, 90184.34, 89981.16, 89992.41, 89951.89, 
    92009.27, 96108.31, 102030.5, 102005.2, 101950.8, 101966.8, 87228.09, 
    77985.49,
  91161.43, 87921.84, 88489.92, 90333.24, 90051.2, 89026.47, 89676.96, 
    91514.6, 95991.48, 102007.2, 102047.6, 102046.5, 101966.6, 86085.5, 
    88250.75,
  94217.47, 89889.77, 89073.73, 90212.16, 89424.94, 87069.47, 88356.62, 
    91079.91, 101509.8, 102044.6, 102034.2, 102036.6, 102007.2, 93844.91, 
    96671.99,
  97357.86, 92722.79, 91265.5, 93719.76, 93997.71, 94154.05, 95216.05, 
    101367, 102014.1, 102077.6, 102068, 102077.8, 102050.9, 99701.09, 100994.2,
  101120, 100758, 97056.59, 94687.65, 94703.08, 93711.62, 91383.79, 91940.04, 
    86031.82, 81355.23, 79054.64, 79318.06, 82347.76, 80932, 91400.63,
  101010.7, 101029.7, 98836.05, 93793.88, 91162.73, 89322.16, 88081.41, 
    88462.25, 83494.85, 80735.46, 79940.41, 80621.05, 82859.54, 81765.77, 
    92905.99,
  92150.74, 88733.65, 93761.05, 92379.12, 85899.57, 84855.42, 87180.7, 
    86470.88, 81545.43, 79304.06, 78351.91, 79075.55, 80510.56, 82112.62, 
    95020.41,
  85977.43, 86179.73, 85299.88, 83740.84, 83501.52, 82054.41, 82959.26, 
    83285.91, 80993.98, 79708.01, 79396.65, 80972.33, 80537.67, 82624.84, 
    88800.34,
  87627.85, 86804.51, 87829.01, 87009.49, 86915.48, 85308.05, 84311.46, 
    83828.29, 82856.55, 84924.44, 100169.3, 100782.1, 90849.09, 91271.91, 
    83751.64,
  88000.9, 86226.04, 88758.7, 89635.66, 88794.06, 88350.88, 87630.23, 
    88021.7, 89658.42, 100913.9, 101887.4, 101829.7, 101593.6, 93391.81, 
    78130.48,
  87225.16, 86480.98, 88661.59, 89942.7, 89748.38, 89807.73, 89737.3, 
    91795.23, 95883.44, 101780.1, 101725.4, 101752.3, 101688.9, 87204.8, 
    77918.52,
  90936.69, 87715.62, 88243.5, 90092.68, 89802.21, 88832.8, 89433.42, 
    91306.2, 95718.33, 101759, 101758.2, 101833.1, 101685.6, 86008.43, 
    88061.43,
  93985.35, 89690.64, 88832.74, 89961.23, 89190.61, 86869.3, 88147.11, 
    90784.72, 101197.8, 101806.7, 101755, 101800.5, 101755.9, 93722.34, 
    96438.38,
  97140.1, 92477.25, 90999.13, 93437.84, 93730.84, 93856.32, 94878.23, 
    101055.7, 101765.9, 101795.9, 101798, 101808.5, 101800.8, 99413.25, 
    100680.4,
  101168.1, 100899.7, 96965.03, 94420.77, 94378.73, 93307.96, 90949.84, 
    91471.77, 85635.31, 81007.95, 78734.02, 79077.94, 82143.47, 80763.98, 
    91224.09,
  101192.8, 101143.1, 98834.91, 93621.44, 90857.93, 88960.07, 87691.68, 
    88049.49, 83101.19, 80395.27, 79635.32, 80345.97, 82600.25, 81519.95, 
    92592.93,
  92066.41, 88566.73, 93616.03, 92159.47, 85576.22, 84549.48, 86853.85, 
    86114.7, 81181.02, 78974.42, 78095.62, 78826.77, 80245, 81853.63, 94710.8,
  85951.72, 86118.21, 85134.61, 83506.73, 83253.29, 81758.53, 82659.44, 
    82980.24, 80669.43, 79415.98, 79091.96, 80660.58, 80345.28, 82387.73, 
    88600.24,
  87572.33, 86655.3, 87670.18, 86830.34, 86698.46, 85068.98, 84033.57, 
    83563.64, 82602.55, 84640.06, 99800.01, 100363, 90488.96, 90956.8, 
    83567.56,
  87926, 86087.09, 88576.69, 89413.41, 88545.97, 88120.63, 87401.11, 
    87745.96, 89375.64, 100430.9, 101358.6, 101323.4, 101130.2, 93078.51, 
    77982.41,
  87075.52, 86326.38, 88456.18, 89726.65, 89519.38, 89560.37, 89477.9, 
    91454.06, 95487.83, 101274.7, 101238.7, 101264.9, 101233.7, 86932.38, 
    77749.72,
  90784.98, 87555.18, 88032.23, 89855.54, 89546.95, 88561.42, 89157.8, 
    90957.42, 95297.62, 101267.4, 101279, 101361.9, 101254.2, 85762.21, 
    87804.91,
  93769.88, 89485.72, 88590.92, 89702.09, 88921.09, 86617.16, 87898.16, 
    90444.98, 100631.1, 101283.6, 101280, 101362.9, 101312.6, 93394.51, 
    96127.36,
  96930.2, 92279.85, 90701.25, 93105.38, 93360.07, 93490.88, 94450.41, 
    100450.7, 101175.7, 101272.4, 101305.4, 101358.4, 101359.3, 99029.82, 
    100322.8,
  101743.1, 101396.4, 97348.81, 94743.12, 94646.45, 93516.65, 91108.92, 
    91648.28, 85692.16, 81109.4, 78823.15, 79192.8, 82274.95, 80828.61, 
    91355.77,
  101643.4, 101537.2, 99301.88, 94056.12, 91171.09, 89209.9, 87941.87, 
    88233.27, 83258.66, 80580.03, 79782.05, 80493.18, 82751.55, 81635.33, 
    92798.59,
  92563.05, 88912.23, 93856.98, 92441.6, 85916.13, 84820.21, 87070.33, 
    86302.7, 81430.65, 79181.67, 78231.75, 78992.14, 80418.98, 82023.2, 
    94908.72,
  86480.2, 86462.27, 85611.43, 83927.09, 83627.93, 82109.23, 82932.7, 
    83227.73, 80935.4, 79627.24, 79325.13, 80875.98, 80489.51, 82564.71, 
    88724.51,
  88099.84, 86917.22, 88013.55, 87186.41, 87025.57, 85389.28, 84319.23, 
    83815.77, 82821.25, 84889.8, 99958.52, 100493.1, 90675.26, 91136.24, 
    83692.38,
  88221.12, 86402.84, 88877.91, 89773.48, 88881.43, 88422.09, 87661.01, 
    88023.55, 89586.61, 100543.4, 101439.8, 101455.3, 101317.5, 93201.94, 
    78159.28,
  87247.41, 86531.4, 88661, 89998.93, 89804.04, 89841.2, 89739.55, 91674.2, 
    95591.62, 101344.9, 101353.5, 101375, 101398, 87088.16, 77959.45,
  90875.16, 87685.98, 88159.17, 90050.16, 89773.95, 88783.08, 89383.16, 
    91172.18, 95363.37, 101268.9, 101321, 101416.1, 101385.6, 85929.15, 
    87977.93,
  93785.73, 89506.35, 88596.98, 89775.88, 89067.2, 86757.63, 88045.16, 
    90584.88, 100586.5, 101216.5, 101269.3, 101378.3, 101390.5, 93549.67, 
    96251.87,
  96908.13, 92266.8, 90621.15, 93056.45, 93398.8, 93566.91, 94542.8, 100482, 
    101111.2, 101161.1, 101230.7, 101331.2, 101402.1, 99138.3, 100396.8,
  101949.7, 101626.1, 97609.16, 95072.41, 94998.04, 93934.09, 91549.91, 
    92098.66, 86174.77, 81600.31, 79296.91, 79613.81, 82639.41, 81167.19, 
    91480.5,
  101791.1, 101783.3, 99497.62, 94320.27, 91465.04, 89577.34, 88350.43, 
    88676.91, 83712.25, 81026.56, 80206.37, 80867.8, 83118.93, 81962.52, 
    92956.29,
  92808.41, 89181.63, 94169.56, 92787.25, 86295.98, 85177.76, 87441.37, 
    86702.55, 81845.51, 79610.39, 78637.91, 79354.74, 80759.77, 82310.12, 
    95048.2,
  86687.3, 86608.95, 85816.73, 84165.19, 83917.29, 82429.41, 83289.92, 
    83582.92, 81299.45, 80021.65, 79746.94, 81289.05, 80805.43, 82886.16, 
    88884.7,
  88340.95, 87073.88, 88199.18, 87379.34, 87264.83, 85664.52, 84632.85, 
    84146.18, 83180.82, 85224.41, 100119.5, 100704.1, 90990.67, 91407.71, 
    83933.12,
  88409.01, 86553.49, 89044.05, 89917.71, 89052.61, 88610.68, 87884.86, 
    88278.15, 89852.41, 100719.8, 101638.7, 101669.3, 101493.4, 93460.87, 
    78420.1,
  87356.05, 86656.84, 88816.91, 90139.48, 89948.88, 89998.02, 89917.46, 
    91874.34, 95790.48, 101481.3, 101519.2, 101573.9, 101568, 87394.88, 
    78225.8,
  90984.32, 87814.3, 88289.41, 90151.45, 89883.23, 88906.19, 89514.3, 
    91356.27, 95550.62, 101392.7, 101435.5, 101568.7, 101519.4, 86212.22, 
    88168.32,
  93951.98, 89669.09, 88772.1, 89913.16, 89211.39, 86903.54, 88201.71, 
    90729.08, 100740.4, 101359.3, 101360.9, 101483.7, 101503.6, 93753.43, 
    96351.67,
  97100.26, 92423.42, 90800.07, 93228.22, 93547.38, 93686.73, 94660.41, 
    100653.3, 101293.9, 101303.1, 101326.6, 101394.3, 101486.7, 99267.4, 
    100444.4,
  101546.4, 101203.4, 97302.44, 94811.26, 94779.73, 93770.61, 91440.73, 
    91941.71, 86116.93, 81531.3, 79254.41, 79520.08, 82455.67, 81033.81, 
    91319.98,
  101348.1, 101406.1, 99136.76, 94002.35, 91239.23, 89385.34, 88161.33, 
    88500.16, 83613.68, 80895.32, 80098.52, 80755.48, 82941.98, 81827.93, 
    92661.2,
  92482.37, 88918.36, 93833.64, 92524.02, 86065.78, 84953.43, 87220.95, 
    86538.54, 81684.73, 79460.2, 78547.35, 79246.91, 80612.96, 82159.51, 
    94744.98,
  86375.52, 86216.88, 85499.45, 83865.3, 83606.85, 82149.66, 83012.62, 
    83330.12, 81086.09, 79865.49, 79521.9, 81056.27, 80685.43, 82679.81, 
    88669.76,
  87918.03, 86644.58, 87809.83, 86958.08, 86882.88, 85295.87, 84289.14, 
    83835.13, 82903.81, 84867.6, 99627.58, 100313.9, 90673.7, 91060.09, 
    83773.61,
  88012.12, 86186.29, 88640.79, 89491.66, 88640.81, 88195.09, 87490, 
    87876.02, 89421.23, 100240.2, 101136.4, 101166.9, 100986.2, 93126.62, 
    78253.17,
  87099.79, 86346.66, 88465.1, 89753.73, 89523.28, 89578.19, 89485.66, 
    91443.64, 95353.42, 100980.2, 100968, 101088.7, 100998, 87133.16, 77980.76,
  90886.69, 87605.38, 88048.12, 89875.47, 89529.42, 88519.75, 89097.14, 
    90940.52, 95126.28, 100919.1, 100903.8, 101043.3, 100937.2, 85934.88, 
    87711.05,
  93898.63, 89508.53, 88598.56, 89688.21, 88905.87, 86547.16, 87813.71, 
    90356.18, 100362.9, 100932.6, 100824.5, 100908.1, 100894.4, 93248.19, 
    95825.8,
  97119.16, 92398.23, 90745.32, 93145.03, 93374.92, 93485.2, 94418.17, 
    100445.5, 101050.9, 100920.5, 100853.2, 100846.4, 100867.6, 98661.64, 
    99828.54,
  101722.2, 101336.6, 97365.87, 94748.77, 94664.55, 93595.46, 91250.59, 
    91690.45, 85934.8, 81288.41, 79012.49, 79298.71, 82195.47, 80828.56, 
    91021.41,
  101600.9, 101466.6, 99204.47, 93987.41, 91146.8, 89206.09, 87931.43, 
    88206.47, 83360.29, 80599.38, 79827.7, 80498.73, 82679.19, 81608.38, 
    92321.98,
  92451.16, 88828.39, 93728.6, 92383.36, 85895.8, 84737.52, 86990.99, 
    86273.34, 81383.88, 79169.54, 78275.55, 78979.31, 80338, 81905.11, 
    94399.78,
  86364.49, 86425.3, 85525.23, 83757.42, 83467.42, 81977.22, 82818.23, 
    83116.18, 80818.34, 79594.45, 79249.68, 80764.55, 80410.32, 82408.42, 
    88343.95,
  87936.86, 86913.09, 87978.08, 87145.28, 86976.79, 85315.23, 84234.97, 
    83728.32, 82745.63, 84754.94, 99997.41, 100750, 90735.91, 90927.23, 
    83578.34,
  88313.04, 86486.41, 88943.76, 89831.61, 88866.34, 88397.76, 87610.83, 
    87957.73, 89579.67, 100907.7, 101827, 101752.3, 101374.4, 93156, 77926.12,
  87475.12, 86714.52, 88812.49, 90125.29, 89846.62, 89865.8, 89746.3, 
    91713.88, 95749.23, 101646.6, 101492.2, 101640.1, 101346.2, 87064.17, 
    77562.74,
  91318.2, 87994.41, 88414.74, 90260.07, 89907.43, 88852.15, 89427.35, 
    91231.5, 95509.84, 101567.2, 101498.7, 101667.6, 101370.8, 85882.73, 
    87347.73,
  94315.61, 89936.82, 88980.11, 90108.97, 89260.93, 86833.21, 88099.33, 
    90699.8, 100997.9, 101524.8, 101430.8, 101489.9, 101344.8, 93464.4, 
    95847.33,
  97525.51, 92837.2, 91167.99, 93585.55, 93823.37, 93973.34, 94862.12, 
    100904.5, 101449.3, 101406.7, 101362.5, 101344.1, 101283.7, 98939.37, 
    99943.15,
  101598.3, 101278.8, 97315.15, 94710.49, 94637.52, 93567.22, 91165.95, 
    91643.21, 85782.12, 81071.01, 78715.33, 78982.59, 81876.19, 80530.29, 
    90624,
  101493.7, 101422.3, 99219.41, 93997.62, 91121.84, 89161.79, 87890.52, 
    88151.48, 83173.48, 80371.95, 79557.24, 80213.42, 82379.43, 81320.56, 
    92045.56,
  92435.3, 88790.64, 93607.55, 92326.38, 85785.39, 84646.95, 86914.8, 
    86187.74, 81232.36, 78965.7, 77982, 78636.16, 80012.53, 81602.92, 94137.45,
  86346.27, 86300.91, 85466.07, 83714.63, 83405.48, 81888.58, 82695.41, 
    83004.06, 80667.77, 79365.71, 79014.37, 80564.06, 80100.41, 82126.48, 
    88113.5,
  87902.43, 86701.23, 87811.06, 86983.71, 86830.05, 85199.39, 84114.48, 
    83592.97, 82575.68, 84596.8, 99675.1, 100344.3, 90440.41, 90745.83, 
    83250.65,
  88115.15, 86294.49, 88759.91, 89652.62, 88700.32, 88222.27, 87430.8, 
    87792.01, 89324.28, 100441.8, 101411.1, 101344.5, 101090.7, 92911.97, 
    77611.44,
  87224.5, 86475.34, 88603.3, 89921.52, 89665.24, 89662.55, 89527.16, 
    91484.59, 95429.56, 101257.5, 101195.6, 101262.4, 101157.2, 86778.8, 
    77340.18,
  91050.88, 87759.08, 88184.77, 90038.14, 89690.89, 88630.34, 89197.61, 
    91001.37, 95248.81, 101234, 101201.1, 101287.3, 101165.8, 85513.2, 
    87379.76,
  94009.8, 89666.4, 88727.23, 89854.04, 89011.02, 86581.76, 87824.61, 
    90441.35, 100709.7, 101219, 101158.5, 101185.2, 101144.6, 93196.02, 
    95801.27,
  97226.29, 92575.95, 90910.04, 93313.82, 93550.11, 93713.16, 94588.62, 
    100619.3, 101162, 101138.6, 101120.8, 101111.8, 101112.8, 98804.8, 99953.7,
  100957.7, 100660.1, 96812.53, 94344.27, 94321.61, 93326.81, 90976.21, 
    91477.48, 85669.67, 80982.88, 78584.02, 78859.34, 81714.71, 80414.59, 
    90525.41,
  100934.8, 100983.2, 98759.75, 93628.75, 90817.83, 88946.11, 87721.41, 
    88027.6, 83092.57, 80311.8, 79498.27, 80151.77, 82310.09, 81212.12, 
    92010.66,
  92027.29, 88492.01, 93320.41, 92046.57, 85655.81, 84520.88, 86781.33, 
    86071.59, 81165.62, 78920.7, 77874.22, 78514.52, 79902.75, 81454.98, 
    94172.27,
  86036.28, 86088.13, 85280.02, 83556.04, 83289.41, 81815.74, 82623.2, 
    82936.38, 80620.02, 79313.99, 78971.34, 80600.88, 80009.19, 82020.96, 
    88051.91,
  87625.28, 86498.23, 87654.91, 86839.37, 86717.53, 85105.11, 84047.73, 
    83555.49, 82539.09, 84590.07, 99741.95, 100348.4, 90416.52, 90710.48, 
    83098.41,
  87895.52, 86111.26, 88640.78, 89531.27, 88591.63, 88150.86, 87378.97, 
    87776.65, 89348.44, 100562.3, 101499.6, 101442.8, 101145.9, 92900.73, 
    77448.13,
  87078.62, 86336.5, 88496.38, 89828, 89587.95, 89619.34, 89524.62, 91521.16, 
    95569.04, 101388.4, 101304.6, 101333.2, 101262.9, 86665.83, 77184.3,
  90870.74, 87650.13, 88116.03, 89971.95, 89668.61, 88624.57, 89215.62, 
    91020.06, 95361.94, 101347.4, 101320.4, 101357.9, 101228.7, 85429.03, 
    87260.17,
  93862.2, 89574.09, 88688.24, 89842.68, 89017.34, 86609.37, 87887.3, 
    90535.89, 100877.1, 101335.7, 101233, 101224.5, 101136.7, 93160.12, 
    95688.24,
  97085.3, 92478.76, 90904.33, 93353.34, 93619.56, 93836.84, 94749.86, 
    100840.4, 101325.2, 101248.9, 101176.1, 101120.8, 101058, 98691.65, 
    99779.66,
  100524.9, 100202.6, 96428.84, 94012.02, 93985.84, 93019.62, 90768.35, 
    91251.56, 85605.7, 80962.85, 78603.63, 78875.17, 81769.44, 80489.35, 
    90708.91,
  100378.3, 100481.7, 98262.03, 93224.69, 90525.02, 88716.42, 87506.43, 
    87834.44, 83043.8, 80259.3, 79473.64, 80120.85, 82325.68, 81244.12, 
    92214.26,
  91682.99, 88183.01, 92991.62, 91746.36, 85432.52, 84321.98, 86568.52, 
    85922.62, 81082.41, 78852.3, 77895.56, 78531.38, 79986.27, 81550.34, 
    94321.38,
  85733.92, 85712.38, 84954.5, 83280.45, 83035.92, 81611.78, 82430.88, 
    82758.07, 80498.52, 79264.03, 78925.94, 80541.21, 80035.27, 82055.16, 
    88130.44,
  87260.12, 86115.91, 87225.78, 86398.03, 86310.78, 84765.9, 83757.71, 
    83313.39, 82387.45, 84404.24, 99601.38, 100233.7, 90368.16, 90747.04, 
    83201.46,
  87481.62, 85683.07, 88100.55, 88997.32, 88129.12, 87714.66, 87031.64, 
    87475.47, 89097.95, 100391.8, 101441.9, 101324.8, 101062.8, 92860.73, 
    77602.49,
  86571.6, 85830.33, 87960.08, 89273.38, 89068.76, 89161.62, 89108.31, 
    91169.61, 95315.15, 101268, 101184.2, 101279.5, 101203.5, 86706.61, 
    77329.05,
  90221.38, 87051.86, 87538.92, 89376.31, 89106.22, 88157.56, 88803.89, 
    90743.84, 95140.09, 101241.6, 101217.1, 101380.3, 101215.7, 85490.23, 
    87361.14,
  93148.23, 88932.34, 88088, 89229.17, 88490.54, 86184.48, 87512.23, 
    90159.63, 100606.2, 101239.6, 101203.7, 101305.4, 101245.4, 93252.16, 
    95910.37,
  96362.06, 91791.19, 90261.29, 92723.98, 93026.57, 93186.79, 94221.82, 
    100433.3, 101153.6, 101204.1, 101239.3, 101284, 101286.3, 98951.93, 
    100104.9,
  100453.6, 100094.2, 96308.01, 93882.12, 93826.41, 92885.72, 90687.81, 
    91169.8, 85568.95, 80986.53, 78724.56, 79006.9, 81834.31, 80534.11, 
    90424.07,
  100291.6, 100356.2, 98096.62, 93034.37, 90363.33, 88592.23, 87380.29, 
    87739.73, 82996.21, 80261.02, 79504.94, 80134.77, 82291.45, 81282.61, 
    91728.95,
  91627.73, 88012.68, 92845.45, 91592.62, 85241.92, 84145.52, 86400.7, 
    85788.82, 80974.7, 78784.66, 77917.16, 78574.78, 79926.59, 81428.34, 
    93698.19,
  85615.13, 85517.12, 84800.32, 83070.19, 82800.52, 81390.23, 82216.45, 
    82543.77, 80285.78, 79118.92, 78745.95, 80222.45, 79907.86, 81853.21, 
    87814.64,
  87171.75, 85965.36, 87132.66, 86220.39, 86108.86, 84505.28, 83459.11, 
    82984.55, 82054.09, 83888.61, 98447.73, 99327.44, 89769.92, 90062.03, 
    82975.73,
  87330.68, 85512.38, 87938.76, 88763.62, 87879.59, 87400.62, 86668.22, 
    87033.12, 88547.01, 99362.02, 100364.6, 100285.8, 99997.57, 92216.64, 
    77432.31,
  86498.48, 85680.3, 87767.97, 89027.77, 88759.75, 88777.68, 88657.24, 
    90586.7, 94551.8, 100212.5, 100105.9, 100169.3, 100052.8, 86221.36, 
    77004.2,
  90266.15, 86966.39, 87418.98, 89190.45, 88826.61, 87788.64, 88356.12, 
    90194.67, 94457.87, 100282.5, 100223, 100267.2, 100076.7, 84894.16, 
    86613.35,
  93247.57, 88893.97, 87977.7, 89042.86, 88232.31, 85849.54, 87081.23, 
    89655.32, 99816.37, 100395.8, 100271, 100320.6, 100199.5, 92359.59, 
    95017.25,
  96449.48, 91808.58, 90175.36, 92591.19, 92865, 92971.38, 93874.34, 
    99872.96, 100444.2, 100390, 100352, 100349.8, 100298.9, 97984.9, 99219.42,
  101357.8, 100978.2, 97024.49, 94456.37, 94375.63, 93341.84, 91053.61, 
    91522.36, 85772.98, 81105.49, 78794.71, 79092.23, 81919.67, 80595.7, 
    90558.17,
  101156, 101164.1, 98865.52, 93642.75, 90851.16, 88961.11, 87719.45, 
    88035.02, 83188.52, 80422.24, 79636.16, 80302.89, 82428.77, 81411.15, 
    91954.72,
  92178.3, 88512.61, 93496.65, 92135.6, 85620.85, 84478.01, 86772.51, 
    86081.59, 81204.34, 78960.61, 78062.42, 78739.02, 80079.38, 81634.65, 
    94022.3,
  86019.44, 85930.38, 85173.69, 83460.23, 83195.77, 81729.68, 82584.2, 
    82890.67, 80614.39, 79387.34, 79063.41, 80537.43, 80192.74, 82140.26, 
    88026.51,
  87591.99, 86402.93, 87546.08, 86675.27, 86571.87, 84961.88, 83925.82, 
    83445.59, 82476.23, 84538.81, 99724.5, 100456.5, 90486.02, 90655.98, 
    83316.18,
  87730.13, 85950.6, 88429.46, 89307.94, 88419.05, 87979.12, 87256.22, 
    87666.08, 89302.73, 100561.4, 101545.2, 101445.8, 101132.7, 92849.04, 
    77715.62,
  86815.03, 86089.27, 88239.11, 89574.52, 89362.07, 89428.81, 89362.78, 
    91403.92, 95497.44, 101381.7, 101262.1, 101365.1, 101147.2, 86762.95, 
    77273.7,
  90587.71, 87312.11, 87812.08, 89675.29, 89379.43, 88405.27, 89036.67, 
    90942.92, 95300.39, 101349.2, 101287.2, 101427.1, 101164, 85535.14, 
    87156.12,
  93540.25, 89222.2, 88317.18, 89471.84, 88724.35, 86402.33, 87714.2, 
    90337.07, 100708.5, 101338.4, 101248.3, 101325.8, 101190.6, 93215.89, 
    95759.52,
  96713.56, 92053.42, 90448.35, 92910.31, 93202.03, 93368.89, 94353.86, 
    100534.3, 101252.5, 101279.7, 101277.8, 101304.9, 101252.9, 98900.98, 
    99958.86,
  101096.8, 100705.5, 96757.85, 94155.95, 94044.5, 93000.7, 90690.2, 
    91150.55, 85415.53, 80721.2, 78443.09, 78776.6, 81746.06, 80463.45, 
    90688.81,
  100937.3, 100868.8, 98572.49, 93318.84, 90491.04, 88570.38, 87243.19, 
    87599.02, 82766.15, 79988.09, 79279.82, 79963.2, 82215.01, 81241.48, 
    91982.73,
  91833.97, 88184.82, 93152.69, 91790.18, 85186.62, 84041.38, 86302.13, 
    85614.06, 80720.34, 78505.08, 77685.64, 78379.47, 79819.94, 81409.89, 
    93914.6,
  85636.45, 85699.77, 84769.85, 83047.08, 82746.85, 81231.04, 82060.84, 
    82353.7, 80079.7, 78935.12, 78578.64, 80087.23, 79883.77, 81821.52, 
    87928.29,
  87221.05, 86242.91, 87281.16, 86402.02, 86229.2, 84543.66, 83448.51, 
    82929.5, 81992.26, 83964.77, 98932.81, 99610.84, 89879.51, 90166.2, 
    83051.69,
  87614.13, 85777.46, 88219.83, 89048.47, 88090.12, 87591.12, 86813.44, 
    87182.84, 88755.98, 99808.02, 100663.1, 100624.5, 100389.7, 92439.34, 
    77458.8,
  86861.09, 86061.8, 88146.27, 89383.38, 89095.47, 89056.38, 88954.35, 
    90909.52, 94890.1, 100590.8, 100467.3, 100542, 100388.9, 86335.94, 
    77117.51,
  90761.77, 87397.73, 87814.09, 89589.63, 89174.88, 88065.74, 88652.08, 
    90461.87, 94759.55, 100647.4, 100532.4, 100624.5, 100495.4, 85170.22, 
    87019.02,
  93859.02, 89409.93, 88465.8, 89525.97, 88598.82, 86136.1, 87389.18, 
    89992.46, 100278.1, 100742, 100613.2, 100639.9, 100560.4, 92758.21, 
    95642.55,
  97174.77, 92404.49, 90789.49, 93161.2, 93337.95, 93403.19, 94255.17, 
    100247.5, 100881.6, 100883.3, 100840.4, 100842.8, 100818.1, 98605.96, 
    99882.25,
  101847.5, 101492.8, 97469.06, 94833.98, 94748.09, 93646.91, 91218.23, 
    91754.47, 85793.59, 81022.8, 78608.45, 78865.69, 81739.56, 80340.28, 
    90433.34,
  101883.4, 101720.1, 99416.7, 94108.27, 91198.97, 89211.87, 87900.76, 
    88169.8, 83130.56, 80331.9, 79468.76, 80136.53, 82287.09, 81167.48, 
    91929.69,
  92553, 88995.35, 93929.52, 92480.62, 85855.25, 84726.59, 86972.73, 
    86166.48, 81154.27, 78893.62, 77894.88, 78579.63, 79894.77, 81443.36, 
    93973.11,
  86490.41, 86605.98, 85597.23, 83870.02, 83544.22, 81979.72, 82780.05, 
    83040.14, 80658.39, 79321.04, 79043.98, 80576.07, 80003.87, 82022.07, 
    87904.12,
  88088.95, 87074.12, 88098.38, 87232.91, 87019.53, 85336.52, 84211.41, 
    83661.56, 82620.64, 84801.29, 100115.5, 100701.8, 90560.57, 90780.84, 
    83021.05,
  88443.44, 86575.77, 89061.65, 89888.2, 88925.26, 88430.48, 87624.53, 
    87993.15, 89609.48, 100830.9, 101664.6, 101619.6, 101294.3, 92936.41, 
    77352.82,
  87630.22, 86824.03, 88926.45, 90188.81, 89914.05, 89884.47, 89759.34, 
    91725.55, 95724.02, 101598.5, 101495.1, 101450.3, 101282.9, 86699.2, 
    77099.87,
  91481.5, 88129.02, 88541.35, 90360.79, 89986.9, 88885.52, 89443.33, 
    91231.62, 95563.27, 101551.8, 101454.1, 101467.6, 101238.6, 85371.16, 
    87232.59,
  94528.52, 90099.04, 89107.34, 90207.08, 89322.72, 86856.83, 88077.44, 
    90740.88, 101013.3, 101539.6, 101415.1, 101396.2, 101214, 93191.09, 
    95830.3,
  97788.59, 93025.35, 91341.83, 93741.16, 93947.32, 94100.59, 94968.95, 
    101017, 101543.3, 101497.2, 101403.2, 101358.7, 101279, 98906.27, 100024.3,
  101899.2, 101511, 97541.72, 94941.66, 94903.9, 93877.9, 91535.95, 92016.2, 
    86165.77, 81386.91, 79030.7, 79323.98, 82225.94, 80853.18, 91024.27,
  101650, 101649.9, 99390.44, 94127.48, 91293.84, 89375.74, 88099.56, 
    88413.03, 83492.73, 80636.31, 79826.43, 80489.48, 82704.74, 81657.27, 
    92424.3,
  92580.06, 88819.14, 93779.23, 92514.38, 85885.37, 84717.71, 87033.05, 
    86375.29, 81389.31, 79091.93, 78182.19, 78869.83, 80254.3, 81847.15, 
    94422.88,
  86353.49, 86221.73, 85396.08, 83657.36, 83318.11, 81843.73, 82670.57, 
    83011.3, 80673.16, 79446.13, 79080.48, 80601.45, 80271.9, 82277.57, 
    88315.25,
  87906.24, 86728.12, 87855.58, 86964.47, 86783.41, 85096.78, 84004.94, 
    83507.35, 82537.26, 84607.23, 99791.63, 100593.5, 90550.55, 90798.53, 
    83433.46,
  88132.74, 86318.17, 88775.14, 89637.8, 88670.86, 88160.77, 87379.38, 
    87762.66, 89445.69, 100716, 101652.7, 101507.7, 101170.8, 93030.45, 
    77715.73,
  87343.14, 86576.73, 88681.14, 89983.07, 89679.39, 89669.52, 89536.2, 
    91579.53, 95693.37, 101565.5, 101414, 101473.9, 101223.3, 86813.89, 
    77257.55,
  91271.27, 87882.12, 88298.8, 90155.73, 89749.97, 88663.44, 89236.94, 
    91129.53, 95485.15, 101509.9, 101408, 101493.6, 101247.7, 85534.53, 
    87117.83,
  94395.55, 89889.19, 88943.34, 90076.99, 89165.33, 86663.78, 87920, 
    90585.55, 101048.4, 101516.2, 101350.2, 101337.4, 101237.1, 93180.86, 
    95739.15,
  97766.76, 92955.78, 91303.84, 93754.12, 93962.7, 94122.26, 94994.08, 
    101120.6, 101589.3, 101444.5, 101341.6, 101267.9, 101214, 98826.5, 
    99933.57,
  101547.4, 101121.6, 97142.22, 94491.57, 94416.98, 93368.64, 91060.38, 
    91478.99, 85718.13, 80902.3, 78657.48, 78946.45, 81927.92, 80639.3, 
    90777.51,
  101550.2, 101429.2, 99078.62, 93726.98, 90855.2, 88941.63, 87637.66, 
    87906.45, 83036.09, 80139.23, 79437.58, 80095.55, 82354.7, 81382.75, 92069,
  92320.3, 88693.36, 93735.05, 92274.06, 85608.8, 84404.97, 86788.85, 
    86019.32, 81003.02, 78683.75, 77852.34, 78546.32, 79994.1, 81591.17, 
    94039.97,
  86204.27, 86357.79, 85406.35, 83596.58, 83294.68, 81744.72, 82619.71, 
    82844.52, 80431, 79203.47, 78931.76, 80401.97, 80062.15, 82055.43, 
    88110.08,
  87945.29, 86959, 88073.47, 87167.02, 86988.05, 85279.64, 84168.09, 
    83653.41, 82616.62, 84873.71, 100444.6, 101083.4, 90702.3, 90814.19, 
    83329.81,
  88390.62, 86551.84, 89177.7, 90005.73, 89020.5, 88527.32, 87753.16, 
    88180.27, 89885.29, 101439.6, 102294, 102158.1, 101836, 93182.23, 77721.52,
  87647.78, 86880.74, 89101.35, 90386.95, 90125.66, 90099.71, 90006.78, 
    92087.09, 96237.27, 102172.5, 101993.7, 102030.8, 101784.9, 86966.04, 
    77296.84,
  91665.73, 88266.41, 88780.72, 90659.38, 90275.98, 89152.08, 89759.73, 
    91631.7, 96088.77, 102175.5, 102047, 102119.8, 101808.5, 85917.5, 87457.17,
  94897.19, 90364.35, 89430.79, 90571.73, 89650.59, 87125.61, 88397.8, 
    91179.3, 101742.2, 102139.9, 101959.7, 101955.4, 101778.2, 93693.24, 
    96297.2,
  98316.42, 93441.22, 91833.26, 94317.59, 94565.84, 94723.7, 95623.19, 
    101787.1, 102198.7, 102090.7, 101961.7, 101888.6, 101802.2, 99423.39, 
    100529.1,
  102259.4, 101943.1, 97783.72, 95110.62, 95035.62, 93876.84, 91377.71, 
    91809.79, 85740.8, 80885.33, 78469.02, 78768.3, 81688.86, 80276.55, 
    90613.22,
  102384.3, 102166.9, 99819.49, 94450.79, 91487.23, 89461.34, 88162.23, 
    88356.25, 83179.29, 80296.69, 79409.94, 80091.95, 82299.31, 81187.84, 
    92197.09,
  92826.2, 89296.27, 94345.09, 92845.42, 86104.77, 84959.33, 87286.1, 
    86431.97, 81333.3, 78973.04, 77915.45, 78606.3, 79946, 81632, 94346.24,
  86695.3, 86903.42, 85862.94, 84111.73, 83816.04, 82224.34, 83085.54, 
    83347.3, 80877.46, 79514.02, 79331.9, 80859.7, 80226.87, 82358.38, 
    88213.25,
  88338.76, 87397.02, 88488.7, 87614.48, 87419.71, 85714.2, 84584.67, 
    84054.7, 82950.1, 85292.64, 101029.9, 101525.4, 91126.68, 91325.88, 
    83292.74,
  88783.9, 86902.24, 89555.5, 90413.95, 89448.63, 88946.5, 88165.12, 
    88570.91, 90293.17, 101832.9, 102598.6, 102561, 102271.1, 93628.84, 
    77678.79,
  87971.68, 87160.94, 89400.07, 90740.39, 90511.2, 90500.78, 90427.25, 
    92470.15, 96630.27, 102608.8, 102493.4, 102474.9, 102259.1, 87311.35, 
    77484.91,
  91910.53, 88517.16, 89032.95, 90917.93, 90598.48, 89491.02, 90112.54, 
    91956.45, 96536.67, 102607.2, 102509.2, 102532.4, 102316.6, 86071.2, 
    87954.7,
  95067.88, 90561.86, 89621.84, 90785.45, 89897, 87423.09, 88729.68, 
    91567.55, 102143.4, 102596.6, 102487.8, 102483, 102337.2, 94053.91, 
    96837.59,
  98409.63, 93567.49, 91939.94, 94428.73, 94689.46, 94885.98, 95841.88, 
    102063.9, 102602.1, 102591.3, 102503.6, 102484.6, 102393, 99968.74, 
    101099.2,
  102318.7, 102027.2, 97987.31, 95433.16, 95458.14, 94370.3, 91922.52, 
    92447.75, 86320.01, 81547.02, 79106.48, 79448, 82364.98, 80978.13, 
    91467.23,
  102412.6, 102320, 99983.62, 94658.46, 91784.07, 89827.25, 88593.1, 
    88906.33, 83712.55, 80942.96, 80072.49, 80788.24, 83011.73, 81848.1, 
    92978.48,
  93007.42, 89429.87, 94542.03, 93102.61, 86417, 85286.34, 87635.37, 
    86864.87, 81822.57, 79496.99, 78433.97, 79144.99, 80530.86, 82149.78, 
    95176.25,
  86750.78, 86972.79, 85971.12, 84236.98, 83972.25, 82433.07, 83301.58, 
    83610.2, 81227.2, 79883.41, 79623.14, 81261.64, 80683, 82763.79, 88898.65,
  88456.3, 87479.02, 88538.69, 87710.62, 87552.38, 85870.98, 84763.4, 
    84233.2, 83189.33, 85357.36, 100951.6, 101572.4, 91377.59, 91737.07, 
    83803.95,
  88812.05, 86911.86, 89492.13, 90372.18, 89449.62, 88983.98, 88206.17, 
    88607.09, 90257.2, 101664.8, 102622.2, 102647.7, 102471.2, 93955.18, 
    78058.66,
  88010.05, 87197.55, 89386.84, 90679.94, 90463.94, 90472.43, 90394.85, 
    92398.93, 96443.22, 102418.5, 102450.1, 102495.5, 102539.2, 87511.5, 
    77836.66,
  91860.52, 88504.83, 88997.21, 90844.23, 90520.96, 89445.73, 90046.31, 
    91866.28, 96278.82, 102367, 102419, 102513.8, 102458, 86259.59, 88251.98,
  94959.16, 90516.11, 89581.81, 90714.25, 89834.59, 87393.7, 88664.26, 
    91394.3, 101796.6, 102350.7, 102341.2, 102412, 102385.6, 94232.54, 
    96857.67,
  98228.45, 93460.71, 91840.3, 94260.73, 94489.59, 94669.66, 95581.8, 101653, 
    102254.3, 102289.9, 102283.5, 102331.4, 102339.4, 99985.67, 101129.9,
  102237.9, 101917.7, 97864.95, 95344.44, 95310.23, 94204.84, 91761.17, 
    92287.2, 86236.62, 81549.12, 79133.49, 79489.77, 82460.02, 81075.58, 
    91564.47,
  102363.4, 102219.7, 99920, 94599.87, 91727.45, 89778.52, 88522.17, 
    88822.23, 83708.95, 80972.76, 80099.44, 80815.84, 83037.59, 81925.68, 
    93029.96,
  92935.22, 89433.35, 94436.58, 92998.37, 86411.43, 85307.15, 87601.26, 
    86825.29, 81870.92, 79575.1, 78575.69, 79301.77, 80684.01, 82297.87, 
    95173.56,
  86897.38, 87058.04, 86033.91, 84351.83, 84075.02, 82533.9, 83395.88, 
    83692.33, 81318.87, 79972.05, 79706.7, 81278.16, 80786.62, 82853.96, 
    88910.93,
  88497.91, 87510.79, 88553.3, 87735.37, 87574.56, 85920.56, 84819.48, 
    84295.45, 83250.85, 85440.1, 100740.9, 101348.1, 91332.77, 91655.52, 
    83932.69,
  88875.74, 86997.66, 89519.57, 90361.43, 89465.38, 89001.08, 88240.14, 
    88631.03, 90254.05, 101389.9, 102277.3, 102303.8, 102085.9, 93812.44, 
    78228.45,
  88018.84, 87235.78, 89373.23, 90641.83, 90430.44, 90442.6, 90375.28, 
    92353.38, 96327.38, 102166.1, 102149.1, 102221.8, 102157.6, 87547.75, 
    77966.39,
  91831.18, 88533.25, 88992.93, 90822.68, 90484.77, 89446.42, 90053.8, 
    91842.67, 96176.85, 102110.2, 102092.7, 102191.3, 102096.8, 86267.83, 
    88097.3,
  94855.77, 90484.81, 89539.25, 90651.55, 89800.7, 87396.64, 88645.18, 
    91323.32, 101535.3, 102061.5, 102030.4, 102072.5, 102022.5, 94036.88, 
    96572.8,
  98099.34, 93374.4, 91743.42, 94133.47, 94362.17, 94531.8, 95438.1, 
    101400.3, 101967.6, 101970.1, 101948, 101962.3, 101966.1, 99638.17, 
    100731.5,
  102476.2, 102121.5, 98086.62, 95552.81, 95507.59, 94429.41, 92002.47, 
    92557.86, 86519.79, 81847.45, 79474.55, 79761.14, 82734.06, 81300.27, 
    91688.86,
  102424.1, 102353.3, 100070.6, 94826.73, 91940.05, 90013.46, 88766.48, 
    89065.51, 83991.34, 81291.67, 80422.41, 81099.52, 83304.4, 82139.27, 
    93126.05,
  93177.15, 89651.98, 94636.73, 93232.4, 86658.45, 85557.41, 87832.76, 
    87064.18, 82144.36, 79853.45, 78789.43, 79509.28, 80899.57, 82487.7, 
    95242.16,
  87025.73, 87184.84, 86228.3, 84556.76, 84280.17, 82763.86, 83605.13, 
    83909.38, 81577.25, 80229.87, 80006.37, 81558.22, 80954.62, 83075.67, 
    89067.85,
  88716.43, 87671.77, 88676.62, 87848.4, 87675.36, 86064.3, 84979.21, 
    84461.98, 83437.07, 85595.34, 100569.4, 101211.5, 91401.62, 91768.04, 
    84064.98,
  88979.46, 87148.17, 89597.67, 90434.88, 89515.98, 89062.6, 88313.54, 
    88706.32, 90281.77, 101213.2, 102126.6, 102227.4, 102040.1, 93864.27, 
    78465.69,
  88079.14, 87329.31, 89418.62, 90685.47, 90452.38, 90457.95, 90368.31, 
    92317.38, 96239.8, 101972.4, 102013.8, 102061.3, 102107.3, 87663.72, 
    78233.68,
  91836.99, 88587.49, 89009.73, 90810.78, 90475.32, 89440.77, 90031.52, 
    91823.7, 96034.05, 101883.7, 101934.2, 102043.3, 102013.4, 86373.32, 
    88288.48,
  94802.84, 90482.55, 89528.06, 90611.19, 89794.97, 87408.13, 88641.12, 
    91225.76, 101324.8, 101860.5, 101853.6, 101933.3, 101932.3, 94069.23, 
    96583.68,
  98013.93, 93319.32, 91665.55, 94011.2, 94241.45, 94387.07, 95277.26, 
    101187.2, 101795.4, 101801.8, 101790.5, 101818.7, 101842.9, 99563.44, 
    100682.8,
  102272.7, 101939.2, 98051.91, 95611.04, 95603.23, 94581.82, 92252.17, 
    92776.02, 86886.78, 82198.99, 79862.27, 80150.1, 83077.12, 81652.98, 
    91864.62,
  102221.8, 102257.3, 99939.77, 94787.42, 92045.89, 90181.28, 88932.27, 
    89259.09, 84316.25, 81570.75, 80748.91, 81406.87, 83594.05, 82470.91, 
    93280.05,
  93213.28, 89729.52, 94710.58, 93351.72, 86805.81, 85727.8, 88022.27, 
    87319.34, 82387.11, 80132.99, 79162.3, 79850.14, 81200.01, 82774.13, 
    95350.94,
  87050.79, 87131, 86284.05, 84650.72, 84392.48, 82919.2, 83781.8, 84094.85, 
    81803.03, 80539.49, 80193.8, 81755.08, 81294.07, 83293.1, 89250.9,
  88695.34, 87646.67, 88707.43, 87896.88, 87771.64, 86176.89, 85132.98, 
    84636.4, 83661.41, 85686.44, 100664.8, 101310.1, 91511.83, 91850.66, 
    84340.16,
  88964.38, 87147.1, 89605.61, 90477.4, 89590.08, 89154.78, 88426.92, 
    88823.37, 90396.74, 101331.1, 102230, 102248.5, 101992.3, 93958.22, 
    78747.91,
  88044.84, 87340.56, 89459.11, 90745.83, 90525.69, 90561.24, 90475.05, 
    92447.44, 96358.35, 102101.8, 102042.6, 102157.3, 102031.6, 87873.47, 
    78455.8,
  91785.85, 88573.08, 89031.23, 90852.81, 90539.48, 89541.07, 90142.17, 
    91977.47, 96177.16, 102066.6, 102016.1, 102167.1, 101991.8, 86610.2, 
    88352.86,
  94742.03, 90463.95, 89565.74, 90671.23, 89886.86, 87533.59, 88789.52, 
    91354.22, 101435.6, 102018.7, 101959.2, 102041.1, 101954.4, 94167.79, 
    96588.34,
  97945.06, 93287.08, 91682.88, 94059.32, 94319.22, 94470.2, 95377.7, 
    101293.8, 101886.9, 101890.5, 101862.5, 101864.9, 101851.3, 99560.22, 
    100578.8,
  101849.9, 101490.7, 97674.25, 95313.91, 95356.38, 94391.48, 92083.48, 
    92622.58, 86764.23, 82142.54, 79811.5, 80120.75, 83031.41, 81620.22, 
    91781.28,
  101840.1, 101831.1, 99533.82, 94487.27, 91832.04, 90021.93, 88799.48, 
    89153.95, 84232.93, 81527.48, 80705.38, 81380.53, 83558.8, 82476.56, 
    93244.09,
  92950.57, 89489.08, 94413.28, 93087.62, 86670.45, 85650.91, 87924.1, 
    87236.59, 82345.11, 80115.91, 79149.54, 79848.62, 81194.02, 82772.28, 
    95291.95,
  86866.16, 87023.05, 86149.6, 84533.74, 84302.66, 82858.66, 83733.39, 
    84054.52, 81779.05, 80520.93, 80204.08, 81757.27, 81295.59, 83300.18, 
    89245.8,
  88473.69, 87548.95, 88580.16, 87786.45, 87677.27, 86106.25, 85090.01, 
    84604, 83636.91, 85671.91, 100615.7, 101238.4, 91512.14, 91831.2, 84352.52,
  88807.63, 87041.7, 89502.2, 90382.37, 89517.48, 89101.15, 88386.78, 
    88790.45, 90374.48, 101287.5, 102159.9, 102150.1, 101957.2, 93948.12, 
    78761.02,
  87950.55, 87252.44, 89368.95, 90678.74, 90485.38, 90530.13, 90456.16, 
    92412.77, 96326.8, 102046.4, 102020.9, 102086, 102049.1, 87840.13, 
    78515.62,
  91666.01, 88493.75, 88960.8, 90797.7, 90507.28, 89532.12, 90142.99, 
    91958.73, 96171.08, 102032.7, 102019.2, 102115.5, 102025.2, 86603.07, 
    88520.41,
  94592.18, 90393.23, 89518.68, 90631.72, 89863.84, 87542.39, 88801.48, 
    91378.61, 101467.8, 101999.5, 101980.7, 102041.8, 101997.4, 94219.02, 
    96765.99,
  97787.13, 93185.81, 91632.48, 94017.66, 94283.24, 94461.18, 95397.02, 
    101331.1, 101928.5, 101939.7, 101939.7, 101963.5, 101962.1, 99685.37, 
    100755.2,
  101437.7, 101136, 97388, 95109.3, 95162.56, 94209.99, 91887.8, 92456.12, 
    86604.15, 82031.35, 79723.54, 80037.7, 82978.93, 81556.62, 91757.92,
  101435.6, 101446.4, 99200.51, 94254.78, 91665.84, 89880.71, 88668.48, 
    89038.39, 84120.78, 81457.59, 80627.16, 81310.55, 83511.73, 82381.17, 
    93179.05,
  92664.12, 89265.39, 94166.42, 92866.58, 86523.52, 85532.99, 87796.27, 
    87118.26, 82263.43, 80051.64, 79092.88, 79800.62, 81161.59, 82726.25, 
    95240.45,
  86627.05, 86820.41, 85949.44, 84387.52, 84174.89, 82765.2, 83651.08, 
    83988.87, 81727.26, 80461.36, 80159.14, 81716.62, 81243.59, 83284.91, 
    89219.04,
  88206.48, 87354.19, 88379.87, 87598.56, 87515.88, 85977.79, 84988.96, 
    84524.02, 83573.4, 85622.93, 100505.9, 101096.9, 91410.7, 91823.41, 
    84317.43,
  88580.02, 86818.63, 89283.53, 90152.92, 89322.99, 88941.13, 88258.55, 
    88682.39, 90269.43, 101141.1, 102048.2, 102030.3, 101860.3, 93868.04, 
    78843.59,
  87736.25, 87046.57, 89171.35, 90459.64, 90293.48, 90359.03, 90333.91, 
    92302.08, 96237.43, 101948.1, 101934.2, 101978.1, 101973.8, 87800.62, 
    78640.8,
  91344.02, 88250.8, 88744.38, 90580.62, 90325.11, 89395.15, 90044.34, 
    91869.41, 96064.45, 101905.8, 101936.8, 102037.5, 101963.4, 86595.84, 
    88609.65,
  94246.43, 90132.98, 89300.9, 90431.37, 89702.34, 87443.96, 88737.28, 
    91308.11, 101317.1, 101881.8, 101912.3, 102021.3, 101977.7, 94240.25, 
    96844.31,
  97410.48, 92877.92, 91379.3, 93786.94, 94076.7, 94262.32, 95241.73, 
    101169.6, 101794.5, 101869, 101916.6, 102001.2, 102030, 99771.55, 100909.9,
  101313.4, 101005.6, 97219.75, 94897.96, 94917.16, 93945.4, 91615.1, 
    92182.86, 86335.01, 81807.8, 79510.81, 79801.47, 82791.73, 81386.35, 
    91642.59,
  101179.7, 101223.6, 98983.99, 94059.92, 91455.3, 89648.57, 88446.76, 
    88807.16, 83891.71, 81249.84, 80419.35, 81105.29, 83310.23, 82212.27, 
    92988.48,
  92431.84, 89081.3, 93962.48, 92658.8, 86330.31, 85333.37, 87586.73, 
    86891.34, 82067.34, 79860.12, 78917.55, 79609.98, 80977.51, 82543.5, 
    95018.62,
  86460.83, 86582.93, 85762.97, 84210.39, 83996.32, 82590.07, 83466.55, 
    83797.08, 81553.55, 80276.54, 79979.56, 81512.91, 81067.3, 83068.09, 
    89025.7,
  88035.49, 87066.61, 88129.51, 87360.23, 87284.26, 85766.34, 84800.67, 
    84347.88, 83394.48, 85427.27, 100265.6, 100845.8, 91190.76, 91592.34, 
    84153.31,
  88342.78, 86571.73, 89008.17, 89867.77, 89064.82, 88698.12, 88043.56, 
    88477.28, 90073.66, 100915.4, 101813.7, 101772.8, 101595.4, 93646.91, 
    78725.04,
  87471.83, 86791.19, 88898.02, 90162.88, 90007.59, 90092.52, 90092.8, 
    92058.22, 96026.65, 101730.6, 101705.6, 101733.7, 101733.2, 87612.62, 
    78508.8,
  91083.85, 87988.14, 88474.59, 90285.63, 90031.27, 89116.53, 89786.23, 
    91618.91, 95879.81, 101731.6, 101740.2, 101822.5, 101750.6, 86397.08, 
    88497.33,
  94001.13, 89883.62, 89030.12, 90151.96, 89430.59, 87207.36, 88518.36, 
    91083.8, 101131.9, 101752.6, 101770.5, 101840.4, 101773.2, 94115.13, 
    96920.49,
  97169.11, 92612.62, 91122.66, 93496.64, 93781.2, 93942.18, 94937.69, 
    100853.1, 101622.9, 101764.2, 101826.9, 101915.9, 101920.3, 99775.71, 
    101116.4,
  101407, 101094.4, 97225.89, 94850.74, 94852.02, 93874.75, 91558.13, 
    92117.23, 86318.27, 81770.43, 79481.6, 79741.62, 82701.09, 81303.35, 
    91710.45,
  101331.3, 101355.8, 99094.4, 94061.59, 91395.45, 89594.64, 88385.13, 
    88729.89, 83852.8, 81188.08, 80371.55, 81018.23, 83211.39, 82066.1, 
    92955.32,
  92557.55, 89093.67, 93944.84, 92649.15, 86304.88, 85287.03, 87517.24, 
    86819.41, 82018.89, 79807.63, 78837.65, 79497.45, 80871.29, 82412.53, 
    94991.41,
  86578.84, 86642.35, 85816.59, 84219.4, 83979.54, 82554.59, 83409.4, 
    83724.04, 81474.98, 80199.34, 79910.65, 81463.78, 80957.61, 82967.47, 
    88942.61,
  88126.45, 87118.01, 88169.49, 87378.89, 87278.55, 85738.27, 84742.78, 
    84272.76, 83321.55, 85340.98, 100113.7, 100668.5, 91071.1, 91442.41, 
    84010.1,
  88423.44, 86638.67, 89073.97, 89915.52, 89071.1, 88671.95, 87984.94, 
    88402.02, 89972.38, 100788.1, 101713.5, 101635.9, 101449.8, 93503.09, 
    78630.65,
  87537.68, 86848.26, 88953.95, 90211.92, 90039.42, 90074.3, 90031.05, 
    91969.61, 95933.77, 101632.7, 101576.1, 101588.1, 101592.5, 87475.45, 
    78383.66,
  91161.7, 88052.47, 88547.99, 90328.42, 90046.34, 89098.87, 89731.34, 
    91534.52, 95811.7, 101654.1, 101619.5, 101689.2, 101606.8, 86249.82, 
    88415.43,
  94053.72, 89941.91, 89100.36, 90185.95, 89423.03, 87156.82, 88439, 
    90991.42, 101113.7, 101694.2, 101653.2, 101700.8, 101599, 93967.1, 
    96863.38,
  97162.87, 92690.56, 91198.85, 93562.3, 93810.6, 93967.06, 94921.76, 
    100894.5, 101662, 101746, 101788.5, 101849, 101807.1, 99701.88, 101095.8,
  101263.6, 100931.1, 97115.23, 94693.09, 94676.29, 93697.52, 91442.45, 
    91978.05, 86271.41, 81716.8, 79448.98, 79716.2, 82667.92, 81274.26, 
    91751.71,
  101104.2, 101161.3, 98937.79, 93912.05, 91245.23, 89456.88, 88245.48, 
    88584.39, 83771.62, 81115.03, 80329.63, 80968.05, 83184.39, 82053.46, 
    93122.12,
  92448.67, 88952.84, 93779.64, 92489.14, 86164.88, 85135.52, 87369.23, 
    86702.7, 81916.78, 79732.05, 78765.57, 79424.03, 80826.38, 82405.48, 
    95241.67,
  86460.04, 86430.95, 85691.1, 84071.98, 83831.91, 82409.68, 83260.45, 
    83597.91, 81359.8, 80109.09, 79815.7, 81393.91, 80899.19, 82944.55, 
    89100.28,
  88005.19, 86866.27, 87985.23, 87174.63, 87103.16, 85565.91, 84584.02, 
    84129.07, 83199.51, 85201.15, 100026.4, 100600.4, 90991.23, 91459.8, 
    84066.19,
  88187.67, 86430.2, 88844.09, 89692.12, 88851.22, 88453.23, 87787.53, 
    88220.22, 89794.03, 100757.1, 101669.4, 101598.2, 101426.8, 93515.89, 
    78618.33,
  87288.38, 86584.52, 88696.17, 89959.04, 89783.01, 89840.73, 89827.93, 
    91817.95, 95884.02, 101556.6, 101498.7, 101524.4, 101567.7, 87444.48, 
    78372.95,
  90903.32, 87765.89, 88269.77, 90065.32, 89784.64, 88845.7, 89521.65, 
    91398.62, 95720.62, 101567.3, 101548.7, 101605.1, 101570.2, 86231.33, 
    88540.05,
  93791.3, 89630.22, 88805.01, 89907.28, 89183.9, 86954.31, 88265.41, 
    90866.35, 101046, 101601.3, 101565.7, 101625.7, 101562, 93959.54, 97008.01,
  96913.42, 92376.8, 90887.38, 93267.77, 93542.67, 93686.15, 94672.6, 
    100771.2, 101603.8, 101667.8, 101722.5, 101801.9, 101784.9, 99772.62, 
    101234.8,
  101595.5, 101206.3, 97298.87, 94707.25, 94599.15, 93519.55, 91183.59, 
    91641.12, 85990.57, 81456.32, 79214.24, 79516.7, 82615.29, 81330.9, 
    91955.2,
  101381.5, 101306.6, 99070.04, 93952.8, 91143.59, 89241.46, 87974.8, 
    88261.08, 83461.09, 80804.74, 80057.75, 80746.88, 83105.55, 82069.84, 
    93412.37,
  92498.07, 88866.49, 93740.42, 92387.61, 85980.89, 84883.38, 87087.84, 
    86381.07, 81609.08, 79455.86, 78561.25, 79251.86, 80765.09, 82419.33, 
    95494.8,
  86478.23, 86474, 85618.95, 83924.42, 83647.62, 82178.46, 82989.59, 
    83276.52, 81036.38, 79819.68, 79521.28, 81083.45, 80726.5, 82911.85, 
    89289.41,
  88047.08, 86964.28, 88019.82, 87153.54, 86995.98, 85414.12, 84390.66, 
    83888.63, 82909.56, 84897.9, 99649.41, 100232.7, 90669.59, 91378.07, 
    84128.56,
  88321.13, 86554.76, 88957.88, 89782.73, 88870.02, 88404.7, 87654.61, 
    88015.72, 89570.91, 100363.4, 101245, 101136.3, 101090.1, 93350.73, 
    78536.98,
  87560.97, 86803, 88840.7, 90086.64, 89830.98, 89815.73, 89709.54, 91594.84, 
    95506.1, 101178.1, 101105.2, 101137.6, 101216.4, 87258.29, 78257.5,
  91309.46, 88053.97, 88481.77, 90266.4, 89898.98, 88854.82, 89414.32, 
    91185.12, 95454.79, 101190.9, 101131.1, 101264.6, 101198.9, 86050.08, 
    88197.7,
  94263.83, 89949.8, 89023.85, 90110.45, 89307.04, 86943.07, 88169.38, 
    90735.99, 100799.6, 101249.4, 101181.2, 101310.3, 101255.3, 93600.85, 
    96591.63,
  97427.63, 92784.83, 91168.92, 93562.81, 93797.79, 93896.83, 94819.32, 
    100802, 101355.7, 101285.7, 101271.3, 101365.9, 101404.2, 99318.65, 
    100830.6,
  101570, 101199.8, 97271.48, 94690.8, 94616.77, 93529.51, 91147.44, 91586.2, 
    85887.53, 81291.56, 79042.65, 79345.56, 82444.2, 81124.8, 91630.62,
  101461.4, 101307.3, 99044.1, 93928.41, 91128.16, 89188.44, 87891.51, 
    88160.05, 83321.89, 80611.8, 79854.31, 80535.84, 82868.12, 81874.04, 
    93034.08,
  92503.89, 88872.66, 93739.88, 92362.23, 85908.78, 84780.46, 86998.12, 
    86258.73, 81425.16, 79244.77, 78404.13, 79089.8, 80567.14, 82207.35, 
    95093.72,
  86476.14, 86527.95, 85612.11, 83858.97, 83588.96, 82100.92, 82925.86, 
    83185.02, 80876.11, 79621.47, 79300.8, 80824.58, 80579.05, 82683.01, 
    88986.63,
  88087.6, 87012.27, 88043.49, 87186.23, 87018.76, 85387.62, 84328.65, 
    83847.2, 82829.45, 84881.44, 100013.8, 100589, 90622.27, 91156.36, 
    83906.88,
  88376.65, 86554.7, 88975.73, 89801.27, 88884.55, 88412.28, 87667.78, 
    88018.8, 89658.87, 100739.1, 101524, 101493.7, 101263.6, 93263.65, 
    78285.92,
  87545.38, 86778.02, 88860.83, 90106.88, 89853.84, 89847.42, 89755.24, 
    91718.01, 95786.86, 101440.7, 101345.9, 101361.8, 101275.6, 87153.48, 
    78020.81,
  91299.89, 88028.22, 88466.7, 90268.22, 89928.91, 88889.95, 89484.4, 
    91281.75, 95618.3, 101438.9, 101352.2, 101388.7, 101303.1, 85908.01, 
    87854.62,
  94256.85, 89936.46, 89014.22, 90117.37, 89312.38, 86934.51, 88199.36, 
    90775.05, 101058.8, 101450.2, 101318.4, 101261.9, 101324.1, 93506.74, 
    96208.12,
  97442.93, 92794.51, 91188.54, 93591.82, 93843.8, 93993.07, 94915.42, 
    100981.8, 101533.1, 101440.2, 101334, 101260.1, 101322.4, 99057.75, 
    100369.6,
  101325.3, 100973.5, 97065.91, 94537.23, 94480.05, 93444.51, 91074.14, 
    91571.76, 85785.4, 81167.8, 78884.01, 79155.17, 82087.7, 80702.43, 
    91068.58,
  101278.1, 101188.7, 98944.51, 93799.24, 91003.78, 89108.09, 87852.52, 
    88147.27, 83203.41, 80494.04, 79708.3, 80395.86, 82630.65, 81513.03, 
    92483.16,
  92291.41, 88721.12, 93618.13, 92248.18, 85791.03, 84722.16, 86983.87, 
    86251.34, 81351.98, 79144.03, 78231.38, 78915.47, 80284.75, 81869.42, 
    94591.3,
  86234.05, 86355.13, 85446.23, 83741.23, 83472.6, 82012.78, 82855.95, 
    83143.95, 80841.98, 79521.49, 79238.38, 80782.89, 80420, 82413.88, 
    88518.18,
  87799.7, 86838.8, 87873.61, 87066.56, 86919.88, 85304.11, 84246.2, 
    83753.02, 82767.92, 84825.29, 100141.6, 100650.9, 90706.39, 91013.48, 
    83572.45,
  88187.84, 86403.57, 88855.53, 89685.3, 88771.52, 88309.66, 87581.37, 
    87969.48, 89606.29, 100839.8, 101611.6, 101595, 101398.9, 93226.95, 
    78009.31,
  87399.46, 86642.06, 88743.42, 90014.6, 89771.54, 89790.53, 89689.59, 
    91735.11, 95823.05, 101598.8, 101496.6, 101533.6, 101414.9, 87054.13, 
    77773.02,
  91198.03, 87931.54, 88386.48, 90224.06, 89868.83, 88841.12, 89438.71, 
    91284.41, 95678.88, 101616.1, 101542.5, 101563, 101433.7, 85829.2, 
    87774.32,
  94217.55, 89898.11, 88977.42, 90090.3, 89253.47, 86866.26, 88154.69, 
    90801.13, 101136.1, 101591.2, 101528.3, 101495.2, 101449.1, 93509.59, 
    96196.32,
  97448.66, 92813.17, 91226.19, 93649.68, 93897.18, 94064.91, 94990.55, 
    101048.4, 101648.1, 101596.1, 101556.6, 101477.3, 101424.9, 99081.76, 
    100273,
  100993.9, 100635.5, 96758.16, 94283.3, 94241.07, 93221.19, 90941.62, 
    91441.3, 85748.34, 81158.34, 78907.91, 79218.98, 82161.2, 80761.55, 
    91054.66,
  100932.5, 100925.3, 98663.91, 93529.26, 90770.49, 88926.51, 87688.19, 
    88015.94, 83195.94, 80498.92, 79731.73, 80433.48, 82659.38, 81558.27, 
    92448.41,
  91983.57, 88481.66, 93400.42, 92074.31, 85626.03, 84571.55, 86851.71, 
    86149.65, 81278.7, 79110.55, 78248.66, 78963.63, 80319.02, 81911.84, 
    94550.22,
  85955.03, 86090.41, 85214.75, 83528.51, 83290.39, 81832.58, 82700.28, 
    83019.29, 80746.02, 79520.63, 79193.23, 80748.64, 80418.89, 82433.62, 
    88490.52,
  87554.34, 86624.48, 87677.65, 86845.15, 86726.23, 85138.08, 84095.91, 
    83612.41, 82648.41, 84655.38, 99819.12, 100407.4, 90528.25, 90947.99, 
    83533.07,
  87976.84, 86201.7, 88688.73, 89534.73, 88619.7, 88168.16, 87453.85, 
    87844.84, 89453.09, 100675, 101541.7, 101459.6, 101225.6, 93103.12, 
    78047.74,
  87205.67, 86453.59, 88598.07, 89877.63, 89637.15, 89668.37, 89565.21, 
    91588.56, 95674.37, 101461.6, 101341.1, 101383.1, 101264.5, 86996.13, 
    77834.13,
  91024.88, 87774.45, 88284.66, 90102.27, 89779.06, 88737.68, 89352.93, 
    91179.09, 95543.74, 101513.4, 101460.7, 101505, 101292.9, 85785.87, 
    87858.55,
  94079.27, 89755.95, 88904.87, 90006.53, 89172.01, 86764.37, 88059.93, 
    90702.5, 101051.2, 101535.7, 101492.9, 101497.5, 101427.5, 93453.14, 
    96242.07,
  97345.38, 92702.09, 91174.86, 93588.16, 93824.21, 94008.62, 94919.73, 
    100983.7, 101580.5, 101556.7, 101550.4, 101530, 101515.3, 99155.95, 
    100332.8,
  101296.9, 100949.3, 97043.45, 94444.54, 94362.88, 93270.05, 90934.91, 
    91372.72, 85665.73, 81092.66, 78867.41, 79196.02, 82127.45, 80849.23, 
    90991.97,
  101317.3, 101182.9, 98930.32, 93757.34, 90962.83, 89055.93, 87794.56, 
    88057.87, 83180.09, 80484.7, 79713.67, 80431.87, 82643.29, 81633.41, 
    92369.47,
  92250.12, 88846.48, 93698.97, 92269.22, 85843.62, 84759.78, 86997.53, 
    86237.76, 81360.19, 79183.61, 78309.52, 79019.88, 80386.75, 81971.92, 
    94455.97,
  86325.24, 86563.02, 85595.79, 83903.53, 83621.39, 82120.14, 82936.73, 
    83223.98, 80922.76, 79640.69, 79383.59, 80908.14, 80534.44, 82525.65, 
    88521.7,
  87924.73, 87050.73, 88105.38, 87294.52, 87129.28, 85499.55, 84414.81, 
    83907.63, 82905.66, 85058.27, 100399.7, 100895.1, 90879.52, 91113.12, 
    83663.59,
  88368.85, 86593.52, 89136.47, 89956.74, 89044.64, 88600.7, 87838.35, 
    88295.6, 89944.16, 101177.8, 101943.3, 101886.7, 101633.9, 93370.53, 
    78163.6,
  87587.75, 86858.62, 89043.33, 90316.3, 90101.13, 90096.45, 90037.12, 
    92079.02, 96147.86, 101929.9, 101828.8, 101811, 101643.4, 87212.02, 
    77926.63,
  91357.34, 88161.12, 88705.41, 90535.86, 90228.32, 89201.4, 89835.69, 
    91650.69, 96028.04, 101954.1, 101888.8, 101870.2, 101668.5, 86020.58, 
    87980.88,
  94380.34, 90141.96, 89305.07, 90436.66, 89587.62, 87198.02, 88497.52, 
    91217.32, 101508.5, 101954, 101882, 101831.2, 101709.1, 93679.41, 96416.71,
  97586.99, 93011.69, 91550.19, 94000.63, 94292.55, 94496.43, 95462.11, 
    101460.9, 101987.3, 101956.4, 101921.5, 101859.3, 101765.4, 99393.52, 
    100479.7,
  101549.5, 101277.1, 97368.08, 94909.27, 94873.98, 93786.53, 91376.22, 
    91860.57, 85944, 81355.22, 79074.71, 79396.52, 82302.42, 80871.3, 91129.82,
  101653.9, 101581, 99302.77, 94204.29, 91418.64, 89527.18, 88311.45, 
    88528.74, 83526.66, 80835.52, 79999.52, 80713.63, 82867.09, 81746.34, 
    92688.06,
  92560.86, 89210.25, 94101.19, 92680.89, 86264.76, 85206.71, 87465.16, 
    86655.6, 81754.21, 79540.69, 78567.06, 79286.59, 80597.73, 82200.16, 
    94777.15,
  86660.09, 86858.95, 85941.12, 84288.04, 84028.74, 82519.02, 83381.73, 
    83668.44, 81302.25, 79965.7, 79762.02, 81323.08, 80789.2, 82897.51, 
    88785.99,
  88226.52, 87336.86, 88427.41, 87636.12, 87509.16, 85908.64, 84853.48, 
    84339.87, 83304.81, 85553.12, 100957.2, 101426, 91362.23, 91686.33, 
    83764.09,
  88616.77, 86870.94, 89439.69, 90276.02, 89421.92, 88999.35, 88302.95, 
    88713.14, 90401.39, 101589.4, 102432.4, 102412.6, 102307.6, 93773.04, 
    78407.78,
  87796.34, 87093.49, 89320.99, 90614.73, 90454.39, 90506.94, 90495.98, 
    92492.59, 96585.06, 102393.1, 102394.1, 102332.9, 102337.9, 87511.32, 
    78251.8,
  91463.73, 88337.26, 88918.01, 90795.67, 90532.27, 89544.81, 90212.53, 
    92020.34, 96492.43, 102377.8, 102361.3, 102404.8, 102251.2, 86450.48, 
    88606.35,
  94424.19, 90288.95, 89488.97, 90669.8, 89872.06, 87536.95, 88857.87, 
    91651.72, 101919.4, 102395, 102337.1, 102367.3, 102301.2, 94264, 96997.53,
  97563.16, 93098.09, 91655.8, 94157.87, 94460.41, 94697.49, 95768.77, 
    101822.7, 102376.4, 102392.1, 102315.2, 102312.7, 102288.8, 99968.19, 
    101100.2,
  100896.3, 100741.3, 97010.98, 94670.52, 94673.82, 93636.37, 91300.9, 
    91854.76, 85983.14, 81444.92, 79208.37, 79568.85, 82606.91, 81119.28, 
    91565.8,
  100922, 101047, 98788.28, 93860.02, 91190.93, 89372.54, 88180.91, 88477.61, 
    83538.27, 80901.33, 80100.43, 80860.58, 83092.98, 81947.37, 93100.29,
  92113.96, 88831.75, 93752.5, 92375.77, 86017.49, 85033.49, 87317.09, 
    86576.55, 81719.53, 79555.34, 78612.64, 79405.96, 80763.69, 82429.06, 
    95185.7,
  86140.28, 86325.99, 85495.1, 83916.9, 83723.57, 82295.68, 83207.84, 
    83531.24, 81238.63, 79962.33, 79717.6, 81347.52, 80889.23, 83024.22, 
    89009.87,
  87736.31, 86849.46, 87949.76, 87180.54, 87116.65, 85567.39, 84597.45, 
    84144.48, 83171.98, 85420.46, 100764.6, 101213.8, 91316.91, 91752.51, 
    83991.38,
  88129.59, 86358.45, 88948.75, 89790.27, 89000.86, 88629.88, 88006.87, 
    88435.78, 90191.91, 101403.4, 102311.7, 102307.3, 102272.1, 93730.7, 
    78616.52,
  87327.49, 86591.75, 88864.86, 90121.55, 90033.37, 90115.35, 90178.01, 
    92231.12, 96406.56, 102203.1, 102238.3, 102213.8, 102315.3, 87552.05, 
    78450.28,
  90921.48, 87795.08, 88444.07, 90291.45, 90065.63, 89150.78, 89870.21, 
    91758.23, 96238.55, 102212.6, 102236.3, 102346.4, 102111.9, 86526.83, 
    88717.73,
  93863.3, 89726.66, 88991.62, 90155.38, 89447.41, 87207.84, 88547.58, 
    91297.3, 101588.1, 102227.7, 102217.2, 102332.2, 102165.1, 94318.38, 
    97009.48,
  97032.34, 92534.2, 91126.19, 93581.45, 93876.99, 94044.89, 95128.9, 
    101258.4, 102109.7, 102219.8, 102235.6, 102302.6, 102262.8, 99980.38, 
    101120.4,
  100511.7, 100133.7, 96324.83, 94001.75, 94013.42, 93099.01, 90890.23, 
    91439.02, 85729.65, 81178.69, 78958.04, 79362.7, 82427.31, 81043.79, 
    91465.39,
  100294.9, 100398, 98136.71, 93189.2, 90629.73, 88888.3, 87701.29, 88093.27, 
    83228.45, 80584.19, 79814.98, 80563.11, 82888.11, 81818.48, 92853.81,
  91550.94, 88343.74, 93165.85, 91845.3, 85537.52, 84550.21, 86838.34, 
    86186.17, 81325.75, 79192.36, 78314.66, 79067.69, 80535.22, 82147.16, 
    94875,
  85563.48, 85779.17, 84917.09, 83426.76, 83194.48, 81806.5, 82722.87, 
    83078.11, 80810.27, 79621.61, 79282.45, 80853.2, 80585.03, 82670.7, 
    88866.27,
  87218.52, 86373.02, 87409.22, 86646.78, 86539.52, 85017.04, 84058.5, 
    83639.34, 82680.66, 84712.14, 99766.47, 100305.6, 90559.04, 91128.16, 
    83846.3,
  87601.82, 85884.55, 88394.45, 89274.38, 88410.58, 88017.53, 87342.08, 
    87765.03, 89438.9, 100554, 101386.8, 101267, 101099.1, 93241.72, 78325.38,
  86784.33, 86125.55, 88326.44, 89605.62, 89405.35, 89486.15, 89478.25, 
    91526.41, 95633.47, 101306.4, 101240.9, 101265.9, 101250.9, 87157.38, 
    78093.57,
  90520.8, 87355.45, 87914.45, 89763.65, 89455.98, 88525.33, 89186.72, 
    91085.07, 95480.12, 101355.1, 101343.9, 101405.4, 101272.8, 85985.29, 
    88109.09,
  93531.16, 89287.23, 88493.95, 89637.99, 88858.2, 86615.02, 87915.55, 
    90610.42, 100783.8, 101390, 101337.7, 101395.4, 101307.1, 93620.45, 
    96470.12,
  96729.09, 92101.28, 90643.21, 93061.91, 93256.97, 93392.8, 94408.86, 
    100484.5, 101335.5, 101402.7, 101415.3, 101471.5, 101468.8, 99315.89, 
    100584.5,
  100506.6, 100194.4, 96324.99, 93798.27, 93738.23, 92707.41, 90395.79, 
    90859.05, 85214.57, 80680.23, 78469.84, 78821.95, 81839.75, 80547.17, 
    90921.75,
  100371.5, 100353.9, 98052.73, 92979.48, 90246.3, 88397.75, 87138.58, 
    87502.15, 82685.95, 80047.97, 79296.2, 80008.58, 82290.98, 81318.62, 
    92283.09,
  91429.5, 87986.23, 92901.88, 91525.41, 85079.1, 84060.19, 86300.27, 
    85602.58, 80791.61, 78658.06, 77824.48, 78552.46, 79990.65, 81620.05, 
    94316.94,
  85413.19, 85577.27, 84621.99, 83036.17, 82784.65, 81347.59, 82213.77, 
    82523.06, 80275.26, 79079.52, 78751.23, 80271.66, 80044.11, 82080.78, 
    88311.16,
  86988.36, 86138.43, 87090.29, 86259.28, 86109.3, 84547.48, 83547.23, 
    83083.68, 82152.45, 84183.03, 99117.81, 99662.27, 89962.16, 90478.13, 
    83340.12,
  87384.84, 85638.55, 88026.58, 88854.19, 87955.61, 87515.09, 86830.09, 
    87260.84, 88892.39, 99833.87, 100613.8, 100571.8, 100473, 92588.4, 
    77802.88,
  86686.38, 85873, 87960.66, 89162.24, 88950, 88984.91, 88974.17, 90995.32, 
    94956.29, 100563.5, 100467.7, 100527.2, 100493.8, 86543.37, 77576.87,
  90523.35, 87158.17, 87652.4, 89387.52, 89049.65, 88089.59, 88739.63, 
    90553.95, 94837.58, 100593.6, 100536.3, 100633.3, 100553, 85403.84, 
    87438.51,
  93543.42, 89133.16, 88294.62, 89335.91, 88497.71, 86209.77, 87487.34, 
    90152.28, 100172.5, 100619.6, 100569.2, 100629, 100602, 92893.55, 95745.76,
  96765.12, 92037.98, 90521.91, 92899.71, 93101.72, 93209.38, 94153.23, 
    100114.6, 100700.8, 100683.7, 100668.1, 100677.9, 100691.1, 98540.06, 
    99852.09,
  100784.8, 100488.9, 96598.57, 94105.77, 94068.57, 93058.58, 90759.28, 
    91255.45, 85501.96, 80916.49, 78649.29, 78979.92, 81889.64, 80580.59, 
    90616.09,
  100697.3, 100713.8, 98431.05, 93302.05, 90553.02, 88700.38, 87447.17, 
    87796.49, 82961.87, 80270.02, 79487.78, 80177.55, 82354.36, 81353.78, 
    91923.11,
  91613.3, 88225.09, 93161.41, 91834.81, 85326.16, 84288.65, 86540.27, 
    85836.41, 80993.86, 78822.41, 77969.5, 78675.06, 80036.26, 81611.96, 
    93930.66,
  85717.97, 85887.34, 84856.32, 83213.19, 82985.17, 81512.12, 82376.61, 
    82725.12, 80486.86, 79236.05, 78901.23, 80420.25, 80117.66, 82090.05, 
    88096.81,
  87313.89, 86405.68, 87374.66, 86494.21, 86355.39, 84752.48, 83718.94, 
    83210.65, 82229.55, 84304.31, 99226.6, 99798.07, 90104.73, 90412.76, 
    83240.4,
  87723.54, 85910.13, 88359.12, 89101.07, 88196.04, 87798.74, 87120.89, 
    87529.62, 89159.66, 100116.9, 100882.6, 100824.4, 100563.4, 92636.43, 
    77792.3,
  87003.86, 86218.65, 88329.69, 89516.2, 89287.34, 89289.11, 89223.06, 
    91184.08, 95152.3, 100735.2, 100636.7, 100643.5, 100525.1, 86602.37, 
    77551.96,
  90789.16, 87533.72, 88014.31, 89754.05, 89398.84, 88398.2, 89034.8, 
    90806.57, 95069.03, 100790.3, 100714.8, 100738.7, 100622.7, 85439.02, 
    87310.34,
  93821.52, 89518.73, 88667.43, 89749.1, 88887.38, 86520.93, 87762.04, 
    90419.16, 100424, 100778.1, 100653.9, 100628.7, 100589.4, 92892.59, 
    95721.45,
  97023.7, 92419.36, 90902.28, 93285.05, 93530.25, 93677.63, 94611.99, 
    100468.3, 100935.4, 100835.9, 100743.6, 100686.4, 100673.6, 98507.23, 
    99821.36,
  101337, 101048.1, 97109.52, 94582.99, 94542.04, 93474.57, 91115.16, 
    91634.88, 85830.5, 81272.52, 78983.84, 79285.05, 82201.08, 80806.27, 
    90847.88,
  101274.7, 101219.2, 98985.22, 93836.85, 91044.19, 89163.42, 87908.5, 
    88211.47, 83304, 80628.83, 79827.09, 80542.73, 82715.4, 81652.99, 92219.72,
  92165.08, 88792.31, 93649.66, 92343.24, 85823.81, 84759.41, 86993.27, 
    86308.33, 81437.27, 79234.54, 78321.91, 79050.89, 80394.62, 81944.04, 
    94222.48,
  86280.6, 86463.41, 85448.47, 83785.61, 83532.89, 82054.35, 82866.32, 
    83187.23, 80909.67, 79656.58, 79342.52, 80869.38, 80505.18, 82488.13, 
    88358.66,
  87857.02, 86903.23, 87941.45, 87121.84, 86953.03, 85344.74, 84300.96, 
    83791.02, 82772.71, 84844.93, 99963.46, 100517.9, 90660.03, 91023.32, 
    83557.98,
  88243.31, 86413.05, 88867.93, 89687.39, 88803.2, 88364.99, 87646, 88055.7, 
    89690.34, 100766.7, 101545.7, 101550, 101323.7, 93157.91, 78146.38,
  87408.96, 86651.29, 88748.73, 89999.81, 89798.16, 89815.17, 89753.91, 
    91722.38, 95722.05, 101426.3, 101342, 101382.1, 101283, 87107.88, 77924.25,
  91072.07, 87889.61, 88397.16, 90182.89, 89862.9, 88878.27, 89490.25, 
    91302.3, 95609.73, 101424.9, 101354.7, 101424.9, 101303.4, 85950.97, 
    87799.63,
  94000.99, 89812.21, 88949.66, 90067.27, 89267.41, 86915.92, 88173.66, 
    90827.23, 100950.8, 101378.2, 101267, 101277.6, 101260.9, 93468.41, 
    96100.85,
  97114.59, 92593.09, 91112.59, 93497.73, 93765.3, 93963.45, 94919.23, 
    100903.5, 101420.5, 101348.7, 101290.8, 101244, 101247.3, 99009.42, 
    100131.3,
  101557.8, 101249.5, 97290.09, 94800.35, 94718.08, 93653.93, 91289.83, 
    91840.34, 85998.41, 81452.91, 79144.3, 79428.38, 82346.43, 80894.46, 
    91046.23,
  101500.6, 101470.6, 99266.45, 94108.26, 91270.98, 89393.22, 88155.11, 
    88431.88, 83505.72, 80848.55, 80033.77, 80721.21, 82899.18, 81778.98, 
    92466.4,
  92520.8, 89054.23, 93917.08, 92526.97, 86143.39, 85074.32, 87285.09, 
    86526.16, 81699.6, 79476.96, 78544.87, 79237.05, 80586.7, 82148.42, 
    94476.22,
  86570.37, 86676.21, 85781.27, 84144.39, 83882.82, 82388.55, 83202.64, 
    83499.23, 81204.75, 79862, 79616.3, 81123.27, 80682.45, 82707.57, 88550.59,
  88162.96, 87101.93, 88136.69, 87332.96, 87193.42, 85625.67, 84579.43, 
    84076.38, 83066.17, 85167.68, 100119.2, 100685.7, 90908.02, 91259.85, 
    83772.6,
  88437.45, 86613.66, 89036.77, 89865.36, 89000.73, 88574.84, 87866.49, 
    88267.27, 89822.59, 100737.9, 101647.3, 101685.6, 101500.8, 93381.02, 
    78323.67,
  87476.36, 86772.28, 88864.51, 90110.77, 89928.97, 89953.73, 89907.23, 
    91836.3, 95745.88, 101541.9, 101550.5, 101609.6, 101559.3, 87295.45, 
    78123.65,
  91017.16, 87944.93, 88430.84, 90238.03, 89942.98, 88973.23, 89603.98, 
    91387.48, 95617.78, 101521.5, 101528.4, 101657.8, 101565.7, 86135.55, 
    88026.33,
  93876.27, 89787.65, 88945.92, 90055.8, 89299.29, 87019.91, 88276.77, 
    90834.44, 100880.7, 101519.8, 101519.5, 101599.9, 101563.9, 93749.1, 
    96340.95,
  96944.07, 92505.07, 91007.16, 93388.01, 93659.54, 93835.37, 94776.14, 
    100750.7, 101453.4, 101508.4, 101520.9, 101562.2, 101573.5, 99317.52, 
    100418.4,
  101232.8, 100952.8, 97135.64, 94711.78, 94659.96, 93640.59, 91296.61, 
    91821.27, 86013.91, 81509.41, 79250.02, 79556.76, 82468.15, 81028.71, 
    91198.62,
  101121.9, 101194.5, 98975.52, 93951.25, 91210.82, 89392.88, 88165.13, 
    88456.61, 83583.38, 80939.04, 80129.02, 80806.62, 82967.22, 81867.2, 
    92540.9,
  92427.24, 88988.22, 93811.3, 92502.83, 86146.66, 85097.47, 87312.14, 
    86582.91, 81772.05, 79573.16, 78627.65, 79331.19, 80677.48, 82227.91, 
    94558.52,
  86443.61, 86467.17, 85710.62, 84081.79, 83842.32, 82391.46, 83224.27, 
    83517.32, 81252.63, 79977.72, 79697.78, 81208.1, 80744.22, 82751.15, 
    88620.52,
  87964.13, 86891.99, 88008.45, 87216.92, 87116.79, 85573.83, 84571.72, 
    84088.62, 83121.64, 85132.91, 99821.4, 100401.6, 90824.21, 91216.74, 
    83832.59,
  88159.12, 86391.86, 88833.03, 89711.02, 88879.98, 88483.33, 87794.23, 
    88197.26, 89739.04, 100449.7, 101351.3, 101344.9, 101161.3, 93258.44, 
    78409.31,
  87239.87, 86553.89, 88655.31, 89951.77, 89794.05, 89864.65, 89805.55, 
    91741.65, 95581.45, 101211.7, 101249.5, 101297.9, 101277.7, 87270.77, 
    78200.59,
  90783.45, 87708.93, 88192.83, 90046.27, 89793.73, 88852.91, 89467.29, 
    91270.95, 95385.34, 101186.7, 101241.1, 101346.1, 101278.9, 86058.04, 
    88020.27,
  93648.33, 89541.16, 88706.34, 89873.01, 89164.27, 86901.97, 88169.79, 
    90683.95, 100565.3, 101194.6, 101232.3, 101342, 101337, 93593.71, 96233.76,
  96660.11, 92244.58, 90736.85, 93172.02, 93483.91, 93634.45, 94573.03, 
    100425.8, 101107.9, 101192.3, 101248.3, 101348.2, 101366.4, 99120.99, 
    100302.5,
  100427.2, 100147, 96523.48, 94271.72, 94304.04, 93335.23, 91061.23, 
    91588.52, 85879.94, 81407.38, 79173.98, 79467.45, 82404.62, 81011.26, 
    91091.46,
  100308.1, 100426.3, 98249.05, 93410.33, 90854.01, 89095.02, 87907.02, 
    88244.04, 83452.29, 80824.65, 80055.17, 80716.66, 82869.26, 81799.06, 
    92362.51,
  91828.9, 88441.81, 93259.3, 92008.64, 85795.05, 84801.11, 87040.84, 
    86383.18, 81620.73, 79444.92, 78562.59, 79257.46, 80613.88, 82159.07, 
    94369.28,
  85847.24, 85869.66, 85183.66, 83628.95, 83429.7, 82067.47, 82947.36, 
    83286.41, 81073.35, 79867.14, 79554.3, 81047.2, 80682.5, 82620.52, 
    88508.75,
  87350.53, 86325.21, 87456.08, 86660.91, 86641.72, 85153.05, 84222.55, 
    83799.31, 82897.72, 84853.72, 99404.09, 100039.3, 90561.35, 90922.93, 
    83749.23,
  87622.3, 85823.22, 88287.81, 89161.38, 88372.41, 87997.82, 87369.79, 
    87807.17, 89380.69, 99993.74, 100893.7, 100875.8, 100712.1, 92979.14, 
    78364.53,
  86770.21, 86082.99, 88153.91, 89416.34, 89260.22, 89360.78, 89350.73, 
    91322.62, 95196.86, 100790.8, 100779.2, 100843.7, 100780.3, 87107.23, 
    78104.29,
  90443.98, 87311.86, 87783.77, 89579.43, 89287.15, 88360.88, 88996.96, 
    90872.21, 95019.48, 100767.2, 100763.5, 100875.3, 100775.7, 85907.83, 
    87757.36,
  93417.78, 89218.91, 88363.49, 89468.49, 88713.51, 86470.98, 87741.92, 
    90268.77, 100204.6, 100767.1, 100737.9, 100828.5, 100827.5, 93261.85, 
    95837.81,
  96537.74, 92004.35, 90438.63, 92851.98, 93114.66, 93222.68, 94178.8, 
    100070.4, 100748.8, 100702.8, 100718.2, 100766.3, 100826.6, 98650.43, 
    99827.82,
  100639.8, 100268.4, 96404.78, 93943.96, 93839.34, 92831.43, 90583.94, 
    91089.83, 85561.26, 81136.62, 78949.24, 79266.16, 82174.26, 80835.33, 
    90864.92,
  100362.3, 100376.6, 98177.19, 93105.22, 90436.38, 88639.84, 87392.95, 
    87769.34, 83092.85, 80520.29, 79785.27, 80476.94, 82649.6, 81621.38, 
    92114.64,
  91685.81, 88065.73, 92926.5, 91662.93, 85330.8, 84278.53, 86521.38, 
    85903.43, 81188.93, 79089.95, 78266.73, 78993.8, 80352.97, 81922.21, 
    94073.37,
  85552.88, 85466.69, 84701.37, 83157.66, 82895.86, 81535.59, 82439.56, 
    82783.2, 80624.95, 79508.59, 79180.21, 80712.31, 80450.85, 82392.4, 
    88313.55,
  87065.71, 86002.88, 87017.31, 86173.34, 86103.62, 84591.21, 83636.04, 
    83254.55, 82420.38, 84297.24, 98800.52, 99432.49, 90088.85, 90529.14, 
    83533.39,
  87199.41, 85456.95, 87818.21, 88698.89, 87867.87, 87460.71, 86824.53, 
    87244.38, 88816.59, 99431.8, 100336.4, 100328.6, 100200.9, 92596.2, 
    78158.34,
  86412.11, 85644.18, 87666.57, 88918.19, 88717.88, 88794.9, 88777.73, 
    90744.32, 94652.05, 100119.1, 100152.9, 100234, 100197, 86734.34, 77907.01,
  90091.49, 86841.2, 87253.6, 89029.16, 88711.53, 87770.5, 88399.76, 
    90279.09, 94418.7, 100125.9, 100181.7, 100273.1, 100211.8, 85569.08, 
    87445.62,
  93065.62, 88712.48, 87774.27, 88826.29, 88037.43, 85793.64, 87100.69, 
    89637.11, 99444.2, 100103, 100123, 100228.9, 100251.3, 92794.61, 95466.26,
  96189.84, 91553.27, 89921.53, 92224.75, 92397.91, 92439.05, 93365.78, 
    99167.51, 99948.22, 100011.4, 100114, 100233.6, 100295, 98167.5, 99361.59,
  100983.9, 100656, 96739.69, 94203.13, 94107.07, 92988.98, 90689.84, 
    91190.06, 85614.18, 81117.53, 78924.02, 79248.71, 82174.96, 80772.01, 
    90840.02,
  100854.7, 100849.9, 98580.98, 93448.15, 90644.08, 88776.45, 87469.18, 
    87792.34, 83079.38, 80476.09, 79761.36, 80453.78, 82667.06, 81605.42, 
    92109.96,
  91928.48, 88392.36, 93308.14, 91966.8, 85510.2, 84405.61, 86621.6, 
    85944.59, 81132.59, 79008.36, 78218.02, 78950.42, 80344.23, 81887.71, 
    94018.32,
  85803.33, 85926.45, 85026.46, 83390.17, 83127.21, 81671.37, 82510.12, 
    82835.22, 80577.76, 79454.7, 79112.3, 80634.61, 80417.61, 82353.14, 
    88249.38,
  87415.09, 86439.24, 87433.52, 86628.77, 86475.26, 84890.52, 83853.2, 
    83366.78, 82460.41, 84354.39, 99000.77, 99634.49, 90130.56, 90480.96, 
    83502.52,
  87672.19, 85885.73, 88287.45, 89127.43, 88254.29, 87825.68, 87115.79, 
    87495.13, 89031.48, 99793.39, 100731, 100648.1, 100389.1, 92646.21, 
    78095.6,
  86849.47, 86115.68, 88167.56, 89411.26, 89176.98, 89188.37, 89112.4, 
    91051.55, 94934.5, 100507.7, 100465.1, 100524.3, 100338.6, 86737.78, 
    77790.72,
  90544.53, 87330.71, 87758.38, 89539.3, 89200.12, 88194.56, 88775.87, 
    90589.81, 94714.21, 100451.2, 100486.3, 100593.8, 100438.9, 85599.3, 
    87344.91,
  93507.95, 89225.11, 88300.34, 89359.72, 88540.75, 86191.74, 87428.98, 
    89963.53, 99861.3, 100427.9, 100420.8, 100469.8, 100477.7, 92827.55, 
    95469.33,
  96624.48, 92032.17, 90421.2, 92723.43, 92937.62, 93057.75, 93931.69, 
    99762.95, 100391.9, 100396.7, 100432.5, 100427.2, 100479.6, 98252.77, 
    99356.27,
  100974.6, 100628.2, 96681.58, 94134.74, 93993.88, 92859.5, 90450.17, 
    91000.46, 85247.38, 80747.38, 78494.67, 78777.66, 81744.26, 80354.17, 
    90539.91,
  100876.8, 100808.9, 98550.29, 93422.62, 90558.94, 88625.46, 87294.41, 
    87627.09, 82782.23, 80140.35, 79339.05, 80033.2, 82235.43, 81188.91, 
    91849.24,
  91932.78, 88383.32, 93266.33, 91873.62, 85425.05, 84343.8, 86507.45, 
    85771.92, 80943.49, 78740.59, 77842.37, 78557.02, 79923.31, 81531.98, 
    93743.68,
  85890.93, 86025.09, 85088.91, 83427.16, 83165.33, 81672.3, 82485.7, 
    82765.5, 80458.82, 79265.52, 78963.93, 80388.86, 80069.38, 82040.81, 
    88009.16,
  87506.84, 86546.79, 87521.55, 86695.56, 86543.85, 84947.07, 83892.54, 
    83379.52, 82405.07, 84462.31, 99196.94, 99761.61, 90019.11, 90307.37, 
    83224.82,
  87792.49, 86007.78, 88412.21, 89231.84, 88345.64, 87910.41, 87191.15, 
    87562.23, 89124.06, 99874.98, 100634.4, 100623.4, 100518.7, 92488.71, 
    77913.41,
  86985.23, 86236.98, 88292, 89522.76, 89302.34, 89320.53, 89248.35, 
    91171.85, 95063.3, 100620.3, 100555, 100559.3, 100465.2, 86559.98, 
    77644.98,
  90662.15, 87462.01, 87910.37, 89683, 89340.7, 88352.84, 88950.28, 90737.04, 
    94906.69, 100614, 100589.1, 100644, 100554.9, 85491.21, 87383.15,
  93573.86, 89346.58, 88442.92, 89517.05, 88721.16, 86405.95, 87660.52, 
    90192.45, 100149.5, 100601.8, 100574.1, 100588.9, 100531.3, 92846.54, 
    95559.74,
  96691.36, 92108.8, 90540.73, 92888.73, 93132.67, 93258.2, 94168.55, 
    100010.7, 100632.9, 100611.1, 100613.5, 100622.8, 100604.5, 98427.48, 
    99537.24,
  101059.8, 100706.6, 96777.1, 94218.01, 94131.19, 93037.16, 90643.56, 
    91142.86, 85392.57, 80794.32, 78485.51, 78758.69, 81629.41, 80150.35, 
    90172.27,
  100867.8, 100823.2, 98553.28, 93437.12, 90632.69, 88721.12, 87426.59, 
    87727.16, 82852.42, 80189.15, 79378.53, 80050.42, 82186.71, 81072.62, 
    91658.72,
  92011.68, 88361.11, 93304.68, 91946.86, 85471.85, 84408.43, 86583.94, 
    85842.59, 81007.57, 78817.09, 77828.7, 78495.05, 79794.48, 81354.26, 
    93637.93,
  85912.52, 85905.16, 85040.62, 83385.49, 83139.01, 81671.27, 82502.67, 
    82785.66, 80495.69, 79205.52, 78950.78, 80498.17, 79959.01, 81944.23, 
    87802.28,
  87475.52, 86457.52, 87486.09, 86629.01, 86500.92, 84905.2, 83875.02, 
    83384.71, 82381.9, 84460.82, 99230.54, 99757.02, 90078.67, 90378.45, 
    82944.45,
  87715.05, 85935.65, 88358.38, 89171.69, 88298.32, 87854.71, 87153.03, 
    87517.38, 89099.4, 99935.51, 100657.7, 100674.3, 100535.5, 92425.47, 
    77644.05,
  86934.78, 86176.09, 88256.56, 89482.04, 89262.57, 89295.54, 89227.55, 
    91169.05, 95103.91, 100662.7, 100582.1, 100595.9, 100495.7, 86398.72, 
    77431.85,
  90639.19, 87423.62, 87869.66, 89631.74, 89300.03, 88296.15, 88939.45, 
    90731.65, 94957.53, 100673, 100609.5, 100647.6, 100503.1, 85222.03, 
    87165.38,
  93610.77, 89346.04, 88453.35, 89519.16, 88728.94, 86431.78, 87706.51, 
    90261.83, 100251.8, 100699, 100633.4, 100622.8, 100544.2, 92729.55, 
    95405.95,
  96759.05, 92129.32, 90573.95, 92945.7, 93168.12, 93265.73, 94272.94, 
    100170.7, 100727, 100719.1, 100696.2, 100658.8, 100645.8, 98353.05, 
    99397.73,
  101105.2, 100748, 96860.88, 94319.1, 94260.98, 93233.98, 90905.3, 91361.52, 
    85631.34, 81021.5, 78736.17, 79006.97, 81895.17, 80450.7, 90521.85,
  100975.6, 100936.5, 98674.52, 93506.97, 90743.43, 88852.44, 87566.21, 
    87905.66, 83053.97, 80345.83, 79542.24, 80232.73, 82395.77, 81288.22, 
    91915.59,
  92031.72, 88386.53, 93356.91, 92012.02, 85514.64, 84434.65, 86662.17, 
    85974.56, 81113.42, 78920.25, 78055.39, 78752.18, 80061.55, 81597.94, 
    93911.98,
  85882.81, 85977.91, 85025.21, 83372.66, 83099.59, 81645.52, 82506.72, 
    82796.85, 80559.64, 79336.49, 78984.28, 80536.43, 80158.34, 82150.63, 
    88003.25,
  87448.96, 86509.12, 87518.7, 86661.81, 86502.1, 84880.66, 83843.37, 
    83378.15, 82415.7, 84377.8, 99304.3, 99807.64, 90152.26, 90558.01, 
    83162.12,
  87783.58, 85973.17, 88410.02, 89226.43, 88312.12, 87865.88, 87143.08, 
    87491.42, 89090.58, 100040.6, 100879.2, 100810.9, 100647.2, 92624.36, 
    77817.71,
  87041.13, 86233.78, 88337.5, 89568.6, 89301.64, 89283.88, 89215.8, 
    91193.55, 95145.36, 100763.4, 100699.6, 100756.8, 100665.5, 86657.27, 
    77587.91,
  90779.8, 87507.14, 87959.15, 89739.11, 89351.61, 88307.36, 88895.45, 
    90706.7, 94959.37, 100762.9, 100745.2, 100815, 100708.3, 85474.78, 
    87350.74,
  93801.3, 89468.62, 88560.99, 89634.41, 88762.47, 86394.12, 87633.41, 
    90271.46, 100266.3, 100744.2, 100722.7, 100733, 100752.1, 92925.18, 
    95679.48,
  96952.05, 92312.16, 90799.86, 93200.12, 93388.86, 93452.41, 94339.59, 
    100242.5, 100763.9, 100743.4, 100740.4, 100709, 100732.2, 98458.2, 
    99647.85,
  101372.2, 101037.7, 97120.7, 94605.91, 94578.07, 93538.95, 91242.62, 
    91683.99, 85954.98, 81312.44, 79074.25, 79342.47, 82308.12, 80896.09, 
    91227.87,
  101305.9, 101270.9, 99001.03, 93846.63, 91060.98, 89176.45, 87906.22, 
    88245.6, 83406.24, 80693.99, 79944.57, 80611.77, 82799.23, 81731.68, 
    92580.14,
  92249.81, 88713.32, 93660.59, 92340.89, 85822.95, 84775.35, 87039.84, 
    86334.57, 81447.9, 79233.31, 78380.62, 79076.23, 80447.43, 82028.83, 
    94549.18,
  86153.12, 86307.46, 85349.54, 83693.95, 83432.17, 81963.55, 82843.57, 
    83155.61, 80889.53, 79691.66, 79363.59, 80884.91, 80577.59, 82530.93, 
    88589.36,
  87752.06, 86812.85, 87809.04, 86972.69, 86839.26, 85217.16, 84198.21, 
    83714.87, 82769.19, 84736.19, 99599.53, 100176, 90467.1, 90896.2, 83671.27,
  88086.59, 86268.96, 88714.2, 89554.76, 88675.69, 88229.37, 87515.99, 
    87882.69, 89457.65, 100359.9, 101290, 101208.2, 100985.7, 93045.63, 
    78193.01,
  87301.76, 86532.68, 88627.81, 89868.48, 89641.62, 89641.01, 89577.23, 
    91541.89, 95477.22, 101091.7, 101049.7, 101089.2, 100935, 87074.95, 
    77934.69,
  91039.57, 87787.93, 88249.81, 90053.15, 89724.16, 88695.13, 89267.31, 
    91051.12, 95272.36, 101114.6, 101107.2, 101202.5, 101040.5, 85916.88, 
    87730.45,
  94040.73, 89738.89, 88828.47, 89915.56, 89082.35, 86721.46, 87983.13, 
    90618.23, 100719.4, 101118.1, 101083.5, 101128.5, 101082.9, 93351.14, 
    96050.34,
  97205.93, 92561.35, 91009.56, 93384.65, 93593.23, 93735.78, 94676.69, 
    100674.6, 101196.1, 101139.3, 101137.7, 101147.8, 101145.2, 98890.23, 
    100035.6,
  101328.1, 100994.8, 97041.66, 94533.92, 94457.74, 93383.65, 91084.02, 
    91599.53, 85851.53, 81273.79, 79006.88, 79310.94, 82260.95, 80817.92, 
    91094.84,
  101223.2, 101237.2, 98939.29, 93776.62, 90972.55, 89115.35, 87858.78, 
    88188.8, 83344.88, 80670.88, 79894.64, 80572.05, 82774.42, 81677.91, 
    92466.27,
  92261.41, 88731.81, 93677.05, 92331.06, 85821.32, 84763.52, 87019.2, 
    86316.66, 81449.48, 79258.14, 78378.68, 79080.29, 80445.55, 82016.45, 
    94487.52,
  86130.34, 86263.82, 85367.73, 83720.69, 83474.47, 82018.63, 82884.66, 
    83205.11, 80932.55, 79712.41, 79374.78, 80899.66, 80580.71, 82542.05, 
    88568.75,
  87742.83, 86796.08, 87810.15, 86997.03, 86864.73, 85273.13, 84249.31, 
    83782.15, 82829.51, 84822.42, 99784.37, 100306.5, 90592.73, 90959.34, 
    83652.9,
  88069.67, 86283.15, 88714.01, 89557.4, 88682.76, 88252.26, 87546.55, 
    87936.52, 89533.61, 100452.9, 101294.1, 101275.8, 101096.3, 93084.03, 
    78282.13,
  87236.12, 86490.38, 88612.95, 89872.39, 89651.8, 89677.07, 89633.72, 
    91614.06, 95551.8, 101209.1, 101146.2, 101206.5, 101071.4, 87104.22, 
    78003.35,
  90968.5, 87744.64, 88215.07, 90031.22, 89696.16, 88702.31, 89316.6, 
    91139.38, 95379.63, 101219.5, 101187.5, 101283.3, 101147.8, 85967.91, 
    87916.73,
  93963.59, 89661.38, 88776.03, 89894.08, 89064.17, 86710.42, 88006.7, 
    90599.39, 100677.7, 101214.2, 101186.6, 101228.9, 101208, 93425.77, 
    96187.88,
  97112.16, 92509.3, 90947.48, 93326.69, 93577.52, 93728.5, 94661.02, 
    100583.3, 101220.3, 101198.3, 101212, 101242.9, 101267.2, 99001.77, 
    100157.4,
  100989.2, 100673.7, 96773.16, 94335.78, 94232.88, 93206.7, 90897.77, 
    91395.55, 85656.74, 81117.6, 78889.95, 79174.66, 82196.71, 80771.86, 
    91147.91,
  101057.8, 100989.4, 98648.52, 93542.32, 90813.39, 88972.21, 87684.94, 
    88048.62, 83188.57, 80528.12, 79749.23, 80442.11, 82708.12, 81588.07, 
    92496.77,
  91981.8, 88539.57, 93521.09, 92114.05, 85630.89, 84631.16, 86864.69, 
    86173.47, 81324.92, 79161.18, 78274.23, 78994.43, 80382.77, 81961.72, 
    94481.33,
  86001.86, 86173.36, 85190.98, 83598.5, 83330.65, 81892.96, 82784.18, 
    83105.02, 80823.52, 79598.17, 79275.73, 80822.99, 80471.84, 82482.85, 
    88559.05,
  87607.79, 86710.95, 87697.77, 86880.73, 86747.73, 85149.48, 84146.88, 
    83678.9, 82722.7, 84764.48, 99752.12, 100204.5, 90495.77, 90926.6, 
    83590.12,
  88002.27, 86212.34, 88650.44, 89459.55, 88600.2, 88157.5, 87476.25, 
    87850.97, 89508.51, 100405.3, 101175.9, 101140.3, 101048.2, 92953.96, 
    78241.35,
  87253.98, 86498.05, 88601.35, 89800.64, 89614.07, 89620.27, 89597.53, 
    91571.05, 95559.39, 101120.3, 101089.1, 101078.3, 101035.6, 87014.44, 
    78026.3,
  91024.95, 87757.86, 88265.47, 90037.45, 89698.8, 88723.89, 89348.75, 
    91136.06, 95413.42, 101157.2, 101137.1, 101144.5, 101014.9, 85883.73, 
    87887.25,
  94030.38, 89714.91, 88870.95, 89925.44, 89139.02, 86795.5, 88088.78, 
    90685.21, 100731.3, 101194.6, 101145.8, 101125.8, 101023, 93364.34, 
    96143.48,
  97209.43, 92552.51, 91055.31, 93433.18, 93660.06, 93817.18, 94766.94, 
    100687.1, 101242.6, 101232.3, 101214.8, 101196.5, 101144, 98950.56, 
    100182.5,
  101123.5, 100817.3, 96902.52, 94384.4, 94288.17, 93239.4, 90915.06, 
    91448.89, 85723.33, 81220.55, 79047.77, 79457.6, 82571.55, 81197.75, 
    91651.37,
  101175.7, 101070.4, 98858.73, 93686.3, 90903.4, 88968.88, 87724.81, 
    88110.31, 83219.2, 80644.16, 79906.77, 80688.43, 83025.05, 81978.19, 
    93068.63,
  92047.21, 88740.41, 93561.02, 92164.35, 85707.39, 84741.4, 86969.37, 
    86214.77, 81378.06, 79300.1, 78451.81, 79239.62, 80678.76, 82340.05, 
    95058.59,
  86322.34, 86483.46, 85452.71, 83843.04, 83536.66, 82041.39, 82894.81, 
    83191.7, 80921.77, 79709.27, 79411.35, 80997.34, 80743.97, 82860.98, 
    89086.8,
  87881.02, 86978.39, 87976.74, 87168.84, 87013.9, 85410.49, 84382.38, 
    83888.01, 82914.58, 85075.77, 100099.7, 100472.1, 90730.85, 91250.19, 
    84036.3,
  88314.12, 86539.02, 89002.88, 89771.13, 88899.67, 88476.6, 87782.68, 
    88155.76, 89869.22, 100696, 101447.4, 101461.6, 101315.5, 93322.17, 
    78581.31,
  87585.91, 86818.2, 88935.44, 90145.02, 89953.55, 89963.87, 89943.53, 
    91885.27, 95884.33, 101425.9, 101383.6, 101346.2, 101341.5, 87322.34, 
    78304.2,
  91293.14, 88102.88, 88595.98, 90356.22, 90038.55, 89050.22, 89703.33, 
    91473.41, 95779.27, 101464.1, 101415.2, 101420.4, 101352.2, 86204.73, 
    88149.96,
  94276.83, 90046.89, 89195.66, 90273.7, 89453.45, 87140.65, 88410.51, 
    91073.81, 101081.6, 101484.4, 101405.9, 101388.1, 101382.3, 93671.12, 
    96340.15,
  97426.4, 92843.15, 91355.2, 93715.27, 93972.98, 94147.38, 95085.08, 
    101038.3, 101554.6, 101504.3, 101451.3, 101412.8, 101406.2, 99156.66, 
    100369.8,
  101178.5, 100891.3, 96982.29, 94461.95, 94430.74, 93390.53, 91096.79, 
    91634.09, 85870.74, 81344.12, 79122.53, 79519.17, 82584.27, 81202.99, 
    91614.11,
  101182.4, 101085.5, 98866.91, 93765.87, 90993.41, 89117.02, 87872.7, 
    88217.16, 83369.61, 80746.74, 79988.45, 80737.49, 83039.27, 82046.99, 
    93011.8,
  92192.25, 88809.95, 93623.57, 92230.85, 85843.42, 84844.71, 87076.68, 
    86365.6, 81540.38, 79359.33, 78506.96, 79254.86, 80712.98, 82386.49, 
    95062.15,
  86356.23, 86513.45, 85532.64, 83915.61, 83629.3, 82164.57, 82990.18, 
    83306.59, 81044.12, 79781.19, 79478.68, 80993.27, 80775.4, 82874.62, 
    89107.34,
  87906.1, 86989.3, 87992.16, 87204.52, 87046.41, 85445.65, 84424.12, 
    83911.22, 82952.88, 85028.51, 100013.3, 100447.9, 90732.4, 91285.15, 
    84087.04,
  88283.54, 86507.52, 88960.24, 89767.29, 88900.73, 88463.89, 87752.13, 
    88125.48, 89790.05, 100652.4, 101424.5, 101416, 101328.5, 93374.46, 
    78589.93,
  87483.38, 86737.61, 88829.66, 90087.89, 89897.33, 89930.45, 89874.16, 
    91796.82, 95778.29, 101378.2, 101324.1, 101350.4, 101362.2, 87293.59, 
    78284.47,
  91107.47, 87974.77, 88453.3, 90244.29, 89948.63, 88973.31, 89598.06, 
    91358.77, 95628.42, 101411.5, 101379.5, 101455.5, 101362.8, 86164.26, 
    88120.12,
  93995.22, 89864.57, 88997.62, 90102.8, 89337.47, 87052.09, 88296.34, 
    90861.44, 100880.3, 101401.1, 101369, 101436.8, 101414.2, 93685.1, 
    96346.93,
  97078.84, 92601.27, 91101.17, 93467.49, 93718.71, 93873.64, 94807.8, 
    100697.7, 101359.9, 101394.1, 101390.3, 101425.6, 101449.8, 99175.23, 
    100341.5,
  101134.9, 100808.2, 96937.71, 94442.38, 94414.09, 93413.95, 91115.16, 
    91612.73, 85850.28, 81332.78, 79061.45, 79364.2, 82380.49, 80932.58, 
    91326.31,
  101027.1, 101016.4, 98785.61, 93713.12, 90970.8, 89110.7, 87886.44, 
    88220.51, 83365.19, 80707.45, 79924.4, 80626.36, 82860.62, 81766.3, 
    92717.2,
  92190.21, 88696.48, 93606.66, 92239.88, 85826.12, 84786.52, 87043.9, 
    86332.55, 81521.66, 79350.54, 78432.23, 79151.11, 80549.96, 82120.87, 
    94650.33,
  86186.47, 86289.1, 85412.14, 83785.01, 83532.92, 82066.3, 82929.93, 
    83259.41, 80975.16, 79761.08, 79409.46, 80953.25, 80580.15, 82645.39, 
    88707.19,
  87785.57, 86839.09, 87855.13, 87028.46, 86889.89, 85303.34, 84274.56, 
    83794.37, 82852.25, 84855.84, 99675.47, 100224.1, 90556.39, 91003.77, 
    83745.53,
  88094.66, 86302.02, 88734.8, 89542.5, 88688.12, 88257.22, 87565.73, 
    87944.74, 89532.96, 100349.2, 101196.6, 101155.8, 100989.1, 93062.22, 
    78346.98,
  87261.56, 86552.59, 88648, 89884.51, 89653.95, 89671.77, 89629.22, 
    91544.72, 95481.06, 101108.5, 101075.7, 101095.2, 101069.1, 87090.15, 
    78095.16,
  90890.52, 87786.05, 88245.34, 90055.61, 89718.98, 88726.16, 89340.04, 
    91125.98, 95317.34, 101102.9, 101114.8, 101180.5, 101085.1, 85909.34, 
    87940.86,
  93787.95, 89668.81, 88839.84, 89917.94, 89117.8, 86827.07, 88110.39, 
    90657.78, 100553.7, 101114.5, 101113.2, 101166.5, 101127.1, 93434.53, 
    96109.11,
  96899.46, 92399.91, 90920.8, 93366.74, 93551.5, 93681.31, 94674.11, 
    100489.7, 101065.3, 101128, 101148.2, 101192.1, 101189.8, 98933.78, 
    100060.9,
  101025.8, 100713.7, 96885.7, 94456.55, 94448.55, 93463.41, 91192.38, 
    91688.02, 85987.02, 81439.41, 79166.74, 79452.03, 82351.9, 80984.41, 
    91142.91,
  100965.7, 100968.7, 98721.09, 93687.47, 90983.78, 89160.76, 87921.16, 
    88268.45, 83453.18, 80786.09, 79987.37, 80659.62, 82846.15, 81776.49, 
    92507.56,
  92242.09, 88702.72, 93579.24, 92259.66, 85887.37, 84840.82, 87067.73, 
    86374.6, 81565.14, 79393.41, 78502.38, 79192.02, 80549.34, 82096.47, 
    94540.73,
  86209.5, 86278.4, 85430.94, 83786.05, 83541.35, 82097.67, 82962.93, 
    83271.77, 81033.88, 79797.23, 79437.81, 80961.2, 80598.8, 82591.65, 
    88613.41,
  87769.59, 86790.05, 87840.64, 87031.48, 86915.16, 85330.2, 84316.93, 
    83832.23, 82889.73, 84842.15, 99656.72, 100196.1, 90555.14, 90969.85, 
    83708.55,
  88077.4, 86303.85, 88741.09, 89561.08, 88706.76, 88259.3, 87577.03, 
    87950.62, 89476.7, 100343.4, 101167.7, 101095.8, 100926.2, 93024.4, 
    78290.44,
  87281.61, 86568.55, 88645.16, 89864.41, 89672.35, 89694.42, 89643.91, 
    91553.95, 95536.49, 101103, 101040.2, 101057.6, 101013.2, 87057.83, 
    78083.91,
  90986.02, 87809.92, 88277.4, 90055.78, 89739.16, 88733.75, 89336.16, 
    91137.85, 95367.88, 101101.8, 101096.4, 101119.5, 101031, 85868.58, 
    87916.23,
  93985.91, 89740.05, 88864.45, 89934.41, 89133.93, 86819.59, 88097.31, 
    90672.34, 100644, 101140.1, 101099.4, 101101.2, 101049, 93375.74, 96018.2,
  97131.61, 92548.25, 91028.27, 93390.93, 93656.15, 93785.23, 94723.29, 
    100608.2, 101170.5, 101156.1, 101136.1, 101125.4, 101079.4, 98840.7, 
    99981.43,
  101391.8, 101085.3, 97126.42, 94698.12, 94695.45, 93704.73, 91446.98, 
    91935.29, 86232, 81686.54, 79417.72, 79708.95, 82568.47, 81174.63, 
    91206.95,
  101265.6, 101254.8, 98956.05, 93893.84, 91230.92, 89425.64, 88174.04, 
    88534.54, 83723.51, 81042.37, 80249.55, 80915.47, 83076.64, 81993.38, 
    92568.61,
  92353.73, 88981.2, 93861.56, 92495.79, 86113.16, 85088.82, 87325, 86652.57, 
    81820.26, 79650.3, 78751.45, 79460.75, 80774.07, 82306.57, 94614.44,
  86345.77, 86534.92, 85595.27, 84042.91, 83797.84, 82366.1, 83223.85, 
    83530.65, 81293.77, 80084.03, 79719.62, 81221.43, 80846.94, 82822.78, 
    88730.44,
  87950.02, 87065.79, 88055.14, 87253.64, 87131.15, 85565.55, 84563.01, 
    84104.12, 83152.59, 85125.09, 99973.3, 100599.1, 90906.56, 91255.75, 
    83885.46,
  88338.98, 86549.76, 89004.34, 89813.7, 88960.75, 88534.77, 87845.94, 
    88224.27, 89807.13, 100719.1, 101600.4, 101494.8, 101306.6, 93357.33, 
    78447.3,
  87572.7, 86820.38, 88924.67, 90125.2, 89930.55, 89952.52, 89896.33, 
    91857.8, 95893.28, 101507.2, 101416.4, 101413.7, 101382.4, 87341.53, 
    78263.17,
  91254.78, 88069.57, 88561.99, 90336.34, 90010.04, 89002.1, 89668.74, 
    91468.97, 95714.47, 101490.3, 101437.3, 101464.9, 101389, 86131.12, 
    88166.98,
  94216.7, 90001.84, 89158.15, 90233.23, 89421.67, 87095.31, 88380.57, 
    90968.46, 101100.7, 101483.1, 101421.1, 101413.7, 101367.2, 93667.19, 
    96268.45,
  97330.74, 92804.04, 91316.98, 93663.51, 93944.21, 94106.87, 95073.55, 
    100988.6, 101518.6, 101474, 101442.2, 101410.2, 101373.8, 99116.41, 
    100207.4,
  101500.3, 101220.3, 97210.02, 94771.97, 94740.88, 93719.13, 91474.16, 
    91972.11, 86280.1, 81767.73, 79535.99, 79869.23, 82781.87, 81381.69, 
    91416.48,
  101518.7, 101437.1, 99156.45, 94039.73, 91299.47, 89492.69, 88229.73, 
    88603.55, 83803.06, 81169.65, 80404.08, 81102.38, 83275.7, 82212.16, 
    92766.61,
  92498.12, 89081.88, 93953.88, 92571.52, 86208.76, 85194.77, 87408.88, 
    86741.84, 81919.91, 79782.04, 78912.52, 79625.89, 80968.07, 82523.4, 
    94782.44,
  86579.25, 86776.4, 85802.88, 84190.11, 83930.54, 82480.55, 83335.95, 
    83651.63, 81416.91, 80228.16, 79886.96, 81395.22, 81079.23, 83013.96, 
    88906.83,
  88180.86, 87221.26, 88236.97, 87435.05, 87294.6, 85724.15, 84700.34, 
    84232.84, 83298.97, 85252.53, 100076.8, 100673.1, 91007.78, 91405.16, 
    84152.83,
  88533.67, 86714.23, 89166.53, 89980.53, 89113.98, 88689.28, 87992.63, 
    88373, 89923.49, 100836.1, 101731.3, 101630, 101416, 93539.62, 78680.12,
  87667.34, 86931.45, 89015.85, 90262.97, 90071.38, 90098.3, 90051.48, 
    91990.3, 95974.79, 101600.3, 101523.2, 101584.7, 101470.4, 87574.77, 
    78464.63,
  91277.93, 88148.12, 88634.84, 90404.06, 90116.64, 89136.45, 89775.87, 
    91549.35, 95783.09, 101595.2, 101580.6, 101661.3, 101538.2, 86366.45, 
    88327.98,
  94160.04, 90038.48, 89173.68, 90268.72, 89497.43, 87198.65, 88473.97, 
    91023.91, 101026.1, 101589.4, 101561, 101602.6, 101579.5, 93855.76, 
    96536.24,
  97260.58, 92759.34, 91266.08, 93612.13, 93878.11, 94034.81, 94995.59, 
    100924.8, 101556.1, 101568.8, 101583.6, 101604.4, 101618.7, 99368.67, 
    100468.6,
  101166.3, 100907.8, 97072.29, 94653.26, 94643.46, 93640.83, 91377.29, 
    91864.42, 86174.84, 81669.52, 79422.02, 79697.77, 82660.45, 81224.74, 
    91303.62,
  101119.3, 101154.6, 98934.84, 93919.06, 91200, 89403.87, 88158.05, 
    88497.82, 83703.29, 81049.95, 80261.37, 80950.54, 83136.34, 82037.79, 
    92650.96,
  92360.99, 88942.62, 93792.88, 92441.92, 86127.02, 85124.2, 87345.76, 
    86629.62, 81841.03, 79681.98, 78797.97, 79491.32, 80830.14, 82391.05, 
    94617.3,
  86413.26, 86514.52, 85702.28, 84081.89, 83851.2, 82398.38, 83240.7, 
    83561.77, 81333.07, 80101.05, 79747.12, 81251.9, 80931.91, 82875.32, 
    88775.81,
  87976, 86932.42, 88031.79, 87248.2, 87141.45, 85598.89, 84596.88, 84117.8, 
    83171.63, 85146.9, 99834.4, 100410.2, 90809.56, 91174.63, 84004.36,
  88285.86, 86457.02, 88900.32, 89747.54, 88916, 88504.91, 87811.46, 
    88220.16, 89768.85, 100459.9, 101347.9, 101305.1, 101123.8, 93303.26, 
    78579.29,
  87369.09, 86676.38, 88770.49, 90031.55, 89866.92, 89920.84, 89863.08, 
    91765.44, 95587.02, 101215.9, 101203.9, 101270, 101163.5, 87381.06, 
    78354.86,
  90963.34, 87854.83, 88337.78, 90141.72, 89870.38, 88925.41, 89550.27, 
    91330.9, 95416.94, 101181.4, 101208.3, 101319.8, 101215.9, 86196.86, 
    88139.94,
  93914.71, 89742.79, 88890.12, 89986.59, 89272.07, 87022.03, 88275.01, 
    90776.75, 100540.1, 101153.5, 101184.2, 101269.5, 101237.9, 93605.44, 
    96284.37,
  97059.22, 92503.88, 90944.77, 93301.81, 93573.62, 93713.3, 94662.05, 
    100441.3, 101036.2, 101124.2, 101187.5, 101257.7, 101291, 99067.17, 
    100197.9,
  100913, 100578.2, 96827.53, 94382.12, 94321.48, 93329.24, 91098.3, 
    91594.05, 85986.51, 81499.12, 79272.12, 79556.01, 82411.26, 81034.61, 
    90928.25,
  100613.4, 100670.7, 98511.58, 93544.3, 90917.69, 89126.27, 87885.32, 
    88237.03, 83499.5, 80868.59, 80096.78, 80765.2, 82899.87, 81840.45, 
    92305.98,
  92020.39, 88493.67, 93360.92, 92073.39, 85793.95, 84769.03, 87012.58, 
    86365.32, 81605.77, 79462.27, 78583.77, 79273.98, 80583.79, 82114.98, 
    94298.75,
  86011.25, 85941.44, 85195.71, 83634.34, 83406.05, 82021.46, 82907.02, 
    83239.11, 81038.23, 79859.79, 79522.73, 81014.68, 80680.46, 82598.74, 
    88452.59,
  87527.3, 86456.91, 87533.59, 86687.73, 86619.45, 85093.03, 84151.63, 
    83741.46, 82848.69, 84760.07, 99224.76, 99872.1, 90440.5, 90835.06, 
    83709.4,
  87773.86, 85996.12, 88407.62, 89216.41, 88377.47, 87972.26, 87317.3, 
    87730.15, 89282.46, 99865.31, 100760.5, 100731.8, 100570, 92900.65, 
    78310.22,
  86987.07, 86257.36, 88306.81, 89537.14, 89310.56, 89357.19, 89317.93, 
    91258.54, 95100.07, 100595.2, 100601.5, 100663.7, 100637.8, 87025.52, 
    78079.34,
  90657.52, 87503.83, 87923.51, 89697.59, 89367.5, 88381.05, 88979.37, 
    90801.59, 94889.84, 100554.8, 100594.3, 100700.5, 100657.3, 85838.98, 
    87762.42,
  93604.13, 89411.24, 88520.09, 89574.93, 88787.72, 86515.91, 87751.77, 
    90261.66, 100039.8, 100564.4, 100564.7, 100653.8, 100698.3, 93124.67, 
    95819.43,
  96740.29, 92167.77, 90633.3, 92990.49, 93221.95, 93341.09, 94257.12, 
    100058, 100590.6, 100532.7, 100585.1, 100641.9, 100720.3, 98523.63, 
    99701.36,
  101300.2, 100920.7, 97081.83, 94579.47, 94497.45, 93470.7, 91184.71, 
    91571.87, 85948.16, 81391.7, 79180.66, 79491.95, 82337.45, 81043.65, 
    90778.04,
  101054.8, 101108.8, 98891.77, 93783.13, 91031.95, 89177.7, 87923.11, 
    88216.37, 83442.42, 80732.52, 79991.41, 80665.05, 82802.68, 81815.28, 
    92089.73,
  92296.07, 88700.73, 93607.61, 92302.32, 85900.56, 84744.66, 87008.05, 
    86329.07, 81499.23, 79311.81, 78460.05, 79164.72, 80489.66, 82030.12, 
    94000.7,
  86152.6, 86100.38, 85323.91, 83690.3, 83430.47, 82005.53, 82853.6, 
    83152.33, 80907.41, 79741.05, 79383.19, 80862.95, 80586.2, 82469.56, 
    88242.64,
  87697.55, 86611.14, 87694.5, 86861.21, 86742.44, 85162.59, 84140.68, 
    83670.39, 82744.09, 84640.65, 99219.9, 99901.47, 90397.33, 90656.38, 
    83615.06,
  87814.88, 86086.95, 88504.16, 89371.05, 88507.88, 88080, 87373.09, 
    87750.83, 89271.27, 99985.25, 100920.8, 100889.9, 100633.7, 92845.83, 
    78184.43,
  86976.71, 86277.98, 88359.55, 89622.09, 89412.77, 89440.28, 89360.77, 
    91290.31, 95133.07, 100690.6, 100652.6, 100741, 100563.2, 86988.04, 
    77868.34,
  90626.7, 87437.88, 87917.91, 89720.95, 89415.77, 88440.37, 89018.39, 
    90803.85, 94892.27, 100644.3, 100627.3, 100744.4, 100568, 85799.52, 
    87366.75,
  93569.18, 89344.81, 88468.52, 89550.48, 88771.96, 86475.73, 87704.31, 
    90223.02, 100095.9, 100633, 100547.6, 100587.9, 100545, 93012.7, 95457.66,
  96677.47, 92101.38, 90568.01, 92918.78, 93161.82, 93289.84, 94206.48, 
    100077.8, 100613.5, 100546.8, 100498.6, 100479.6, 100496.8, 98316.48, 
    99379.88,
  101354.1, 101000.9, 97128.89, 94632.97, 94550.86, 93526.38, 91268.62, 
    91669.64, 86048, 81505.04, 79264.18, 79576.77, 82397.48, 81102.02, 
    90912.73,
  101260.1, 101231.3, 98967.69, 93853.69, 91114.77, 89257.52, 88010.41, 
    88317.82, 83557.42, 80849.44, 80111.82, 80778.03, 82904.12, 81920.06, 
    92244.73,
  92338.85, 88823.97, 93731.77, 92394.26, 85969.38, 84877.62, 87136.24, 
    86456.16, 81631.12, 79443.12, 78578.36, 79276.55, 80602.08, 82157.78, 
    94220.13,
  86254.02, 86363.17, 85437.43, 83821.41, 83562.73, 82133.36, 82990.15, 
    83297.1, 81048.14, 79869.17, 79510.86, 80992.98, 80692.32, 82600.77, 
    88419.19,
  87853.04, 86903.74, 87889.57, 87066.21, 86911.52, 85333.55, 84310.86, 
    83851.62, 82897.19, 84863.12, 99561.8, 100231.6, 90619, 90899.41, 83756.76,
  88128.95, 86326.59, 88760.62, 89591.88, 88712.85, 88276.16, 87562.94, 
    87939.45, 89515.03, 100343.7, 101186.5, 101137.5, 100877.4, 93079.77, 
    78256.84,
  87338.67, 86588.87, 88666.22, 89906.05, 89683.45, 89702.02, 89632.84, 
    91602.45, 95494.62, 101080.9, 100970, 101037.5, 100878.6, 87132.86, 
    77944.56,
  91055.88, 87804.12, 88271.25, 90046.5, 89704.79, 88715.57, 89326.84, 
    91126.38, 95300.54, 101062.2, 100989.4, 101046.1, 100895.3, 85913.17, 
    87613.87,
  94047.16, 89767.21, 88901.33, 89966.31, 89112.89, 86775.36, 88041.68, 
    90643.38, 100671.2, 101054.9, 100934.3, 100944, 100876.2, 93265.27, 
    95787.59,
  97205.17, 92614.19, 91065.91, 93436.27, 93676.52, 93840.56, 94755.55, 
    100629, 101095.7, 101013.9, 100948.7, 100908.6, 100874.8, 98652.2, 
    99725.25,
  101570, 101217, 97288.81, 94733.47, 94605.93, 93486.72, 91134.61, 91639.05, 
    85886.21, 81366.9, 79096.78, 79408.19, 82342.45, 80973.71, 91049.95,
  101543.7, 101401.3, 99193.41, 94047.91, 91219.27, 89292.97, 88022.35, 
    88303.73, 83406.2, 80764.3, 79964.58, 80712.3, 82878.7, 81733.52, 92487.19,
  92451.54, 89071.41, 93889.87, 92484.29, 86074.23, 84997.25, 87206.56, 
    86456.53, 81606.27, 79434.66, 78503.38, 79188.16, 80564.1, 82134.52, 
    94557.2,
  86588.23, 86794.75, 85787.57, 84138.34, 83873.52, 82360.2, 83168.87, 
    83455.77, 81151.58, 79882.52, 79591.99, 81097.16, 80648.12, 82653.25, 
    88483.53,
  88166.37, 87247.12, 88274.62, 87443.54, 87257.95, 85652.51, 84613.93, 
    84100.71, 83099.08, 85235.23, 100265.8, 100721.9, 90885.5, 91152.2, 
    83741.43,
  88582.2, 86770.42, 89258.21, 90052.17, 89146.52, 88703.77, 87984.77, 
    88381.56, 90028.12, 101020.9, 101731.8, 101651.2, 101366.9, 93280.45, 
    78274.87,
  87810.57, 87028.46, 89140.9, 90378.67, 90170.77, 90176.52, 90148.62, 
    92129.94, 96126.12, 101771.9, 101666.4, 101621.8, 101455.7, 87277.02, 
    78117.02,
  91509.77, 88295.31, 88807.11, 90578.39, 90276.75, 89238.29, 89880.27, 
    91654.62, 96005.02, 101777.6, 101687.6, 101672.2, 101521.3, 86060.15, 
    87999.73,
  94482.27, 90247.79, 89382.47, 90490.47, 89665.73, 87312.43, 88591.1, 
    91253.07, 101366.8, 101781.8, 101675.8, 101651.7, 101530.2, 93710.68, 
    96314.3,
  97665.5, 93073.2, 91555.28, 93928.76, 94191.59, 94384.16, 95319.84, 
    101298.7, 101817.9, 101782.3, 101701, 101646.4, 101573, 99277.54, 100337.1,
  101783.8, 101410, 97494.16, 94965.77, 94874.59, 93814.3, 91453.61, 91964.8, 
    86175.56, 81656.43, 79372.43, 79714.59, 82648.95, 81194.32, 91309.97,
  101682.6, 101626.6, 99415.52, 94300.79, 91484.08, 89592.53, 88333.93, 
    88598.98, 83688.95, 81046.55, 80261.91, 80949.02, 83105.01, 81981.96, 
    92798.16,
  92723.12, 89299.41, 94117.11, 92734.55, 86340.02, 85274.07, 87482.1, 
    86715.93, 81881.07, 79706.89, 78765.13, 79486.51, 80808.12, 82386.15, 
    94788.99,
  86805.98, 86926.4, 85997.85, 84342.76, 84076.45, 82586.35, 83405.84, 
    83697.27, 81391.27, 80113.34, 79819.43, 81387.98, 80914.84, 82965.77, 
    88821.03,
  88439.17, 87372.01, 88368.95, 87577.63, 87426.73, 85851.49, 84806.13, 
    84302.09, 83298.4, 85386.01, 100363.3, 100905.8, 91115.23, 91530.31, 
    83970.68,
  88675.14, 86881.23, 89272.71, 90099.73, 89233.85, 88816.48, 88105.31, 
    88490.26, 90076.61, 100961.2, 101870.1, 101878.6, 101735.4, 93600.78, 
    78516.8,
  87794.07, 87066.4, 89110.04, 90350.66, 90160.08, 90191.42, 90147.09, 
    92080.9, 95974.09, 101713.7, 101754.9, 101780.7, 101798.1, 87500.73, 
    78356.54,
  91404.95, 88263.53, 88701.91, 90482.86, 90167.88, 89187.62, 89814.5, 
    91621.3, 95788.32, 101645.5, 101704.8, 101815.4, 101748.8, 86344.55, 
    88329.88,
  94271.69, 90114.85, 89227.44, 90310.16, 89544.28, 87239.8, 88493.45, 
    91026.34, 100953.3, 101592.9, 101633.9, 101735.2, 101731.4, 93934.31, 
    96551.32,
  97372.94, 92861.59, 91293.31, 93631.29, 93882.06, 94039.34, 94960.4, 
    100834, 101455.5, 101525.5, 101584.7, 101650.8, 101715.8, 99489.5, 
    100621.3,
  101664.1, 101309.6, 97429.44, 94913.45, 94838.35, 93782.18, 91468.16, 
    91961.23, 86271.82, 81736.48, 79471.57, 79746.48, 82628.02, 81265.55, 
    91294.37,
  101562.8, 101472.5, 99309.66, 94251.96, 91452.29, 89568.93, 88327.91, 
    88601.95, 83782.58, 81099.16, 80305.59, 80968.24, 83137.29, 82059.05, 
    92622.28,
  92683.66, 89191.05, 93966.18, 92667.26, 86316.23, 85243.94, 87437.17, 
    86723.45, 81920.61, 79734.68, 78813.9, 79485.98, 80817.83, 82364.26, 
    94663.04,
  86778.08, 86851.15, 85931.03, 84283.1, 84006.61, 82546.94, 83344.08, 
    83644.6, 81380.59, 80130.89, 79789.66, 81282.73, 80892.97, 82838.07, 
    88731.56,
  88366.08, 87323.36, 88275.34, 87476, 87288.27, 85725.96, 84685.48, 84199.2, 
    83235.73, 85237.02, 99859.19, 100467.7, 90873.91, 91192.48, 83958.64,
  88594.96, 86822.31, 89192.08, 90011.42, 89117.34, 88672.49, 87934.55, 
    88310.34, 89842.54, 100531.4, 101356.1, 101331.4, 101097.6, 93303.31, 
    78504.21,
  87764.88, 87036.48, 89057.93, 90269.09, 90039.76, 90045.02, 89957.55, 
    91865.57, 95717.73, 101269.3, 101241.1, 101301.7, 101172.4, 87386.15, 
    78228.82,
  91423.92, 88249.66, 88671.45, 90425.66, 90096.7, 89089.46, 89666.05, 
    91413.41, 95560.25, 101237.1, 101216.8, 101312.5, 101182.6, 86181.55, 
    87985.46,
  94305.59, 90119.8, 89208.74, 90271.84, 89451.17, 87122.19, 88336.88, 
    90897.59, 100752.3, 101220.8, 101184.9, 101251.9, 101223.4, 93585.48, 
    96193.69,
  97426.47, 92895.9, 91324.92, 93633.76, 93839.49, 94028.58, 94903.11, 
    100683.6, 101202.3, 101189.8, 101171.2, 101201.1, 101237.1, 99055.3, 
    100190.6,
  101507.9, 101158.8, 97318.73, 94856.22, 94764.37, 93734.64, 91450.86, 
    91961.22, 86239.05, 81733.38, 79471.62, 79757.35, 82634.04, 81251.16, 
    91273.52,
  101436, 101408, 99186.88, 94144.4, 91381.04, 89548.36, 88315.75, 88603.48, 
    83775.43, 81124.51, 80332.09, 80995.03, 83163.27, 82062.09, 92704.96,
  92629.9, 89178.59, 93973.29, 92635.55, 86314.34, 85275.85, 87476.09, 
    86755.06, 81949.73, 79782.74, 78851.26, 79547.31, 80881.2, 82417.55, 
    94753.46,
  86757.45, 86834.27, 85947.63, 84297.41, 84056.12, 82599.27, 83416.09, 
    83715.91, 81457.93, 80179.8, 79878.86, 81454.67, 80951.71, 82990.34, 
    88796.7,
  88316.23, 87293.12, 88301.72, 87490.08, 87347.81, 85794.89, 84781.33, 
    84297.71, 83334.23, 85371.82, 100205.1, 100715.2, 91115.97, 91448.95, 
    83992.38,
  88600.77, 86823.67, 89222.6, 90048.05, 89177.98, 88753.85, 88053.45, 
    88452.33, 90012.48, 100803.9, 101647.2, 101654, 101456.8, 93507.2, 
    78564.48,
  87726.85, 87013.68, 89083.41, 90325.3, 90130.55, 90161.41, 90109.28, 
    92027.42, 95910.4, 101551.3, 101527.2, 101589.6, 101541.3, 87508.45, 
    78378.16,
  91321.23, 88209.01, 88683.53, 90465.41, 90160.44, 89193.93, 89814.35, 
    91598.4, 95744.41, 101491.3, 101500.2, 101598.8, 101519.9, 86288.82, 
    88254.18,
  94187.34, 90071.34, 89212.04, 90306.83, 89543.91, 87265.23, 88515.55, 
    91061.16, 100930.5, 101463.6, 101456.9, 101515.8, 101486.7, 93824.31, 
    96369.4,
  97260.59, 92804.98, 91298.68, 93654.69, 93901.02, 94049.77, 94980.34, 
    100812.6, 101386, 101408.2, 101424.4, 101446.5, 101456.7, 99238.34, 
    100316.4,
  101458.7, 101134.8, 97317.84, 94856.2, 94775.22, 93752.88, 91467.77, 
    91965.13, 86280.11, 81781.77, 79530.03, 79824.09, 82709.63, 81355.02, 
    91361.48,
  101373.1, 101345.9, 99175.53, 94165.59, 91414.11, 89569.16, 88338.79, 
    88619.9, 83824.38, 81162.96, 80371.18, 81042.64, 83206.11, 82148.46, 
    92716.92,
  92659.11, 89175.88, 93908.13, 92617.24, 86312.07, 85267.16, 87464.1, 
    86761.02, 81974.37, 79797.61, 78894.73, 79582.91, 80921.17, 82468.09, 
    94744.77,
  86749, 86773.21, 85945.5, 84307.82, 84047.27, 82596.69, 83406.1, 83693.91, 
    81449.71, 80204.87, 79876.99, 81366.76, 81000.27, 82948.95, 88869.66,
  88250.78, 87199.47, 88212.46, 87414.33, 87268.36, 85734.6, 84716.47, 
    84238.75, 83288.76, 85264.46, 99882.34, 100459.5, 90924.32, 91300.7, 
    84070.06,
  88498.32, 86744.07, 89113.68, 89930.77, 89063.51, 88648.29, 87941.91, 
    88326.4, 89859.63, 100497.7, 101349, 101331.1, 101156.5, 93390.47, 
    78627.17,
  87602.83, 86910.73, 88949.13, 90188.53, 89993.19, 90024.76, 89954, 
    91859.07, 95674.44, 101246.2, 101243, 101319.5, 101253, 87466.05, 78391.99,
  91233.56, 88118.15, 88571.21, 90334.03, 90024.52, 89056.36, 89655.81, 
    91418.05, 95503.15, 101202.9, 101233.5, 101349.8, 101281, 86250.68, 
    88153.34,
  94120.91, 89978.53, 89110.51, 90180.75, 89416.65, 87125.68, 88352.4, 
    90852.25, 100613.5, 101151.5, 101201.4, 101294.4, 101315.2, 93666.42, 
    96343.66,
  97220.08, 92733.54, 91193.29, 93508.8, 93753.64, 93903.2, 94801.84, 
    100562.7, 101096.8, 101116, 101179.9, 101251, 101332.9, 99115.68, 100265.9,
  101291.6, 100917.5, 97142.84, 94686.15, 94624.8, 93613.73, 91357.35, 
    91843.99, 86235.2, 81748.58, 79522.95, 79817.82, 82648.36, 81274.41, 
    91178.9,
  101239.8, 101192.5, 98996.19, 93991.66, 91271.55, 89434.45, 88220.71, 
    88506.08, 83767.87, 81101.62, 80330.75, 80995.19, 83150.78, 82102.05, 
    92565.25,
  92480.88, 89032.23, 93800.46, 92493.87, 86199.11, 85160.74, 87363.23, 
    86676.8, 81914.86, 79748.29, 78859.91, 79544.91, 80864.26, 82389.05, 
    94571.59,
  86631, 86718.52, 85822.75, 84185.34, 83936.36, 82499.1, 83318.18, 83612.66, 
    81384, 80164.96, 79816.1, 81308.31, 80947.54, 82886.36, 88693.89,
  88174.06, 87220.3, 88192.03, 87397.51, 87235.67, 85694.94, 84672.38, 
    84192.3, 83228.91, 85211.33, 99866.18, 100467.2, 90878.09, 91202.59, 
    83978.62,
  88497.43, 86749.89, 89114.85, 89943.9, 89068.5, 88640.23, 87927.95, 
    88310.48, 89854.36, 100601.1, 101341.6, 101290.2, 101057.9, 93287.16, 
    78555,
  87676.76, 86960.43, 89002.44, 90235.07, 90021.26, 90036.34, 89957.83, 
    91884.98, 95781.9, 101322.8, 101204.6, 101244.1, 101083, 87401.19, 
    78292.22,
  91337.55, 88192.08, 88654.48, 90408.61, 90091.54, 89105.86, 89703.8, 
    91481.88, 95615.18, 101313.6, 101233.7, 101282.4, 101121.4, 86200.91, 
    87972.8,
  94195.74, 90063.1, 89197.43, 90278.73, 89493.45, 87164, 88399.55, 90952.41, 
    100888.6, 101312.8, 101206.9, 101209.8, 101145.1, 93550.43, 96087.48,
  97300.88, 92821.88, 91314.87, 93641.48, 93901.61, 94103.39, 95009.35, 
    100854.5, 101343.7, 101268.7, 101203.3, 101169.5, 101148.1, 98938.62, 
    100019.1,
  100674.1, 100399, 96705.87, 94334.66, 94259.97, 93242.87, 91018.32, 
    91479.55, 85893.57, 81455.7, 79267.96, 79611.56, 82481.34, 81200.34, 
    91036.4,
  100663.5, 100705.3, 98510.34, 93586.62, 90922.66, 89142.83, 87927.05, 
    88196, 83447.14, 80821.23, 80080.23, 80779.84, 82942.38, 81965.19, 
    92354.48,
  92051.68, 88674.34, 93426.37, 92151.68, 85872.32, 84866.61, 87080.13, 
    86386.18, 81628.71, 79484.13, 78634.02, 79343.29, 80684.27, 82239.24, 
    94372.08,
  86168.95, 86309.68, 85459.51, 83849.37, 83613.02, 82198.12, 83036.77, 
    83343.97, 81115.5, 79911.39, 79563.5, 81052.95, 80756.46, 82693.59, 
    88566.1,
  87717.2, 86787.57, 87789.71, 86993.97, 86878.75, 85358.67, 84361.48, 
    83903.7, 82971.52, 84931.82, 99673.91, 100249.5, 90647.34, 91008.83, 
    83847.28,
  88073.45, 86321.72, 88697.64, 89518.29, 88676.67, 88283.2, 87595.72, 
    88001.9, 89542.45, 100355.6, 101200, 101180.7, 100978.2, 93152.48, 
    78407.29,
  87241.09, 86538.45, 88605.97, 89835.89, 89659.97, 89689.03, 89624.38, 
    91560.3, 95457.02, 101098.4, 101047.4, 101144.8, 100989.3, 87225.69, 
    78154.95,
  90861.57, 87766.16, 88233.43, 90000.46, 89699.43, 88739.71, 89362.74, 
    91161.02, 95295.89, 101106.4, 101085.7, 101223.5, 101048.4, 86058.18, 
    87889.63,
  93730.46, 89633.59, 88768.44, 89853.66, 89085.44, 86808.05, 88060.37, 
    90574.55, 100470, 101088.5, 101069, 101152.7, 101097.1, 93456.14, 96011.83,
  96768.55, 92355.36, 90844.29, 93184.47, 93420.44, 93584.7, 94514.7, 
    100383.1, 101017.7, 101066.6, 101086.8, 101134.4, 101144, 98925.93, 
    100013.1,
  100029.8, 99705.31, 95945.45, 93537.3, 93461.03, 92527.98, 90409, 90930.11, 
    85433.17, 80988.72, 78827.95, 79174.98, 82060.13, 80752.25, 90565.26,
  100089.7, 99975.21, 97735.12, 92801.02, 90164.25, 88415.03, 87251.62, 
    87623.05, 82960.55, 80360.66, 79634.63, 80333.86, 82500.25, 81515.29, 
    91828.2,
  91488.35, 88030.2, 92771.38, 91471.64, 85233, 84207.69, 86416.23, 85770.41, 
    81040.84, 78927.88, 78112, 78833.16, 80199.12, 81756.22, 93748.11,
  85699.12, 85744.22, 84869.65, 83246.07, 83031.57, 81593.81, 82446.43, 
    82749.96, 80525.01, 79358.84, 79030.95, 80511.41, 80257.48, 82179.55, 
    88026.58,
  87219.25, 86239.73, 87248.37, 86432.3, 86299.02, 84748.7, 83748.43, 
    83297.84, 82393.48, 84309.18, 98748.02, 99382.55, 89939.76, 90304.89, 
    83322.48,
  87533.73, 85792.47, 88160.51, 88970.46, 88100.3, 87661.77, 86955.41, 
    87325.89, 88862.12, 99473.82, 100447.5, 100348.9, 100097.6, 92441.63, 
    77937.12,
  86724.2, 86006.91, 88028.77, 89255.33, 89044.73, 89064.84, 88971.12, 
    90879.01, 94739.55, 100269.1, 100200.5, 100239.6, 100110.4, 86587.4, 
    77670.07,
  90348.35, 87219.7, 87655.84, 89410.7, 89081.02, 88095.69, 88676.52, 
    90451.81, 94538.94, 100271.9, 100240.4, 100334.8, 100202.2, 85427.52, 
    87251.24,
  93202.45, 89061.33, 88180.09, 89250.54, 88483.17, 86187.7, 87409.39, 
    89910.64, 99734.53, 100289, 100241.5, 100264.8, 100221.1, 92671.36, 
    95345.02,
  96290.34, 91807.5, 90249, 92559.41, 92819.59, 92951.56, 93867.9, 99651.63, 
    100211.1, 100255, 100281.6, 100277.5, 100287.2, 98104.27, 99257.91,
  100107.7, 99720.89, 95962.04, 93514.36, 93469.83, 92491.79, 90299.65, 
    90788.72, 85243.88, 80768.1, 78550.55, 78849.9, 81662.35, 80375.43, 
    90131.15,
  99917.58, 99887.63, 97699.77, 92719.24, 90064.66, 88292.05, 87092.29, 
    87440.96, 82747.42, 80099.71, 79350.24, 80022.12, 82136.87, 81176.52, 
    91423.61,
  91236.12, 87741.13, 92510.22, 91262.7, 84996.97, 83965.66, 86190.93, 
    85558.59, 80820.12, 78690.23, 77844.06, 78536.38, 79865.03, 81407.36, 
    93320.8,
  85331.73, 85376.42, 84502.56, 82887.73, 82650.35, 81270.53, 82122.74, 
    82450.14, 80266.59, 79087.82, 78749.99, 80227.05, 79961.82, 81848.42, 
    87634.9,
  86826.88, 85913.3, 86903.34, 86083.03, 85939.8, 84391.35, 83410.52, 
    82972.95, 82085.81, 84000.02, 98475.78, 99067.13, 89647.69, 89945.33, 
    82976.83,
  87247.91, 85482.45, 87842.29, 88633.98, 87739.92, 87318.36, 86612.54, 
    87011.8, 88548.41, 99170.66, 100078.8, 100041, 99809.61, 92128.08, 
    77619.66,
  86513.33, 85752.15, 87769.4, 88967.39, 88722.7, 88746.89, 88655.05, 
    90583.99, 94456.2, 99946.2, 99861.88, 99927.3, 99810.55, 86277.99, 77312.2,
  90222.62, 86991.88, 87431.88, 89155.23, 88796.52, 87800.77, 88399.66, 
    90194.39, 94300.02, 99966.52, 99928.5, 100019.6, 99885.72, 85126.78, 
    86870.63,
  93156.34, 88899.45, 87978.12, 89047.74, 88242.65, 85926.2, 87175.69, 
    89712.53, 99563.94, 99996.67, 99941.59, 99960.19, 99937.55, 92360.85, 
    95003.92,
  96255.48, 91693.59, 90117.58, 92423.35, 92635.09, 92762.48, 93683.74, 
    99496.65, 99996.5, 99978.99, 99969.31, 99948.66, 99958.84, 97764.51, 
    98864.32,
  100574, 100259.3, 96396.79, 93899.82, 93813.94, 92731.27, 90447.48, 
    90883.41, 85284.79, 80796.42, 78612.89, 78981.84, 81875.95, 80597.02, 
    90420.44,
  100516, 100370.7, 98199.29, 93165.66, 90396.57, 88517.82, 87233.73, 
    87548.77, 82776.84, 80160.85, 79429.81, 80140.4, 82331.44, 81371.56, 
    91703.98,
  91617.66, 88250.75, 93008.78, 91633.12, 85264.36, 84213.69, 86385.31, 
    85676.52, 80895.76, 78774.28, 77962.38, 78686.26, 80081.97, 81626.43, 
    93631.64,
  85816.88, 85990.37, 84976.27, 83328.45, 83032.09, 81553.48, 82348.95, 
    82643.47, 80384.88, 79186.88, 78852.2, 80348.06, 80155.36, 82078.32, 
    87949.04,
  87397.65, 86474, 87442.16, 86618.12, 86408.08, 84783.37, 83744.01, 83231.1, 
    82255.41, 84276.66, 98980.74, 99521.34, 89922.31, 90225.46, 83253.47,
  87820.58, 86014.66, 88395.55, 89176.26, 88241.29, 87774.34, 87048.84, 
    87393.11, 88974.65, 99682.87, 100435.4, 100453.9, 100195.7, 92439.42, 
    77897.26,
  87071.98, 86271.37, 88311.54, 89515.09, 89235.98, 89238.3, 89121.08, 
    91067.68, 94955.29, 100430.6, 100263.4, 100342.5, 100171.3, 86520.99, 
    77599.52,
  90798.99, 87534.71, 87953.02, 89714.55, 89355.41, 88336.59, 88911.57, 
    90698.16, 94853.19, 100507.2, 100402.9, 100417.9, 100272.3, 85391.99, 
    87224.26,
  93738.09, 89457.72, 88549.7, 89590.97, 88749.57, 86426.91, 87657.02, 
    90245.38, 100131.4, 100530.7, 100451.2, 100397.3, 100359.9, 92739.77, 
    95419.19,
  96878.02, 92292.31, 90734.61, 93030.47, 93239.61, 93417.1, 94274.82, 
    100109.5, 100577.2, 100549.5, 100507.9, 100440.2, 100439, 98204.95, 
    99334.45,
  101435.5, 101131.4, 97250.41, 94733.55, 94680.11, 93653.59, 91316.91, 
    91853.72, 86082.91, 81547.77, 79260.18, 79553.32, 82379.9, 80997.88, 
    90845.68,
  101392.1, 101319.9, 99129.8, 94047.9, 91251.09, 89368.5, 88117.91, 88415.7, 
    83570.84, 80914.45, 80111.7, 80808.48, 82927.46, 81872.16, 92256.8,
  92435.38, 89078.33, 93848.66, 92461.73, 86128.61, 85066.68, 87282.88, 
    86544.14, 81726.55, 79559.67, 78622.64, 79321.26, 80610.22, 82136.41, 
    94187.7,
  86610.04, 86765.41, 85821.94, 84193.08, 83914.91, 82391.93, 83232.1, 
    83495.98, 81216.39, 79907.84, 79626.24, 81131.91, 80696.75, 82651.21, 
    88379.94,
  88154.45, 87222.9, 88238.12, 87439.89, 87279.8, 85662.32, 84623.08, 
    84100.4, 83115.38, 85218.76, 100048.6, 100572.9, 90774.36, 91104.67, 
    83661.95,
  88526.62, 86746.06, 89199.03, 89995.26, 89106.45, 88660.94, 87924.86, 
    88303.81, 89904.27, 100710.3, 101438.8, 101393.6, 101197.2, 93219.66, 
    78272.33,
  87710.7, 86975.62, 89064, 90280.77, 90091.16, 90094.9, 90009.75, 91940.89, 
    95850.84, 101432.3, 101358, 101294.4, 101203.3, 87165.76, 78048.66,
  91344.06, 88196.7, 88691.8, 90438.23, 90153.86, 89142.4, 89751.83, 
    91494.42, 95711.56, 101408.9, 101353.6, 101306, 101192.6, 85953.91, 
    87914.42,
  94226.39, 90074.45, 89219.29, 90313.91, 89511.64, 87201.6, 88433.84, 
    91019.73, 100945.7, 101400.4, 101331.6, 101281.1, 101200.3, 93486.12, 
    96089.55,
  97316.22, 92819.48, 91323.67, 93665.69, 93905.21, 94103.25, 95010.38, 
    100835, 101380.7, 101368.2, 101325.9, 101272.1, 101212.9, 98957.48, 
    100000.9,
  101607.6, 101282.1, 97450.21, 95046.57, 95006.4, 93974.97, 91665.37, 
    92201.48, 86445.95, 81935.59, 79662.45, 79977.65, 82876.6, 81471.45, 
    91477.88,
  101554, 101565.8, 99356.39, 94328.39, 91594, 89771.71, 88556.35, 88840.88, 
    83964.94, 81341.73, 80557.48, 81241.74, 83397.59, 82294.36, 92907.64,
  92788.61, 89364.04, 94186.12, 92824.16, 86515.86, 85485.63, 87694.87, 
    86946.98, 82168.87, 79995.41, 79041.98, 79738.14, 81086.46, 82643.95, 
    94893.23,
  86837.33, 86912.07, 86114.05, 84502.58, 84250.85, 82795.76, 83630.23, 
    83935.16, 81688.6, 80376.33, 80108.14, 81607.44, 81163.49, 83185.87, 
    88988.81,
  88411.32, 87350.44, 88386.82, 87622.42, 87515.03, 85986.97, 84969.59, 
    84484.18, 83504.4, 85571.43, 100223.1, 100806.6, 91234.26, 91600.93, 
    84261.16,
  88668.89, 86891.05, 89271.54, 90116.06, 89271.62, 88879.7, 88195.07, 
    88609.7, 90160.61, 100836.6, 101759.8, 101762.3, 101608.5, 93691.24, 
    78810.94,
  87715.87, 87042.09, 89119.47, 90362.69, 90194.89, 90253.3, 90217.47, 
    92131.66, 95947.07, 101586.6, 101645.4, 101686.9, 101687.3, 87705.48, 
    78600.91,
  91218.73, 88180.2, 88677.96, 90455.17, 90183.95, 89254.27, 89886.52, 
    91668.15, 95763.58, 101512.8, 101591.9, 101719.2, 101677.9, 86514.41, 
    88458.51,
  94030.19, 89978.28, 89172, 90273.14, 89559.82, 87338.11, 88598.24, 
    91108.76, 100860.8, 101456.9, 101534.8, 101643, 101660.3, 93995.95, 
    96583.47,
  97068.41, 92646.66, 91147.69, 93514.6, 93808.91, 93972.94, 94914.2, 
    100670.1, 101272.3, 101383.6, 101484.9, 101576.3, 101642.8, 99445.8, 
    100534.1,
  101230.6, 100966.2, 97332.42, 94996.48, 94977.27, 93988.32, 91690.23, 
    92234.48, 86495.7, 82068.53, 79836.66, 80165.34, 83061.51, 81625.66, 
    91658.3,
  101157.4, 101262.1, 99083.28, 94211.91, 91598.6, 89823.47, 88617.12, 
    88915.85, 84094.78, 81528.33, 80718.11, 81424.27, 83572.98, 82462.73, 
    93078.45,
  92662.68, 89338.21, 94115.66, 92829.41, 86578.26, 85580.94, 87789.23, 
    87069.78, 82323.29, 80170.32, 79198.74, 79936.77, 81259.13, 82848.16, 
    95019.84,
  86746.77, 86815.02, 86101.68, 84522.51, 84301.83, 82893.84, 83737.27, 
    84053.3, 81830.12, 80565.39, 80309.71, 81826.08, 81326.84, 83378.8, 
    89163.33,
  88267.4, 87230.55, 88360.36, 87581.25, 87509.86, 86008.94, 85055.5, 
    84608.29, 83669.09, 85663.85, 100157.2, 100669.9, 91273.52, 91703.77, 
    84401.13,
  88508.32, 86739.17, 89176.39, 90049.34, 89260.93, 88876.3, 88219.8, 
    88634.78, 90195.27, 100728.4, 101608.8, 101611, 101497.6, 93694.09, 
    79080.45,
  87558.89, 86900.09, 89006.39, 90299.12, 90169.79, 90251.95, 90225.23, 
    92138.44, 95965.17, 101472.1, 101518.2, 101547.6, 101605.3, 87799.96, 
    78871.83,
  91005.27, 87991.12, 88532.3, 90353.82, 90140.27, 89239.85, 89889.77, 
    91695.04, 95765.19, 101411.2, 101495.9, 101595.9, 101587.9, 86644.27, 
    88667.35,
  93870.86, 89815.2, 89037.75, 90157.67, 89495.93, 87320.98, 88616.15, 
    91112.84, 100797.9, 101357, 101440.4, 101547.8, 101603.3, 94038.48, 
    96675.64,
  96969.95, 92529.05, 91038.53, 93426.83, 93723.92, 93889.45, 94844.98, 
    100598.1, 101209.6, 101259.7, 101390.4, 101489.5, 101602.7, 99448.54, 
    100619,
  101119.7, 100809.1, 97189.12, 94881.49, 94885.83, 93917.41, 91679.7, 
    92220.89, 86556.87, 82197.33, 80000.76, 80373.68, 83266.82, 81869.95, 
    91913.56,
  101037.5, 101099.1, 98915.53, 94128.48, 91562.06, 89799.59, 88609.31, 
    88931.8, 84194.73, 81662.73, 80866.53, 81614.41, 83748.13, 82698.16, 
    93257.13,
  92648.91, 89334.9, 94067.5, 92760.19, 86582.68, 85634.84, 87828.12, 
    87123.38, 82410.54, 80319.88, 79407.36, 80172.34, 81483.96, 83082.91, 
    95216.22,
  86747.02, 86793.94, 86078.2, 84568.74, 84343.9, 82966.7, 83815.21, 
    84145.38, 81931.7, 80716.02, 80403.2, 81938.06, 81544.68, 83587.27, 
    89400.05,
  88294.52, 87236.95, 88351.31, 87574.01, 87521.18, 86048.18, 85120.33, 
    84709.16, 83766.6, 85767.96, 100195.7, 100660, 91302.3, 91800.54, 84617.86,
  88522.28, 86764.16, 89162.93, 90005.38, 89230.17, 88868.38, 88254.72, 
    88682.96, 90237.19, 100740.9, 101570.7, 101581.7, 101471.2, 93764.2, 
    79342.56,
  87656.45, 86958.19, 89017.95, 90268.93, 90113.48, 90223.6, 90226.18, 
    92170.16, 95988.62, 101478.6, 101516.6, 101547.3, 101557.4, 87949.62, 
    79115.17,
  91284.97, 88165.38, 88620.84, 90423.28, 90134.22, 89236.2, 89894.97, 
    91732.65, 95800.45, 101456.2, 101504.1, 101598.9, 101559, 86812.94, 
    88802.78,
  94275.44, 90086.99, 89207.95, 90300.77, 89589.55, 87398.39, 88696.98, 
    91208.24, 100835.8, 101432.5, 101478.5, 101572.2, 101609.4, 94105.59, 
    96744.91,
  97425.81, 92842.59, 91274.78, 93605.94, 93876.87, 93976.54, 94947.51, 
    100678.9, 101326.4, 101370.8, 101454.1, 101540.1, 101628.6, 99475.03, 
    100657.3,
  101232, 100858.6, 97168.55, 94855.8, 94882.02, 93930, 91720.78, 92251.93, 
    86585.76, 82226.43, 80053.46, 80440.3, 83351.15, 81933, 91994.87,
  101073.6, 101102.3, 98909.77, 94104.59, 91572.99, 89835.35, 88660.9, 
    88984.78, 84242.05, 81706.43, 80905.37, 81653.2, 83793.1, 82749.89, 
    93290.94,
  92693.02, 89335.47, 94054.64, 92745.75, 86611.76, 85659.85, 87860.38, 
    87186.41, 82457.14, 80362.69, 79469.01, 80231.83, 81551.59, 83139.52, 
    95236.8,
  86898.71, 86912.95, 86119.98, 84600.14, 84400.45, 83024.45, 83864, 
    84201.41, 81986.87, 80769.6, 80432.44, 81972.98, 81594, 83627.54, 89443.9,
  88452.48, 87433.84, 88437.55, 87662.09, 87603.72, 86131.11, 85186.69, 
    84744.58, 83805.2, 85829.28, 100390.4, 100843.6, 91405.41, 91833.48, 
    84683.74,
  88751.71, 86994.16, 89399.2, 90204.24, 89370.16, 89017.81, 88386.39, 
    88790.83, 90424.36, 101013.6, 101762.3, 101726.4, 101576.8, 93801.74, 
    79408.95,
  87972.02, 87301.88, 89360.26, 90588.39, 90347.62, 90410.38, 90417.61, 
    92390.91, 96314.66, 101785.7, 101683.1, 101626.9, 101589.2, 87992.91, 
    79166.76,
  91682.38, 88558.91, 89052.3, 90790.57, 90441.02, 89504.51, 90153.13, 
    92029.12, 96191.98, 101767.6, 101670.2, 101666.1, 101551.7, 86844.91, 
    88800.09,
  94716.39, 90522.23, 89687.8, 90792, 89968.77, 87686.22, 88993.58, 91613.86, 
    101425.7, 101810.8, 101678.1, 101631.9, 101608.8, 94093.93, 96696.84,
  97877.01, 93375.13, 91846.78, 94239.54, 94537.98, 94668.62, 95592.05, 
    101438.9, 101946.4, 101805.1, 101700.6, 101616.9, 101641.2, 99467.55, 
    100547.8,
  101218.3, 100884.6, 97122.95, 94753.64, 94758.52, 93832.07, 91630.09, 
    92173.79, 86522.28, 82170.6, 79984.11, 80343.37, 83239.9, 81820.19, 
    91832.25,
  101065.8, 101101.8, 98870.93, 94020.36, 91484.68, 89740.95, 88565.8, 
    88902.23, 84180.7, 81621.16, 80833.73, 81565.3, 83722.23, 82681.84, 
    93161.77,
  92690.09, 89200.62, 93996.95, 92681.98, 86526.83, 85552.2, 87759.91, 
    87084.3, 82373.73, 80288.2, 79424.23, 80166.82, 81484.37, 83054.5, 
    95088.66,
  86828.54, 86785.22, 86017.64, 84480.95, 84271.51, 82897.84, 83770.26, 
    84098.78, 81911.23, 80691.58, 80353.2, 81902.75, 81564.7, 83560.59, 
    89342.61,
  88332.44, 87355.35, 88349.39, 87557.61, 87513.06, 86025.72, 85087.89, 
    84661.56, 83722.41, 85742.23, 100582.7, 101031.5, 91452.98, 91828.62, 
    84614.02,
  88588.69, 86884.3, 89319.54, 90141.13, 89315.98, 88950.09, 88311.49, 
    88751.09, 90449.05, 101272.8, 102068.7, 102046, 101851.3, 93916.41, 
    79319.59,
  87858.85, 87196.52, 89283.74, 90526.72, 90332.7, 90437.05, 90461.85, 
    92489.31, 96505.88, 102036.8, 101895.7, 101885.6, 101841.6, 87980.58, 
    79093.12,
  91540.01, 88433.02, 88947.88, 90728.61, 90449.95, 89557.58, 90230.67, 
    92110.38, 96366.37, 102044.8, 101911.4, 101914.7, 101829.2, 86864.97, 
    88818.09,
  94591.48, 90425.94, 89627.22, 90710.45, 89896.73, 87654.58, 89013.26, 
    91670.13, 101686.8, 102083.1, 101948, 101875.7, 101858.8, 94193.11, 
    96844.32,
  97808.7, 93309.55, 91857.93, 94252.43, 94525.98, 94668.83, 95674.61, 
    101637.7, 102236.3, 102137.6, 102055.3, 101954.1, 101922.7, 99662.68, 
    100760.7,
  101098.5, 100719, 96904.28, 94558.78, 94554.62, 93632.07, 91417.06, 
    91927.04, 86317.37, 81922.24, 79743.34, 80066.23, 82998.57, 81594.55, 
    91538.1,
  100883.8, 100903.8, 98702.37, 93826.48, 91272.38, 89530.74, 88329.84, 
    88662.49, 83959.67, 81382.8, 80626.63, 81286.12, 83462.02, 82424.44, 
    92862.38,
  92433.94, 88982.45, 93737.23, 92443.85, 86289.18, 85294.65, 87526.87, 
    86858.04, 82145.77, 80016.91, 79191.59, 79904.76, 81238.78, 82776.7, 
    94792.27,
  86483.6, 86556.2, 85753.6, 84204.63, 84017.12, 82644.98, 83520.53, 
    83842.23, 81663.95, 80486.24, 80133.11, 81635.36, 81337.04, 83272.26, 
    89057.93,
  88045.57, 87094.76, 88098.62, 87274.61, 87216.53, 85760.13, 84835.05, 
    84419.31, 83491.09, 85455.16, 100218.1, 100741.2, 91134.02, 91525.42, 
    84365.77,
  88367.6, 86696.7, 89130.13, 89913.28, 89043.38, 88667.99, 88035.05, 
    88498.39, 90175.42, 100999.4, 101784.2, 101754.4, 101511.7, 93622.1, 
    79066.06,
  87697.02, 86990.93, 89078.69, 90314.69, 90131.75, 90224.45, 90237.38, 
    92248.76, 96222.33, 101740.6, 101572.1, 101619.8, 101491.3, 87772.41, 
    78827.74,
  91368.7, 88265.15, 88788.49, 90550.56, 90227.65, 89305.99, 89981.99, 
    91852.76, 96083.92, 101755.9, 101644.4, 101697.4, 101543.3, 86636.98, 
    88451.62,
  94419.7, 90253.01, 89465.7, 90547.97, 89729.67, 87464.04, 88793.14, 
    91451.23, 101414.8, 101798.9, 101695.8, 101663.9, 101587.9, 93987.07, 
    96652.93,
  97604.74, 93089.98, 91688.31, 94073.02, 94336.72, 94474.66, 95454.47, 
    101363.6, 101908.6, 101858.5, 101791.9, 101737.1, 101687.7, 99478.03, 
    100569,
  101140.4, 100801.7, 96903.22, 94413.54, 94392.49, 93409.09, 91194.1, 
    91711.27, 86126.78, 81758.95, 79589.49, 79907.02, 82790.35, 81407.48, 
    91281.51,
  100918.6, 100905.3, 98681.02, 93699.03, 91098.88, 89327.58, 88123.25, 
    88466.4, 83765.05, 81187.8, 80435.3, 81121.84, 83280.88, 82237.45, 92580.2,
  92239.52, 88891.84, 93677.09, 92315.15, 86116.61, 85128.5, 87337.73, 
    86658.76, 81960.4, 79857.21, 79028.2, 79721.79, 81065.99, 82605.03, 
    94533.16,
  86360.96, 86407.91, 85571.02, 84100.21, 83877.81, 82493.83, 83372.48, 
    83694.93, 81503.07, 80311.91, 79995.73, 81493.85, 81162.48, 83106.99, 
    88836.99,
  87864.2, 86980.55, 87976.94, 87205.74, 87128.67, 85642.16, 84701.67, 
    84272.34, 83373.16, 85408.84, 100208, 100720.3, 91076.22, 91423.13, 
    84210.48,
  88302.35, 86593.04, 89010.02, 89812.86, 88991.63, 88643.53, 88025.43, 
    88473.89, 90141.66, 100923.7, 101658.1, 101639.9, 101457.1, 93516.05, 
    78868.48,
  87578.11, 86886.84, 89003.45, 90231.36, 90070.23, 90159.41, 90169.77, 
    92177.24, 96126.91, 101617.1, 101492.3, 101536.2, 101448.6, 87633.08, 
    78654.73,
  91248.79, 88164.75, 88672.09, 90461.88, 90170.18, 89271.77, 89952.21, 
    91802.37, 96027.75, 101661.3, 101575.3, 101608.4, 101468.9, 86470.46, 
    88412.91,
  94271.05, 90138.67, 89343.18, 90438.34, 89651.85, 87420.62, 88748.49, 
    91399.62, 101294.9, 101703.6, 101615.5, 101597.9, 101473.2, 93940.33, 
    96576.27,
  97439.34, 92969.16, 91581.43, 93957.66, 94212.2, 94366.89, 95395.18, 
    101266.2, 101791.4, 101761.9, 101711.5, 101697.7, 101629.9, 99430.55, 
    100491.4,
  101175, 100840.2, 96949.84, 94363.99, 94275.77, 93250.58, 91025.4, 
    91463.98, 85933.92, 81580.75, 79448.62, 79806.62, 82740.23, 81392.39, 
    91339.73,
  101016.5, 100968.3, 98716.15, 93682.68, 90963.09, 89140.38, 87913.19, 
    88230.73, 83560.72, 81004.4, 80305.75, 80986.68, 83184.52, 82167.73, 
    92608.8,
  92216.74, 88852.52, 93640.08, 92206.98, 85952.2, 84964.02, 87161.61, 
    86470.62, 81774.81, 79701.57, 78894.3, 79604.58, 80980.8, 82525.18, 
    94540.22,
  86313.77, 86375.58, 85494.45, 83994.24, 83738.14, 82339.07, 83191.52, 
    83505.16, 81309.05, 80140.17, 79845.44, 81336.36, 81051.41, 83004.83, 
    88856.37,
  87879.12, 86997.78, 87966.96, 87175.51, 87081.65, 85550.34, 84595.88, 
    84165.48, 83255.45, 85312.92, 100083.2, 100540.6, 90916.26, 91317.94, 
    84160.57,
  88259.16, 86548.65, 88982.64, 89808.2, 88989.98, 88604.1, 87958.98, 
    88359.2, 90058.16, 100729.4, 101464.2, 101454.9, 101320.8, 93357.73, 
    78809.98,
  87544.64, 86842.44, 88942.95, 90169.81, 90015.7, 90086.93, 90103.44, 
    92068.71, 96005.3, 101432.7, 101353.8, 101383.9, 101366.6, 87507.91, 
    78636.78,
  91202.14, 88111.27, 88641.03, 90429.17, 90153.15, 89237.39, 89888.92, 
    91697.25, 95934.09, 101514, 101434.5, 101429.5, 101249.4, 86368.95, 
    88433.54,
  94218.82, 90077.4, 89280.46, 90374.04, 89600.4, 87368.93, 88677.79, 
    91336.22, 101164.5, 101590.4, 101506.4, 101491.6, 101375.1, 93897.86, 
    96550.5,
  97360.77, 92911.91, 91523.52, 93875.07, 94127.62, 94280.98, 95303.45, 
    101136.4, 101672, 101663.3, 101610.9, 101584.4, 101501.6, 99314.45, 
    100420.1,
  101107.7, 100791.9, 96928.23, 94407.15, 94278.5, 93203.33, 90950.02, 
    91390.19, 85865.68, 81442.27, 79254.72, 79584.85, 82399.02, 81148.24, 
    91051.9,
  101001.4, 100980.9, 98714.54, 93669, 90915.02, 89022.5, 87780.5, 88071.42, 
    83389.46, 80789.62, 80056.18, 80750.05, 82885.91, 81908.27, 92298.78,
  92143.39, 88766.82, 93596.09, 92223.49, 85879.03, 84825.07, 86993.96, 
    86302.12, 81571.19, 79461.42, 78637.52, 79336.42, 80681.7, 82215.88, 
    94196.59,
  86204.38, 86378.43, 85432.8, 83841.21, 83578.18, 82139.39, 82996.41, 
    83268.5, 81049.43, 79856.21, 79535.37, 81021.12, 80763.4, 82670.87, 
    88542.98,
  87804.2, 86899.56, 87880.3, 87115.18, 87029.15, 85471.43, 84480.12, 
    84006.4, 83045.54, 85032.88, 99685.71, 100204.4, 90594.13, 90878.32, 
    83864.06,
  88211.15, 86460.21, 88902.04, 89680.02, 88853.8, 88447.83, 87766.03, 
    88136.27, 89732.44, 100411.4, 101151, 101133, 100920, 93053.62, 78516.98,
  87451.97, 86721.05, 88856.42, 90073.71, 89913.45, 89961.9, 89940.81, 
    91870.48, 95704.93, 101047.3, 100906.4, 100936.8, 100878.4, 87184.2, 
    78306.67,
  91087.69, 87991.22, 88504.73, 90273.38, 89979.31, 89021.77, 89654.88, 
    91389.94, 95598.88, 101075.9, 100938.7, 100941, 100897.3, 86019.39, 
    87915.71,
  94039.71, 89933.55, 89118.36, 90207.48, 89417.26, 87166.08, 88436.34, 
    91083.42, 100832.1, 101154.9, 100982, 100905.1, 100848.9, 93371.7, 
    96058.17,
  97148.98, 92718.7, 91309.41, 93644.31, 93892.8, 94055.13, 95028.69, 
    100817.3, 101325, 101277.2, 101137.8, 101051, 100960.9, 98815.23, 99939.34,
  101229.1, 100899.2, 97063.84, 94574.34, 94482.31, 93408.99, 91156.49, 
    91594.84, 86027.27, 81576.45, 79365.34, 79670.23, 82444.63, 81075.51, 
    90800.77,
  101183.2, 101168.2, 98885.42, 93814.91, 91077.77, 89207.45, 87983.37, 
    88265.34, 83557.16, 80940.11, 80181.51, 80860.72, 82969.88, 81936.54, 
    92162.73,
  92288.69, 88892.33, 93769.57, 92396.45, 85993.02, 84972.24, 87154.75, 
    86446.8, 81707.55, 79591.79, 78739.56, 79437.29, 80737.38, 82256.98, 
    94149.52,
  86356.58, 86491.3, 85545.55, 83969.16, 83741.64, 82242.16, 83104.76, 
    83429.62, 81205.59, 79987.68, 79656.6, 81149.78, 80827.6, 82766.47, 
    88475.66,
  87919.3, 86996.79, 87986.37, 87171.29, 87055.64, 85516.36, 84522.41, 
    84011.85, 83063.51, 85123.46, 99803.25, 100363.4, 90722.59, 91059.34, 
    83836.78,
  88296.01, 86518.92, 88955.85, 89758.35, 88914.5, 88497.74, 87823.19, 
    88205.42, 89837.32, 100526.7, 101244.6, 101239.8, 101032.2, 93224.44, 
    78491.75,
  87505.02, 86777.75, 88863.62, 90093.62, 89914.02, 89947.96, 89916.83, 
    91838.88, 95737.22, 101187, 101048.9, 101077.6, 100999.6, 87309.55, 
    78237.18,
  91125.51, 88027.98, 88514.25, 90266.24, 89991.27, 89040.34, 89670.61, 
    91432.89, 95645.32, 101187.2, 101062.1, 101099.6, 100994.6, 86078.45, 
    87880.32,
  94039.84, 89937.68, 89106.12, 90180.91, 89383.93, 87125.2, 88379.63, 
    90960.8, 100830, 101202.1, 101065.1, 101047.4, 101022.8, 93467.21, 
    96038.79,
  97130.56, 92694.34, 91258.77, 93583.13, 93837.9, 94005.86, 94962.33, 
    100781.7, 101293.7, 101240.5, 101120.1, 101048.5, 101034.9, 98847.55, 
    99948.29,
  101376.3, 101036.5, 97167.45, 94676.34, 94575.34, 93522.27, 91250.15, 
    91744.18, 86140.05, 81706.62, 79495.39, 79795.85, 82602.73, 81225.49, 
    91044.23,
  101342.2, 101307.5, 99046.99, 93978.78, 91203.64, 89365.48, 88125.7, 
    88429.26, 83684.8, 81088.34, 80319.76, 81005.93, 83121.09, 82062.68, 
    92436.56,
  92413.8, 89013.65, 93900.12, 92542.82, 86159.73, 85162.09, 87322.65, 
    86611.65, 81873.77, 79782.46, 78911.75, 79624.16, 80924.16, 82451.91, 
    94446.38,
  86569.92, 86745.31, 85766.52, 84141.34, 83931.21, 82481.84, 83353, 
    83655.24, 81417.74, 80184.19, 79867.5, 81416.46, 80987.21, 83003.77, 
    88728.27,
  88137.76, 87251.02, 88243.45, 87435.59, 87294.38, 85715.21, 84731.88, 
    84239.45, 83300.75, 85443.38, 100233.7, 100719.8, 91047.73, 91432.09, 
    84005.61,
  88524.91, 86759.63, 89189.59, 89987.02, 89147.23, 88738.38, 88068.92, 
    88470.09, 90151, 100840.3, 101574.9, 101553.8, 101415.6, 93478.05, 
    78653.05,
  87760.13, 87022.38, 89107.82, 90326.31, 90153.59, 90182.63, 90173.44, 
    92103.24, 96048.3, 101532.8, 101510.4, 101481.2, 101507.6, 87455.41, 
    78527.38,
  91379.3, 88256.16, 88746.27, 90501.48, 90229.3, 89275.3, 89942.64, 91697.4, 
    95949.94, 101566.6, 101517.1, 101533.2, 101429.3, 86309.86, 88406.04,
  94296.23, 90177.3, 89329.66, 90406.38, 89626.83, 87375.8, 88661.15, 
    91256.95, 101153, 101585.6, 101509.9, 101522.4, 101442.8, 93905.05, 
    96465.98,
  97353.51, 92884.52, 91448.27, 93779.25, 94046.81, 94198.46, 95177.99, 
    101048, 101623.4, 101617.8, 101564.2, 101545.5, 101482.8, 99297.74, 
    100382.5,
  101360.8, 100996.3, 97152.62, 94666.05, 94513.69, 93428.48, 91197.45, 
    91727.27, 86128.56, 81714.01, 79511.02, 79845.34, 82742.59, 81373.69, 
    91297.01,
  101289.1, 101235.1, 99029.69, 93947.78, 91200.01, 89354.55, 88109.74, 
    88425.84, 83704.38, 81136.04, 80356.93, 81057.35, 83240.24, 82202.24, 
    92730.3,
  92417, 89047.72, 93896.88, 92530.45, 86161.37, 85169.35, 87340.72, 
    86640.08, 81912.44, 79829.14, 78964.64, 79690.03, 81004.41, 82574.66, 
    94729.8,
  86621.11, 86789.6, 85823.85, 84205.44, 83952.34, 82521.85, 83377.19, 
    83678.98, 81453.24, 80239.51, 79906.62, 81478.2, 81088.67, 83156.1, 
    88959.98,
  88183.27, 87287.28, 88284.72, 87460.75, 87321.56, 85750.89, 84751.62, 
    84269.54, 83330.02, 85419, 100203.3, 100661, 91029.64, 91514.54, 84119.73,
  88584.66, 86829.38, 89243.12, 90025.49, 89172.78, 88757.34, 88090.03, 
    88467.76, 90109.98, 100818, 101601.7, 101585.4, 101515.7, 93456.7, 
    78922.56,
  87848.51, 87098.77, 89168.41, 90363.16, 90180.32, 90209.39, 90187.32, 
    92103.37, 96039.44, 101523.9, 101519.7, 101513.1, 101560.9, 87535.34, 
    78772.63,
  91503.36, 88346.89, 88815.77, 90565.4, 90266.66, 89305.7, 89938.39, 
    91692.43, 95910.92, 101552.5, 101524.2, 101592.2, 101441.7, 86551.73, 
    88611.08,
  94426.14, 90255.12, 89402.47, 90474.61, 89696.23, 87424.68, 88678.02, 
    91264.04, 101114.8, 101581.1, 101529.7, 101583.2, 101471.2, 93986.34, 
    96700.06,
  97479.7, 92993.3, 91510.83, 93818.84, 94063.03, 94205.75, 95120.4, 
    100974.7, 101595.1, 101618.9, 101594.3, 101621.5, 101605.7, 99484.34, 
    100646.7,
  101138, 100788.2, 96977.37, 94477.88, 94374, 93280.12, 91003.01, 91502.7, 
    85947.83, 81551.39, 79355.85, 79653.98, 82586.54, 81220.84, 91185.36,
  101041.6, 100980.6, 98808.34, 93773.38, 91042.43, 89207.44, 87941.07, 
    88225.65, 83525.41, 80951.77, 80174.85, 80882.89, 83054.15, 82032.16, 
    92550.08,
  92284.49, 88928.89, 93674.96, 92310.23, 86021.62, 85019.28, 87185.17, 
    86469.89, 81733.06, 79626.22, 78766.16, 79484.16, 80824.29, 82390.77, 
    94535.77,
  86499.32, 86670.88, 85722.82, 84092.3, 83830.44, 82377.78, 83195.17, 
    83496.42, 81272.69, 80051.12, 79701.62, 81221.49, 80903.62, 82895.42, 
    88759.66,
  88081.72, 87163.96, 88167.93, 87357.89, 87214.73, 85632.93, 84599.95, 
    84100.45, 83130.86, 85149.07, 99873.46, 100335.2, 90745.62, 91176.49, 
    83990.62,
  88481.16, 86716.53, 89112.41, 89889.58, 89021.71, 88604.72, 87914.18, 
    88276.98, 89869.34, 100534.2, 101263.4, 101241, 101056.6, 93195.38, 
    78664.46,
  87758.66, 87000.83, 89050.1, 90244.87, 90041.5, 90024.59, 89983.12, 
    91862.84, 95725.1, 101216.1, 101170.5, 101170.2, 101064.9, 87347.38, 
    78500.89,
  91441.22, 88252.77, 88725.12, 90457.3, 90130.04, 89149.34, 89751.29, 
    91483.76, 95606.38, 101244.8, 101210.9, 101223.8, 101099.6, 86214.65, 
    88159.1,
  94377.74, 90174.75, 89312.07, 90375.89, 89555.7, 87257.79, 88488.78, 
    91047.91, 100809.5, 101237.1, 101190.8, 101179.5, 101162.3, 93564.28, 
    96232.91,
  97470.38, 92977.15, 91469.3, 93788.3, 94037.03, 94203.36, 95102.75, 
    100808.8, 101281.9, 101235.8, 101189.4, 101166.2, 101176.5, 98979.91, 
    100119,
  101008.9, 100669.7, 96876.7, 94398.72, 94289.79, 93267.27, 91007.02, 
    91482.36, 85893.8, 81462.67, 79270.14, 79570.59, 82449.19, 81085.43, 
    90971.73,
  100948.4, 100889.7, 98680.11, 93681.66, 90981.31, 89142.95, 87901.56, 
    88196.52, 83444.96, 80874.12, 80092.98, 80779.3, 82912.5, 81868.57, 
    92318.04,
  92228.66, 88861.22, 93636.9, 92246.66, 85965.51, 84964.26, 87146.71, 
    86413.98, 81665.94, 79572.59, 78703.42, 79401.21, 80705.02, 82235.4, 
    94347.47,
  86434.73, 86595.02, 85655.23, 84052.77, 83813, 82371.34, 83196.09, 
    83480.78, 81228.61, 80018.88, 79718.74, 81223.9, 80817.66, 82783.62, 
    88554.11,
  88017.5, 87159.41, 88154.83, 87356.77, 87224.58, 85644.04, 84643.25, 
    84148.19, 83189.76, 85272.7, 99984.35, 100436.5, 90839.59, 91183.55, 
    83803.24,
  88438.51, 86695.71, 89139.55, 89922.85, 89083.42, 88670.77, 87983.98, 
    88347.3, 89967.54, 100596.2, 101308, 101294.2, 101159.1, 93223.09, 
    78500.91,
  87741.91, 87021.91, 89124.27, 90315.76, 90125.23, 90134.62, 90104.01, 
    92001.61, 95858.4, 101297.3, 101259.3, 101223.9, 101189.8, 87252.65, 
    78369.57,
  91423.87, 88293.45, 88809.09, 90562.03, 90250.01, 89270.16, 89877.38, 
    91613.04, 95780.02, 101318.5, 101259.1, 101247.7, 101158.1, 86154.26, 
    88153.79,
  94422.97, 90255.13, 89442.06, 90521.23, 89702.41, 87425.92, 88662.62, 
    91269.22, 101003, 101341.3, 101252.3, 101224.4, 101151.2, 93587.02, 
    96164.85,
  97553.8, 93068.94, 91656.8, 94040.65, 94298.44, 94447.37, 95387.58, 
    101083.7, 101474.2, 101377.6, 101299.4, 101244.7, 101174.6, 98971.91, 
    100047.4,
  100995.4, 100685.9, 96851.57, 94366.45, 94282.55, 93274.84, 91036.79, 
    91508.38, 85918.95, 81496.51, 79299.82, 79594.27, 82461.68, 81107.84, 
    90997.71,
  101031.2, 100907.1, 98717.12, 93699.95, 91013.61, 89184.92, 87950.73, 
    88262.28, 83497.21, 80895.56, 80119.93, 80801.8, 82927.34, 81896.91, 
    92326.53,
  92212.5, 88892.22, 93652.19, 92276.72, 85992.95, 85003.51, 87190.08, 
    86451.73, 81685.79, 79615.17, 78740.12, 79454.87, 80767.35, 82276.05, 
    94399.96,
  86480.2, 86655.76, 85694.99, 84104.68, 83845.44, 82427.98, 83256.97, 
    83564.97, 81315.26, 80077.01, 79748.37, 81280.99, 80883.25, 82803.84, 
    88591.35,
  88011.96, 87170.06, 88168.42, 87381.36, 87231.78, 85655.1, 84664.88, 
    84178.92, 83193.91, 85293.88, 100071.9, 100519.6, 90891.41, 91229.45, 
    83822.42,
  88446.69, 86722.67, 89172.23, 89962.95, 89122.48, 88703.07, 88010.55, 
    88402.08, 90046.56, 100717.4, 101383, 101356.1, 101301.2, 93249.05, 
    78589.62,
  87694.51, 86985.05, 89109.27, 90325.14, 90143.32, 90166.65, 90133.72, 
    92046.49, 95948.62, 101407.9, 101315.5, 101256.4, 101242.1, 87323.12, 
    78442.49,
  91342.45, 88230.6, 88751.66, 90534.44, 90245.06, 89267.04, 89914.28, 
    91677.29, 95872.45, 101442.9, 101316.4, 101287.2, 101230.4, 86230.39, 
    88179.59,
  94300.89, 90160.88, 89362.63, 90460.74, 89662.35, 87402.42, 88655.72, 
    91277.14, 101122.2, 101472.6, 101348.6, 101276.3, 101187.5, 93619.43, 
    96320.2,
  97408.89, 92946.59, 91528.78, 93921.59, 94195.52, 94346.57, 95319.09, 
    101126.5, 101594.4, 101533.7, 101436.5, 101365.5, 101297.3, 99101.64, 
    100207.9,
  101046.8, 100708.4, 96894.34, 94384.28, 94320.85, 93294.45, 91010.64, 
    91492.99, 85866.45, 81481.59, 79293.43, 79634.73, 82509.12, 81148.46, 
    91025.33,
  101028.4, 100909.2, 98721.74, 93727.98, 91044.49, 89211.73, 87998.35, 
    88275.7, 83492.49, 80939.39, 80163.82, 80867.89, 82972.93, 81951.01, 
    92389.53,
  92292.18, 88959.06, 93671.89, 92296.72, 86076.56, 85073.14, 87231.09, 
    86475.38, 81749.62, 79672.7, 78784.04, 79514.28, 80804.92, 82369.57, 
    94406.21,
  86542.89, 86722.61, 85785.21, 84170.99, 83913.96, 82479.7, 83307.51, 
    83611.66, 81355.95, 80099.55, 79812.94, 81357.55, 80890.23, 82892.52, 
    88599.45,
  88091.43, 87199.87, 88205.21, 87409.93, 87280.59, 85728.73, 84721.39, 
    84231.24, 83257.95, 85413.98, 100145.2, 100617.9, 90964.36, 91330.65, 
    83922.36,
  88481.25, 86740.33, 89146.55, 89964.67, 89122.45, 88716.74, 88052.19, 
    88449.72, 90093.27, 100753.4, 101489.5, 101469.8, 101325.1, 93368.3, 
    78573.52,
  87690.79, 86976.14, 89034.73, 90294.66, 90123.3, 90180.17, 90126.28, 
    92054.98, 95986.83, 101492.8, 101427.3, 101369.8, 101357.3, 87375.9, 
    78449.86,
  91269.09, 88187.28, 88666.89, 90457.22, 90176.27, 89257.4, 89887.95, 
    91693.86, 95884.23, 101491.3, 101420.6, 101400.1, 101349.5, 86275.95, 
    88239.82,
  94146.48, 90069.27, 89228.48, 90341.49, 89593.15, 87348.05, 88613.43, 
    91202.46, 101119.1, 101502.2, 101415.4, 101371.1, 101317.9, 93665.52, 
    96308.41,
  97194.38, 92798.98, 91340.84, 93728.22, 93985.86, 94135.33, 95154.59, 
    101081.7, 101572.1, 101520.7, 101440.7, 101384.4, 101324.3, 99089.25, 
    100176,
  101213.8, 100855.1, 97079.73, 94571.62, 94484.66, 93443.25, 91153.04, 
    91615.71, 86000.01, 81651.33, 79484.82, 79840.99, 82718.95, 81382.06, 
    91328.59,
  101115, 101081.2, 98868.4, 93892.95, 91210.29, 89383.07, 88151.97, 
    88397.31, 83657.05, 81109.75, 80342.06, 81056.45, 83214.09, 82151.26, 
    92700.73,
  92522.22, 89116.06, 93860.49, 92481.3, 86265.61, 85221.44, 87390.24, 
    86634.09, 81898.94, 79815.94, 78962.92, 79691.78, 81008.32, 82569.04, 
    94709.7,
  86725.6, 86803.59, 85969.4, 84322.55, 84072.55, 82623.02, 83433.02, 
    83707.58, 81474.97, 80268, 79959.55, 81516.88, 81070.1, 83135.85, 88851.05,
  88297.3, 87247.4, 88308.3, 87505.16, 87379.55, 85839.88, 84828.2, 84352.76, 
    83376.87, 85451.9, 100166.2, 100664.4, 91073.87, 91512.8, 84100.95,
  88527.16, 86803.92, 89182.45, 90009.46, 89170.64, 88753.98, 88072.12, 
    88472.38, 90069.74, 100801.4, 101617, 101618.1, 101491.3, 93485.55, 
    78813.59,
  87687.34, 86988.01, 89035.28, 90292.79, 90113.75, 90175.89, 90133.11, 
    92056.3, 95978.92, 101531, 101498.8, 101515.3, 101536.7, 87572.3, 78679.08,
  91242.11, 88159.41, 88629.18, 90408.09, 90121.81, 89188.73, 89825.22, 
    91629.28, 95795.5, 101531.6, 101519.3, 101581.2, 101476.5, 86438.62, 
    88488.72,
  94116.97, 89996.32, 89141.05, 90229.72, 89506.7, 87292.51, 88571.52, 
    91079.21, 100948.6, 101510.3, 101491, 101529.3, 101502, 93907.52, 96541.16,
  97211.35, 92703.95, 91178.31, 93534.45, 93801.87, 93924.95, 94880.77, 
    100702, 101421.4, 101473, 101499.5, 101510.3, 101526.7, 99315.6, 100416.2,
  101272.9, 100908.4, 97152.59, 94703.73, 94603.74, 93581.73, 91317.66, 
    91751.13, 86184.3, 81782.3, 79606.79, 79983.66, 82911.88, 81574.91, 
    91501.14,
  101142.1, 101140.9, 98943.48, 94002.43, 91314.9, 89515.2, 88278.7, 
    88525.03, 83807.26, 81236.45, 80495.72, 81177.77, 83368.23, 82323.02, 
    92837.52,
  92648.32, 89140.62, 93902.23, 92583.94, 86357.59, 85314.45, 87489.34, 
    86766.97, 82030.62, 79910.51, 79089.95, 79785.07, 81140.25, 82688.59, 
    94824.29,
  86764.01, 86758.82, 85972.13, 84352.51, 84114.77, 82702.2, 83518.91, 
    83798.28, 81582.12, 80373.5, 80033.48, 81513.85, 81219.76, 83183.21, 
    89051.12,
  88290.85, 87236.26, 88282.79, 87473.73, 87339.88, 85826.1, 84845.36, 
    84388.74, 83455.37, 85411.8, 99921.08, 100487.8, 90942.84, 91385.58, 
    84324.82,
  88492.92, 86784.02, 89132.62, 89949.48, 89093.93, 88676.73, 88014.59, 
    88432.33, 89970.55, 100556.4, 101396.2, 101423.8, 101168.6, 93470.12, 
    78957.19,
  87690.59, 86996.54, 89012.94, 90248.32, 90050.53, 90091.6, 90043, 91957.47, 
    95760.02, 101301.3, 101261.8, 101351.3, 101202.9, 87658.98, 78732.73,
  91346.81, 88229.23, 88674.79, 90417.88, 90099.87, 89160.38, 89768.35, 
    91565.77, 95614.01, 101286.3, 101311.7, 101417.8, 101283.5, 86490.2, 
    88327.43,
  94295.23, 90112.55, 89224.4, 90299.57, 89539.56, 87275.61, 88532.14, 
    91018.38, 100724, 101268.4, 101293.8, 101353.1, 101338.7, 93783.28, 
    96409.79,
  97433.38, 92888.54, 91337.49, 93653.98, 93901.19, 94020.85, 94923.8, 
    100731.4, 101288.9, 101257, 101315.6, 101358.7, 101399.9, 99191.26, 
    100334.8,
  101244.6, 100874.6, 97125.68, 94679.74, 94593.54, 93544.91, 91320.22, 
    91759.23, 86191.99, 81782.48, 79589.98, 79931.3, 82841.46, 81515.18, 
    91378.27,
  101183.2, 101116.9, 98922.88, 93983.76, 91299.82, 89484.05, 88260.93, 
    88522.43, 83803.45, 81203.62, 80457.35, 81137.32, 83298.02, 82286.78, 
    92654.32,
  92592.73, 89137.9, 93871.75, 92521.4, 86313.78, 85306.48, 87465.17, 
    86767.66, 82033.95, 79912.45, 79077.23, 79762.9, 81079.77, 82613.56, 
    94684.02,
  86723.45, 86872.41, 86001.24, 84367.92, 84116.62, 82696.47, 83519.97, 
    83804.27, 81580.77, 80381.23, 80069.98, 81540.3, 81194.77, 83119.14, 
    88929.48,
  88248.45, 87365.98, 88364.46, 87578.25, 87425.47, 85892.69, 84883.62, 
    84420.02, 83480.58, 85486.02, 100084, 100558.5, 91082.36, 91368.5, 
    84250.87,
  88607.55, 86908.07, 89307.58, 90137.64, 89272.66, 88828.42, 88127.46, 
    88504.73, 90095.55, 100796.2, 101495, 101484, 101252.7, 93472.1, 78910.53,
  87862.32, 87180.13, 89221.3, 90468.03, 90253.12, 90251.71, 90201.27, 
    92135.56, 96047, 101542.3, 101403.9, 101443, 101253.4, 87607.76, 78694.78,
  91507.84, 88419.55, 88889.52, 90638.72, 90338.53, 89365.24, 89959.73, 
    91735.35, 95900.26, 101554.1, 101460.8, 101484.7, 101289.2, 86466.99, 
    88401.34,
  94444.3, 90307.36, 89453.46, 90537.66, 89745.93, 87455.61, 88690.76, 
    91238.82, 101140, 101569.3, 101469.2, 101449.4, 101358.9, 93812.91, 
    96378.34,
  97548.23, 93050.25, 91581.04, 93895.8, 94138.43, 94324.83, 95239.03, 
    101052.1, 101609.6, 101550, 101492.6, 101452.2, 101402.9, 99209.8, 
    100207.2,
  101141.2, 100810, 97070.69, 94614.91, 94538.9, 93521.86, 91251.55, 
    91685.62, 86127.42, 81733.19, 79529.3, 79915.77, 82824.9, 81499.89, 
    91397.16,
  101152.3, 101056, 98845.8, 93916.62, 91275.83, 89459.03, 88224.04, 
    88469.86, 83746, 81187.68, 80448.7, 81161.52, 83308.77, 82301.88, 92733.42,
  92485.48, 89152.86, 93872.95, 92525.53, 86339.29, 85341.75, 87481.01, 
    86729.71, 82009.23, 79925.33, 79084.39, 79788.99, 81111.42, 82697.24, 
    94757.29,
  86755.62, 86951.18, 86022.25, 84433.73, 84184.45, 82758.33, 83576.27, 
    83845.06, 81618.91, 80425.15, 80127.61, 81638.65, 81273.77, 83256.61, 
    88958.1,
  88280.75, 87442.23, 88425.45, 87651.04, 87521.25, 85985.9, 84983.2, 
    84491.76, 83525.38, 85645.61, 100389.4, 100837.1, 91230.34, 91592.68, 
    84273.73,
  88696.89, 86978.92, 89413.8, 90204.43, 89358.9, 88955.05, 88289.78, 
    88660.17, 90318.39, 101018.3, 101780.7, 101787.3, 101622.5, 93618.66, 
    79001.11,
  87950.15, 87257.88, 89319.55, 90545.06, 90362.59, 90378.96, 90372.79, 
    92286.27, 96234.3, 101747.6, 101707.5, 101702.4, 101608.3, 87735.64, 
    78858.71,
  91549.77, 88501.88, 88992.21, 90733.24, 90456.34, 89504.38, 90129.83, 
    91879.8, 96059.69, 101775.4, 101752.3, 101767.2, 101603.6, 86603.98, 
    88643.57,
  94463.11, 90400.27, 89562.16, 90657.05, 89868.52, 87598.75, 88850.47, 
    91417.39, 101247.6, 101773.5, 101745.9, 101742.8, 101682.5, 94033.2, 
    96665.79,
  97513.55, 93104.32, 91666.84, 93964.75, 94218.83, 94408.11, 95349.42, 
    101129.1, 101724.4, 101765, 101751.5, 101739.3, 101707.2, 99494.95, 
    100519.4,
  101125.7, 100810.4, 97040.07, 94644.48, 94573.43, 93525.1, 91271.5, 
    91746.03, 86153.9, 81785.62, 79577.49, 79919.14, 82839, 81479.98, 91422.91,
  101196.5, 101088.3, 98860.02, 93991.81, 91331.66, 89497.61, 88293.67, 
    88548.98, 83789.34, 81236.12, 80491.48, 81206.38, 83337.18, 82318.83, 
    92831.34,
  92535.74, 89286.98, 93963.85, 92588.84, 86394.63, 85405.97, 87525.54, 
    86784.27, 82089.16, 80002.65, 79110.19, 79811.23, 81150.22, 82706.53, 
    94809.4,
  86921, 87081.2, 86138.16, 84570.14, 84301.31, 82871.37, 83673.46, 83940.68, 
    81681.23, 80457.24, 80206.27, 81724.88, 81306.17, 83311.73, 89045.73,
  88446.03, 87587.3, 88572.08, 87799.41, 87665.89, 86112.09, 85101.7, 
    84599.99, 83595.03, 85851.71, 100450.7, 100897.3, 91343.26, 91679.77, 
    84327.36,
  88860.34, 87143.42, 89574.37, 90347.2, 89515.84, 89105.5, 88441.82, 
    88800.3, 90462.05, 101023.2, 101839.4, 101863.1, 101733.8, 93628.85, 
    79114.35,
  88133.4, 87423.62, 89496.89, 90695.27, 90522.24, 90532.5, 90516.32, 
    92382.31, 96308.85, 101819.3, 101823.5, 101769.4, 101689.5, 87796.57, 
    78956.3,
  91745.28, 88683, 89170.05, 90901.28, 90609.52, 89657.39, 90280.37, 
    91992.35, 96174.16, 101837.5, 101824.7, 101851.8, 101643.8, 86679.95, 
    88692.01,
  94644.24, 90585.31, 89756.2, 90829.92, 90031.41, 87766.18, 88993.79, 
    91579.11, 101311.7, 101854.8, 101820.6, 101837.8, 101714.5, 94154.63, 
    96738.52,
  97688.17, 93312.71, 91870.77, 94160.91, 94411.16, 94595.81, 95503.95, 
    101224.1, 101796.7, 101865.6, 101840.5, 101841.5, 101792.1, 99520.01, 
    100582.8,
  101023.1, 100742.2, 96986.91, 94631.59, 94577.15, 93522.06, 91264.4, 
    91768.34, 86141.71, 81796.68, 79633.84, 79932.16, 82796.46, 81439.07, 
    91424.9,
  101162.7, 101050.9, 98855.27, 93997.48, 91352.98, 89534.95, 88352.45, 
    88591.23, 83823.5, 81285.17, 80535.43, 81264.65, 83429.16, 82312.29, 
    92901.61,
  92509.22, 89306.91, 93971.04, 92595.23, 86419.18, 85469.09, 87596.87, 
    86849.22, 82147.23, 80047.55, 79112.22, 79812.86, 81175.51, 82705.53, 
    94961.36,
  86934.73, 87103.4, 86168.09, 84614.09, 84348.75, 82939.02, 83760.12, 
    84031.06, 81739.2, 80467.84, 80324.95, 81852.57, 81336.56, 83389.06, 
    89165.87,
  88474.33, 87633.67, 88628.87, 87871.83, 87737.27, 86196.28, 85189.88, 
    84701.95, 83691.12, 85972.98, 100469.8, 100919, 91445.12, 91747.91, 
    84264.2,
  88885.46, 87215, 89645.39, 90426.62, 89607.97, 89206.61, 88547.74, 
    88910.47, 90565.95, 101071.9, 101924.9, 101924.4, 101799.6, 93672.38, 
    79105.18,
  88207.94, 87508.92, 89594.88, 90789.95, 90631.01, 90645.05, 90639.98, 
    92509.91, 96411.74, 101900.7, 101894.7, 101790.7, 101805.1, 87795.6, 
    78922.67,
  91844.52, 88797.62, 89298.65, 91044.97, 90752.4, 89808.95, 90429.34, 
    92130.47, 96325.51, 101903.6, 101874.7, 101856, 101693.7, 86696.92, 88740,
  94770.44, 90721.62, 89912.59, 90991.07, 90180.27, 87912.42, 89152.16, 
    91796.35, 101507.4, 101945.6, 101859.3, 101844.2, 101731.3, 94183.53, 
    96676.12,
  97860.36, 93486.15, 92085.85, 94421.83, 94698.46, 94892.15, 95813.79, 
    101492.5, 101975.1, 101955.7, 101863, 101819.8, 101744.1, 99526.73, 
    100526.2,
  100940.2, 100646.2, 96889, 94542.56, 94470.23, 93404.34, 91141.11, 
    91631.92, 86016, 81698.4, 79549.35, 79902.32, 82835.08, 81426.16, 91335.02,
  101044.3, 100959.2, 98742.77, 93888.82, 91238.86, 89417.96, 88244.7, 
    88484.41, 83741.98, 81241.87, 80485.56, 81201.77, 83310.59, 82216.95, 
    92824.34,
  92418.64, 89200.64, 93876.46, 92490.27, 86322.67, 85360.74, 87493.89, 
    86739.37, 82058.08, 79966.8, 79042.29, 79783.57, 81112.02, 82659.27, 
    94756.98,
  86808.75, 86969.88, 86049.38, 84473.86, 84216.7, 82814.41, 83648.55, 
    83935.32, 81691.12, 80415.99, 80251.68, 81739.27, 81197.87, 83222.04, 
    88940.17,
  88354.06, 87522.12, 88534.23, 87767.05, 87628.91, 86090.44, 85073.29, 
    84599.62, 83618.1, 85815.83, 100438.3, 100902.2, 91366.59, 91655.54, 
    84238.41,
  88744.32, 87091.26, 89530, 90328.99, 89503.31, 89116.81, 88454.98, 
    88842.95, 90487.71, 101124.8, 101860.1, 101867.7, 101662.6, 93699.9, 
    78877.15,
  88059.34, 87372.66, 89478.14, 90690.27, 90525.52, 90556.61, 90566.86, 
    92489.3, 96403.91, 101893.7, 101815.7, 101766.5, 101709, 87767.47, 
    78690.97,
  91694.11, 88651.68, 89167.02, 90933.57, 90644.59, 89714.84, 90360.3, 
    92092.66, 96321.88, 101920.8, 101825.2, 101826.9, 101698.8, 86556.67, 
    88527.51,
  94629.16, 90579.27, 89780, 90868.96, 90062.66, 87776.42, 89039.12, 
    91723.42, 101573.7, 101956.7, 101845.8, 101822.6, 101712.4, 94099.88, 
    96589.61,
  97744.62, 93368.14, 91971.23, 94314.41, 94599.08, 94796.69, 95765.06, 
    101540.6, 102021, 102002.1, 101900.4, 101848.3, 101766.4, 99505.63, 
    100517.9,
  100810.2, 100516.8, 96719.14, 94354.88, 94307.29, 93286.22, 91031.65, 
    91480.95, 85941.47, 81583.78, 79464.88, 79823.61, 82721.7, 81395.23, 
    91300.72,
  100809.5, 100790.5, 98565.72, 93683.57, 91054.88, 89257.94, 88076.85, 
    88328.55, 83618.18, 81082.99, 80366.63, 81046.79, 83208.81, 82182.62, 
    92685.35,
  92258.62, 88934.62, 93624.59, 92263.96, 86140.48, 85165.48, 87308.58, 
    86579.66, 81867.3, 79787.42, 78931.38, 79656.86, 81009.8, 82557.27, 
    94682.42,
  86591.72, 86702.68, 85818.66, 84207.84, 83956.51, 82579.44, 83410.52, 
    83690.65, 81479.39, 80259.8, 79998.19, 81535.05, 81073.97, 83080.22, 
    88875.44,
  88105.49, 87255.65, 88270.27, 87483.17, 87344.55, 85806.19, 84803.79, 
    84332.41, 83382.45, 85484.8, 100241.7, 100732.5, 91141.44, 91504.91, 
    84152.38,
  88468.05, 86808.46, 89231.94, 90040.48, 89190.16, 88789.48, 88137.98, 
    88540.63, 90155.67, 100931.3, 101725.1, 101720.3, 101507.7, 93560.35, 
    78742.18,
  87776.97, 87072.23, 89164.23, 90385.7, 90203.05, 90244.11, 90227.03, 
    92161.32, 96109.33, 101678.1, 101614.6, 101628.1, 101565.1, 87620.91, 
    78556.02,
  91402.84, 88344.67, 88833.94, 90600.11, 90312.89, 89369.84, 89996.81, 
    91763.78, 95946.63, 101677.1, 101632.9, 101678.4, 101555.8, 86415.61, 
    88327.8,
  94337.4, 90274.83, 89452.03, 90536.52, 89732.32, 87433.36, 88696.01, 
    91292.99, 101184.8, 101663.9, 101607.9, 101612.6, 101528.5, 93937.27, 
    96439.19,
  97454.48, 93065.95, 91628.98, 93955.66, 94213.52, 94396.63, 95322.58, 
    101100.3, 101636.9, 101641.1, 101601.7, 101578.8, 101530.7, 99305.8, 
    100335.2,
  100667, 100299.8, 96580.37, 94173.52, 94124.28, 93102.78, 90934.9, 
    91371.24, 85881.23, 81493.18, 79298.7, 79610.32, 82426.61, 81143.2, 
    90946.8,
  100580.8, 100581.2, 98392.38, 93491.59, 90878.69, 89084.33, 87910.91, 
    88163.45, 83502.13, 80883.38, 80143.35, 80794.98, 82901.44, 81894.1, 
    92277.98,
  92050.65, 88722, 93403.41, 92081.99, 85992.97, 84992.08, 87147.09, 
    86433.17, 81720.58, 79611.2, 78766.13, 79455.37, 80753.48, 82281.62, 
    94323.64,
  86346.04, 86512.13, 85641.15, 84033.02, 83781.8, 82418.64, 83255.09, 
    83519.34, 81301.72, 80102.68, 79810.07, 81304.67, 80882.63, 82797.13, 
    88556.64,
  87899.91, 87063.71, 88079.29, 87290.2, 87174.28, 85643.77, 84651.8, 
    84181.95, 83236.83, 85311.59, 100004, 100553.5, 90942.94, 91172.27, 
    83963.38,
  88294.16, 86637.14, 89049.07, 89852.26, 89005.01, 88630.56, 87967.45, 
    88382.86, 89979.12, 100725.2, 101504.2, 101489.3, 101240.7, 93317.19, 
    78529.64,
  87605.27, 86930.29, 89015.76, 90230.25, 90021.8, 90087.7, 90068.94, 
    92025.31, 95925.32, 101469.9, 101347.2, 101432.8, 101266, 87413.16, 
    78239.91,
  91249.66, 88204.16, 88718.01, 90486.7, 90175.16, 89231.98, 89873.59, 
    91640.18, 95787.65, 101477.3, 101401, 101479.7, 101279.2, 86224.95, 
    87917.93,
  94188.04, 90141.88, 89344.37, 90434.78, 89630.96, 87331.55, 88582.67, 
    91198.2, 101093, 101498, 101400.3, 101401.4, 101277.8, 93668.55, 96154.52,
  97336.21, 92943.71, 91530.38, 93879.69, 94151.52, 94351.05, 95284.49, 
    101086.1, 101545.7, 101503.4, 101438.3, 101384.4, 101309.1, 99054.78, 
    100078.8,
  100759.4, 100430.5, 96645.39, 94190.73, 94114.54, 93123.16, 90950.77, 
    91363.95, 85889.68, 81541.88, 79371.11, 79739.33, 82546.53, 81296.23, 
    91116.55,
  100688.6, 100673.9, 98453.44, 93534.53, 90893.45, 89107.17, 87921.12, 
    88200.91, 83563.93, 80978.61, 80256.8, 80947.07, 83045.97, 82062.54, 
    92487.28,
  92131.07, 88792.98, 93485.12, 92142.02, 86015.16, 85036.33, 87185.12, 
    86479.47, 81794.55, 79690.7, 78858.2, 79554.48, 80867.71, 82408.08, 
    94524.01,
  86400.34, 86549.34, 85662.23, 84060.35, 83816.3, 82450.02, 83278.81, 
    83555.03, 81348.66, 80162.22, 79875.5, 81378.82, 80987.28, 82919.84, 
    88684.97,
  87926.59, 87098.38, 88119.84, 87340.25, 87206.84, 85659.85, 84687.3, 
    84217.34, 83294.52, 85368.17, 100134.8, 100647.8, 91054.04, 91307.41, 
    84057.99,
  88309.12, 86634.8, 89083.22, 89894.84, 89066.09, 88669.72, 88006.12, 
    88425.65, 90043.61, 100870.3, 101663.7, 101660.6, 101378.8, 93432.9, 
    78595.5,
  87588.35, 86890.65, 89027.73, 90254.95, 90077.77, 90143.81, 90109.7, 
    92109.08, 96043.93, 101671.9, 101543.9, 101616.8, 101427.9, 87528.38, 
    78289.45,
  91185.38, 88157.62, 88676.23, 90464.47, 90198.93, 89267.82, 89891.25, 
    91701.14, 95890.01, 101679.6, 101584.8, 101670.3, 101448.9, 86306.27, 
    87960.77,
  94133.97, 90101.1, 89314.75, 90422.64, 89621.37, 87334.95, 88608.31, 
    91236.94, 101210.1, 101680.1, 101574.2, 101578, 101420.8, 93788.24, 
    96176.53,
  97287.52, 92862.14, 91478.1, 93864.52, 94151.26, 94355.1, 95300.98, 
    101167.1, 101673.1, 101636.4, 101555.7, 101516.6, 101429.9, 99156.06, 
    100143.3,
  100966.3, 100606.6, 96831.2, 94388.42, 94345.27, 93329.58, 91097.43, 
    91530.8, 85978.37, 81620.45, 79424.96, 79783.36, 82621.98, 81317.27, 
    91251.73,
  100834.4, 100815.2, 98633.45, 93707.05, 91101.73, 89293.62, 88118.09, 
    88377.98, 83671.12, 81097.24, 80368.05, 81057.02, 83144.35, 82143.82, 
    92678.3,
  92313.77, 88935.78, 93635.33, 92297.95, 86209.51, 85211.16, 87379.04, 
    86656.52, 81949.07, 79858.21, 78986.89, 79695.78, 81004.8, 82584.61, 
    94730.29,
  86531.95, 86677.05, 85812.99, 84212.13, 84006.53, 82650.86, 83495.57, 
    83791.01, 81595.98, 80341.55, 80110.83, 81636.94, 81148.84, 83131.97, 
    88863.61,
  88090.38, 87282.3, 88308.74, 87524.71, 87414.52, 85880.79, 84914.38, 
    84444.58, 83504.62, 85680.06, 100603.5, 101054.9, 91405.88, 91641.5, 
    84228.75,
  88481.54, 86800.64, 89262.91, 90097.01, 89305.95, 88939.03, 88292.8, 
    88740.12, 90418.3, 101302.4, 102050.6, 102056.8, 101798.2, 93732.72, 
    78764.71,
  87762.67, 87063.76, 89230.68, 90468.36, 90333.2, 90419.76, 90442.04, 
    92451.9, 96423, 102065, 101988.3, 102012.1, 101871.6, 87738.67, 78514.76,
  91297.56, 88299.56, 88851.49, 90672.16, 90422.03, 89530.88, 90229.34, 
    92024.14, 96326.09, 102102.3, 102021.5, 102080.4, 101876.6, 86480.26, 
    88386.45,
  94258.1, 90233.28, 89473.07, 90601.2, 89842.52, 87594.37, 88910.75, 
    91622.91, 101655, 102120.7, 102044.2, 102061.3, 101914.9, 94199.66, 
    96701.48,
  97379.62, 92996.57, 91647.31, 94047.84, 94362.17, 94577.56, 95649.48, 
    101568, 102116.2, 102140.5, 102083, 102064.4, 101983.9, 99657.2, 100682.1,
  101031, 100702, 96876.6, 94496.02, 94428.98, 93443.77, 91246.45, 91675.7, 
    86128.96, 81768.61, 79575.91, 80061.84, 83005.69, 81706.77, 91818.27,
  100953.4, 100943.7, 98691.59, 93780.8, 91174.38, 89413.89, 88233.98, 
    88516.61, 83809.91, 81257.06, 80555.38, 81263.72, 83468.49, 82462.88, 
    93124.01,
  92371.81, 89032.54, 93786.52, 92447.68, 86282.67, 85290.81, 87464.91, 
    86757.48, 82020.05, 79966.09, 79160.94, 79886, 81268.71, 82857.75, 
    95178.46,
  86617.4, 86764.37, 85860.53, 84279.85, 84054.62, 82708.93, 83561.6, 
    83865.34, 81669.33, 80467.97, 80186.41, 81751.1, 81333.68, 83361.45, 
    89244.49,
  88176.14, 87363.62, 88370.44, 87584.21, 87464.38, 85919.66, 84972.5, 
    84505.82, 83581.52, 85726.27, 100730.5, 101202.8, 91459.7, 91884, 84460.31,
  88524.63, 86870.43, 89329.59, 90154.91, 89342.74, 88964.7, 88333.25, 
    88750.09, 90488.65, 101421.2, 102242.5, 102208.8, 102042.8, 93934.52, 
    79067.88,
  87804.99, 87130.67, 89297.47, 90527.22, 90384.06, 90462.19, 90493.05, 
    92502.77, 96551.81, 102158, 102144.9, 102123.3, 102129.5, 87892.26, 
    78921.59,
  91386.11, 88354.02, 88896.4, 90705.59, 90448.44, 89532.12, 90236.45, 
    92059.04, 96424.32, 102225.2, 102204.2, 102224.8, 102030.2, 86770.62, 
    88876.91,
  94311.59, 90256.28, 89487.12, 90601.78, 89863.84, 87622.07, 88940.34, 
    91607.9, 101709, 102248.5, 102210.1, 102268.4, 102140.9, 94477.2, 97161.69,
  97403.01, 93021.27, 91626.38, 94005.29, 94276.38, 94420.34, 95479.98, 
    101470.8, 102190.3, 102266.5, 102258.8, 102288.1, 102244.6, 100005.9, 
    101142.2,
  101048.7, 100714.8, 96921.98, 94564.77, 94489, 93479.73, 91310.91, 
    91756.32, 86267.63, 81900.33, 79706.28, 80074.44, 83097.09, 81802.44, 
    91932.22,
  100981.3, 100964.5, 98727.45, 93844.96, 91225.69, 89445.55, 88269.91, 
    88559.79, 83909.52, 81316.42, 80606.66, 81333.82, 83583.51, 82549.55, 
    93253.89,
  92430.19, 89103.47, 93803.59, 92478.21, 86327.82, 85356.93, 87470.7, 
    86796.88, 82092.8, 80005.15, 79211.03, 79930.47, 81339.25, 82882.85, 
    95256.55,
  86707.14, 86856.02, 85929.45, 84338.1, 84084.1, 82745.31, 83573.74, 
    83871.08, 81653.58, 80468.67, 80167.88, 81687.52, 81398.22, 83407.09, 
    89424.25,
  88266.12, 87428.51, 88432.96, 87650.25, 87499.49, 85926.46, 84945.22, 
    84468.16, 83516.69, 85598.83, 100346.8, 100836.7, 91194.77, 91661.26, 
    84566.49,
  88594.7, 86888.36, 89347.07, 90138.62, 89304.97, 88899.18, 88229.13, 
    88636.96, 90267.4, 101055.1, 101937.1, 101915.7, 101654.8, 93739.6, 
    79190.95,
  87863.45, 87145.88, 89276.87, 90502.66, 90312.75, 90367.77, 90338, 
    92294.16, 96256.67, 101835.9, 101753.7, 101786.2, 101682.7, 87838.64, 
    78953.47,
  91420.11, 88366.48, 88846.45, 90655.53, 90375.22, 89406.53, 90071.39, 
    91863.48, 96087.98, 101856.1, 101801.5, 101857, 101728.2, 86699.87, 
    88637.44,
  94356.48, 90263.21, 89445.28, 90545.25, 89812.96, 87543.79, 88800.9, 
    91348.31, 101310.5, 101854.3, 101789.4, 101826.5, 101756.4, 94119.1, 
    96770.43,
  97435.44, 93002.01, 91561.3, 93908.67, 94181.38, 94327.04, 95263.95, 
    101120.4, 101818.8, 101854.9, 101846.2, 101852.2, 101811.2, 99577.76, 
    100797.3,
  100976.6, 100630, 96896.3, 94488.85, 94403.79, 93403.49, 91231.33, 
    91694.16, 86188.35, 81857.34, 79658.47, 79987.41, 82923.68, 81607.81, 
    91561.23,
  100850.9, 100848, 98633.12, 93759.05, 91154.19, 89375.29, 88223.38, 
    88516.49, 83854.71, 81289.23, 80558.04, 81235.45, 83414.73, 82387.2, 
    92884.48,
  92359.12, 89027.45, 93733.85, 92442.98, 86289.15, 85318.23, 87419.07, 
    86757.08, 82084.31, 80003.97, 79171.34, 79866.18, 81241.43, 82763.66, 
    94914.45,
  86601.18, 86701, 85788.62, 84229.56, 84001.22, 82679.96, 83515.79, 
    83852.97, 81663.12, 80455.26, 80123.55, 81621.03, 81269.41, 83237.3, 
    89110.5,
  88196.25, 87276.3, 88248.94, 87449.11, 87302.14, 85799.24, 84858.02, 
    84432.58, 83500.39, 85497.55, 100131.5, 100643.8, 91134.17, 91508.93, 
    84362.74,
  88460.24, 86734.84, 89148.63, 89970.66, 89142.95, 88734.2, 88094.65, 
    88537.77, 90115.09, 100833.8, 101669.1, 101654.8, 101415.3, 93548.37, 
    79025.82,
  87746.37, 87026.34, 89094.9, 90309.09, 90119.5, 90202.62, 90170.52, 
    92141.33, 96025.57, 101580.6, 101508.3, 101553.6, 101468.2, 87685, 
    78869.67,
  91361.71, 88233.34, 88734.62, 90515.08, 90224.95, 89296.95, 89932.75, 
    91705.59, 95871.2, 101591.4, 101575.9, 101630.9, 101439.1, 86529.01, 
    88578.97,
  94309.15, 90158.69, 89359.78, 90456.91, 89706.9, 87463.59, 88716.45, 
    91229.48, 101095.7, 101599.5, 101560.4, 101595.7, 101533.9, 93939.66, 
    96511.89,
  97419.83, 92968.77, 91504.42, 93831.44, 94086.48, 94239.68, 95174.83, 
    101030.3, 101592.3, 101620.7, 101599.9, 101598.9, 101539.9, 99261.74, 
    100383.5,
  100777.4, 100418.1, 96702.27, 94263.05, 94156.2, 93108.71, 90919.3, 
    91428.38, 85944.34, 81614.87, 79427.77, 79759.53, 82666.6, 81343.84, 
    91244.16,
  100634, 100633.8, 98438.86, 93537.75, 90900.38, 89071.41, 87924.2, 
    88235.52, 83609.61, 81059.91, 80330.84, 81005.48, 83179.09, 82145.35, 
    92551.49,
  92095.85, 88775.98, 93478.56, 92192.69, 85995.2, 85027.34, 87144.83, 
    86490.38, 81863.93, 79787.02, 78954.73, 79654.81, 81004.76, 82535.2, 
    94562.31,
  86335.27, 86416.8, 85545.93, 83993.48, 83753.03, 82425.6, 83263.48, 
    83611.5, 81431.9, 80223.66, 79904.93, 81406.74, 81067.44, 83011.36, 
    88812.95,
  87958.67, 87005.28, 87980.99, 87174.89, 87038.71, 85536.06, 84604.56, 
    84187.5, 83253.44, 85263.85, 99871.95, 100347.1, 90857.51, 91274.02, 
    84119.88,
  88229.9, 86544.67, 88947.12, 89727.47, 88867.03, 88475.56, 87835.04, 
    88257.26, 89886.41, 100559.1, 101358.3, 101335.1, 101112.9, 93284.09, 
    78833.59,
  87534.48, 86842.62, 88918.14, 90097.88, 89890.78, 89946.63, 89959.34, 
    91906.23, 95813.46, 101291.3, 101219.3, 101243.9, 101172.3, 87439.84, 
    78664.14,
  91144.49, 88091.91, 88591.91, 90329.59, 90025.77, 89082.31, 89720.74, 
    91478.55, 95667.16, 101314.5, 101266.2, 101296.9, 101117.6, 86331.55, 
    88374.7,
  94121.75, 89997.98, 89196.23, 90269.64, 89493.88, 87252.56, 88523.59, 
    91059.35, 100878.6, 101328.7, 101252.1, 101269.5, 101167.1, 93722.16, 
    96302.32,
  97234.66, 92805.76, 91352.92, 93672.52, 93929.52, 94056.73, 94983.04, 
    100822.6, 101357.5, 101351.1, 101278.7, 101250.8, 101194.8, 99057.04, 
    100238.3,
  100636, 100290.9, 96517.62, 94068.22, 93919.16, 92841.17, 90667.62, 
    91142.4, 85676.31, 81348.07, 79165.78, 79499.65, 82409.2, 81089.68, 
    90970.75,
  100474.7, 100487.6, 98276.09, 93386.22, 90698.25, 88884.8, 87689.55, 
    87980.93, 83339.32, 80783.72, 80054.82, 80714.77, 82902.2, 81866.52, 
    92261.95,
  91943.31, 88607.05, 93269.26, 91959.85, 85789.84, 84829.65, 86926.71, 
    86243.87, 81614.05, 79540.12, 78690.16, 79370.77, 80719.18, 82240.45, 
    94217.98,
  86185.55, 86255.96, 85379.52, 83788.13, 83536.95, 82205.19, 83048.8, 
    83362.93, 81165.27, 79951.25, 79628.99, 81144.84, 80761.95, 82711.37, 
    88541.04,
  87773.87, 86829.55, 87809.52, 87030.84, 86892.02, 85361.88, 84393.76, 
    83943.63, 83020.43, 85017.33, 99607.93, 100057.9, 90614.96, 90975.26, 
    83832.12,
  88041.82, 86329.47, 88698.3, 89516.36, 88661.95, 88276.47, 87627, 88044.84, 
    89629.32, 100262.7, 101020.5, 101019.5, 100820.3, 92996.24, 78539.43,
  87285.48, 86593.32, 88656.92, 89889.83, 89669.81, 89729.48, 89703.08, 
    91649.28, 95513.92, 100967.8, 100884.3, 100921.9, 100852.4, 87170.87, 
    78360.57,
  90908.24, 87830.38, 88312.51, 90076.4, 89784.11, 88825.9, 89463.11, 
    91235.14, 95390.62, 100978.2, 100914.4, 100967.4, 100845.3, 86046.23, 
    88030.8,
  93850.2, 89736.38, 88935.02, 90008.89, 89249, 87010.81, 88281.72, 90805.2, 
    100578.7, 100973.4, 100898.2, 100910.5, 100815.4, 93416.2, 95983.86,
  96945.3, 92535.52, 91083.65, 93408.82, 93662.6, 93798.31, 94736.8, 
    100532.1, 101038.1, 100987.3, 100944.9, 100951.4, 100917.5, 98804.18, 
    99940.16,
  100538.7, 100185.7, 96444.77, 93989.87, 93828.2, 92765.09, 90626.8, 
    91075.11, 85575.58, 81223.2, 79033.8, 79355.14, 82185.73, 80884.36, 90760,
  100345.9, 100374.3, 98200.6, 93279.48, 90598.61, 88782.73, 87631.41, 
    87897.09, 83253.16, 80678.65, 79930.92, 80583.16, 82715.55, 81668.95, 
    92017.02,
  91825.77, 88465.3, 93157.8, 91904.34, 85739.52, 84726.63, 86867.6, 
    86172.62, 81513.81, 79409.07, 78524.73, 79193.33, 80500.06, 82021.45, 
    94019.48,
  86054.51, 86115.13, 85244.84, 83660.35, 83449.66, 82119.44, 82977.09, 
    83280.88, 81073.78, 79845.96, 79580.88, 81070.13, 80619.45, 82541.26, 
    88288.44,
  87601.53, 86689.66, 87708.07, 86938.27, 86830.44, 85326.39, 84360.6, 
    83900.85, 82972.05, 85019.35, 99522.4, 99980.35, 90535.7, 90850.11, 
    83614.23,
  87888.02, 86223.93, 88638.01, 89449.72, 88634.7, 88269.05, 87619.28, 
    88061.84, 89667.95, 100222.2, 100923, 100909.2, 100719.2, 92899.24, 
    78283.77,
  87211.08, 86520.95, 88616.17, 89838.22, 89670.12, 89753.66, 89752.95, 
    91679.47, 95549.12, 100923.7, 100826.4, 100813.2, 100789.4, 87018.3, 
    78151.58,
  90815.25, 87757.88, 88276.09, 90047.86, 89768.93, 88861.03, 89515.51, 
    91304.13, 95484.06, 100999, 100884.8, 100872.6, 100734.7, 85876.41, 
    87909.41,
  93766.6, 89690.01, 88907.54, 89989.34, 89233.2, 87022.7, 88320.66, 
    90966.12, 100697.9, 101083.6, 100980.9, 100945.6, 100786.6, 93380.88, 
    95875.83,
  96886.78, 92474.67, 91077.23, 93420.13, 93670.36, 93843.3, 94875.55, 
    100681.6, 101197.8, 101201.6, 101153.2, 101128.7, 101016.7, 98836.55, 
    99941.79 ;

 sftlf =
  0.0008770345, 0.4596241, 0.9892928, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.01035247, 0.004304647, 0.6546783, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.8534847, 0.8118016, 0.9951549, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9894952, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4452189, 0.3028796, 0.7140614, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9903189, 0.3150955, 0.0007410151, 0, 0.02645395, 
    0.9012984, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.681631, 0, 0, 0, 0.004980796, 0.7708192, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5536854, 0, 0, 0, 0.004666397, 0.9395298, 1,
  1, 1, 1, 1, 1, 1, 1, 0.9995009, 0.3626226, 0, 0, 0, 0, 0.8367797, 1,
  1, 1, 1, 1, 1, 0.8451425, 0.7016711, 0.3953246, 0, 0, 0, 0, 0.006316811, 
    0.8673657, 1 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0.2038203, 25.08469, 362.922, 581.3585, 583.7158, 677.0037, 892.3406, 
    840.3151, 1394.918, 1845.667, 2078.668, 2048.803, 1746.472, 1895.031, 
    903.5963,
  0.04938461, 3.284697, 202.5217, 654.3141, 903.2668, 1076.606, 1196.302, 
    1163.293, 1639.916, 1906.256, 1988.945, 1916.741, 1695.228, 1807.269, 
    774.2457,
  790.1076, 1114.346, 653.3495, 780.126, 1392.106, 1491.591, 1273.753, 
    1344.373, 1825.463, 2046.944, 2142.644, 2067.535, 1930.862, 1770.506, 
    591.146,
  1359.809, 1341.669, 1435.043, 1594.124, 1615.893, 1763.274, 1677.539, 
    1645.991, 1875.931, 2003.645, 2040.039, 1879.801, 1919.839, 1717.029, 
    1138.974,
  1205.389, 1290.31, 1192.454, 1271.409, 1283.839, 1439.06, 1538.882, 
    1587.552, 1685.139, 1482.705, 108.3495, 67.86669, 940.4369, 898.4109, 
    1612.947,
  1168.617, 1342.769, 1106.133, 1029.211, 1110.353, 1151.071, 1218.088, 
    1182.275, 1031.226, 58.02261, 0, 0, 7.641389, 710.6758, 2161.482,
  1244.873, 1316.863, 1112.963, 998.5415, 1017.03, 1014.576, 1020.14, 
    838.6226, 484.287, 0, 0, 0, 0, 1273.715, 2180.106,
  896.0552, 1198.27, 1151.006, 981.8504, 1010.922, 1103.887, 1045.003, 
    880.1057, 498.0692, 0, 0, 0, 0, 1386.297, 1186.975,
  625.923, 1015.673, 1096.604, 994.0698, 1069.039, 1288.357, 1166.806, 
    927.0013, 34.64387, 0, 0, 0, 0, 678.2806, 439.0615,
  346.5426, 755.811, 896.7624, 677.1516, 656.058, 642.5463, 557.833, 
    41.91994, 0, 0, 0, 0, 0, 191.3587, 93.07086 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
