netcdf \00010101.atmos_daily.tile6.pr {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pr(time, grid_yt, grid_xt) ;
		pr:_FillValue = 1.e+20f ;
		pr:missing_value = 1.e+20f ;
		pr:units = "kg m-2 s-1" ;
		pr:long_name = "Precipitation" ;
		pr:cell_methods = "time: mean" ;
		pr:cell_measures = "area: area" ;
		pr:time_avg_info = "average_T1,average_T2,average_DT" ;
		pr:standard_name = "precipitation_flux" ;
		pr:interp_method = "conserve_order1" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:11 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile6.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile6.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pr =
  4.935544e-06, 8.669232e-06, 7.880827e-06, 9.642461e-06, 9.401841e-06, 
    7.358928e-06, 6.497738e-06, 7.129477e-06, 8.335194e-06, 6.89705e-06, 
    7.903425e-06, 6.231838e-06, 8.873928e-06, 6.634148e-06, 4.472528e-06,
  4.072285e-06, 6.69937e-06, 6.587232e-06, 6.769203e-06, 7.658098e-06, 
    7.454943e-06, 7.065874e-06, 6.650766e-06, 7.472097e-06, 6.549661e-06, 
    7.419354e-06, 7.858023e-06, 8.520199e-06, 5.096533e-06, 5.500795e-06,
  7.18965e-06, 5.09165e-06, 5.582237e-06, 7.474494e-06, 6.444301e-06, 
    5.820695e-06, 8.533938e-06, 6.890264e-06, 3.992357e-06, 5.518267e-06, 
    6.061213e-06, 7.61206e-06, 5.96662e-06, 4.954127e-06, 7.506804e-06,
  8.295286e-06, 6.156186e-06, 6.921537e-06, 5.763321e-06, 7.159228e-06, 
    7.547847e-06, 7.498587e-06, 7.066327e-06, 3.900836e-06, 6.365308e-06, 
    5.990045e-06, 6.550981e-06, 4.628474e-06, 6.702026e-06, 8.486608e-06,
  1.210464e-05, 9.303099e-06, 8.229322e-06, 7.226047e-06, 4.630325e-06, 
    6.541086e-06, 5.542287e-06, 7.05038e-06, 5.303815e-06, 5.342267e-06, 
    6.093222e-06, 6.185023e-06, 8.141426e-06, 6.601173e-06, 8.758681e-06,
  1.13243e-05, 9.405739e-06, 9.505738e-06, 6.755864e-06, 6.133313e-06, 
    3.709512e-06, 5.707478e-06, 4.959293e-06, 6.364463e-06, 3.173879e-06, 
    3.663628e-06, 6.119421e-06, 8.614092e-06, 8.10389e-06, 9.546279e-06,
  1.568661e-05, 1.092151e-05, 1.125675e-05, 8.77475e-06, 6.803327e-06, 
    7.231684e-06, 5.999937e-06, 5.408805e-06, 3.942196e-06, 4.308752e-06, 
    3.052419e-06, 6.108362e-06, 7.925044e-06, 7.381254e-06, 9.957332e-06,
  1.814334e-05, 1.703472e-05, 1.374231e-05, 1.05557e-05, 9.245543e-06, 
    8.305958e-06, 7.129302e-06, 5.150614e-06, 4.095245e-06, 7.039715e-06, 
    4.41356e-06, 5.713365e-06, 9.011726e-06, 7.631253e-06, 1.002147e-05,
  2.109248e-05, 1.820515e-05, 1.510357e-05, 1.101098e-05, 1.235277e-05, 
    1.050718e-05, 8.800232e-06, 6.573062e-06, 5.884405e-06, 3.682753e-06, 
    6.406504e-06, 4.899152e-06, 7.875115e-06, 7.526164e-06, 9.505437e-06,
  2.719414e-05, 2.298024e-05, 1.597636e-05, 1.461397e-05, 1.296648e-05, 
    1.138221e-05, 1.023421e-05, 6.482797e-06, 5.88911e-06, 3.780231e-06, 
    5.352351e-06, 6.363538e-06, 6.091254e-06, 8.036482e-06, 9.271093e-06,
  6.356047e-06, 4.979139e-06, 4.154731e-06, 3.869193e-06, 4.051995e-06, 
    6.26994e-06, 7.186257e-06, 6.361599e-06, 6.513287e-06, 4.817141e-06, 
    2.809482e-06, 2.482078e-06, 2.624655e-06, 2.803319e-06, 1.473691e-06,
  6.985473e-06, 7.114739e-06, 3.636911e-06, 4.438356e-06, 3.749375e-06, 
    5.079718e-06, 5.087345e-06, 7.203395e-06, 6.677275e-06, 5.088484e-06, 
    4.000296e-06, 4.99371e-06, 3.594169e-06, 2.293325e-06, 6.4738e-07,
  8.061549e-06, 7.715169e-06, 8.423547e-07, 2.909505e-06, 3.602898e-06, 
    3.927464e-06, 6.040739e-06, 6.224293e-06, 5.159824e-06, 3.618379e-06, 
    5.028022e-06, 2.757093e-06, 3.830882e-06, 2.103137e-06, 8.875623e-07,
  8.663998e-06, 6.131322e-06, 5.087109e-06, 3.354871e-06, 3.738197e-06, 
    3.679872e-06, 6.075106e-06, 5.827237e-06, 5.506994e-06, 6.775172e-06, 
    3.669207e-06, 4.945294e-06, 3.071293e-06, 2.358404e-06, 1.067548e-06,
  4.573321e-06, 5.376243e-06, 7.121745e-06, 6.218807e-06, 3.371749e-06, 
    5.516461e-06, 8.55724e-06, 6.355394e-06, 5.498176e-06, 4.798328e-06, 
    4.30111e-06, 2.991139e-06, 6.655673e-06, 2.429497e-06, 7.742067e-07,
  7.233455e-06, 6.899063e-06, 7.146499e-06, 5.115976e-06, 6.459179e-06, 
    9.526439e-06, 5.725004e-06, 4.194063e-06, 3.75343e-06, 4.526625e-06, 
    3.846133e-06, 5.234845e-06, 5.40661e-06, 2.087812e-06, 2.778024e-07,
  1.059153e-05, 8.761326e-06, 5.823259e-06, 3.86886e-06, 1.296187e-05, 
    1.054575e-05, 7.898468e-06, 3.059461e-06, 2.806587e-06, 4.837052e-06, 
    6.137193e-06, 5.457128e-06, 4.313153e-06, 1.188654e-06, 3.365813e-07,
  1.041195e-05, 9.087723e-06, 8.414342e-06, 4.973987e-06, 7.015959e-06, 
    9.963303e-06, 4.824841e-06, 4.339869e-06, 3.265771e-06, 2.429326e-06, 
    2.300251e-06, 6.204073e-06, 3.731389e-06, 2.591327e-06, 2.736714e-07,
  1.582719e-05, 1.178565e-05, 8.337133e-06, 6.370266e-06, 7.529473e-06, 
    1.068943e-05, 5.828334e-06, 4.338912e-06, 4.601746e-06, 4.231068e-06, 
    3.983792e-06, 5.926589e-06, 3.167979e-06, 2.065702e-06, 1.204727e-06,
  1.470237e-05, 1.215216e-05, 1.015181e-05, 5.868306e-06, 5.683103e-06, 
    8.237042e-06, 8.340332e-06, 3.457004e-06, 5.622464e-06, 3.188527e-06, 
    2.475417e-06, 4.484701e-06, 3.560335e-06, 1.136922e-06, 2.633564e-06,
  3.233854e-06, 1.75515e-06, 1.878002e-06, 1.073448e-06, 2.150406e-06, 
    1.644166e-06, 2.419905e-06, 4.144854e-06, 8.286862e-06, 2.334795e-05, 
    4.477989e-05, 7.300486e-05, 0.000121737, 0.0002393822, 0.0005103793,
  3.901941e-06, 1.22153e-06, 1.18089e-06, 1.109753e-06, 1.06624e-06, 
    1.657034e-06, 2.896925e-06, 2.217325e-06, 5.000121e-06, 1.692718e-05, 
    3.194766e-05, 4.570654e-05, 8.224472e-05, 0.0001774821, 0.0003947448,
  2.875284e-06, 2.396631e-06, 1.018814e-06, 2.289757e-06, 1.415737e-06, 
    1.230066e-06, 1.585873e-06, 2.183009e-06, 3.746751e-06, 1.031262e-05, 
    2.667152e-05, 4.014086e-05, 6.536125e-05, 0.0001353094, 0.000315355,
  4.241237e-06, 2.548818e-06, 1.628605e-06, 5.39059e-06, 4.468136e-06, 
    2.473141e-06, 2.591796e-06, 3.134122e-06, 2.948234e-06, 7.184445e-06, 
    2.544378e-05, 4.729993e-05, 7.71495e-05, 0.000128361, 0.0002790236,
  6.21481e-06, 5.103796e-06, 4.774666e-06, 3.055298e-06, 2.619365e-06, 
    4.157848e-06, 2.315787e-06, 2.437318e-06, 2.542811e-06, 3.338991e-06, 
    1.874186e-05, 5.811371e-05, 9.754212e-05, 0.0001585698, 0.0002975493,
  1.187745e-05, 9.628849e-06, 5.555378e-06, 3.932878e-06, 1.663272e-06, 
    2.428698e-06, 5.016575e-06, 5.274133e-06, 6.061477e-06, 3.134596e-06, 
    4.661444e-06, 3.538987e-05, 9.419942e-05, 0.0001833705, 0.0003276168,
  1.666018e-05, 9.886649e-06, 8.848587e-06, 7.103989e-06, 6.211805e-06, 
    4.049461e-06, 3.951436e-06, 3.122648e-06, 3.233807e-06, 3.595846e-06, 
    3.925115e-06, 8.105868e-06, 3.331426e-05, 0.0001561189, 0.0002981648,
  1.462785e-05, 1.228245e-05, 6.209044e-06, 5.536641e-06, 7.38464e-06, 
    7.710951e-06, 5.387607e-06, 3.249815e-06, 4.758218e-06, 7.276697e-06, 
    1.260419e-05, 1.177377e-05, 2.991296e-05, 9.648456e-05, 0.0001968876,
  1.199602e-05, 1.281447e-05, 8.094448e-06, 7.808166e-06, 8.382853e-06, 
    9.108713e-06, 8.348042e-06, 7.895704e-06, 3.985369e-06, 3.856328e-06, 
    6.992674e-06, 1.069801e-05, 3.271376e-05, 8.079591e-05, 0.0001267952,
  1.057258e-05, 1.115268e-05, 6.368955e-06, 1.276956e-05, 8.028337e-06, 
    3.549318e-06, 6.394523e-06, 6.022131e-06, 6.2174e-06, 3.631638e-06, 
    2.321391e-06, 4.252056e-06, 5.297831e-06, 2.853929e-05, 6.670409e-05,
  3.345399e-06, 4.532988e-06, 4.497263e-06, 2.05168e-06, 1.260828e-05, 
    9.29178e-05, 0.0002482043, 0.0004087228, 0.0005550707, 0.0005871432, 
    0.0006321421, 0.0005507109, 0.0004019248, 0.0002226593, 6.811127e-05,
  2.311882e-06, 2.478574e-06, 4.185862e-06, 5.338048e-06, 1.142507e-05, 
    3.821807e-05, 0.0001464093, 0.0003259385, 0.0005212168, 0.0006405628, 
    0.0006932605, 0.0006178681, 0.0004901646, 0.0003289565, 0.0001563755,
  2.039864e-06, 1.134997e-06, 2.26534e-06, 6.008051e-06, 7.00323e-06, 
    1.65345e-05, 7.07685e-05, 0.0002165035, 0.0004340021, 0.0006146263, 
    0.0006970704, 0.0007195451, 0.0005399333, 0.0003897213, 0.0002616538,
  2.331762e-06, 1.747807e-06, 3.781228e-06, 6.170901e-06, 8.895321e-06, 
    8.935805e-06, 1.695948e-05, 0.0001093675, 0.0002822443, 0.0004781014, 
    0.0006446604, 0.0007264635, 0.00060045, 0.0004412161, 0.0003376643,
  1.781066e-06, 1.032751e-06, 3.112182e-06, 2.921895e-06, 7.091294e-06, 
    6.262204e-06, 7.666378e-06, 2.916789e-05, 0.0001378203, 0.0003066271, 
    0.0005153639, 0.0006718185, 0.0007033007, 0.0005051963, 0.0003961688,
  3.590395e-06, 1.842581e-06, 1.120791e-06, 2.024385e-06, 2.220062e-06, 
    2.655067e-06, 5.948832e-06, 1.338275e-05, 4.745631e-05, 0.0001383992, 
    0.0002781691, 0.0005392462, 0.0006936874, 0.0006441587, 0.000474121,
  5.807914e-06, 4.682592e-06, 2.174415e-06, 2.863323e-06, 1.113922e-06, 
    1.845598e-06, 2.724149e-06, 5.744247e-06, 2.308986e-05, 5.380779e-05, 
    0.0001183682, 0.000244638, 0.0005565084, 0.0006678237, 0.0006155418,
  6.664087e-06, 5.411518e-06, 3.730459e-06, 2.865791e-06, 3.761346e-06, 
    3.749208e-06, 2.512935e-06, 3.193924e-06, 1.39234e-05, 3.621988e-05, 
    5.747988e-05, 9.016284e-05, 0.0001799884, 0.0004846463, 0.0006408201,
  9.257805e-06, 6.720708e-06, 4.119096e-06, 3.173384e-06, 2.952441e-06, 
    3.514763e-06, 2.174835e-06, 1.139169e-06, 2.29967e-06, 1.273536e-05, 
    4.247064e-05, 7.398419e-05, 9.139907e-05, 0.0001610968, 0.0003505635,
  7.594565e-06, 3.612586e-06, 4.139747e-06, 3.15338e-06, 2.097484e-06, 
    1.016048e-06, 2.824387e-07, 2.432676e-07, 4.794366e-07, 7.277594e-07, 
    8.884838e-06, 3.616308e-05, 7.843574e-05, 0.0001088289, 0.0001587153,
  0.0001700033, 0.0002101425, 0.0002624586, 0.0003099173, 0.0003257402, 
    0.0002276821, 7.568435e-05, 8.009257e-06, 2.336618e-06, 3.667829e-06, 
    8.462347e-06, 2.330431e-05, 3.815981e-05, 5.495098e-05, 8.474416e-05,
  0.0001687791, 0.0002439392, 0.0002993704, 0.0003403911, 0.000367846, 
    0.0003430962, 0.0001835864, 4.834805e-05, 5.515263e-06, 3.256872e-06, 
    7.544428e-06, 2.163996e-05, 4.401683e-05, 6.22244e-05, 8.300431e-05,
  0.0001119514, 0.0002392125, 0.0002945686, 0.0003218249, 0.0003552249, 
    0.0003718663, 0.0002754025, 0.0001307251, 2.892381e-05, 3.14164e-06, 
    3.749544e-06, 1.216454e-05, 3.686613e-05, 5.814129e-05, 7.524656e-05,
  4.368388e-05, 0.0001680907, 0.0002437371, 0.0002492139, 0.0002668854, 
    0.0003080943, 0.0003286284, 0.0001999619, 9.801763e-05, 2.035925e-05, 
    2.643418e-06, 4.837689e-06, 1.762066e-05, 4.14203e-05, 6.162921e-05,
  4.926e-06, 4.849603e-05, 0.0001324955, 0.0001648975, 0.000174206, 
    0.0002059138, 0.000270661, 0.0002792739, 0.0001568796, 7.912341e-05, 
    1.665776e-05, 3.004192e-06, 6.37968e-06, 2.273397e-05, 4.867755e-05,
  7.697403e-06, 1.471743e-05, 3.311401e-05, 6.630511e-05, 8.622459e-05, 
    0.0001026429, 0.0001688935, 0.0002471145, 0.0002388762, 0.0001375768, 
    7.953657e-05, 2.180489e-05, 4.228928e-06, 7.128434e-06, 2.762091e-05,
  6.913115e-06, 3.048542e-05, 4.382518e-05, 6.438397e-05, 4.835547e-05, 
    4.612398e-05, 6.860614e-05, 0.0001653124, 0.0002652121, 0.0002404808, 
    0.000140069, 8.606545e-05, 2.747159e-05, 5.392594e-06, 1.016413e-05,
  5.498181e-06, 2.376728e-05, 5.878049e-05, 8.413338e-05, 8.259862e-05, 
    5.836795e-05, 4.208031e-05, 5.448856e-05, 0.0001846294, 0.0002757625, 
    0.0002473514, 0.0001526164, 9.170536e-05, 3.828474e-05, 7.021531e-06,
  4.271481e-06, 3.511946e-06, 1.035082e-05, 3.617893e-05, 6.393273e-05, 
    8.19359e-05, 8.253165e-05, 7.309119e-05, 5.2948e-05, 0.0001795426, 
    0.0002688495, 0.0002503263, 0.000166189, 0.0001033908, 4.787582e-05,
  5.917962e-06, 8.324124e-06, 5.564859e-06, 1.826759e-06, 3.322999e-06, 
    6.533734e-06, 2.981709e-05, 5.675916e-05, 5.580837e-05, 4.671121e-05, 
    0.0001513705, 0.0002461055, 0.0002490725, 0.0001786536, 0.0001250132,
  1.592049e-05, 1.933219e-05, 2.089553e-05, 2.412236e-05, 4.718097e-05, 
    7.41331e-05, 9.245671e-05, 9.295202e-05, 8.049682e-05, 6.478302e-05, 
    4.913731e-05, 2.871959e-05, 2.139101e-05, 2.030456e-05, 2.861802e-05,
  4.232459e-05, 3.157437e-05, 2.441598e-05, 1.907204e-05, 5.080636e-05, 
    8.548661e-05, 0.0001067592, 0.0001177348, 0.0001088092, 8.282581e-05, 
    5.538671e-05, 3.633185e-05, 2.234902e-05, 2.413262e-05, 3.184492e-05,
  0.0001272675, 5.507827e-05, 2.268527e-05, 9.237636e-06, 2.641946e-05, 
    6.550259e-05, 9.522842e-05, 0.0001058577, 0.0001058525, 7.580435e-05, 
    4.609582e-05, 4.368532e-05, 2.981974e-05, 2.009986e-05, 3.402364e-05,
  0.000256362, 0.0001510142, 5.107635e-05, 1.373047e-05, 1.176321e-05, 
    2.673485e-05, 7.342823e-05, 0.0001067441, 0.0001148947, 8.128874e-05, 
    4.22329e-05, 3.111756e-05, 2.433419e-05, 2.817536e-05, 2.994558e-05,
  0.000198983, 0.0002127786, 0.0001197809, 4.215106e-05, 1.729478e-05, 
    9.134854e-06, 2.855229e-05, 9.872386e-05, 0.0001355104, 0.0001098432, 
    6.195041e-05, 3.092536e-05, 1.975575e-05, 2.071421e-05, 1.870815e-05,
  0.0001101104, 9.426031e-05, 8.752591e-05, 6.140608e-05, 4.436243e-05, 
    2.48368e-05, 1.170909e-05, 3.737324e-05, 0.000121037, 0.0001458288, 
    9.566391e-05, 4.251307e-05, 2.682726e-05, 1.669148e-05, 2.258192e-05,
  0.0001996021, 0.0001664161, 0.0001342435, 7.944641e-05, 5.248112e-05, 
    4.928648e-05, 3.281709e-05, 1.328339e-05, 4.182227e-05, 0.0001417055, 
    0.0001355439, 7.961501e-05, 4.468039e-05, 3.136816e-05, 2.136447e-05,
  0.0003237118, 0.0003022891, 0.0002760142, 0.0002219461, 0.000118947, 
    6.980451e-05, 5.410711e-05, 3.885909e-05, 1.788149e-05, 2.345675e-05, 
    0.0001132388, 0.0001172326, 6.257609e-05, 4.107742e-05, 3.403414e-05,
  0.0002530107, 0.0002563643, 0.0003059705, 0.0003150484, 0.0002672667, 
    0.0001994921, 0.0001402348, 9.241774e-05, 5.68757e-05, 2.760821e-05, 
    2.037355e-05, 6.451849e-05, 8.135125e-05, 5.155688e-05, 3.945762e-05,
  9.927136e-05, 0.0001181028, 0.0001609327, 0.0002164645, 0.0002414731, 
    0.0002355414, 0.0002312044, 0.0002222387, 0.0001788946, 0.0001119108, 
    6.041845e-05, 4.6275e-05, 4.205098e-05, 4.943215e-05, 4.274381e-05,
  5.019445e-05, 6.072061e-05, 6.469595e-05, 4.770034e-05, 2.139583e-05, 
    2.357364e-05, 2.837866e-05, 3.396636e-05, 3.545289e-05, 2.965389e-05, 
    2.331216e-05, 2.052158e-05, 1.711352e-05, 1.264686e-05, 1.251875e-05,
  2.989564e-05, 6.438301e-05, 0.0001071415, 9.091455e-05, 3.924458e-05, 
    2.026314e-05, 2.555213e-05, 4.059887e-05, 4.91739e-05, 4.70742e-05, 
    3.869643e-05, 3.099974e-05, 2.335247e-05, 1.60142e-05, 1.549171e-05,
  1.738826e-05, 3.312478e-05, 9.346049e-05, 0.0001291094, 7.033814e-05, 
    3.182098e-05, 2.390025e-05, 3.431454e-05, 4.562272e-05, 5.558e-05, 
    6.169559e-05, 6.05301e-05, 4.744008e-05, 3.271757e-05, 2.082685e-05,
  3.414884e-05, 1.409157e-05, 4.870803e-05, 0.0001139567, 0.0001148451, 
    6.182405e-05, 3.696336e-05, 2.76085e-05, 3.232918e-05, 4.550565e-05, 
    5.934514e-05, 6.0873e-05, 5.596539e-05, 4.021599e-05, 3.131698e-05,
  6.371542e-05, 2.890402e-05, 2.234309e-05, 7.579738e-05, 0.0001180831, 
    8.821456e-05, 7.369334e-05, 4.123109e-05, 3.783372e-05, 2.497761e-05, 
    3.376575e-05, 3.837926e-05, 4.326055e-05, 4.091397e-05, 3.709532e-05,
  9.633353e-05, 5.270487e-05, 4.012807e-05, 4.549661e-05, 9.158099e-05, 
    9.531753e-05, 5.843345e-05, 7.957056e-05, 6.527207e-05, 2.349926e-05, 
    1.632484e-05, 2.229325e-05, 2.400422e-05, 3.147328e-05, 3.50684e-05,
  0.000247955, 0.0001108286, 5.033232e-05, 4.39776e-05, 5.247762e-05, 
    0.0001179781, 9.589988e-05, 7.24272e-05, 0.000114827, 0.0001006112, 
    2.808692e-05, 1.965821e-05, 2.453302e-05, 3.132614e-05, 1.784754e-05,
  0.0002814569, 0.0002408939, 0.00013735, 6.908051e-05, 5.626192e-05, 
    8.290654e-05, 0.0001407928, 0.0001241431, 8.818909e-05, 0.0001231036, 
    0.000136762, 0.00010258, 4.730156e-05, 7.992442e-05, 7.472136e-05,
  0.0002464348, 0.0002787677, 0.0002470758, 0.0001539372, 7.498698e-05, 
    5.799828e-05, 8.773544e-05, 0.0001313033, 0.0001164568, 8.233768e-05, 
    9.831871e-05, 0.0001422035, 0.0001926259, 0.0002638064, 0.0002503224,
  0.0002256185, 0.0002906702, 0.0003235613, 0.0002657978, 0.0001652832, 
    0.0001007488, 6.625133e-05, 7.091487e-05, 9.710754e-05, 0.0001072863, 
    7.336382e-05, 5.468506e-05, 0.0001409101, 0.0002551615, 0.0003171577,
  3.25039e-05, 2.928869e-05, 2.069474e-05, 1.830361e-05, 1.901857e-05, 
    1.966172e-05, 1.793927e-05, 1.465007e-05, 1.62519e-05, 1.252302e-05, 
    8.613229e-06, 6.172019e-06, 4.627828e-06, 3.137577e-06, 1.341642e-06,
  2.747853e-05, 2.483464e-05, 2.828819e-05, 3.66879e-05, 2.629876e-05, 
    3.077903e-05, 2.612766e-05, 2.14741e-05, 1.654121e-05, 1.21608e-05, 
    1.07067e-05, 8.58513e-06, 7.138821e-06, 4.83647e-06, 2.932304e-06,
  1.712756e-05, 1.828955e-05, 2.292237e-05, 3.324509e-05, 4.286396e-05, 
    3.826172e-05, 4.059078e-05, 3.659731e-05, 2.22604e-05, 1.368648e-05, 
    1.197127e-05, 1.134351e-05, 8.923147e-06, 6.907361e-06, 5.112033e-06,
  1.18242e-05, 1.575842e-05, 2.433358e-05, 2.786728e-05, 4.082331e-05, 
    3.757735e-05, 4.021233e-05, 2.423423e-05, 1.599579e-05, 1.313032e-05, 
    1.225609e-05, 1.032099e-05, 7.875071e-06, 8.035417e-06, 6.349588e-06,
  8.405719e-06, 1.064947e-05, 2.272859e-05, 2.091472e-05, 3.505468e-05, 
    4.437812e-05, 3.066318e-05, 2.548298e-05, 2.172266e-05, 2.970973e-05, 
    2.795957e-05, 1.631423e-05, 7.751512e-06, 7.788557e-06, 6.530613e-06,
  3.311837e-06, 4.997334e-06, 1.423214e-05, 2.453676e-05, 2.781796e-05, 
    3.064302e-05, 2.502902e-05, 1.890218e-05, 4.465362e-05, 0.0001141441, 
    0.0001276864, 0.0001098673, 3.986676e-05, 9.16175e-06, 7.390939e-06,
  2.990209e-06, 2.914066e-06, 6.257232e-06, 1.778999e-05, 3.181159e-05, 
    2.684522e-05, 1.391501e-05, 1.786037e-05, 5.430863e-05, 0.00015078, 
    0.0001444954, 0.0001673114, 0.0001425797, 5.608058e-05, 1.001543e-05,
  8.72571e-06, 7.87887e-06, 7.988315e-06, 9.782349e-06, 2.160442e-05, 
    1.726374e-05, 1.261142e-05, 9.056744e-06, 2.074622e-05, 5.636853e-05, 
    8.926999e-05, 0.0001237297, 0.0001775355, 0.0001113678, 1.455597e-05,
  6.462414e-05, 1.579655e-05, 8.215252e-06, 1.479118e-05, 1.474344e-05, 
    1.689813e-05, 8.637475e-06, 3.94359e-06, 7.333587e-06, 9.022229e-06, 
    2.209533e-05, 3.793146e-05, 0.0001314255, 0.0001669196, 4.484804e-05,
  0.000151334, 3.425794e-05, 1.096215e-05, 7.09897e-06, 1.099433e-05, 
    1.101365e-05, 9.983313e-06, 4.70912e-06, 5.350518e-06, 2.815155e-06, 
    3.565131e-06, 1.479499e-05, 4.606425e-05, 0.0001515638, 0.0001082572,
  4.710621e-06, 2.662739e-06, 2.837665e-06, 1.852286e-06, 1.733597e-06, 
    1.591967e-06, 1.012668e-06, 6.093331e-07, 1.841993e-07, 4.462463e-08, 
    7.093283e-08, 7.813223e-07, 5.439783e-07, 3.668322e-06, 4.933361e-06,
  8.19271e-06, 5.629518e-06, 5.15482e-06, 5.727355e-06, 5.176e-06, 
    3.391614e-06, 2.190782e-06, 1.47865e-06, 1.090984e-06, 4.762198e-07, 
    1.187629e-07, 3.461592e-07, 1.116335e-06, 8.808622e-07, 3.265896e-06,
  1.201842e-05, 8.701005e-06, 1.068805e-05, 8.323482e-06, 6.82521e-06, 
    6.866014e-06, 4.801653e-06, 5.222545e-06, 2.30088e-06, 2.362014e-06, 
    1.279128e-06, 8.086987e-07, 2.713075e-07, 1.00385e-06, 2.045029e-06,
  1.780441e-05, 1.508937e-05, 2.232921e-05, 1.243016e-05, 9.045511e-06, 
    9.241307e-06, 9.353166e-06, 5.919783e-06, 4.36284e-06, 4.135558e-06, 
    3.057567e-06, 2.118416e-06, 1.614153e-06, 1.273176e-06, 2.895816e-06,
  1.98389e-05, 2.00809e-05, 1.694763e-05, 1.968303e-05, 1.544287e-05, 
    1.165481e-05, 9.707967e-06, 7.96544e-06, 5.281972e-06, 4.263322e-06, 
    4.367832e-06, 3.648819e-06, 3.129476e-06, 1.3171e-06, 6.403044e-07,
  2.128363e-05, 1.45562e-05, 1.582083e-05, 2.077778e-05, 2.16981e-05, 
    1.732033e-05, 1.370104e-05, 1.225234e-05, 6.364566e-06, 6.476941e-06, 
    4.057016e-06, 3.855764e-06, 3.17324e-06, 3.568075e-06, 4.679295e-06,
  1.756462e-05, 1.220116e-05, 2.102612e-05, 1.554702e-05, 1.938075e-05, 
    2.399921e-05, 2.375757e-05, 2.072367e-05, 1.503408e-05, 8.81845e-06, 
    6.568144e-06, 6.911612e-06, 1.678315e-06, 1.999291e-06, 2.323087e-06,
  1.109245e-05, 1.622477e-05, 2.841843e-05, 1.756008e-05, 1.450767e-05, 
    1.386485e-05, 1.870155e-05, 1.892174e-05, 2.023537e-05, 2.013577e-05, 
    1.625771e-05, 9.700232e-06, 6.111883e-06, 2.91907e-06, 3.397514e-06,
  8.802924e-06, 1.326486e-05, 7.953134e-06, 1.340518e-05, 8.927806e-06, 
    8.485286e-06, 1.392655e-05, 2.173572e-05, 2.587624e-05, 2.654919e-05, 
    2.481253e-05, 2.507027e-05, 1.606411e-05, 6.087537e-06, 5.42929e-06,
  1.258311e-05, 1.176765e-05, 1.016621e-05, 1.022822e-05, 1.627362e-05, 
    4.806062e-06, 6.363077e-06, 1.84203e-05, 2.051015e-05, 2.293916e-05, 
    1.944616e-05, 2.283012e-05, 2.719806e-05, 3.055658e-05, 1.410849e-05,
  2.54693e-07, 1.609546e-07, 1.793441e-07, 9.073005e-09, 2.739156e-07, 
    1.830418e-06, 4.468879e-06, 7.876664e-06, 1.210519e-05, 1.79235e-05, 
    1.55874e-05, 1.572984e-05, 1.322001e-05, 1.191318e-05, 9.192834e-06,
  1.256543e-06, 6.364693e-07, 4.101188e-07, 2.451292e-07, 9.928376e-08, 
    3.722054e-06, 9.497519e-06, 8.800496e-06, 1.394026e-05, 1.956917e-05, 
    1.983357e-05, 1.699302e-05, 1.89032e-05, 2.205602e-05, 2.140746e-05,
  3.667513e-06, 2.588062e-06, 1.451868e-06, 1.096568e-06, 7.07024e-07, 
    1.583e-06, 1.291204e-05, 1.455297e-05, 1.89911e-05, 2.299354e-05, 
    2.654994e-05, 2.536887e-05, 2.897394e-05, 3.351191e-05, 3.521989e-05,
  5.977935e-06, 4.223391e-06, 2.710994e-06, 2.061882e-06, 9.774019e-07, 
    5.83138e-07, 1.028691e-05, 2.362569e-05, 2.472556e-05, 3.182273e-05, 
    3.346575e-05, 3.940981e-05, 5.021285e-05, 6.271955e-05, 7.012442e-05,
  6.510736e-06, 5.105298e-06, 4.078434e-06, 3.380376e-06, 2.018544e-06, 
    2.015763e-06, 7.952748e-06, 3.225745e-05, 4.55085e-05, 4.929003e-05, 
    5.60361e-05, 7.759828e-05, 0.000115169, 0.0001321348, 0.000125366,
  7.000815e-06, 4.715669e-06, 4.791092e-06, 2.796736e-06, 3.081258e-06, 
    2.349126e-06, 5.983717e-06, 2.783491e-05, 6.280661e-05, 7.389866e-05, 
    9.001768e-05, 0.0001349356, 0.000187742, 0.0002039697, 0.0001665174,
  1.180495e-05, 7.074197e-06, 5.542922e-06, 4.029402e-06, 3.256769e-06, 
    3.270603e-06, 5.711253e-06, 1.910295e-05, 5.49989e-05, 0.0001036471, 
    0.0001331435, 0.0001749049, 0.0002268821, 0.0002370786, 0.0001904962,
  1.644102e-05, 1.257663e-05, 1.071319e-05, 8.920842e-06, 5.620059e-06, 
    3.680404e-06, 4.154801e-06, 1.150601e-05, 2.944705e-05, 8.3417e-05, 
    0.0001418625, 0.0001912426, 0.0002229135, 0.0002304837, 0.0002179023,
  1.5472e-05, 1.333111e-05, 1.204421e-05, 1.131292e-05, 1.089842e-05, 
    8.303875e-06, 5.205102e-06, 4.217701e-06, 9.392079e-06, 3.481848e-05, 
    8.805721e-05, 0.0001522832, 0.0001911066, 0.0002021841, 0.0002343024,
  1.745961e-05, 1.15769e-05, 1.166484e-05, 9.356733e-06, 8.763414e-06, 
    8.757211e-06, 1.064876e-05, 7.172374e-06, 3.766344e-06, 3.747954e-06, 
    1.455279e-05, 4.306766e-05, 9.050985e-05, 0.0001342644, 0.0001915431,
  6.627716e-06, 6.1625e-06, 8.364368e-06, 1.288197e-05, 7.680229e-06, 
    4.318675e-06, 9.081712e-07, 7.48964e-08, 1.286347e-07, 7.399459e-08, 
    6.352985e-08, 8.61707e-08, 7.575227e-08, 1.101117e-08, 3.584584e-07,
  7.157467e-06, 8.940407e-06, 1.358728e-05, 1.085485e-05, 1.171402e-05, 
    1.003696e-05, 1.248214e-06, 2.522407e-07, 1.639642e-07, 3.175255e-07, 
    1.410448e-07, 1.303535e-07, 6.380506e-08, 4.187489e-07, 1.112452e-08,
  8.427728e-06, 7.941847e-06, 1.13506e-05, 1.302499e-05, 1.374871e-05, 
    1.42195e-05, 5.677552e-06, 9.267358e-07, 6.241573e-07, 5.297218e-07, 
    6.378492e-07, 4.377659e-07, 4.850961e-07, 3.041718e-07, 3.165598e-07,
  4.890082e-06, 8.863901e-06, 9.699534e-06, 7.127283e-06, 1.088253e-05, 
    2.248493e-05, 1.769597e-05, 3.113123e-06, 1.908611e-06, 1.809724e-06, 
    2.413787e-06, 1.74354e-06, 1.025354e-06, 5.89657e-07, 4.246746e-07,
  5.92923e-06, 5.986669e-06, 7.474458e-06, 1.089476e-05, 1.694179e-05, 
    2.367883e-05, 2.944911e-05, 1.46327e-05, 5.812905e-06, 6.606675e-06, 
    6.082416e-06, 4.478137e-06, 2.523157e-06, 2.106045e-06, 7.049719e-07,
  4.317226e-06, 7.063052e-06, 9.771354e-06, 1.651381e-05, 2.325493e-05, 
    2.919041e-05, 3.37337e-05, 3.434213e-05, 1.983393e-05, 1.453671e-05, 
    8.55581e-06, 1.481755e-05, 1.370696e-05, 8.556266e-06, 4.969102e-06,
  5.145903e-06, 1.221352e-05, 1.057714e-05, 1.149392e-05, 2.173547e-05, 
    2.873564e-05, 3.799089e-05, 5.285001e-05, 4.040104e-05, 2.814475e-05, 
    2.561284e-05, 2.920298e-05, 2.353771e-05, 2.37006e-05, 2.783721e-05,
  3.613568e-06, 7.736796e-06, 1.489017e-05, 1.384566e-05, 1.682993e-05, 
    2.774243e-05, 3.926328e-05, 4.554956e-05, 5.470087e-05, 4.404298e-05, 
    2.85582e-05, 2.59938e-05, 2.544464e-05, 3.824372e-05, 9.237946e-05,
  3.530681e-06, 4.197112e-06, 1.089305e-05, 1.291211e-05, 1.778168e-05, 
    1.528869e-05, 3.25515e-05, 4.87813e-05, 5.033845e-05, 5.530774e-05, 
    4.154432e-05, 3.308917e-05, 2.273274e-05, 3.292902e-05, 9.147456e-05,
  2.577468e-06, 3.78092e-06, 7.877338e-06, 9.41824e-06, 1.86731e-05, 
    1.90413e-05, 2.082909e-05, 2.909712e-05, 6.05287e-05, 5.798074e-05, 
    5.725895e-05, 4.765935e-05, 4.568962e-05, 7.348884e-05, 0.000202286,
  7.311012e-13, 1.297437e-10, 1.787194e-09, 8.558591e-09, 1.97274e-08, 
    1.283209e-07, 4.56487e-07, 1.415436e-06, 3.475966e-06, 4.041068e-06, 
    4.329151e-06, 3.008443e-06, 5.783275e-06, 5.101562e-06, 7.216333e-06,
  2.632012e-09, 1.634238e-08, 5.581565e-09, 1.436244e-08, 8.726927e-09, 
    3.802342e-07, 4.565828e-07, 2.245602e-06, 2.155308e-06, 2.634087e-06, 
    4.871253e-06, 6.161826e-06, 6.621324e-06, 7.60543e-06, 6.384219e-06,
  8.264972e-09, 2.20774e-07, 6.874507e-07, 9.003471e-07, 1.297742e-06, 
    2.099758e-06, 1.902394e-06, 1.636801e-06, 1.206882e-06, 2.746166e-06, 
    4.365445e-06, 5.165781e-06, 6.088566e-06, 5.123458e-06, 2.410982e-06,
  1.380989e-08, 1.490722e-07, 2.158196e-07, 1.495332e-07, 1.137795e-08, 
    4.610997e-07, 4.528016e-07, 5.394487e-07, 7.890077e-07, 1.744985e-06, 
    2.272834e-06, 3.260177e-06, 4.467914e-06, 3.61227e-06, 5.463744e-06,
  7.924043e-10, 3.221512e-09, 1.452735e-08, 6.00857e-09, 5.445027e-07, 
    7.869106e-07, 1.16002e-06, 1.749457e-06, 1.558187e-06, 2.604257e-06, 
    2.257837e-06, 1.080623e-06, 1.959884e-06, 2.299369e-06, 4.844335e-06,
  2.462598e-09, 5.054884e-09, 1.539872e-09, 9.273484e-07, 1.100928e-06, 
    3.126988e-06, 2.666074e-06, 2.878041e-06, 2.337835e-06, 2.474303e-06, 
    2.862124e-06, 2.693805e-06, 2.425425e-06, 4.499035e-06, 3.407039e-06,
  4.199247e-07, 1.147157e-09, 8.45683e-07, 9.797494e-07, 2.980696e-06, 
    4.092998e-06, 4.524169e-06, 4.174442e-06, 3.617093e-06, 3.295603e-06, 
    5.200564e-06, 3.97345e-06, 1.835816e-06, 3.541803e-06, 5.228126e-06,
  9.833968e-07, 1.459265e-08, 6.460093e-07, 2.969153e-06, 4.883098e-06, 
    5.546539e-06, 6.682052e-06, 6.517837e-06, 5.731462e-06, 9.89019e-06, 
    5.023363e-06, 2.544585e-06, 2.730196e-06, 4.022603e-06, 3.88934e-06,
  1.961523e-06, 6.000094e-08, 1.025845e-06, 3.976301e-06, 6.31751e-06, 
    7.185882e-06, 6.824727e-06, 6.709045e-06, 7.601953e-06, 3.138426e-06, 
    5.631373e-06, 7.943587e-06, 5.455865e-06, 3.501336e-06, 4.830974e-06,
  1.994931e-06, 5.341722e-07, 2.10603e-06, 4.333821e-06, 7.31734e-06, 
    9.244123e-06, 9.524249e-06, 7.273435e-06, 6.88358e-06, 5.76326e-06, 
    8.97579e-06, 7.809177e-06, 5.728317e-06, 4.250131e-06, 3.555376e-06,
  9.81878e-08, 2.988748e-08, 1.203974e-07, 2.356517e-08, 8.129986e-07, 
    6.100075e-07, 3.46082e-06, 1.069737e-06, 9.592566e-07, 2.474653e-06, 
    4.915672e-06, 6.051267e-06, 7.76214e-06, 4.56071e-06, 1.806329e-05,
  2.151644e-08, 6.100994e-08, 5.763249e-08, 5.301762e-08, 2.042039e-06, 
    1.528917e-06, 1.570435e-06, 1.814135e-06, 1.002954e-06, 2.248207e-07, 
    2.430026e-06, 3.508714e-06, 9.723668e-06, 7.919858e-06, 2.988068e-05,
  1.801183e-08, 1.24767e-07, 6.164978e-08, 1.731382e-07, 1.565982e-07, 
    5.177146e-07, 2.620599e-06, 4.48153e-06, 1.283455e-06, 5.546573e-07, 
    3.805806e-07, 2.578197e-06, 7.428626e-06, 8.235475e-06, 3.852626e-05,
  7.369953e-07, 1.39019e-07, 3.138362e-08, 1.017433e-07, 4.926207e-08, 
    5.222106e-07, 3.857755e-06, 6.013753e-06, 3.176987e-06, 6.692188e-07, 
    5.583137e-08, 8.429814e-07, 2.754746e-06, 4.990198e-06, 3.90964e-05,
  1.381356e-06, 7.645806e-08, 1.213989e-07, 1.013655e-06, 2.175124e-06, 
    1.406057e-06, 4.796393e-06, 6.714839e-06, 5.894208e-06, 3.073143e-06, 
    1.064069e-07, 1.233507e-07, 7.660338e-07, 2.37274e-06, 4.420322e-05,
  2.055409e-07, 5.115198e-08, 3.500369e-07, 1.303341e-06, 1.787551e-06, 
    1.376541e-06, 2.924241e-06, 5.479035e-06, 7.052689e-06, 1.876438e-06, 
    7.470888e-07, 6.382677e-08, 1.023941e-07, 6.422631e-07, 4.330004e-05,
  8.821287e-09, 1.418146e-07, 2.286526e-07, 1.095775e-06, 4.302902e-07, 
    1.055524e-06, 1.79687e-06, 2.404407e-06, 3.194591e-06, 1.982459e-06, 
    5.462473e-07, 6.242971e-07, 5.574844e-07, 1.149239e-06, 5.027801e-05,
  2.235178e-08, 2.351323e-06, 3.18248e-07, 1.462381e-06, 5.44423e-07, 
    5.491524e-07, 1.762414e-06, 8.60823e-07, 3.277678e-06, 2.600912e-06, 
    4.153818e-07, 2.592936e-06, 2.495855e-06, 2.095692e-06, 6.430256e-05,
  4.096604e-08, 7.092243e-07, 8.048855e-07, 1.831437e-06, 1.042243e-06, 
    6.342341e-07, 8.083371e-07, 1.040551e-06, 2.081395e-06, 1.213675e-06, 
    1.26149e-06, 2.094281e-06, 3.355613e-06, 4.836251e-06, 8.362115e-05,
  4.767657e-07, 1.747912e-06, 1.433392e-06, 1.080747e-06, 8.684332e-07, 
    8.345277e-07, 1.011371e-06, 9.359806e-07, 9.808535e-07, 1.473343e-06, 
    2.475429e-06, 6.232413e-07, 2.234499e-06, 1.998345e-05, 0.0001028845,
  2.384863e-05, 1.482446e-05, 1.189337e-05, 4.472237e-06, 1.233138e-06, 
    1.327289e-06, 3.47242e-06, 3.573507e-06, 1.122303e-05, 1.345451e-05, 
    9.213256e-06, 5.206125e-06, 6.061822e-06, 1.094445e-05, 9.318254e-06,
  2.910284e-05, 2.702437e-05, 2.154841e-05, 1.038444e-05, 5.877737e-06, 
    1.781603e-06, 2.655e-06, 4.341551e-06, 3.758962e-06, 9.073964e-06, 
    9.59833e-06, 5.391855e-06, 3.739657e-06, 5.770928e-06, 6.573191e-06,
  3.000409e-05, 2.984927e-05, 1.888794e-05, 1.454744e-05, 7.66334e-06, 
    3.011135e-06, 2.590665e-06, 3.38406e-06, 6.464253e-07, 5.290372e-06, 
    1.008206e-05, 5.686405e-06, 4.891381e-06, 4.775024e-06, 7.537936e-06,
  2.896389e-05, 1.336598e-05, 9.285495e-06, 9.255123e-06, 4.715324e-06, 
    3.029342e-06, 2.442667e-06, 3.922316e-06, 1.117924e-07, 1.749504e-06, 
    5.208751e-06, 3.350479e-06, 4.253944e-06, 5.786513e-06, 6.313766e-06,
  8.461651e-06, 2.963453e-06, 3.941123e-06, 5.394106e-06, 4.129049e-06, 
    6.587668e-06, 8.907494e-06, 7.781626e-06, 1.663076e-07, 2.279084e-09, 
    2.998183e-06, 2.731051e-06, 3.832647e-06, 3.693772e-06, 6.328691e-06,
  2.187425e-06, 1.821114e-06, 3.27006e-06, 4.520094e-06, 7.039518e-06, 
    6.926967e-06, 1.112123e-05, 1.198736e-05, 2.169818e-06, 3.184683e-09, 
    1.155836e-06, 1.1406e-06, 2.336269e-06, 2.558812e-06, 1.515907e-05,
  2.556841e-06, 3.154381e-06, 5.260963e-06, 3.450808e-06, 5.230718e-06, 
    7.598546e-06, 1.137818e-05, 9.760543e-06, 1.96956e-06, 1.1237e-09, 
    7.619319e-07, 6.398924e-07, 1.363028e-06, 1.328009e-06, 4.270038e-05,
  5.255833e-06, 4.08766e-06, 4.533736e-06, 6.81747e-06, 3.536652e-06, 
    4.479831e-06, 6.903571e-06, 9.728094e-06, 5.628318e-06, 3.393979e-07, 
    8.890486e-08, 4.044053e-07, 1.881053e-06, 3.525324e-06, 0.0001091435,
  3.790448e-06, 3.995569e-06, 3.832096e-06, 8.732826e-06, 7.26476e-06, 
    3.297505e-06, 5.183654e-06, 5.235907e-06, 5.318801e-06, 1.478595e-06, 
    2.66747e-09, 2.345362e-07, 3.948302e-06, 3.722204e-05, 0.0002198142,
  2.886309e-06, 2.715109e-06, 5.604245e-06, 3.525942e-06, 2.466955e-06, 
    1.605649e-06, 4.774602e-06, 3.809378e-06, 1.31566e-06, 1.259977e-06, 
    1.494933e-09, 1.159909e-08, 5.228989e-06, 5.582192e-05, 0.0002933239,
  6.223028e-06, 1.126559e-05, 1.682072e-05, 1.797479e-05, 6.019281e-06, 
    1.249099e-06, 1.229255e-06, 9.942451e-05, 0.0001820136, 0.0001844435, 
    0.0001824014, 0.0001777128, 0.0001605226, 0.0001003859, 3.298422e-05,
  8.577564e-07, 7.973334e-06, 1.426581e-05, 1.394143e-05, 8.359146e-06, 
    3.357139e-06, 1.494759e-06, 8.733891e-05, 0.0002312113, 0.0002897131, 
    0.000322856, 0.0003027547, 0.0002307318, 0.0001134125, 3.074278e-05,
  1.383485e-06, 3.420065e-07, 7.494262e-06, 9.379352e-06, 1.489718e-05, 
    8.669743e-06, 4.790799e-06, 3.262251e-05, 0.0001903656, 0.0003347444, 
    0.0003884406, 0.0003795056, 0.0002743105, 0.0001123951, 2.397172e-05,
  2.283004e-06, 4.858691e-07, 2.334422e-06, 5.17841e-06, 1.715347e-05, 
    2.149611e-05, 3.506208e-06, 5.286116e-06, 7.9578e-05, 0.0002516485, 
    0.0003521022, 0.0003608541, 0.0002579849, 9.176401e-05, 2.016979e-05,
  2.689941e-06, 1.506759e-06, 3.881084e-06, 6.363428e-06, 7.886311e-06, 
    1.242576e-05, 3.461957e-06, 1.163823e-06, 1.232409e-05, 7.817594e-05, 
    0.0001991968, 0.0002652275, 0.0001935155, 5.783137e-05, 1.246059e-05,
  2.922661e-06, 3.617875e-06, 2.801486e-06, 1.189317e-06, 2.070859e-06, 
    6.120212e-06, 7.183069e-06, 2.879259e-06, 1.049281e-06, 1.217854e-05, 
    2.88694e-05, 8.642924e-05, 0.0001083976, 4.159964e-05, 1.463193e-05,
  6.304402e-06, 5.541965e-06, 4.73022e-06, 2.422171e-06, 3.742679e-06, 
    4.618297e-06, 4.22693e-06, 2.308489e-06, 1.640404e-07, 2.225108e-06, 
    6.182646e-06, 2.403786e-05, 9.386456e-05, 5.999869e-05, 2.087023e-05,
  3.090911e-06, 7.790986e-06, 6.736526e-06, 6.011384e-06, 4.095378e-06, 
    4.95169e-06, 3.577568e-06, 3.197875e-06, 8.233903e-07, 7.490248e-07, 
    3.062e-06, 2.456124e-05, 0.0001051526, 8.97158e-05, 2.748022e-05,
  4.825073e-06, 5.1904e-06, 4.761855e-06, 8.215909e-06, 5.256511e-06, 
    4.426446e-06, 5.038401e-06, 5.785024e-06, 1.336899e-06, 6.29379e-08, 
    6.373139e-07, 2.598759e-05, 0.0001162518, 0.0001142495, 2.901785e-05,
  5.741799e-06, 6.426628e-06, 2.829019e-06, 5.402327e-06, 6.428394e-06, 
    4.618329e-06, 6.651683e-06, 4.434055e-06, 9.507997e-07, 9.293775e-09, 
    4.702605e-07, 2.161306e-05, 0.0001356658, 0.0001440574, 4.148939e-05,
  2.487465e-06, 2.397567e-07, 6.287343e-08, 4.158636e-06, 8.651869e-06, 
    4.358459e-06, 3.241845e-05, 6.266328e-05, 8.001766e-06, 3.905282e-06, 
    3.232054e-06, 7.783946e-06, 1.85169e-05, 2.367553e-05, 2.688107e-05,
  2.844484e-06, 6.335061e-07, 3.490128e-07, 2.025362e-06, 7.435295e-06, 
    1.291558e-05, 3.218296e-05, 3.259911e-05, 2.422126e-05, 1.371853e-05, 
    9.393303e-06, 6.43884e-06, 8.397132e-06, 4.24531e-05, 4.241627e-05,
  2.390005e-06, 3.547975e-07, 1.127847e-07, 3.668446e-06, 3.179088e-06, 
    9.114395e-06, 7.266317e-06, 1.895558e-05, 1.801952e-05, 1.155794e-05, 
    6.173927e-06, 1.046053e-05, 5.168325e-05, 8.92969e-05, 5.162938e-05,
  1.734934e-06, 1.222027e-06, 1.082496e-07, 5.89571e-08, 4.900518e-07, 
    9.941915e-06, 3.408974e-06, 1.111082e-05, 1.187489e-05, 6.627756e-06, 
    2.480592e-06, 1.064917e-05, 9.177716e-05, 0.0001203594, 3.9874e-05,
  2.611437e-06, 2.155659e-06, 7.828655e-07, 9.321512e-08, 3.996688e-06, 
    9.64554e-06, 5.76409e-06, 1.211309e-05, 1.68963e-05, 7.908731e-06, 
    6.779251e-06, 4.030869e-05, 0.0001565665, 0.000116971, 1.634657e-05,
  1.869455e-06, 3.536355e-06, 4.292067e-06, 1.217065e-06, 3.12184e-06, 
    5.750655e-06, 7.917012e-06, 1.323171e-05, 1.691007e-05, 1.066111e-05, 
    7.966182e-06, 0.000154482, 0.0002455467, 8.747616e-05, 6.779996e-06,
  2.535606e-06, 1.660768e-06, 2.623241e-06, 1.117851e-06, 4.086146e-07, 
    6.054338e-06, 8.674267e-06, 1.293748e-05, 1.009136e-05, 7.760649e-06, 
    5.929502e-05, 0.0002355186, 0.0002565087, 2.765934e-05, 5.527852e-06,
  4.734025e-06, 5.16239e-06, 4.495384e-06, 4.382128e-06, 2.364396e-06, 
    5.695368e-06, 1.002274e-05, 1.236732e-05, 9.265012e-06, 5.884959e-06, 
    8.36844e-05, 0.0002207989, 0.0001275209, 8.764273e-06, 5.157898e-06,
  2.647994e-06, 3.959497e-06, 5.258891e-06, 5.026253e-06, 2.22775e-06, 
    3.920855e-06, 1.001925e-05, 1.369298e-05, 9.153014e-06, 9.458045e-06, 
    5.920994e-05, 0.0001031902, 1.458868e-05, 8.614369e-06, 5.852259e-06,
  5.083168e-06, 3.699036e-06, 4.761931e-06, 4.793094e-06, 4.104025e-06, 
    3.898423e-06, 7.783655e-06, 1.405476e-05, 9.814148e-06, 9.124463e-06, 
    1.571653e-05, 1.73842e-05, 2.420875e-05, 9.749439e-06, 7.021213e-06,
  4.486198e-06, 3.853991e-06, 4.126079e-06, 5.539747e-06, 3.293952e-06, 
    1.801813e-06, 1.353284e-06, 1.094917e-06, 1.206951e-07, 1.637349e-06, 
    4.144809e-05, 0.0001057701, 7.984052e-05, 2.547149e-05, 8.450508e-06,
  5.333735e-06, 3.685377e-06, 3.633259e-06, 5.739984e-06, 2.345103e-06, 
    1.759152e-06, 2.955625e-06, 9.469724e-07, 1.001355e-06, 4.380898e-08, 
    1.214318e-05, 4.848031e-05, 4.395132e-05, 2.323451e-05, 1.567304e-05,
  4.985263e-06, 3.021007e-06, 1.181676e-06, 2.985483e-06, 3.360387e-06, 
    3.923314e-06, 3.330222e-06, 2.192499e-06, 2.185103e-07, 8.067298e-07, 
    1.861393e-06, 1.880751e-05, 2.79979e-05, 3.303853e-05, 2.388351e-05,
  3.435967e-06, 3.103005e-06, 2.279678e-06, 3.051785e-06, 2.969965e-06, 
    3.280865e-06, 4.531973e-06, 9.453402e-07, 1.486224e-07, 6.247064e-07, 
    7.411713e-07, 4.868406e-06, 1.636773e-05, 3.985009e-05, 3.250166e-05,
  3.754887e-06, 4.356673e-06, 3.235531e-06, 5.363042e-06, 3.023447e-06, 
    2.752239e-06, 1.105063e-06, 4.415683e-06, 4.357797e-07, 1.275586e-06, 
    1.651229e-06, 4.576381e-06, 1.004434e-05, 4.080658e-05, 3.982496e-05,
  3.33713e-06, 5.90307e-06, 5.50624e-06, 4.367992e-06, 3.119859e-06, 
    2.713391e-06, 1.438409e-06, 4.040868e-06, 6.455282e-06, 1.508866e-06, 
    2.552909e-06, 6.125815e-06, 5.254782e-06, 2.739382e-05, 4.198836e-05,
  4.157127e-06, 4.217029e-06, 5.562416e-06, 4.97794e-06, 3.103405e-06, 
    2.660599e-06, 9.442551e-07, 4.448421e-06, 8.275506e-06, 4.498919e-06, 
    3.215056e-06, 6.806308e-06, 5.042661e-06, 1.307475e-05, 4.314888e-05,
  4.653389e-06, 3.143718e-06, 2.885398e-06, 5.44892e-06, 2.133319e-06, 
    1.164557e-06, 2.211819e-06, 4.954692e-06, 7.121111e-06, 9.434848e-06, 
    5.780356e-06, 1.38576e-05, 9.695148e-06, 6.166095e-06, 3.915546e-05,
  2.785401e-06, 5.368121e-06, 2.97412e-06, 2.397402e-06, 1.294229e-06, 
    5.958883e-07, 2.283223e-06, 6.441357e-06, 8.475009e-06, 1.21181e-05, 
    1.309515e-05, 3.064393e-05, 9.698224e-06, 6.637897e-06, 3.203048e-05,
  2.493359e-06, 3.631925e-06, 2.093369e-06, 2.201326e-06, 6.436121e-07, 
    1.246054e-06, 2.902547e-06, 6.354106e-06, 6.119355e-06, 1.685259e-05, 
    2.392756e-05, 1.736245e-05, 8.497758e-06, 7.679772e-06, 1.98106e-05,
  2.610382e-06, 2.754109e-06, 2.520697e-06, 3.552184e-06, 3.955085e-06, 
    1.777598e-06, 2.592636e-06, 2.145432e-06, 1.599532e-06, 4.166945e-07, 
    7.444208e-07, 2.374694e-06, 4.378635e-06, 2.978746e-06, 3.052518e-06,
  2.297476e-06, 3.159212e-06, 3.333256e-06, 3.789162e-06, 4.799561e-06, 
    3.285239e-06, 3.970201e-06, 1.238031e-06, 1.112417e-06, 9.21003e-07, 
    2.31183e-07, 1.636405e-06, 6.5727e-06, 5.798498e-06, 8.374587e-07,
  2.997011e-06, 2.438751e-06, 2.524697e-06, 3.755766e-06, 3.835039e-06, 
    4.704256e-06, 4.805873e-06, 3.517332e-06, 3.535726e-06, 3.485589e-06, 
    1.113894e-06, 1.334713e-06, 8.822477e-06, 6.953886e-06, 1.485412e-06,
  4.141237e-06, 3.004154e-06, 2.908616e-06, 2.293481e-06, 3.321878e-06, 
    3.271076e-06, 1.927777e-06, 5.334437e-06, 3.679519e-06, 1.012535e-06, 
    6.495557e-07, 2.865602e-06, 9.026359e-06, 9.715022e-06, 3.774892e-06,
  3.373234e-06, 3.439713e-06, 2.161262e-06, 2.65137e-06, 2.94366e-06, 
    3.577819e-06, 4.224129e-06, 3.651538e-06, 3.334212e-06, 1.248013e-06, 
    2.642012e-07, 2.94115e-06, 8.099318e-06, 9.927689e-06, 3.698143e-06,
  2.103237e-06, 3.860095e-06, 2.91218e-06, 1.758888e-06, 4.791808e-06, 
    4.104611e-06, 5.590618e-06, 3.810999e-06, 4.146832e-06, 1.720454e-06, 
    1.572159e-07, 2.008082e-06, 6.700183e-06, 7.204157e-06, 5.792177e-06,
  3.310861e-06, 3.047028e-06, 4.255841e-06, 3.856053e-06, 4.110733e-06, 
    6.73048e-06, 4.323094e-06, 2.556967e-06, 2.348616e-06, 4.022668e-07, 
    4.109445e-08, 9.784048e-07, 5.08116e-06, 6.242627e-06, 7.215475e-06,
  4.056217e-06, 3.651896e-06, 6.001262e-06, 4.494261e-06, 5.843361e-06, 
    7.445806e-06, 5.43949e-06, 1.929569e-06, 1.082541e-06, 3.824318e-07, 
    2.129562e-08, 3.712268e-07, 5.429587e-06, 4.60791e-06, 6.162408e-06,
  5.503282e-06, 4.040241e-06, 2.904656e-06, 2.885764e-06, 2.859676e-06, 
    3.005322e-06, 5.791365e-06, 2.086605e-06, 1.160984e-06, 5.25976e-07, 
    2.588727e-08, 1.637183e-07, 7.161898e-06, 8.114715e-06, 7.315192e-06,
  8.145248e-06, 2.87458e-06, 2.075466e-06, 2.803894e-06, 3.276567e-06, 
    2.260928e-06, 3.425386e-06, 1.606565e-06, 9.021691e-07, 2.21377e-06, 
    1.696521e-07, 7.762448e-07, 8.211214e-06, 1.051917e-05, 5.868509e-06,
  5.033479e-06, 3.740497e-06, 2.794433e-06, 3.044718e-06, 2.525501e-06, 
    2.200783e-06, 1.265649e-06, 1.15929e-06, 1.35459e-06, 2.942317e-06, 
    5.518261e-06, 4.446173e-06, 9.243091e-07, 2.810526e-07, 3.256579e-07,
  4.327069e-06, 2.475814e-06, 1.763751e-06, 3.877029e-06, 4.229347e-06, 
    2.235785e-06, 1.627326e-06, 1.509642e-06, 1.63514e-06, 1.437436e-06, 
    2.844637e-06, 3.163221e-06, 2.237314e-07, 9.863071e-08, 5.712108e-07,
  2.843553e-06, 2.729721e-06, 2.88289e-06, 2.890781e-06, 3.240407e-06, 
    2.365415e-06, 2.045312e-06, 2.004379e-06, 1.499095e-06, 1.73869e-06, 
    1.135377e-06, 1.194424e-06, 1.965398e-07, 1.302426e-07, 9.992657e-07,
  3.423532e-06, 2.580237e-06, 1.199482e-06, 2.792194e-06, 3.270784e-06, 
    2.670268e-06, 1.4553e-06, 2.037604e-06, 2.579306e-06, 7.169445e-07, 
    1.512557e-06, 1.792235e-07, 3.729404e-08, 1.040163e-07, 8.896076e-07,
  6.124586e-06, 3.179412e-06, 2.292585e-06, 2.41826e-06, 2.584515e-06, 
    3.020794e-06, 2.456581e-06, 1.57822e-06, 1.875993e-06, 2.484302e-06, 
    3.217221e-06, 6.889407e-08, 8.584515e-08, 6.658995e-08, 7.570866e-07,
  5.872982e-06, 6.776691e-06, 5.001647e-06, 6.430597e-06, 4.986605e-06, 
    4.041126e-06, 2.845522e-06, 1.615233e-06, 9.952297e-07, 7.083112e-07, 
    4.126252e-07, 9.263348e-08, 1.646074e-07, 1.506087e-07, 2.720431e-06,
  6.061056e-06, 6.189383e-06, 5.849001e-06, 6.37194e-06, 8.159095e-06, 
    7.58615e-06, 4.890776e-06, 3.028918e-06, 2.440379e-06, 4.407149e-06, 
    6.731596e-06, 2.613907e-07, 2.041381e-07, 1.584257e-07, 4.81996e-06,
  6.986781e-06, 4.000258e-06, 3.164784e-06, 3.819842e-06, 6.564739e-06, 
    7.572578e-06, 7.766233e-06, 4.681819e-06, 4.745755e-06, 6.683642e-06, 
    9.334153e-06, 5.350456e-06, 9.297589e-08, 2.185761e-07, 8.192591e-06,
  4.635593e-06, 2.639367e-06, 1.711739e-06, 4.069083e-06, 2.608846e-06, 
    2.520891e-06, 4.744528e-06, 6.094906e-06, 7.08873e-06, 7.532441e-06, 
    9.509345e-06, 8.09262e-06, 2.286284e-06, 3.903145e-07, 1.212927e-05,
  3.240569e-06, 2.655145e-06, 1.917345e-06, 3.628407e-06, 8.53512e-06, 
    6.766562e-06, 3.776741e-06, 2.74375e-06, 8.71637e-06, 7.402836e-06, 
    7.342574e-06, 9.221384e-06, 6.22372e-06, 2.075793e-07, 1.596892e-05,
  0.0001006313, 0.0001085342, 7.099135e-05, 5.178458e-05, 3.578777e-05, 
    8.690673e-06, 4.154547e-06, 3.72556e-06, 4.953563e-07, 2.103215e-06, 
    1.68673e-05, 9.312746e-06, 4.743206e-06, 9.060371e-06, 8.996401e-06,
  0.0001122679, 0.0001229403, 0.000100842, 9.399316e-05, 7.904023e-05, 
    1.282067e-05, 5.515232e-06, 5.719953e-06, 3.236906e-07, 2.294739e-06, 
    9.731789e-06, 7.472513e-06, 5.477143e-06, 4.405952e-06, 1.864126e-05,
  0.000107065, 0.0001220714, 0.0001201718, 0.0001144498, 0.0001160278, 
    2.997795e-05, 8.849805e-06, 5.822543e-06, 2.63374e-06, 3.575472e-06, 
    8.739862e-06, 8.118246e-06, 4.919397e-06, 1.615188e-05, 4.3549e-05,
  5.947268e-05, 7.632373e-05, 0.0001089768, 0.0001460507, 0.00014545, 
    4.808017e-05, 7.417727e-06, 6.466434e-06, 2.921761e-06, 3.136202e-06, 
    7.420389e-06, 5.465929e-06, 1.363285e-05, 3.915519e-05, 4.56313e-05,
  1.3793e-05, 2.261496e-05, 7.046606e-05, 0.0001515636, 0.0001461601, 
    5.225583e-05, 9.002603e-06, 8.034138e-06, 3.915436e-06, 4.885304e-06, 
    5.93008e-06, 7.611998e-06, 4.324276e-05, 4.237118e-05, 3.908927e-05,
  4.350983e-06, 4.933522e-06, 3.344781e-05, 0.0001348043, 0.0001374105, 
    4.334625e-05, 4.832459e-06, 7.070212e-06, 2.76528e-06, 8.265281e-06, 
    7.359843e-06, 1.480137e-05, 4.673182e-05, 3.356615e-05, 2.920247e-05,
  3.510227e-06, 3.095689e-06, 1.70443e-05, 0.0001004171, 0.0001116645, 
    2.738101e-05, 7.417998e-06, 9.180654e-06, 2.845494e-06, 7.427429e-06, 
    9.104317e-06, 3.539303e-05, 4.213254e-05, 3.184003e-05, 2.150577e-05,
  5.649052e-06, 5.268945e-06, 4.135924e-06, 6.262607e-05, 8.66055e-05, 
    1.424959e-05, 6.30355e-06, 9.438391e-06, 2.428934e-06, 7.425734e-06, 
    1.216038e-05, 5.372805e-05, 3.596783e-05, 3.387362e-05, 1.977955e-05,
  1.006256e-05, 6.435389e-06, 6.045964e-06, 3.046951e-05, 4.261938e-05, 
    7.806072e-06, 5.924299e-06, 9.726845e-06, 3.596578e-06, 7.383712e-06, 
    1.661838e-05, 5.898398e-05, 3.473392e-05, 3.129851e-05, 2.100789e-05,
  9.653276e-06, 9.061723e-06, 1.152214e-05, 7.838796e-06, 9.479627e-06, 
    5.369684e-06, 6.231263e-06, 9.13382e-06, 4.337757e-06, 8.005339e-06, 
    2.413716e-05, 6.097303e-05, 4.047053e-05, 3.111355e-05, 2.435291e-05,
  3.380741e-05, 4.319881e-05, 1.996123e-05, 8.315487e-06, 8.251241e-06, 
    8.499421e-06, 1.007114e-05, 7.400447e-06, 1.09489e-05, 9.472701e-06, 
    7.298588e-06, 3.535719e-06, 2.313932e-06, 2.759823e-06, 3.145179e-06,
  3.614269e-05, 5.23525e-05, 2.835202e-05, 1.182117e-05, 1.071492e-05, 
    6.149473e-06, 6.664505e-06, 6.098944e-06, 9.021536e-06, 7.07655e-06, 
    3.791662e-06, 1.683043e-06, 1.422141e-06, 1.971407e-06, 2.342927e-06,
  4.995757e-05, 6.166242e-05, 3.594363e-05, 1.992446e-05, 1.786847e-05, 
    5.745806e-06, 6.253022e-06, 7.563626e-06, 7.817613e-06, 5.727597e-06, 
    1.386615e-06, 6.473257e-07, 7.184e-07, 1.248138e-06, 1.654348e-06,
  5.660149e-05, 6.557427e-05, 5.277984e-05, 3.97444e-05, 3.080112e-05, 
    1.10328e-05, 6.987135e-06, 7.825484e-06, 5.794293e-06, 6.468085e-06, 
    1.384404e-06, 7.765179e-07, 1.666883e-06, 1.523222e-06, 2.450406e-06,
  5.050682e-05, 5.493384e-05, 7.19882e-05, 7.048098e-05, 5.408892e-05, 
    1.71305e-05, 6.682547e-06, 5.900743e-06, 4.634942e-06, 3.591355e-06, 
    1.057702e-06, 9.285946e-07, 1.824404e-06, 2.406681e-06, 2.901717e-06,
  1.585447e-05, 4.106e-05, 7.316258e-05, 8.848817e-05, 7.642592e-05, 
    2.152059e-05, 5.548718e-06, 4.764271e-06, 5.16562e-06, 3.238919e-06, 
    5.633965e-07, 7.716015e-07, 1.636176e-06, 2.495979e-06, 3.815058e-06,
  3.524217e-05, 2.73561e-05, 5.942116e-05, 0.0001010735, 9.89792e-05, 
    2.665991e-05, 6.584212e-06, 5.918046e-06, 3.93253e-06, 2.102135e-06, 
    7.860691e-07, 9.300703e-07, 1.296886e-06, 2.214065e-06, 2.434096e-06,
  0.0001258592, 2.972485e-05, 4.52745e-05, 0.0001135748, 0.0001347812, 
    3.874239e-05, 6.446154e-06, 3.964987e-06, 4.108594e-06, 2.765121e-06, 
    8.381604e-07, 1.240835e-06, 1.20789e-06, 1.85488e-06, 2.339373e-06,
  0.0002670483, 7.128644e-05, 4.252748e-05, 0.0001330866, 0.0001807868, 
    5.136428e-05, 6.071512e-06, 4.97655e-06, 4.569292e-06, 4.868757e-06, 
    1.249153e-06, 1.955368e-06, 1.736015e-06, 1.959271e-06, 2.161386e-06,
  0.00044707, 0.0001940407, 8.851204e-05, 0.0001385137, 0.0002195992, 
    7.23729e-05, 6.371133e-06, 6.829498e-06, 5.175444e-06, 7.973374e-06, 
    1.951531e-06, 1.940285e-06, 2.052364e-06, 1.899198e-06, 2.550894e-06,
  1.660534e-05, 6.061765e-06, 9.074879e-06, 8.428432e-06, 9.801245e-06, 
    1.230778e-05, 1.174536e-05, 1.030835e-05, 1.313144e-05, 1.026168e-05, 
    9.804092e-06, 1.074201e-05, 8.027073e-06, 7.626728e-06, 4.566917e-06,
  7.375225e-06, 6.317509e-06, 1.053461e-05, 1.248684e-05, 8.145535e-06, 
    1.124957e-05, 1.101725e-05, 1.122229e-05, 1.200084e-05, 9.583632e-06, 
    1.086851e-05, 1.135226e-05, 9.765783e-06, 7.57223e-06, 5.765051e-06,
  8.171171e-06, 7.553189e-06, 1.071911e-05, 1.141138e-05, 1.163811e-05, 
    9.517237e-06, 1.109398e-05, 1.297417e-05, 1.132693e-05, 9.42734e-06, 
    1.146768e-05, 1.251793e-05, 1.260322e-05, 9.883792e-06, 6.035172e-06,
  5.761791e-06, 9.974729e-06, 1.06853e-05, 1.085462e-05, 1.091084e-05, 
    1.250247e-05, 1.303685e-05, 1.312303e-05, 9.168029e-06, 8.003975e-06, 
    1.103129e-05, 8.58325e-06, 1.012436e-05, 7.113542e-06, 4.821833e-06,
  5.570747e-06, 1.058925e-05, 1.128525e-05, 1.584653e-05, 1.243168e-05, 
    1.305711e-05, 1.444642e-05, 1.304656e-05, 8.403782e-06, 8.103503e-06, 
    7.50028e-06, 6.218252e-06, 8.460469e-06, 5.004883e-06, 4.642653e-06,
  6.477131e-06, 9.883039e-06, 1.109618e-05, 1.204041e-05, 1.40795e-05, 
    1.15801e-05, 1.197324e-05, 1.352748e-05, 1.064192e-05, 6.82362e-06, 
    6.756896e-06, 6.754997e-06, 7.850266e-06, 5.252401e-06, 3.708271e-06,
  6.913892e-06, 8.709846e-06, 1.134181e-05, 1.035012e-05, 1.391123e-05, 
    1.100991e-05, 8.477574e-06, 1.133843e-05, 1.214944e-05, 1.069471e-05, 
    9.588201e-06, 8.769729e-06, 8.014583e-06, 6.742653e-06, 3.118192e-06,
  5.321673e-06, 4.555267e-06, 9.979348e-06, 7.704019e-06, 1.211807e-05, 
    8.30621e-06, 6.910839e-06, 7.725566e-06, 8.034041e-06, 1.000725e-05, 
    9.8598e-06, 8.946502e-06, 8.707385e-06, 6.662331e-06, 3.022526e-06,
  3.502909e-06, 1.302994e-06, 6.344982e-06, 4.573518e-06, 8.867429e-06, 
    1.131222e-05, 7.379565e-06, 6.88618e-06, 6.487717e-06, 1.0648e-05, 
    1.155956e-05, 1.067173e-05, 1.181184e-05, 6.935561e-06, 5.85375e-06,
  9.152949e-07, 2.433201e-06, 3.144995e-06, 4.182662e-06, 7.786717e-06, 
    7.70336e-06, 6.961543e-06, 7.306458e-06, 7.92737e-06, 6.41661e-06, 
    7.780603e-06, 1.111365e-05, 1.060439e-05, 9.103708e-06, 6.493143e-06,
  9.82431e-06, 1.078315e-05, 9.182424e-06, 9.978467e-06, 8.715984e-06, 
    1.178313e-05, 1.2675e-05, 1.467194e-05, 1.430353e-05, 1.190822e-05, 
    9.320353e-06, 8.66474e-06, 8.334881e-06, 9.770383e-06, 8.114302e-06,
  1.381356e-05, 1.136648e-05, 1.040995e-05, 1.082283e-05, 1.101068e-05, 
    1.066085e-05, 1.250405e-05, 1.283885e-05, 1.210835e-05, 1.115578e-05, 
    8.828077e-06, 8.002914e-06, 6.470607e-06, 6.209122e-06, 6.195959e-06,
  1.250251e-05, 1.137466e-05, 1.131263e-05, 1.125126e-05, 1.279777e-05, 
    1.10013e-05, 1.245852e-05, 1.192939e-05, 1.151477e-05, 1.018356e-05, 
    9.492741e-06, 6.765822e-06, 6.206151e-06, 5.22023e-06, 4.900241e-06,
  1.453124e-05, 1.211462e-05, 1.131957e-05, 1.087139e-05, 9.35897e-06, 
    1.103119e-05, 1.318908e-05, 1.219887e-05, 1.022532e-05, 9.075113e-06, 
    7.661835e-06, 5.686281e-06, 5.362328e-06, 3.905234e-06, 5.034317e-06,
  1.425056e-05, 1.280872e-05, 1.19273e-05, 1.184278e-05, 1.023985e-05, 
    1.193761e-05, 1.244839e-05, 1.151194e-05, 9.032178e-06, 7.859542e-06, 
    7.494619e-06, 5.27495e-06, 5.521473e-06, 4.750987e-06, 5.355833e-06,
  1.239452e-05, 1.411693e-05, 1.102714e-05, 1.133372e-05, 1.038054e-05, 
    1.104093e-05, 1.191245e-05, 1.028997e-05, 8.613185e-06, 8.438677e-06, 
    6.460242e-06, 5.097815e-06, 4.658454e-06, 5.89034e-06, 9.738805e-06,
  1.092222e-05, 1.42794e-05, 1.049305e-05, 1.049013e-05, 1.1961e-05, 
    1.133373e-05, 1.306707e-05, 8.857606e-06, 8.386283e-06, 6.485116e-06, 
    5.325121e-06, 4.78971e-06, 4.078361e-06, 7.596522e-06, 1.192277e-05,
  1.237412e-05, 1.192648e-05, 1.050914e-05, 9.78404e-06, 1.092126e-05, 
    1.226953e-05, 1.136408e-05, 8.334838e-06, 6.545527e-06, 7.934898e-06, 
    6.432572e-06, 5.935983e-06, 5.566323e-06, 7.461561e-06, 1.002723e-05,
  1.019127e-05, 1.082299e-05, 1.163597e-05, 8.250988e-06, 1.355223e-05, 
    1.299413e-05, 1.055215e-05, 7.565908e-06, 8.372586e-06, 7.791275e-06, 
    8.29042e-06, 8.253432e-06, 7.47533e-06, 9.804507e-06, 9.638415e-06,
  1.265579e-05, 1.229807e-05, 8.666628e-06, 8.238262e-06, 1.213014e-05, 
    1.056903e-05, 1.098526e-05, 8.131391e-06, 1.045642e-05, 1.03586e-05, 
    1.128891e-05, 9.58665e-06, 9.778231e-06, 1.184208e-05, 8.501349e-06,
  1.074307e-05, 1.145919e-05, 1.181531e-05, 1.303241e-05, 1.301078e-05, 
    1.098936e-05, 1.150249e-05, 9.339513e-06, 8.613682e-06, 6.531718e-06, 
    4.791436e-06, 1.175281e-05, 1.332442e-05, 1.294314e-05, 1.304977e-05,
  1.050417e-05, 1.118936e-05, 1.124606e-05, 1.213653e-05, 1.418881e-05, 
    1.274619e-05, 1.144627e-05, 9.270566e-06, 8.713579e-06, 5.985706e-06, 
    6.237582e-06, 8.788051e-06, 1.118937e-05, 1.372391e-05, 1.129627e-05,
  1.109197e-05, 1.143478e-05, 1.064637e-05, 1.404929e-05, 1.496535e-05, 
    1.256622e-05, 1.096356e-05, 1.114167e-05, 1.006929e-05, 8.820033e-06, 
    8.260046e-06, 7.137132e-06, 8.379535e-06, 1.041912e-05, 8.490206e-06,
  1.37057e-05, 1.244886e-05, 1.140777e-05, 1.427202e-05, 1.308165e-05, 
    1.313018e-05, 1.267674e-05, 1.315693e-05, 1.081768e-05, 1.114945e-05, 
    8.860579e-06, 7.427731e-06, 1.032058e-05, 6.832072e-06, 7.115884e-06,
  1.373153e-05, 1.201036e-05, 1.19624e-05, 1.328551e-05, 1.496667e-05, 
    1.347772e-05, 1.359734e-05, 1.320052e-05, 1.448597e-05, 1.29455e-05, 
    9.913552e-06, 8.317508e-06, 9.352944e-06, 5.668864e-06, 5.800702e-06,
  1.212479e-05, 1.211617e-05, 1.326226e-05, 1.455543e-05, 1.537737e-05, 
    1.528843e-05, 1.528588e-05, 1.409737e-05, 1.467104e-05, 1.316016e-05, 
    1.033102e-05, 9.868431e-06, 8.558996e-06, 8.915405e-06, 6.266121e-06,
  1.127662e-05, 1.072386e-05, 1.208849e-05, 1.36679e-05, 1.512492e-05, 
    1.288924e-05, 1.45528e-05, 1.602618e-05, 1.41762e-05, 1.358191e-05, 
    1.214451e-05, 9.249656e-06, 9.158181e-06, 9.994616e-06, 8.891122e-06,
  9.236202e-06, 1.152397e-05, 1.095493e-05, 1.257834e-05, 1.408741e-05, 
    9.987379e-06, 1.581603e-05, 1.680524e-05, 1.498803e-05, 1.713649e-05, 
    1.440898e-05, 1.221581e-05, 9.249246e-06, 1.195824e-05, 1.332183e-05,
  9.381728e-06, 8.076301e-06, 8.98857e-06, 1.285471e-05, 1.340689e-05, 
    1.520274e-05, 1.785121e-05, 1.583667e-05, 1.595974e-05, 1.787045e-05, 
    1.547973e-05, 1.46218e-05, 1.434327e-05, 1.352235e-05, 1.585804e-05,
  8.162914e-06, 9.443228e-06, 1.120621e-05, 9.93876e-06, 1.26429e-05, 
    1.492377e-05, 1.46838e-05, 1.477334e-05, 1.516906e-05, 1.789169e-05, 
    2.147219e-05, 1.314549e-05, 1.715776e-05, 1.423688e-05, 1.224888e-05,
  1.447733e-05, 1.381168e-05, 1.217802e-05, 1.098542e-05, 9.333036e-06, 
    7.872514e-06, 9.109916e-06, 9.302894e-06, 6.987225e-06, 6.288072e-06, 
    6.385273e-06, 6.359037e-06, 5.258303e-06, 8.389102e-06, 6.848727e-06,
  1.641189e-05, 1.604383e-05, 1.418732e-05, 1.205583e-05, 1.058187e-05, 
    8.846873e-06, 8.796796e-06, 9.130074e-06, 7.290836e-06, 5.713895e-06, 
    6.318704e-06, 6.73252e-06, 6.833065e-06, 6.632382e-06, 7.563614e-06,
  2.180204e-05, 1.785404e-05, 1.782013e-05, 1.571709e-05, 1.225906e-05, 
    1.098946e-05, 8.710732e-06, 9.487359e-06, 8.178207e-06, 5.051931e-06, 
    6.91581e-06, 6.715905e-06, 6.19413e-06, 3.760334e-06, 3.51066e-06,
  2.206242e-05, 1.94673e-05, 1.970141e-05, 1.756665e-05, 1.453684e-05, 
    1.188769e-05, 9.7477e-06, 9.778077e-06, 9.141314e-06, 5.199747e-06, 
    7.49564e-06, 8.601702e-06, 7.495753e-06, 4.921179e-06, 4.381548e-06,
  2.011614e-05, 2.146813e-05, 2.202394e-05, 1.954593e-05, 1.675964e-05, 
    1.325408e-05, 1.152726e-05, 7.830266e-06, 8.698163e-06, 6.281184e-06, 
    7.561684e-06, 8.472102e-06, 7.024664e-06, 6.414184e-06, 6.205167e-06,
  2.008525e-05, 2.006797e-05, 2.191806e-05, 2.197574e-05, 1.810457e-05, 
    1.343071e-05, 1.26719e-05, 9.46058e-06, 9.5818e-06, 6.996534e-06, 
    6.075929e-06, 7.808162e-06, 6.995719e-06, 5.683105e-06, 6.043894e-06,
  1.793132e-05, 2.033355e-05, 2.076745e-05, 2.331113e-05, 2.050209e-05, 
    1.538157e-05, 1.205997e-05, 1.047699e-05, 9.190963e-06, 6.720071e-06, 
    6.112013e-06, 7.121754e-06, 6.702489e-06, 6.214666e-06, 7.14244e-06,
  1.629338e-05, 1.925746e-05, 1.958084e-05, 2.115377e-05, 2.108205e-05, 
    1.522712e-05, 1.366443e-05, 1.118932e-05, 8.499997e-06, 7.889119e-06, 
    7.505712e-06, 8.526464e-06, 7.903708e-06, 7.916874e-06, 7.823075e-06,
  1.694775e-05, 1.675587e-05, 1.825782e-05, 2.048495e-05, 1.844388e-05, 
    1.721535e-05, 1.463336e-05, 1.151889e-05, 7.745182e-06, 8.380331e-06, 
    7.570994e-06, 8.426286e-06, 5.929843e-06, 7.476521e-06, 9.917175e-06,
  1.785363e-05, 1.639409e-05, 1.683486e-05, 1.826364e-05, 2.045101e-05, 
    1.686483e-05, 1.303747e-05, 1.102438e-05, 8.294186e-06, 8.747666e-06, 
    8.442615e-06, 9.619785e-06, 7.630813e-06, 7.991979e-06, 9.632779e-06,
  7.437973e-06, 6.982293e-06, 6.35936e-06, 7.053842e-06, 7.001276e-06, 
    6.566044e-06, 4.945765e-06, 4.636252e-06, 4.38474e-06, 5.5153e-06, 
    7.497852e-06, 6.731144e-06, 6.321072e-06, 7.438676e-06, 7.201897e-06,
  8.651516e-06, 8.101733e-06, 7.135694e-06, 7.759241e-06, 7.450706e-06, 
    7.564078e-06, 6.041905e-06, 6.051994e-06, 5.087313e-06, 6.674923e-06, 
    1.032218e-05, 7.872696e-06, 6.399113e-06, 8.211461e-06, 9.89054e-06,
  1.139548e-05, 9.299342e-06, 7.672315e-06, 7.645604e-06, 7.275356e-06, 
    7.223935e-06, 6.939317e-06, 6.044352e-06, 7.447773e-06, 7.530814e-06, 
    9.867287e-06, 9.925167e-06, 8.372883e-06, 1.078778e-05, 8.410479e-06,
  1.52588e-05, 1.163323e-05, 8.388254e-06, 8.010636e-06, 9.916604e-06, 
    8.461953e-06, 5.589638e-06, 5.270704e-06, 8.035214e-06, 7.347518e-06, 
    7.345704e-06, 7.474852e-06, 6.380677e-06, 7.963473e-06, 5.529916e-06,
  1.919057e-05, 1.502512e-05, 1.359663e-05, 1.007982e-05, 9.197268e-06, 
    9.951293e-06, 7.314464e-06, 6.153587e-06, 6.284958e-06, 5.298301e-06, 
    5.185735e-06, 5.82404e-06, 7.132509e-06, 9.597012e-06, 6.930585e-06,
  2.15625e-05, 2.124669e-05, 1.710916e-05, 1.513429e-05, 1.169584e-05, 
    1.027552e-05, 1.016839e-05, 7.72884e-06, 7.096329e-06, 7.871077e-06, 
    7.961597e-06, 8.574462e-06, 1.36466e-05, 9.484178e-06, 7.592711e-06,
  2.377003e-05, 2.570478e-05, 2.298466e-05, 2.441133e-05, 2.620462e-05, 
    1.924073e-05, 1.403813e-05, 9.492245e-06, 9.089644e-06, 8.633214e-06, 
    7.555935e-06, 9.462647e-06, 1.35237e-05, 1.137162e-05, 8.523113e-06,
  2.282397e-05, 2.418908e-05, 2.445775e-05, 2.933247e-05, 4.03835e-05, 
    3.619519e-05, 3.095554e-05, 2.044529e-05, 1.147923e-05, 9.949575e-06, 
    9.29417e-06, 1.229148e-05, 1.155544e-05, 1.238045e-05, 1.161524e-05,
  2.52923e-05, 2.457849e-05, 2.568413e-05, 2.304386e-05, 2.894945e-05, 
    4.006916e-05, 5.103655e-05, 4.973616e-05, 3.711778e-05, 1.67221e-05, 
    1.213925e-05, 1.104744e-05, 7.276819e-06, 1.012324e-05, 1.292132e-05,
  2.736452e-05, 2.426733e-05, 2.494473e-05, 2.443567e-05, 2.478584e-05, 
    3.025449e-05, 3.903978e-05, 5.300258e-05, 6.850365e-05, 6.562188e-05, 
    2.828617e-05, 1.160355e-05, 1.101257e-05, 1.056087e-05, 9.301919e-06,
  6.391115e-06, 6.602481e-06, 6.302148e-06, 6.884165e-06, 8.315621e-06, 
    8.35193e-06, 4.78328e-06, 6.260119e-06, 7.065987e-06, 8.639591e-06, 
    1.605445e-05, 2.190969e-05, 2.323677e-05, 2.127433e-05, 2.012428e-05,
  7.45402e-06, 7.722248e-06, 7.375134e-06, 8.4358e-06, 1.022799e-05, 
    9.360859e-06, 6.006247e-06, 6.991116e-06, 5.837766e-06, 9.683225e-06, 
    1.33195e-05, 2.296661e-05, 2.414369e-05, 2.187302e-05, 2.198628e-05,
  1.44902e-05, 1.495299e-05, 1.193933e-05, 8.958809e-06, 1.106095e-05, 
    6.047211e-06, 6.309868e-06, 8.927644e-06, 7.705393e-06, 9.827313e-06, 
    1.669883e-05, 2.977492e-05, 3.138706e-05, 2.448233e-05, 3.04145e-05,
  2.784128e-05, 3.068385e-05, 2.057499e-05, 1.670893e-05, 1.214708e-05, 
    8.988634e-06, 8.287884e-06, 8.561715e-06, 1.018601e-05, 1.102969e-05, 
    1.364737e-05, 2.358697e-05, 2.749077e-05, 3.877064e-05, 3.353008e-05,
  3.525338e-05, 3.471331e-05, 3.192789e-05, 2.864054e-05, 2.461571e-05, 
    2.015439e-05, 1.396021e-05, 1.307114e-05, 1.29104e-05, 9.602588e-06, 
    1.18609e-05, 1.7561e-05, 3.136684e-05, 4.883579e-05, 4.35274e-05,
  2.430765e-05, 2.740284e-05, 3.422662e-05, 3.30716e-05, 3.312854e-05, 
    3.258163e-05, 2.730308e-05, 2.022322e-05, 1.171533e-05, 1.126902e-05, 
    1.343666e-05, 1.482999e-05, 2.864482e-05, 4.940865e-05, 7.402306e-05,
  2.720091e-05, 2.482316e-05, 3.817261e-05, 2.444777e-05, 3.043029e-05, 
    3.34622e-05, 3.071088e-05, 3.420822e-05, 2.646391e-05, 1.59495e-05, 
    1.133157e-05, 1.316765e-05, 1.674419e-05, 3.914277e-05, 8.127615e-05,
  4.272973e-05, 3.360215e-05, 3.050499e-05, 2.629865e-05, 2.666564e-05, 
    2.595732e-05, 2.128839e-05, 2.972595e-05, 2.263061e-05, 2.579347e-05, 
    1.554534e-05, 9.519718e-06, 1.100292e-05, 1.303813e-05, 2.720045e-05,
  4.009406e-05, 2.907404e-05, 2.766706e-05, 2.595259e-05, 2.37871e-05, 
    1.638551e-05, 1.831376e-05, 1.593114e-05, 2.411046e-05, 2.588204e-05, 
    1.96639e-05, 1.14389e-05, 6.815295e-06, 6.650618e-06, 9.886603e-06,
  2.581736e-05, 2.834142e-05, 2.939485e-05, 2.21288e-05, 1.750132e-05, 
    1.551384e-05, 1.163775e-05, 1.129612e-05, 1.493863e-05, 2.526934e-05, 
    2.24875e-05, 1.592526e-05, 1.166954e-05, 6.634397e-06, 5.652578e-06,
  3.538281e-06, 1.996467e-06, 4.112547e-06, 6.768454e-06, 1.380506e-05, 
    2.139671e-05, 2.739645e-05, 3.705532e-05, 5.470754e-05, 5.387615e-05, 
    5.313582e-05, 4.790358e-05, 4.799032e-05, 3.167111e-05, 1.240249e-05,
  3.668591e-06, 4.156671e-06, 4.911591e-06, 8.708086e-06, 1.248547e-05, 
    1.87698e-05, 1.968416e-05, 2.290094e-05, 3.473356e-05, 4.974553e-05, 
    5.329548e-05, 4.318588e-05, 4.063502e-05, 3.283057e-05, 1.252508e-05,
  5.912397e-06, 6.87838e-06, 8.835647e-06, 9.423811e-06, 1.319701e-05, 
    1.440797e-05, 1.518251e-05, 1.860202e-05, 2.269032e-05, 2.921173e-05, 
    4.427291e-05, 4.644787e-05, 3.748711e-05, 3.179357e-05, 1.617296e-05,
  7.702502e-06, 7.774872e-06, 1.100833e-05, 1.007811e-05, 9.667338e-06, 
    9.304817e-06, 9.354262e-06, 8.068503e-06, 8.18946e-06, 1.092556e-05, 
    1.398356e-05, 2.968275e-05, 3.586505e-05, 2.374268e-05, 1.886527e-05,
  2.170746e-06, 3.255357e-06, 4.219439e-06, 8.283157e-06, 1.068099e-05, 
    1.12599e-05, 9.914778e-06, 4.584796e-06, 4.450524e-06, 3.424013e-06, 
    7.544733e-06, 1.185537e-05, 1.218839e-05, 1.906962e-05, 1.247442e-05,
  1.767699e-06, 6.037314e-07, 1.960625e-06, 2.261869e-06, 7.945833e-06, 
    1.19061e-05, 9.453795e-06, 7.239012e-06, 3.83667e-06, 3.072201e-06, 
    1.768995e-06, 5.216471e-06, 5.578667e-06, 9.895856e-06, 1.012708e-05,
  1.808319e-06, 1.695734e-06, 1.8827e-06, 1.637645e-06, 3.780327e-06, 
    6.389065e-06, 8.900092e-06, 1.315807e-05, 1.005377e-05, 5.936439e-06, 
    6.040167e-06, 6.959638e-06, 7.255919e-06, 8.162853e-06, 6.991441e-06,
  2.369179e-06, 2.574986e-06, 2.280123e-06, 2.083318e-06, 2.805201e-06, 
    3.68243e-06, 1.015237e-05, 1.215245e-05, 1.420614e-05, 1.223705e-05, 
    1.249118e-05, 6.167601e-06, 8.636584e-06, 8.050248e-06, 8.963163e-06,
  2.189868e-06, 2.267361e-06, 2.857584e-06, 2.587609e-06, 3.552024e-06, 
    2.677612e-06, 1.771029e-06, 3.858007e-06, 1.141502e-05, 1.49798e-05, 
    1.95552e-05, 1.151626e-05, 1.098917e-05, 8.172611e-06, 8.683286e-06,
  3.817692e-06, 4.492476e-06, 5.818868e-06, 5.970069e-06, 4.526113e-06, 
    3.872129e-06, 2.571506e-06, 1.489488e-06, 2.837147e-06, 1.164296e-05, 
    1.619697e-05, 1.732608e-05, 1.374524e-05, 8.786897e-06, 9.689002e-06,
  6.885621e-06, 4.812013e-06, 8.154281e-06, 1.167252e-05, 1.156391e-05, 
    8.282613e-06, 7.454158e-06, 7.113118e-06, 7.080141e-06, 7.525121e-06, 
    8.908772e-06, 6.938123e-06, 6.63274e-06, 6.756129e-06, 6.905587e-06,
  1.246822e-05, 8.577714e-06, 8.951787e-06, 8.54773e-06, 7.143745e-06, 
    9.019752e-06, 8.095407e-06, 8.177037e-06, 8.500111e-06, 9.651451e-06, 
    9.220569e-06, 8.132217e-06, 7.26911e-06, 6.95238e-06, 5.803329e-06,
  1.568926e-05, 1.111744e-05, 9.102518e-06, 5.963421e-06, 4.879011e-06, 
    7.694549e-06, 9.441619e-06, 9.486467e-06, 1.116034e-05, 1.047925e-05, 
    8.757087e-06, 8.545727e-06, 6.500062e-06, 6.575867e-06, 6.70769e-06,
  1.19904e-05, 1.450946e-05, 1.047537e-05, 4.960099e-06, 5.145077e-06, 
    9.165259e-06, 1.059856e-05, 1.186204e-05, 1.305198e-05, 9.503156e-06, 
    9.175906e-06, 9.004633e-06, 8.526089e-06, 7.766242e-06, 6.983123e-06,
  5.061149e-06, 1.091789e-05, 1.166844e-05, 7.108784e-06, 6.525269e-06, 
    9.942881e-06, 1.172419e-05, 1.26116e-05, 1.270264e-05, 8.928728e-06, 
    9.266497e-06, 7.742015e-06, 8.19361e-06, 7.406582e-06, 7.335071e-06,
  1.993458e-06, 1.930238e-06, 4.694627e-06, 6.245597e-06, 9.453875e-06, 
    1.270988e-05, 1.311222e-05, 1.388566e-05, 1.380436e-05, 8.184206e-06, 
    7.198154e-06, 8.057271e-06, 7.435877e-06, 6.19618e-06, 6.939246e-06,
  1.627022e-06, 1.173512e-06, 2.441799e-06, 8.108189e-06, 1.332533e-05, 
    1.339701e-05, 1.007589e-05, 1.250107e-05, 1.21427e-05, 9.288849e-06, 
    6.393794e-06, 6.952349e-06, 6.85356e-06, 6.537506e-06, 6.482749e-06,
  2.98689e-06, 1.820571e-06, 3.763678e-06, 8.011229e-06, 1.247211e-05, 
    1.240996e-05, 1.085194e-05, 1.170107e-05, 1.119679e-05, 6.625356e-06, 
    5.325998e-06, 4.909051e-06, 7.871111e-06, 7.322407e-06, 7.05341e-06,
  3.428209e-06, 2.915605e-06, 3.415516e-06, 5.672956e-06, 9.353756e-06, 
    1.172834e-05, 1.393486e-05, 9.575284e-06, 9.809683e-06, 6.727566e-06, 
    5.877905e-06, 8.482541e-06, 7.554575e-06, 8.33865e-06, 1.075409e-05,
  4.385223e-06, 3.219162e-06, 3.191057e-06, 2.817379e-06, 3.991823e-06, 
    6.689159e-06, 1.445481e-05, 1.55142e-05, 9.906754e-06, 9.410322e-06, 
    8.459124e-06, 5.816972e-06, 6.874249e-06, 7.432961e-06, 8.399334e-06,
  5.195996e-06, 6.20141e-06, 6.970431e-06, 8.091851e-06, 6.412581e-06, 
    5.4053e-06, 4.038511e-06, 4.339803e-06, 6.025863e-06, 5.666851e-06, 
    5.290478e-06, 6.371226e-06, 6.296115e-06, 2.772375e-06, 3.373523e-06,
  6.258155e-06, 6.193897e-06, 7.253643e-06, 8.0027e-06, 7.547695e-06, 
    4.885232e-06, 4.629572e-06, 4.005748e-06, 5.198548e-06, 5.37751e-06, 
    5.125405e-06, 6.459829e-06, 6.269296e-06, 2.978124e-06, 2.791751e-06,
  9.254086e-06, 7.898791e-06, 8.28486e-06, 8.649867e-06, 6.565909e-06, 
    4.874155e-06, 4.032026e-06, 4.465601e-06, 5.546704e-06, 6.364435e-06, 
    6.98865e-06, 6.931668e-06, 3.814941e-06, 4.097277e-06, 3.537108e-06,
  1.184342e-05, 9.742733e-06, 9.886799e-06, 8.999584e-06, 7.956701e-06, 
    6.493208e-06, 4.823069e-06, 5.329829e-06, 5.954494e-06, 5.91265e-06, 
    5.75493e-06, 4.803553e-06, 3.790867e-06, 4.840232e-06, 4.148553e-06,
  1.316256e-05, 1.081349e-05, 1.303834e-05, 1.19641e-05, 9.433315e-06, 
    6.026194e-06, 5.889343e-06, 5.119932e-06, 4.341606e-06, 4.848167e-06, 
    4.596486e-06, 3.91519e-06, 4.609353e-06, 4.486788e-06, 6.090983e-06,
  1.699578e-05, 1.454187e-05, 1.609392e-05, 1.574154e-05, 9.607214e-06, 
    7.277558e-06, 5.61441e-06, 4.790341e-06, 4.915742e-06, 4.981997e-06, 
    5.76345e-06, 5.736443e-06, 4.071276e-06, 4.387088e-06, 8.000677e-06,
  2.166752e-05, 2.255993e-05, 1.968306e-05, 1.701637e-05, 1.076405e-05, 
    8.390083e-06, 6.453026e-06, 4.955888e-06, 5.434091e-06, 5.368045e-06, 
    5.751719e-06, 5.248302e-06, 5.580221e-06, 4.989411e-06, 4.69832e-06,
  2.305159e-05, 2.204211e-05, 2.167883e-05, 2.142588e-05, 1.367508e-05, 
    8.47261e-06, 7.38515e-06, 5.973014e-06, 6.201956e-06, 5.38669e-06, 
    4.587048e-06, 4.755154e-06, 7.964777e-06, 3.476827e-06, 2.615805e-06,
  2.123415e-05, 1.946085e-05, 2.322074e-05, 2.077104e-05, 1.625343e-05, 
    1.091697e-05, 8.625692e-06, 7.738461e-06, 5.691591e-06, 6.375639e-06, 
    5.990872e-06, 5.249064e-06, 3.907298e-06, 4.446636e-06, 3.902689e-06,
  1.706977e-05, 2.083209e-05, 2.354175e-05, 9.578069e-06, 1.76665e-05, 
    1.31462e-05, 9.96064e-06, 8.912711e-06, 7.197618e-06, 7.756627e-06, 
    5.952169e-06, 5.138955e-06, 3.505276e-06, 3.488888e-06, 5.002094e-06,
  2.84191e-06, 5.008202e-06, 5.89233e-06, 6.823815e-06, 7.093372e-06, 
    5.071212e-06, 7.05006e-06, 5.986864e-06, 4.966741e-06, 6.545067e-06, 
    9.821883e-06, 9.170137e-06, 1.439605e-05, 1.482486e-05, 1.084835e-05,
  2.801915e-06, 5.539169e-06, 7.900651e-06, 7.083213e-06, 7.56074e-06, 
    6.593486e-06, 5.40598e-06, 4.645336e-06, 4.230446e-06, 5.569563e-06, 
    1.010877e-05, 1.546179e-05, 1.344274e-05, 1.002708e-05, 8.287429e-06,
  5.739031e-06, 7.41102e-06, 8.199582e-06, 8.156494e-06, 5.96826e-06, 
    5.986104e-06, 6.535195e-06, 4.540211e-06, 4.687952e-06, 8.6829e-06, 
    1.695897e-05, 2.126225e-05, 1.922799e-05, 1.45267e-05, 1.164041e-05,
  4.486245e-06, 6.229697e-06, 8.07932e-06, 9.221774e-06, 7.348782e-06, 
    4.460076e-06, 4.624131e-06, 6.023075e-06, 9.607256e-06, 1.762533e-05, 
    2.358906e-05, 2.726477e-05, 2.036326e-05, 1.149135e-05, 1.164235e-05,
  3.503421e-06, 5.624255e-06, 7.984257e-06, 7.544294e-06, 7.038349e-06, 
    4.349838e-06, 5.594529e-06, 9.496044e-06, 1.705694e-05, 2.46235e-05, 
    2.919037e-05, 2.10552e-05, 1.14445e-05, 1.034336e-05, 1.55415e-05,
  4.506316e-06, 4.567472e-06, 5.823085e-06, 6.528754e-06, 4.859176e-06, 
    4.795412e-06, 8.05786e-06, 1.613283e-05, 1.936455e-05, 2.359738e-05, 
    2.048661e-05, 1.153637e-05, 8.631258e-06, 1.050378e-05, 1.401286e-05,
  4.495677e-06, 5.608552e-06, 4.849515e-06, 5.223979e-06, 6.382413e-06, 
    7.828675e-06, 1.085479e-05, 1.594063e-05, 1.456394e-05, 1.731987e-05, 
    1.259303e-05, 9.216613e-06, 9.933649e-06, 1.117154e-05, 9.958771e-06,
  4.977918e-06, 5.953339e-06, 5.855941e-06, 6.13838e-06, 7.272552e-06, 
    9.739131e-06, 1.228637e-05, 1.319407e-05, 1.267046e-05, 1.525923e-05, 
    1.363734e-05, 1.265931e-05, 1.453154e-05, 1.29309e-05, 1.520693e-05,
  4.229705e-06, 6.359161e-06, 6.230422e-06, 7.882848e-06, 8.125762e-06, 
    1.04893e-05, 1.247517e-05, 1.196142e-05, 1.71685e-05, 1.873063e-05, 
    1.571893e-05, 1.818672e-05, 2.057905e-05, 2.089032e-05, 2.784132e-05,
  5.088156e-06, 6.006173e-06, 8.723641e-06, 8.288035e-06, 9.501206e-06, 
    1.148842e-05, 1.397795e-05, 1.727878e-05, 2.236466e-05, 2.155837e-05, 
    2.230467e-05, 2.375629e-05, 2.709819e-05, 2.478479e-05, 3.122506e-05,
  6.605359e-06, 5.883175e-06, 6.567411e-06, 7.067428e-06, 6.758168e-06, 
    1.0829e-05, 2.576055e-05, 1.833676e-05, 1.189302e-05, 5.83433e-06, 
    6.26531e-06, 6.182359e-06, 6.72271e-06, 5.942192e-06, 5.187095e-06,
  6.202981e-06, 4.312957e-06, 6.786237e-06, 1.000294e-05, 8.962928e-06, 
    1.612728e-05, 2.474816e-05, 1.366188e-05, 7.495712e-06, 7.425209e-06, 
    8.322511e-06, 8.886266e-06, 7.377133e-06, 7.709045e-06, 8.555235e-06,
  6.647664e-06, 6.71948e-06, 8.139414e-06, 9.128387e-06, 1.545801e-05, 
    2.653451e-05, 2.054263e-05, 1.133757e-05, 8.669313e-06, 1.049102e-05, 
    1.157006e-05, 1.102249e-05, 1.034614e-05, 8.939543e-06, 9.743749e-06,
  6.056453e-06, 8.469916e-06, 1.07564e-05, 1.410879e-05, 1.782135e-05, 
    3.505436e-05, 1.372171e-05, 8.759572e-06, 1.125989e-05, 1.41462e-05, 
    1.429927e-05, 1.415201e-05, 1.379904e-05, 1.508085e-05, 1.458048e-05,
  9.264037e-06, 8.95533e-06, 1.378768e-05, 2.315024e-05, 2.604762e-05, 
    2.235982e-05, 1.155176e-05, 7.701356e-06, 1.49628e-05, 1.712163e-05, 
    1.629281e-05, 1.981303e-05, 2.136935e-05, 2.10313e-05, 2.164822e-05,
  9.475921e-06, 1.194752e-05, 1.488484e-05, 2.899218e-05, 2.812499e-05, 
    1.58839e-05, 1.23809e-05, 1.16637e-05, 1.689991e-05, 2.422357e-05, 
    2.404934e-05, 2.492846e-05, 2.649352e-05, 2.673895e-05, 3.065555e-05,
  1.106687e-05, 1.472173e-05, 2.018027e-05, 3.243724e-05, 3.037514e-05, 
    2.040722e-05, 1.334112e-05, 1.507572e-05, 2.738911e-05, 2.713702e-05, 
    3.04758e-05, 3.392647e-05, 3.173244e-05, 3.784389e-05, 3.807967e-05,
  1.591336e-05, 1.587028e-05, 2.3712e-05, 3.760948e-05, 3.40891e-05, 
    2.156843e-05, 1.713413e-05, 2.164813e-05, 3.088614e-05, 3.476642e-05, 
    3.161396e-05, 3.330483e-05, 4.013565e-05, 4.259626e-05, 4.044155e-05,
  1.267992e-05, 1.824001e-05, 3.112842e-05, 4.050641e-05, 4.161309e-05, 
    2.6075e-05, 1.892045e-05, 3.204603e-05, 4.604702e-05, 3.687431e-05, 
    4.2773e-05, 4.428589e-05, 3.968645e-05, 4.188087e-05, 4.649321e-05,
  1.830845e-05, 2.134176e-05, 3.597575e-05, 5.174385e-05, 4.01953e-05, 
    3.077588e-05, 2.653526e-05, 4.050565e-05, 4.908596e-05, 7.378736e-05, 
    6.691929e-05, 5.153513e-05, 4.680461e-05, 6.911075e-05, 4.822647e-05,
  1.635455e-05, 1.993967e-05, 1.964763e-05, 2.336802e-05, 2.561802e-05, 
    2.647443e-05, 2.384633e-05, 2.468465e-05, 2.944087e-05, 2.431285e-05, 
    2.47548e-05, 2.402177e-05, 2.086633e-05, 2.106606e-05, 1.624779e-05,
  1.987634e-05, 2.273011e-05, 2.576375e-05, 3.057503e-05, 3.722795e-05, 
    3.443259e-05, 4.346653e-05, 3.2115e-05, 4.032426e-05, 3.183535e-05, 
    2.767069e-05, 2.489761e-05, 2.159438e-05, 1.969152e-05, 1.859312e-05,
  2.584668e-05, 3.23605e-05, 4.141071e-05, 5.681102e-05, 6.691881e-05, 
    5.390992e-05, 4.712676e-05, 4.829778e-05, 4.201403e-05, 4.409291e-05, 
    3.309039e-05, 2.393004e-05, 2.263286e-05, 1.912681e-05, 2.058057e-05,
  3.25923e-05, 4.842186e-05, 5.521656e-05, 8.436671e-05, 7.394433e-05, 
    6.299739e-05, 6.845046e-05, 5.275887e-05, 6.271909e-05, 4.457531e-05, 
    3.993668e-05, 3.312947e-05, 2.900243e-05, 2.240583e-05, 1.634576e-05,
  3.071338e-05, 4.951608e-05, 8.017123e-05, 8.17295e-05, 8.695692e-05, 
    6.455679e-05, 6.08712e-05, 6.229679e-05, 6.076592e-05, 5.068547e-05, 
    4.740836e-05, 4.519976e-05, 3.4622e-05, 2.500509e-05, 2.057218e-05,
  3.22075e-05, 5.104526e-05, 8.748494e-05, 8.613885e-05, 9.266409e-05, 
    8.597306e-05, 6.496556e-05, 6.788242e-05, 5.412708e-05, 5.000042e-05, 
    5.008634e-05, 4.393215e-05, 3.02943e-05, 3.12232e-05, 2.20319e-05,
  3.488662e-05, 5.977214e-05, 9.62195e-05, 9.859374e-05, 0.0001002759, 
    7.380731e-05, 6.605998e-05, 6.546084e-05, 5.835593e-05, 4.038116e-05, 
    3.125489e-05, 3.363026e-05, 2.814599e-05, 2.791437e-05, 2.357358e-05,
  3.537066e-05, 6.784448e-05, 0.0001111757, 0.000105139, 8.647778e-05, 
    8.971382e-05, 7.426868e-05, 6.618474e-05, 5.252418e-05, 4.068936e-05, 
    3.065e-05, 3.126116e-05, 2.425119e-05, 2.11856e-05, 1.962197e-05,
  3.588909e-05, 8.040226e-05, 0.0001155537, 0.0001095877, 0.0001009206, 
    8.246744e-05, 6.348094e-05, 5.503525e-05, 5.479521e-05, 2.374405e-05, 
    2.265922e-05, 2.158511e-05, 1.754153e-05, 1.648556e-05, 1.569378e-05,
  2.133801e-05, 7.397844e-05, 0.0001225021, 0.0001192237, 9.845754e-05, 
    8.385882e-05, 5.650293e-05, 4.408767e-05, 3.392537e-05, 2.574714e-05, 
    2.50814e-05, 2.544479e-05, 2.242911e-05, 1.612589e-05, 1.426198e-05,
  2.559672e-05, 2.278377e-05, 1.750602e-05, 9.537897e-06, 4.943145e-06, 
    3.446511e-06, 2.509127e-06, 3.415332e-06, 3.688533e-06, 4.09922e-06, 
    2.231428e-06, 3.978412e-06, 2.872664e-06, 1.901022e-06, 6.629072e-06,
  3.307249e-05, 1.701172e-05, 2.482541e-05, 9.12371e-06, 4.640989e-06, 
    4.975268e-06, 4.900014e-06, 4.045543e-06, 4.377397e-06, 3.829157e-06, 
    5.352708e-06, 4.293001e-06, 3.630494e-06, 2.99372e-06, 5.567959e-06,
  2.837849e-05, 1.571023e-05, 1.058127e-05, 4.444043e-06, 3.566554e-06, 
    5.052315e-06, 5.402161e-06, 6.018937e-06, 4.817885e-06, 4.761982e-06, 
    4.878987e-06, 3.816181e-06, 4.642655e-06, 2.189221e-06, 4.553668e-06,
  4.464659e-05, 2.871236e-05, 1.126517e-05, 4.09252e-06, 4.922519e-06, 
    5.636581e-06, 6.033116e-06, 6.01999e-06, 5.911339e-06, 6.840619e-06, 
    5.22825e-06, 5.437397e-06, 6.046145e-06, 3.810195e-06, 3.583649e-06,
  5.515493e-05, 3.136681e-05, 5.398079e-06, 3.833299e-06, 5.247477e-06, 
    6.130966e-06, 6.666261e-06, 6.823946e-06, 7.448232e-06, 7.242127e-06, 
    6.709823e-06, 6.197904e-06, 6.023396e-06, 6.408018e-06, 5.049934e-06,
  3.073393e-05, 1.663023e-05, 1.026344e-05, 3.72874e-06, 4.840297e-06, 
    6.806432e-06, 7.126825e-06, 6.65208e-06, 9.322433e-06, 8.93385e-06, 
    8.543969e-06, 7.990139e-06, 7.093203e-06, 6.544874e-06, 8.279121e-06,
  3.476431e-05, 2.730329e-05, 1.010628e-05, 3.326573e-06, 5.333495e-06, 
    6.537293e-06, 6.80809e-06, 8.390476e-06, 1.100588e-05, 1.163712e-05, 
    8.161272e-06, 8.959542e-06, 1.115881e-05, 7.130311e-06, 1.124397e-05,
  3.978487e-05, 2.425338e-05, 8.265338e-06, 4.117418e-06, 4.485878e-06, 
    5.119202e-06, 5.952725e-06, 8.621174e-06, 9.194072e-06, 9.820295e-06, 
    1.177778e-05, 1.06718e-05, 1.171372e-05, 9.074682e-06, 1.075974e-05,
  5.294154e-05, 3.177109e-05, 1.336569e-05, 2.940333e-06, 5.124261e-06, 
    5.916166e-06, 8.294134e-06, 8.92428e-06, 8.880258e-06, 9.98186e-06, 
    1.281817e-05, 1.452126e-05, 1.158304e-05, 1.213544e-05, 1.227866e-05,
  4.69899e-05, 3.760617e-05, 1.686963e-05, 4.654813e-06, 5.502209e-06, 
    7.374577e-06, 8.315726e-06, 1.11113e-05, 1.135888e-05, 1.128038e-05, 
    1.422643e-05, 1.66494e-05, 1.53784e-05, 1.456394e-05, 1.585053e-05,
  5.662572e-06, 5.763882e-06, 5.294641e-06, 5.756087e-06, 6.164966e-06, 
    4.948184e-06, 4.946303e-06, 7.084302e-06, 5.95748e-06, 5.782872e-06, 
    4.913935e-06, 4.389346e-06, 5.601878e-06, 6.164858e-06, 7.14372e-06,
  6.308681e-06, 6.763687e-06, 6.721386e-06, 6.91026e-06, 5.953577e-06, 
    6.239297e-06, 7.048372e-06, 6.623207e-06, 7.447336e-06, 7.60767e-06, 
    7.271417e-06, 5.40128e-06, 6.407492e-06, 6.315709e-06, 7.199252e-06,
  7.648235e-06, 7.602652e-06, 7.47286e-06, 7.852294e-06, 8.189888e-06, 
    8.435036e-06, 7.500371e-06, 7.403602e-06, 7.651364e-06, 9.469727e-06, 
    6.489207e-06, 5.276936e-06, 6.430679e-06, 6.596718e-06, 6.202828e-06,
  9.599753e-06, 1.001302e-05, 9.577812e-06, 9.914855e-06, 9.4516e-06, 
    8.324413e-06, 6.733464e-06, 8.263851e-06, 8.844214e-06, 8.352235e-06, 
    7.930497e-06, 8.735242e-06, 6.413117e-06, 6.253691e-06, 6.262655e-06,
  1.110729e-05, 1.061848e-05, 1.019072e-05, 1.096794e-05, 9.413418e-06, 
    9.628868e-06, 7.646401e-06, 9.40201e-06, 6.477249e-06, 7.181484e-06, 
    9.583264e-06, 5.555135e-06, 5.858296e-06, 5.544034e-06, 5.734229e-06,
  1.141593e-05, 1.277706e-05, 1.00491e-05, 1.212899e-05, 1.012857e-05, 
    9.669227e-06, 1.027243e-05, 8.12824e-06, 7.218489e-06, 7.559037e-06, 
    6.49097e-06, 5.155723e-06, 5.587655e-06, 5.270688e-06, 5.815125e-06,
  1.196722e-05, 1.409957e-05, 1.371689e-05, 1.281126e-05, 1.358116e-05, 
    1.203501e-05, 9.624907e-06, 8.143917e-06, 6.977555e-06, 6.933161e-06, 
    6.867158e-06, 6.785511e-06, 5.282326e-06, 4.617337e-06, 5.495656e-06,
  1.227424e-05, 1.399514e-05, 1.455158e-05, 1.46161e-05, 1.414026e-05, 
    1.378798e-05, 1.197089e-05, 1.069825e-05, 9.174648e-06, 6.962945e-06, 
    7.655625e-06, 6.636738e-06, 5.364081e-06, 4.233088e-06, 3.46338e-06,
  1.35465e-05, 1.469442e-05, 1.328433e-05, 1.510472e-05, 1.594228e-05, 
    1.410923e-05, 1.373713e-05, 1.318485e-05, 9.323848e-06, 6.349043e-06, 
    8.25849e-06, 6.43172e-06, 7.200982e-06, 4.584326e-06, 4.187229e-06,
  1.020048e-05, 1.175789e-05, 1.561809e-05, 1.443265e-05, 1.7956e-05, 
    1.431513e-05, 1.659815e-05, 1.215092e-05, 8.384071e-06, 8.559598e-06, 
    9.566211e-06, 6.886767e-06, 5.746477e-06, 5.186672e-06, 4.011187e-06,
  4.711659e-06, 4.505951e-06, 3.674388e-06, 1.067215e-06, 2.763807e-06, 
    2.305399e-06, 1.312572e-06, 1.776399e-06, 2.153749e-06, 2.088856e-06, 
    3.47526e-06, 4.091192e-06, 4.31026e-06, 5.338996e-06, 6.654971e-06,
  3.680962e-06, 2.88282e-06, 2.049467e-06, 1.683224e-06, 8.743359e-07, 
    4.634357e-07, 3.740645e-07, 6.102829e-07, 2.785364e-07, 1.088592e-06, 
    1.745387e-06, 1.738985e-06, 2.71766e-06, 1.969342e-06, 5.061856e-06,
  3.384732e-06, 3.14004e-06, 8.513039e-07, 7.805272e-07, 3.686418e-08, 
    6.961508e-11, 7.273777e-09, 2.02529e-07, 3.852112e-07, 5.435614e-07, 
    2.152086e-06, 3.034795e-06, 1.397416e-06, 1.476758e-06, 2.138752e-06,
  3.080708e-06, 1.452629e-06, 3.672389e-07, 2.179464e-07, 1.658144e-08, 
    1.204521e-08, 1.426322e-09, 1.63235e-07, 2.425726e-07, 7.572704e-07, 
    4.918393e-07, 6.370361e-07, 1.712323e-06, 1.111207e-06, 1.664318e-06,
  3.127811e-06, 1.529743e-06, 6.45768e-08, 2.153243e-08, 6.222602e-09, 
    9.882068e-09, 8.347627e-08, 1.216074e-07, 2.948008e-07, 1.666109e-07, 
    4.63092e-08, 2.783553e-07, 2.545453e-07, 9.178113e-07, 2.467333e-06,
  3.898196e-06, 1.001543e-06, 2.826536e-07, 1.291767e-07, 1.733304e-07, 
    5.307718e-08, 4.380427e-09, 2.011285e-07, 3.371563e-07, 2.298163e-07, 
    4.650452e-08, 1.906536e-07, 1.061969e-06, 1.203555e-06, 1.395603e-06,
  3.529687e-06, 7.013084e-07, 7.661181e-07, 2.289864e-07, 3.9071e-07, 
    3.099512e-07, 1.387402e-08, 1.698918e-07, 2.883542e-07, 1.65448e-07, 
    2.925006e-07, 3.540796e-07, 1.16155e-06, 1.587424e-06, 1.713625e-06,
  1.796304e-06, 5.238138e-07, 6.200879e-07, 1.884635e-07, 5.146278e-08, 
    4.051565e-08, 2.198318e-08, 2.475649e-08, 4.162323e-07, 2.34072e-07, 
    2.397602e-07, 4.464434e-07, 1.309618e-06, 1.550853e-06, 2.052844e-06,
  2.309637e-06, 7.879394e-07, 1.081862e-06, 1.7041e-06, 6.521407e-07, 
    2.905337e-07, 5.842071e-07, 9.328893e-08, 4.972924e-07, 4.81056e-07, 
    4.248556e-07, 4.520835e-07, 9.327067e-07, 1.921054e-06, 6.670961e-06,
  3.341354e-06, 1.538119e-06, 1.204681e-06, 1.541116e-06, 1.64077e-06, 
    4.968376e-07, 4.957619e-07, 2.046121e-06, 2.763217e-06, 1.70802e-06, 
    4.471702e-07, 3.229404e-07, 5.8117e-07, 3.593096e-06, 8.42693e-06,
  2.620211e-07, 7.359373e-08, 1.953029e-06, 3.155249e-06, 4.165704e-06, 
    5.908835e-06, 6.203654e-06, 6.300085e-06, 6.952667e-06, 5.742438e-06, 
    6.346012e-06, 3.774564e-06, 4.794691e-06, 4.474807e-06, 3.264918e-06,
  7.593602e-07, 3.740681e-07, 1.090623e-06, 2.262261e-06, 6.361381e-06, 
    8.601326e-06, 6.838166e-06, 7.127125e-06, 6.064212e-06, 7.265986e-06, 
    7.179471e-06, 6.790947e-06, 5.910607e-06, 3.99571e-06, 3.20619e-06,
  1.26676e-06, 1.367601e-07, 1.02495e-06, 3.177578e-06, 5.332632e-06, 
    1.077376e-05, 9.729335e-06, 1.085465e-05, 6.993035e-06, 5.911819e-06, 
    7.072537e-06, 7.076724e-06, 6.47272e-06, 3.833024e-06, 4.296611e-06,
  2.870929e-06, 5.737772e-07, 1.765137e-06, 3.208252e-06, 7.42662e-06, 
    1.377969e-05, 8.691346e-06, 5.754615e-06, 6.576371e-06, 6.681736e-06, 
    6.692058e-06, 4.224858e-06, 3.632315e-06, 3.573724e-06, 5.794614e-06,
  4.975836e-07, 1.178097e-06, 3.630169e-06, 3.349769e-06, 9.04654e-06, 
    1.08202e-05, 6.671285e-06, 6.276091e-06, 6.137423e-06, 6.447543e-06, 
    4.015689e-06, 4.81674e-06, 5.656373e-06, 7.410818e-06, 9.084633e-06,
  6.652283e-07, 1.005951e-06, 2.752307e-06, 4.099367e-06, 9.657369e-06, 
    8.827183e-06, 4.199238e-06, 5.296802e-06, 3.727105e-06, 3.758956e-06, 
    3.305692e-06, 5.678568e-06, 9.646167e-06, 1.086891e-05, 1.558973e-05,
  2.194968e-06, 1.25703e-06, 4.178731e-06, 6.706958e-06, 9.601281e-06, 
    7.025881e-06, 2.196039e-06, 3.83194e-06, 2.459704e-06, 4.184565e-06, 
    3.875856e-06, 8.663535e-06, 2.02526e-05, 2.959128e-05, 3.790742e-05,
  2.68659e-06, 2.468942e-06, 3.143447e-06, 6.658935e-06, 1.257507e-05, 
    7.875926e-06, 4.540032e-06, 4.871923e-06, 7.342177e-06, 1.059563e-05, 
    2.118963e-05, 3.800977e-05, 4.813707e-05, 5.289389e-05, 6.013347e-05,
  3.051762e-06, 4.227619e-06, 5.807019e-06, 7.557512e-06, 1.036279e-05, 
    1.179121e-05, 7.270513e-06, 1.086367e-05, 2.107256e-05, 4.304395e-05, 
    6.289101e-05, 7.512597e-05, 7.532963e-05, 7.157534e-05, 6.531579e-05,
  4.910351e-06, 5.309004e-06, 6.049516e-06, 7.062225e-06, 1.251059e-05, 
    1.363535e-05, 2.231863e-05, 5.626881e-05, 7.901062e-05, 8.681827e-05, 
    8.439994e-05, 7.540188e-05, 5.858502e-05, 4.409423e-05, 3.335948e-05,
  2.586799e-06, 7.021888e-06, 1.068154e-05, 1.075987e-05, 4.488063e-06, 
    1.826308e-06, 2.399196e-06, 3.056633e-06, 2.695183e-06, 2.410068e-06, 
    2.449943e-06, 1.45665e-06, 8.770371e-07, 1.316882e-06, 1.370658e-06,
  3.335536e-06, 5.320127e-06, 5.754025e-06, 6.962669e-06, 3.963731e-06, 
    3.479618e-06, 2.89077e-06, 2.854791e-06, 3.025465e-06, 2.914649e-06, 
    2.721125e-06, 2.949226e-06, 3.211572e-06, 1.527356e-06, 8.178723e-07,
  1.948918e-06, 5.261681e-06, 6.932607e-06, 5.881516e-06, 3.760666e-06, 
    2.899733e-06, 2.660653e-06, 2.552906e-06, 3.200248e-06, 2.967485e-06, 
    3.506252e-06, 4.463655e-06, 3.799514e-06, 2.135508e-06, 2.091057e-06,
  3.165654e-06, 8.232201e-06, 7.654515e-06, 7.15935e-06, 4.392814e-06, 
    1.791176e-06, 2.001184e-06, 2.427097e-06, 3.641734e-06, 4.251585e-06, 
    4.851523e-06, 5.767617e-06, 6.910837e-06, 1.183185e-05, 1.001608e-05,
  6.383325e-06, 1.190905e-05, 8.823805e-06, 4.819291e-06, 2.844779e-06, 
    1.974208e-06, 2.594419e-06, 3.267081e-06, 4.782543e-06, 6.188853e-06, 
    1.062036e-05, 1.309563e-05, 1.036376e-05, 1.004255e-05, 1.121535e-05,
  8.888173e-06, 1.052844e-05, 6.955713e-06, 4.160812e-06, 3.397519e-06, 
    4.396029e-06, 5.47543e-06, 6.810892e-06, 9.503128e-06, 1.273511e-05, 
    2.034255e-05, 2.391852e-05, 2.599738e-05, 1.697046e-05, 1.275899e-05,
  1.277614e-05, 8.079602e-06, 7.593983e-06, 5.234311e-06, 8.060838e-06, 
    8.379838e-06, 9.254221e-06, 7.1747e-06, 7.742196e-06, 1.135966e-05, 
    1.78909e-05, 2.317429e-05, 2.669096e-05, 2.330364e-05, 2.038942e-05,
  1.09615e-05, 7.69639e-06, 7.116277e-06, 7.977979e-06, 8.372523e-06, 
    9.320491e-06, 5.977467e-06, 4.100146e-06, 1.619207e-06, 7.939141e-07, 
    3.576832e-06, 6.063006e-06, 7.962775e-06, 1.12853e-05, 1.113643e-05,
  1.145186e-05, 8.116534e-06, 6.575555e-06, 5.838853e-06, 8.932831e-06, 
    5.210311e-06, 5.377634e-06, 3.047295e-06, 3.23287e-06, 1.91629e-06, 
    2.236971e-06, 2.231323e-06, 2.420006e-06, 2.302719e-06, 4.73949e-06,
  1.199642e-05, 1.139064e-05, 9.839233e-06, 6.624257e-06, 5.449642e-06, 
    3.968199e-06, 1.588483e-06, 5.777701e-07, 1.168234e-06, 1.105448e-06, 
    1.15298e-06, 1.3682e-06, 1.229741e-06, 8.96204e-07, 1.308346e-06,
  7.509945e-06, 1.087572e-05, 6.344956e-06, 3.227417e-06, 3.955977e-06, 
    3.023703e-06, 3.408161e-06, 2.13345e-06, 2.262195e-06, 2.502314e-06, 
    1.559738e-06, 1.661399e-06, 1.421892e-06, 1.581282e-06, 2.669599e-06,
  5.835218e-06, 5.080335e-06, 3.865127e-06, 3.100456e-06, 2.811201e-06, 
    1.244201e-06, 2.249373e-06, 2.362238e-06, 2.507522e-06, 2.451045e-06, 
    2.787097e-06, 2.683251e-06, 1.782178e-06, 1.324221e-06, 9.921073e-07,
  7.148778e-06, 4.679654e-06, 3.017713e-06, 2.031283e-06, 1.917341e-06, 
    1.208614e-06, 9.726594e-07, 1.505753e-06, 2.615091e-06, 2.779217e-06, 
    3.140942e-06, 2.242833e-06, 2.976913e-06, 2.863165e-06, 4.183052e-06,
  4.162814e-06, 3.037934e-06, 1.975855e-06, 2.187566e-06, 2.487693e-06, 
    1.268224e-06, 1.14071e-06, 3.488856e-06, 4.484214e-06, 3.980338e-06, 
    5.011719e-06, 2.358652e-06, 6.475696e-06, 7.719036e-06, 7.14959e-06,
  7.437254e-07, 1.636043e-06, 1.274572e-06, 2.917845e-06, 2.807527e-06, 
    5.261283e-06, 1.377797e-06, 1.156932e-05, 6.585837e-06, 5.616799e-06, 
    3.937919e-06, 4.496546e-06, 4.959174e-06, 6.562691e-06, 9.369394e-06,
  2.013591e-06, 3.12151e-06, 6.490052e-06, 5.464556e-06, 4.041477e-06, 
    1.262155e-06, 6.661703e-06, 7.101243e-06, 9.519807e-06, 9.308423e-06, 
    5.256838e-06, 7.5313e-06, 6.681083e-06, 6.872124e-06, 6.799567e-06,
  5.655039e-06, 7.470261e-06, 1.162097e-05, 1.262866e-05, 6.198881e-06, 
    4.082036e-06, 4.483987e-06, 9.532434e-06, 1.608643e-05, 1.365158e-05, 
    9.780585e-06, 9.600192e-06, 8.192345e-06, 7.460185e-06, 9.653282e-06,
  8.468754e-06, 1.258323e-05, 1.168084e-05, 9.909519e-06, 9.209222e-06, 
    5.068521e-06, 4.992173e-08, 8.366394e-06, 1.652582e-05, 2.099992e-05, 
    1.8225e-05, 1.684279e-05, 1.085921e-05, 1.615201e-05, 1.329346e-05,
  7.775522e-06, 8.218531e-06, 4.635646e-06, 5.956571e-06, 8.519759e-06, 
    8.143395e-06, 5.159123e-06, 2.857754e-06, 5.051775e-06, 9.449882e-06, 
    1.248287e-05, 1.654308e-05, 1.463257e-05, 1.516763e-05, 1.076379e-05,
  3.900293e-06, 3.253787e-06, 3.013339e-06, 3.023408e-06, 4.810701e-06, 
    8.212146e-06, 9.276033e-06, 7.030494e-06, 4.920947e-06, 6.966693e-06, 
    9.768655e-06, 1.209659e-05, 9.293284e-06, 8.900663e-06, 8.403851e-06,
  6.272885e-06, 6.279182e-06, 4.747043e-06, 2.927929e-06, 1.941603e-06, 
    3.772874e-06, 6.037522e-06, 5.066514e-06, 4.820091e-06, 2.750767e-06, 
    2.206424e-06, 1.445626e-06, 8.745566e-07, 4.539116e-07, 1.292756e-06,
  7.49288e-06, 5.489647e-06, 3.7649e-06, 1.679454e-06, 2.813994e-06, 
    4.057916e-06, 5.764085e-06, 7.902235e-06, 7.672256e-06, 3.402677e-06, 
    3.954186e-06, 3.472404e-06, 3.893478e-06, 2.441336e-06, 1.637356e-06,
  6.148873e-06, 7.583751e-06, 2.244784e-06, 6.627253e-07, 1.646677e-06, 
    3.614345e-06, 7.597102e-06, 1.407096e-05, 1.236053e-05, 1.19389e-05, 
    1.117834e-05, 8.037548e-06, 5.909141e-06, 5.98099e-06, 3.268705e-06,
  5.399437e-06, 5.401624e-06, 2.225519e-06, 5.432122e-07, 9.625494e-07, 
    7.75936e-06, 1.892749e-05, 2.217517e-05, 1.511768e-05, 1.263958e-05, 
    9.773038e-06, 9.417851e-06, 8.754781e-06, 1.03177e-05, 1.13642e-05,
  3.789801e-06, 4.580205e-06, 2.592813e-06, 1.576913e-06, 3.35885e-06, 
    1.798669e-05, 2.2896e-05, 2.089942e-05, 4.647679e-06, 4.824306e-06, 
    6.911485e-06, 7.029232e-06, 5.048472e-06, 6.574338e-06, 9.84098e-06,
  4.247977e-06, 5.327981e-06, 3.435731e-06, 2.484497e-06, 3.914568e-06, 
    1.543177e-05, 2.012785e-05, 9.83457e-06, 2.814814e-06, 8.678005e-06, 
    9.058811e-06, 1.003672e-05, 6.24236e-06, 8.301441e-06, 6.609318e-06,
  1.732323e-05, 1.566958e-05, 1.076922e-05, 4.723567e-06, 3.649619e-06, 
    1.534068e-05, 1.770192e-05, 8.06357e-06, 6.056522e-06, 8.079828e-06, 
    7.012672e-06, 7.437394e-06, 9.377669e-06, 1.083584e-05, 6.941681e-06,
  2.267049e-05, 2.366712e-05, 2.12254e-05, 7.513632e-06, 1.543845e-06, 
    1.503399e-05, 1.259628e-05, 1.055013e-05, 5.974484e-06, 9.723399e-06, 
    1.159027e-05, 1.494944e-05, 1.196101e-05, 1.065205e-05, 8.209188e-06,
  9.608531e-06, 3.729065e-06, 6.406661e-06, 6.423835e-06, 1.736105e-06, 
    6.229828e-06, 1.559333e-05, 1.171467e-05, 1.151269e-05, 1.325084e-05, 
    1.482043e-05, 1.383963e-05, 1.352641e-05, 5.156314e-06, 1.040642e-05,
  1.884634e-06, 2.665167e-06, 7.574448e-06, 5.435607e-06, 4.237771e-06, 
    3.610085e-06, 1.541933e-05, 1.932978e-05, 1.082477e-05, 1.8433e-05, 
    1.721433e-05, 6.9996e-06, 7.093495e-06, 5.719193e-06, 1.048372e-05,
  3.344212e-06, 2.199086e-06, 4.482278e-06, 6.441544e-06, 9.912318e-06, 
    9.728917e-06, 8.658498e-06, 8.250929e-06, 6.183911e-06, 5.242248e-06, 
    2.084558e-06, 1.988616e-06, 2.46686e-06, 2.186457e-06, 4.070481e-06,
  4.030818e-06, 3.060192e-06, 3.987673e-06, 6.384942e-06, 5.386194e-06, 
    4.962346e-06, 7.071912e-06, 8.90067e-06, 3.753899e-06, 4.188038e-06, 
    3.381509e-06, 3.980541e-06, 4.119421e-06, 1.454444e-06, 2.874402e-06,
  3.345972e-06, 3.210235e-06, 3.770306e-06, 6.166413e-06, 4.857434e-06, 
    6.924165e-06, 3.875772e-06, 4.655285e-06, 3.702802e-06, 2.074686e-06, 
    2.551674e-06, 2.809812e-06, 3.291281e-06, 1.95025e-06, 2.462594e-06,
  3.380989e-06, 2.001035e-06, 2.918757e-06, 4.985737e-06, 3.280531e-06, 
    4.545363e-06, 3.76404e-06, 3.617532e-06, 3.047129e-06, 3.974531e-06, 
    3.474306e-06, 1.450629e-06, 3.989211e-06, 3.555007e-06, 3.532259e-06,
  3.338242e-06, 3.518764e-06, 2.26919e-06, 5.516079e-06, 5.541842e-06, 
    5.578466e-06, 4.77682e-06, 4.376262e-06, 4.210738e-06, 2.647863e-06, 
    3.234074e-06, 1.498765e-06, 2.378067e-06, 3.632627e-06, 4.809328e-06,
  6.002183e-06, 4.564103e-06, 4.702291e-06, 5.322724e-06, 8.584367e-06, 
    8.194825e-06, 5.357669e-06, 4.050588e-06, 5.633156e-06, 6.596958e-06, 
    5.340653e-06, 3.171374e-06, 3.626502e-07, 2.244412e-06, 4.076183e-06,
  1.40816e-05, 1.180938e-05, 6.214132e-06, 4.596391e-06, 8.667083e-06, 
    8.215255e-06, 4.966028e-06, 4.350271e-06, 5.346442e-06, 5.162664e-06, 
    4.160363e-06, 5.070359e-06, 4.780076e-06, 1.969726e-06, 1.148642e-07,
  1.451951e-05, 1.316508e-05, 8.169632e-06, 6.966981e-06, 8.88663e-06, 
    7.97185e-06, 6.136997e-06, 4.740135e-06, 5.082684e-06, 4.409158e-06, 
    7.382623e-06, 7.567494e-06, 7.499893e-06, 3.319511e-06, 2.661104e-07,
  7.327432e-06, 6.136593e-06, 3.753793e-06, 8.898553e-06, 1.739534e-05, 
    9.780716e-06, 7.997177e-06, 6.009016e-06, 5.387912e-06, 4.42106e-06, 
    6.298811e-06, 6.40889e-06, 6.546939e-06, 6.451482e-06, 4.064063e-06,
  1.680088e-06, 8.9008e-07, 5.38651e-06, 1.026666e-05, 1.179793e-05, 
    7.935178e-06, 9.157719e-06, 8.408747e-06, 6.090633e-06, 3.565981e-06, 
    4.646306e-06, 5.227694e-06, 6.099385e-06, 6.91419e-06, 6.418155e-06,
  5.91656e-06, 4.906312e-06, 3.306375e-06, 4.987246e-06, 1.227693e-06, 
    2.350386e-06, 2.233038e-06, 1.45866e-06, 5.848422e-07, 1.659769e-06, 
    3.098987e-06, 3.900012e-06, 3.91302e-06, 2.89625e-06, 5.625001e-08,
  6.373164e-06, 4.40925e-06, 3.683803e-06, 3.048867e-06, 1.068975e-06, 
    1.422985e-06, 2.237288e-06, 2.544303e-06, 9.920363e-07, 1.48738e-07, 
    1.691199e-06, 3.075131e-06, 4.56048e-06, 3.704763e-06, 2.430733e-06,
  5.978249e-06, 3.646538e-06, 4.886508e-06, 3.296421e-06, 1.915499e-06, 
    2.088035e-06, 2.539305e-06, 2.916199e-06, 2.509703e-06, 4.204462e-07, 
    1.633738e-06, 8.797221e-07, 4.981617e-06, 9.84798e-06, 6.434459e-06,
  6.240115e-06, 7.02016e-06, 5.764735e-06, 4.508923e-06, 3.174891e-06, 
    2.95356e-06, 3.707795e-06, 3.045498e-06, 2.662276e-06, 2.940281e-06, 
    9.386451e-07, 3.543181e-07, 9.189335e-06, 2.350824e-05, 1.579883e-05,
  7.903715e-06, 8.883551e-06, 1.061192e-05, 8.903107e-06, 7.628797e-06, 
    6.915261e-06, 6.215574e-06, 3.779545e-06, 2.952015e-06, 2.583263e-06, 
    1.628119e-06, 4.038295e-07, 1.396911e-05, 5.495684e-05, 3.876148e-05,
  7.670051e-06, 8.778522e-06, 8.32606e-06, 9.389324e-06, 9.070341e-06, 
    9.606275e-06, 6.799962e-06, 3.732245e-06, 2.62068e-06, 5.149357e-06, 
    1.885363e-06, 1.182234e-06, 1.73118e-05, 7.049152e-05, 7.330482e-05,
  6.999749e-06, 8.637752e-06, 9.685933e-06, 1.018856e-05, 9.275917e-06, 
    7.296791e-06, 4.942423e-06, 3.943871e-06, 3.228168e-06, 6.035049e-06, 
    6.378684e-06, 3.644131e-06, 7.345773e-06, 6.08712e-05, 0.0001028648,
  8.149193e-06, 1.128942e-05, 1.248454e-05, 9.083478e-06, 4.735667e-06, 
    7.016451e-06, 3.444365e-06, 2.481052e-06, 3.591388e-06, 1.031063e-05, 
    7.902025e-06, 6.938767e-06, 5.743378e-06, 3.853985e-05, 0.0001242448,
  9.051173e-06, 1.169389e-05, 8.72804e-06, 7.47453e-06, 6.189103e-06, 
    3.075978e-06, 7.325519e-06, 4.609277e-06, 5.411388e-06, 1.007808e-05, 
    1.321891e-05, 9.961673e-06, 1.262688e-05, 3.27474e-05, 0.0001538958,
  1.07138e-05, 1.201651e-05, 7.601637e-06, 4.042565e-06, 4.182096e-06, 
    6.665721e-07, 5.537164e-06, 6.826984e-06, 4.840394e-06, 6.400261e-06, 
    8.587574e-06, 9.906594e-06, 1.048068e-05, 3.596005e-05, 0.0001516696,
  3.190635e-06, 4.461288e-06, 5.804058e-06, 6.03029e-06, 6.429078e-06, 
    5.194946e-06, 6.827847e-06, 9.305717e-06, 2.095385e-05, 5.367117e-05, 
    1.374324e-05, 5.912299e-05, 2.810755e-05, 8.543153e-06, 4.599973e-06,
  3.819811e-06, 5.703049e-06, 4.495718e-06, 7.368703e-06, 4.822696e-06, 
    3.481799e-06, 4.267975e-06, 8.305635e-06, 5.874743e-06, 1.758949e-05, 
    5.902499e-06, 6.179231e-05, 4.649494e-05, 7.841318e-06, 1.437736e-05,
  4.463222e-06, 2.542803e-06, 6.063513e-06, 3.941253e-06, 4.879829e-06, 
    4.499182e-06, 3.689258e-06, 7.971921e-06, 5.506053e-06, 5.287771e-06, 
    1.981614e-06, 5.933123e-05, 7.122522e-05, 5.673639e-06, 4.923855e-06,
  5.139185e-06, 5.698114e-06, 4.956452e-06, 5.713325e-06, 5.964072e-06, 
    5.780689e-06, 4.376293e-06, 9.909459e-06, 4.472426e-06, 4.208533e-06, 
    1.621517e-06, 3.004255e-05, 0.0001056901, 8.689694e-06, 5.495994e-06,
  8.081406e-06, 8.051811e-06, 7.657068e-06, 5.108289e-06, 7.230995e-06, 
    7.555266e-06, 4.59886e-06, 6.836479e-06, 4.013771e-06, 2.703651e-06, 
    9.996218e-07, 1.568408e-05, 0.0001197802, 4.357349e-05, 7.872879e-06,
  9.204106e-06, 1.094394e-05, 8.894691e-06, 6.309905e-06, 5.523576e-06, 
    4.519442e-06, 3.812963e-06, 5.486831e-06, 4.61731e-06, 3.260552e-06, 
    1.090094e-06, 6.949625e-06, 9.860902e-05, 0.0001171704, 2.199165e-05,
  1.177264e-05, 9.246382e-06, 7.713697e-06, 7.277053e-06, 5.318328e-06, 
    1.381794e-06, 1.109474e-06, 4.184767e-06, 1.002513e-06, 5.743827e-07, 
    6.367518e-07, 1.159045e-06, 6.048208e-05, 0.0001738027, 0.0001340921,
  1.167378e-05, 9.092072e-06, 7.218929e-06, 5.584857e-06, 4.340081e-06, 
    5.804763e-06, 4.294381e-06, 2.682746e-07, 7.906652e-07, 6.554423e-07, 
    1.294007e-06, 5.307511e-07, 4.51733e-05, 0.0002085964, 0.0003026571,
  1.013591e-05, 1.073902e-05, 9.383403e-06, 6.863142e-06, 8.230933e-06, 
    9.428175e-06, 5.257577e-06, 2.843245e-06, 8.364649e-07, 1.466707e-06, 
    4.965781e-06, 1.923988e-06, 3.042306e-05, 0.0001758212, 0.0003998532,
  1.237636e-05, 1.198937e-05, 1.100865e-05, 1.010845e-05, 5.162767e-06, 
    7.884597e-06, 8.663611e-06, 4.959745e-06, 6.119064e-06, 3.721122e-06, 
    2.926329e-06, 3.606219e-06, 1.808002e-05, 0.000103679, 0.0004010977,
  4.389474e-06, 4.87621e-06, 4.577911e-06, 5.337796e-06, 5.738305e-06, 
    6.047242e-06, 8.473366e-05, 0.0001278968, 0.0001192323, 0.0001927798, 
    0.000188964, 7.644414e-05, 3.271489e-05, 1.939448e-05, 1.216892e-05,
  5.00542e-06, 4.258064e-06, 4.808629e-06, 4.59171e-06, 5.469546e-06, 
    3.526418e-06, 7.442804e-06, 4.895716e-05, 3.836884e-05, 9.684332e-05, 
    0.0001475135, 0.0001085052, 4.195494e-05, 1.546176e-05, 1.256014e-05,
  5.080237e-06, 4.239453e-06, 3.52083e-06, 5.177419e-06, 4.470761e-06, 
    3.208403e-06, 4.74234e-06, 1.457127e-05, 2.180227e-05, 4.961266e-05, 
    0.0001310868, 0.0001327374, 5.041822e-05, 8.804784e-06, 1.260489e-05,
  5.471425e-06, 5.301026e-06, 6.401276e-06, 5.345772e-06, 5.995098e-06, 
    4.032367e-06, 3.755996e-06, 5.066045e-06, 1.757446e-05, 2.843959e-05, 
    0.0001203705, 0.0001526651, 5.27447e-05, 5.100682e-06, 1.437682e-05,
  7.130781e-06, 6.742235e-06, 5.450173e-06, 5.288715e-06, 4.738391e-06, 
    3.543341e-06, 2.390241e-06, 3.943145e-06, 6.728471e-06, 1.972076e-05, 
    0.0001047423, 0.0001332894, 3.803311e-05, 2.578606e-06, 3.887572e-05,
  8.091734e-06, 6.398001e-06, 4.79473e-06, 7.336297e-06, 5.860288e-06, 
    3.491132e-06, 1.953168e-06, 4.558053e-06, 3.502974e-06, 9.904505e-06, 
    6.202778e-05, 9.693688e-05, 3.671651e-05, 8.11507e-06, 7.401502e-05,
  6.513247e-06, 7.328934e-06, 8.316586e-06, 1.241151e-05, 5.796211e-06, 
    3.7109e-06, 1.632432e-06, 6.69715e-07, 6.27368e-07, 2.905843e-06, 
    2.970126e-05, 7.363223e-05, 3.090044e-05, 4.526946e-05, 0.000127277,
  5.725198e-06, 5.447228e-06, 6.415163e-06, 4.190656e-06, 4.707529e-06, 
    5.3467e-06, 4.098762e-06, 3.686056e-07, 9.630738e-07, 2.772468e-07, 
    1.750991e-05, 6.59537e-05, 4.473179e-05, 0.0001262942, 0.0001753533,
  4.160461e-06, 4.190634e-06, 8.320501e-06, 5.821182e-06, 8.306846e-06, 
    1.022274e-05, 4.19804e-06, 1.936443e-06, 9.737512e-08, 4.018752e-08, 
    9.368589e-06, 6.202593e-05, 7.627192e-05, 0.0001832371, 0.0001996422,
  4.438255e-06, 3.79678e-06, 8.080432e-06, 1.200946e-05, 9.024279e-06, 
    1.05848e-05, 1.018798e-05, 5.408671e-06, 3.189574e-06, 2.910563e-08, 
    6.282818e-06, 5.29148e-05, 7.839489e-05, 0.0001791993, 0.0002013015,
  3.964486e-06, 4.00607e-06, 4.556964e-06, 5.062129e-06, 3.70466e-06, 
    3.129874e-06, 2.782325e-06, 7.936512e-06, 2.401578e-05, 4.200299e-05, 
    6.064101e-05, 9.318486e-05, 9.040356e-05, 0.000168276, 0.0002281974,
  4.563138e-06, 5.078747e-06, 4.205613e-06, 4.848958e-06, 3.825844e-06, 
    2.798604e-06, 2.826015e-06, 2.250781e-06, 3.037839e-06, 1.525236e-05, 
    1.507872e-05, 1.569505e-05, 2.771631e-05, 8.901704e-05, 0.0001510263,
  5.061819e-06, 3.977782e-06, 4.303698e-06, 3.780587e-06, 4.358163e-06, 
    4.987131e-06, 3.327264e-06, 2.086219e-06, 2.396139e-06, 2.255638e-06, 
    6.087869e-07, 9.95051e-07, 6.30039e-06, 3.384266e-05, 6.166815e-05,
  7.180271e-06, 6.918239e-06, 6.259228e-06, 5.319952e-06, 7.738297e-06, 
    6.57446e-06, 3.019876e-06, 5.647092e-06, 2.766084e-06, 2.471692e-06, 
    1.623629e-06, 2.684952e-06, 3.833956e-06, 5.954309e-06, 1.096426e-05,
  1.08422e-05, 9.811754e-06, 8.69002e-06, 7.216157e-06, 8.477713e-06, 
    5.832972e-06, 5.172179e-06, 3.571549e-06, 4.752748e-06, 4.182768e-06, 
    2.36918e-06, 5.371294e-06, 8.957847e-06, 8.674714e-06, 7.350945e-06,
  1.056118e-05, 1.357306e-05, 8.981868e-06, 6.820452e-06, 6.566554e-06, 
    7.648656e-06, 6.091221e-06, 3.138311e-06, 1.891637e-06, 1.945066e-06, 
    1.038205e-06, 3.31566e-06, 6.438522e-06, 6.898075e-06, 7.319912e-06,
  1.262708e-05, 1.084121e-05, 9.621635e-06, 9.397965e-06, 4.103131e-06, 
    5.887461e-06, 6.966299e-06, 1.194702e-06, 9.819204e-07, 4.607148e-07, 
    3.4039e-07, 5.962958e-07, 2.702923e-06, 6.573577e-06, 4.072483e-06,
  1.297883e-05, 1.421277e-05, 1.29099e-05, 1.066029e-05, 8.335091e-06, 
    5.417082e-06, 4.587363e-06, 9.064187e-07, 5.109603e-07, 1.83367e-08, 
    5.159284e-08, 9.82195e-08, 1.21705e-06, 6.394893e-06, 1.002513e-05,
  1.181062e-05, 1.537906e-05, 1.784454e-05, 1.554115e-05, 9.82544e-06, 
    5.729501e-06, 4.818977e-06, 9.676471e-07, 1.357272e-06, 1.686721e-08, 
    1.762592e-08, 6.06659e-08, 6.00885e-07, 7.992428e-06, 1.063575e-05,
  1.371703e-05, 1.677949e-05, 1.577001e-05, 1.415594e-05, 1.395509e-05, 
    7.441053e-06, 4.717311e-06, 3.54287e-06, 1.243755e-06, 2.531831e-07, 
    3.250335e-07, 1.40792e-07, 5.720424e-07, 1.302032e-05, 1.068428e-05,
  4.628378e-06, 4.784125e-06, 4.989231e-06, 6.609581e-06, 5.171783e-06, 
    6.923688e-06, 5.510551e-06, 4.380927e-06, 4.403457e-06, 4.819788e-06, 
    2.808537e-06, 1.108985e-06, 2.764482e-07, 2.562735e-06, 4.364833e-05,
  5.397096e-06, 5.846234e-06, 5.170921e-06, 5.689429e-06, 6.527906e-06, 
    5.169425e-06, 5.0413e-06, 6.085e-06, 4.187641e-06, 4.326445e-06, 
    3.750473e-06, 2.159132e-06, 1.925716e-06, 1.898941e-06, 7.330065e-06,
  5.443085e-06, 5.556545e-06, 5.619359e-06, 5.643271e-06, 6.547916e-06, 
    5.590109e-06, 5.550969e-06, 7.599121e-06, 5.287513e-06, 4.116539e-06, 
    3.608366e-06, 2.504637e-06, 1.749033e-06, 1.605958e-06, 5.627186e-07,
  6.010024e-06, 5.748625e-06, 7.009289e-06, 6.34323e-06, 6.91463e-06, 
    7.306523e-06, 6.810159e-06, 5.848821e-06, 7.765202e-06, 4.105332e-06, 
    2.807431e-06, 2.445091e-06, 1.000891e-06, 1.239511e-06, 1.384621e-07,
  6.338339e-06, 5.085798e-06, 5.283934e-06, 5.448921e-06, 6.308288e-06, 
    8.297273e-06, 7.852717e-06, 6.487575e-06, 9.235574e-06, 5.593913e-06, 
    2.658236e-06, 1.807664e-06, 7.275917e-07, 7.804748e-07, 3.179037e-07,
  7.299587e-06, 6.230675e-06, 3.559219e-06, 6.790188e-06, 8.964821e-06, 
    5.862359e-06, 8.899916e-06, 5.35254e-06, 3.679847e-06, 2.996286e-06, 
    1.734626e-06, 2.302245e-06, 2.975054e-07, 3.521378e-07, 6.448498e-08,
  5.353036e-06, 6.540095e-06, 7.540989e-06, 5.689124e-06, 6.926873e-06, 
    1.074801e-05, 1.270782e-05, 1.019345e-05, 7.510632e-06, 3.809471e-06, 
    1.225352e-06, 6.369941e-07, 2.318119e-07, 2.054547e-07, 4.192986e-07,
  5.84817e-06, 6.127718e-06, 6.275138e-06, 1.088308e-05, 1.095302e-05, 
    7.318723e-06, 8.424527e-06, 6.809429e-06, 6.933236e-06, 4.588409e-06, 
    1.415919e-06, 1.684968e-06, 2.647416e-07, 3.346739e-06, 6.063674e-06,
  6.099086e-06, 9.658112e-06, 1.153573e-05, 1.557071e-05, 1.202764e-05, 
    1.020278e-05, 8.423311e-06, 8.238617e-06, 6.127965e-06, 4.764776e-06, 
    2.758796e-06, 2.095972e-06, 6.257105e-07, 1.99979e-06, 7.641133e-06,
  9.399213e-06, 9.998735e-06, 1.301357e-05, 1.583473e-05, 1.237047e-05, 
    1.337198e-05, 9.187224e-06, 6.006352e-06, 5.810672e-06, 3.125757e-06, 
    2.068798e-06, 8.240622e-07, 7.923697e-07, 3.1334e-06, 8.665881e-06,
  5.283291e-06, 4.892528e-06, 4.591052e-06, 4.792329e-06, 4.572083e-06, 
    3.70949e-06, 4.959596e-06, 3.684028e-06, 2.31417e-06, 2.448809e-06, 
    8.635031e-07, 1.051546e-07, 5.342329e-07, 3.062992e-07, 1.748045e-06,
  5.991204e-06, 5.194846e-06, 4.569901e-06, 4.466877e-06, 4.580104e-06, 
    3.301423e-06, 3.981801e-06, 4.04349e-06, 3.224369e-06, 2.71764e-06, 
    1.52077e-06, 3.154406e-07, 3.718421e-07, 1.709301e-06, 1.081903e-06,
  4.833405e-06, 3.67923e-06, 4.246512e-06, 4.722688e-06, 4.602428e-06, 
    3.485491e-06, 2.978244e-06, 4.573497e-06, 4.137981e-06, 3.529507e-06, 
    2.374963e-06, 9.642665e-07, 1.211892e-06, 3.927054e-06, 1.176309e-06,
  5.039103e-06, 3.606375e-06, 3.730394e-06, 3.768587e-06, 4.01968e-06, 
    4.530687e-06, 3.079004e-06, 3.878203e-06, 4.270436e-06, 4.328437e-06, 
    4.381691e-06, 3.389129e-06, 2.43098e-06, 1.197123e-06, 6.226034e-07,
  5.050669e-06, 4.502052e-06, 5.189709e-06, 6.212175e-06, 5.635187e-06, 
    6.946229e-06, 6.545334e-06, 6.114566e-06, 4.856286e-06, 4.156776e-06, 
    3.425149e-06, 4.46454e-06, 1.115807e-06, 4.437887e-07, 3.678115e-08,
  6.577114e-06, 7.330362e-06, 5.888057e-06, 8.831233e-06, 7.923403e-06, 
    7.652438e-06, 6.784656e-06, 5.958146e-06, 4.853314e-06, 3.399758e-06, 
    3.006014e-06, 2.863493e-06, 1.78048e-06, 8.548371e-07, 1.010574e-08,
  8.057125e-06, 8.010608e-06, 5.8878e-06, 9.848835e-06, 8.812087e-06, 
    7.695957e-06, 7.615532e-06, 5.575494e-06, 6.337075e-06, 4.244726e-06, 
    2.104132e-06, 3.260069e-06, 1.741702e-07, 9.205126e-09, 7.317627e-07,
  6.790593e-06, 8.676989e-06, 1.255254e-05, 6.981651e-06, 1.094755e-05, 
    1.21071e-05, 1.034224e-05, 1.540203e-05, 9.613285e-06, 6.521312e-06, 
    3.811576e-06, 3.156159e-06, 5.630551e-06, 1.526679e-06, 1.003296e-07,
  7.933051e-06, 7.985552e-06, 1.080958e-05, 1.112879e-05, 1.112943e-05, 
    1.215152e-05, 1.292565e-05, 9.161708e-06, 7.306995e-06, 5.351644e-06, 
    5.292516e-06, 5.748396e-06, 7.729954e-06, 5.124009e-06, 1.546004e-06,
  1.004757e-05, 9.681102e-06, 1.224595e-05, 8.662506e-06, 1.078528e-05, 
    1.137174e-05, 1.201079e-05, 1.087936e-05, 1.001682e-05, 8.715248e-06, 
    7.536618e-06, 6.037018e-06, 7.705897e-06, 3.47401e-06, 3.70083e-06,
  5.394319e-06, 5.182296e-06, 4.130917e-06, 2.366319e-06, 1.921824e-06, 
    4.417479e-06, 4.05395e-06, 4.030646e-06, 3.608895e-06, 2.884521e-06, 
    2.326105e-06, 2.105886e-06, 2.804802e-06, 2.226028e-06, 5.848889e-07,
  6.290515e-06, 5.096071e-06, 3.490471e-06, 2.192881e-06, 1.960681e-06, 
    2.729972e-06, 6.054797e-06, 3.974951e-06, 2.805476e-06, 2.551852e-06, 
    2.726039e-06, 2.075803e-06, 2.220837e-06, 3.282067e-06, 5.901339e-07,
  6.680512e-06, 5.330629e-06, 4.392021e-06, 3.402858e-06, 4.197141e-06, 
    6.996575e-06, 7.224858e-06, 5.871565e-06, 3.811784e-06, 3.277819e-06, 
    2.105088e-06, 1.696717e-06, 2.028982e-06, 2.711279e-06, 2.311537e-06,
  7.582381e-06, 8.036909e-06, 5.966595e-06, 5.716044e-06, 7.423195e-06, 
    5.792903e-06, 6.673589e-06, 6.769759e-06, 6.448774e-06, 5.277817e-06, 
    3.35258e-06, 2.719582e-06, 1.467282e-06, 2.577154e-06, 2.068761e-06,
  8.665279e-06, 7.767502e-06, 7.795252e-06, 5.673523e-06, 5.63192e-06, 
    6.189886e-06, 8.999332e-06, 9.2254e-06, 7.1619e-06, 4.668128e-06, 
    4.087128e-06, 2.594825e-06, 1.765004e-06, 2.039785e-06, 1.74916e-06,
  8.189062e-06, 6.108364e-06, 5.491292e-06, 6.240322e-06, 6.151326e-06, 
    5.411354e-06, 5.744949e-06, 8.897993e-06, 1.08506e-05, 7.639559e-06, 
    3.58293e-06, 1.460597e-06, 1.527512e-06, 2.188624e-06, 1.143686e-06,
  4.495323e-06, 4.362599e-06, 3.717265e-06, 5.283952e-06, 7.422493e-06, 
    1.012187e-05, 5.951081e-06, 6.939034e-06, 6.678063e-06, 6.656313e-06, 
    4.127256e-06, 3.42084e-06, 2.21628e-06, 2.318012e-06, 1.267259e-06,
  5.926728e-06, 4.510982e-06, 4.030667e-06, 3.478799e-06, 4.092515e-06, 
    6.877428e-06, 1.024062e-05, 1.02836e-05, 8.985849e-06, 1.064635e-05, 
    8.634058e-06, 2.657597e-06, 2.144041e-06, 1.530599e-07, 1.347278e-06,
  5.428199e-06, 5.864516e-06, 6.807371e-06, 5.382786e-06, 5.305161e-06, 
    6.022439e-06, 7.357272e-06, 1.391881e-05, 1.446423e-05, 9.156038e-06, 
    1.144144e-05, 5.458645e-06, 3.135859e-06, 3.80579e-06, 2.898649e-06,
  8.190695e-06, 8.649097e-06, 6.55909e-06, 8.658032e-06, 9.653424e-06, 
    9.081823e-06, 4.551342e-06, 6.286783e-06, 1.09713e-05, 1.28188e-05, 
    8.664048e-06, 7.259478e-06, 3.544395e-06, 5.247228e-06, 4.754477e-06,
  5.055473e-06, 4.552486e-06, 4.490986e-06, 4.208358e-06, 2.836325e-06, 
    3.551217e-06, 4.046767e-06, 5.042861e-06, 2.357234e-06, 2.013742e-06, 
    1.662435e-06, 8.557407e-07, 2.923883e-06, 1.012975e-06, 4.905762e-07,
  3.507366e-06, 3.384893e-06, 3.666629e-06, 3.850754e-06, 2.336299e-06, 
    3.124652e-06, 5.475181e-06, 5.135414e-06, 3.460153e-06, 2.801786e-06, 
    1.698253e-06, 4.650366e-06, 4.061675e-06, 2.674031e-06, 9.661682e-07,
  2.975769e-06, 3.110783e-06, 3.547075e-06, 2.971554e-06, 3.126921e-06, 
    3.222998e-06, 4.088359e-06, 3.72596e-06, 2.439961e-06, 3.303026e-06, 
    3.672302e-06, 3.337859e-06, 4.297136e-06, 3.95663e-06, 3.684031e-06,
  5.009465e-06, 4.193422e-06, 3.155606e-06, 3.824886e-06, 3.983444e-06, 
    2.705291e-06, 2.02689e-06, 2.743211e-06, 3.03286e-06, 4.18894e-06, 
    3.423613e-06, 3.208063e-06, 6.045856e-06, 4.824753e-06, 1.657689e-06,
  4.936797e-06, 5.711332e-06, 3.7407e-06, 4.045417e-06, 5.007419e-06, 
    3.761824e-06, 2.620106e-06, 2.052773e-06, 2.994046e-06, 3.931353e-06, 
    3.345471e-06, 2.614736e-06, 4.500895e-06, 4.803582e-06, 1.324387e-06,
  6.994757e-06, 6.486896e-06, 3.470115e-06, 6.656053e-06, 4.514407e-06, 
    4.39194e-06, 3.029106e-06, 2.468707e-06, 2.218515e-06, 3.507503e-06, 
    2.963899e-06, 3.212885e-06, 2.767112e-06, 1.719237e-06, 7.963691e-07,
  7.866475e-06, 6.504145e-06, 5.642525e-06, 7.999955e-06, 7.378162e-06, 
    7.345947e-06, 5.106459e-06, 3.967276e-06, 2.369881e-06, 1.869608e-06, 
    2.447511e-06, 1.054639e-06, 7.902182e-07, 8.237601e-07, 5.941436e-07,
  8.274797e-06, 5.739358e-06, 8.696289e-06, 1.013788e-05, 8.333925e-06, 
    9.134483e-06, 7.386258e-06, 6.600966e-06, 3.10217e-06, 3.216192e-06, 
    1.125025e-06, 1.353782e-06, 1.848775e-06, 1.642448e-06, 6.187058e-07,
  6.258376e-06, 5.247871e-06, 7.042989e-06, 1.059463e-05, 1.46061e-05, 
    1.129505e-05, 7.506372e-06, 7.502165e-06, 5.02601e-06, 3.204512e-06, 
    6.692102e-07, 1.726392e-06, 5.247397e-06, 4.374579e-06, 3.544192e-07,
  4.969653e-06, 5.808364e-06, 7.461911e-06, 1.10697e-05, 1.144543e-05, 
    1.314724e-05, 1.003237e-05, 8.509266e-06, 9.084132e-06, 5.209886e-06, 
    5.731423e-06, 9.412187e-06, 9.950722e-06, 7.6593e-06, 1.852652e-06,
  6.340596e-06, 7.604877e-06, 7.178384e-06, 7.503903e-06, 1.199487e-05, 
    9.598699e-06, 8.673561e-06, 9.626345e-06, 8.962368e-06, 6.249147e-06, 
    5.039378e-06, 3.661938e-06, 2.592354e-06, 1.234074e-06, 1.406361e-07,
  7.295741e-06, 7.886959e-06, 7.042714e-06, 5.623397e-06, 4.877837e-06, 
    5.458437e-06, 4.025017e-06, 6.851456e-06, 3.459934e-06, 4.210695e-06, 
    2.561252e-06, 1.245073e-06, 1.486983e-06, 1.698353e-06, 7.542308e-07,
  5.971946e-06, 7.145562e-06, 6.85978e-06, 6.679971e-06, 5.827291e-06, 
    4.958254e-06, 5.091383e-06, 4.817013e-06, 3.933213e-06, 3.715848e-06, 
    2.666665e-06, 3.572203e-06, 1.759324e-06, 2.67581e-06, 9.195605e-07,
  6.443263e-06, 5.064738e-06, 7.579176e-06, 6.261682e-06, 5.007995e-06, 
    4.795557e-06, 4.952296e-06, 5.512079e-06, 3.83106e-06, 3.175147e-06, 
    2.502735e-06, 3.756197e-06, 1.811584e-06, 2.571406e-06, 2.684709e-06,
  5.511859e-06, 5.039886e-06, 3.804608e-06, 5.20272e-06, 4.983408e-06, 
    4.785907e-06, 5.101201e-06, 5.132801e-06, 4.416484e-06, 3.937597e-06, 
    2.909826e-06, 2.324216e-06, 3.570428e-06, 2.612684e-06, 3.155472e-07,
  5.516661e-06, 4.461867e-06, 3.823231e-06, 3.995909e-06, 5.066207e-06, 
    5.807046e-06, 4.026938e-06, 4.280492e-06, 3.789891e-06, 2.859853e-06, 
    2.96149e-06, 2.741023e-06, 2.024583e-06, 9.772228e-07, 5.707963e-06,
  5.186041e-06, 4.761081e-06, 4.613614e-06, 3.344337e-06, 3.76772e-06, 
    3.443624e-06, 2.973277e-06, 4.107331e-06, 4.094092e-06, 4.003155e-06, 
    3.616911e-06, 2.807e-06, 2.053599e-06, 2.040176e-06, 9.665096e-06,
  6.05888e-06, 5.940573e-06, 4.0108e-06, 1.827211e-06, 4.525081e-06, 
    5.731205e-06, 3.850219e-06, 3.717495e-06, 3.778636e-06, 2.822796e-06, 
    2.34596e-06, 2.421338e-06, 2.48458e-06, 1.037321e-06, 7.979454e-06,
  5.698686e-06, 5.016032e-06, 4.10073e-06, 2.566914e-06, 5.103071e-06, 
    5.316189e-06, 4.119371e-06, 4.028841e-06, 5.85354e-06, 3.378691e-06, 
    2.747282e-06, 2.647222e-06, 1.253278e-06, 3.296423e-06, 9.45276e-06,
  6.162472e-06, 4.583184e-06, 4.153943e-06, 5.720122e-06, 5.010805e-06, 
    4.178772e-06, 5.949509e-06, 6.574507e-06, 8.197935e-06, 1.023257e-05, 
    5.291953e-06, 3.669601e-06, 3.348383e-06, 8.29634e-06, 9.071423e-06,
  3.757969e-06, 8.318254e-06, 2.066544e-05, 6.140209e-05, 0.0001135573, 
    0.0001427636, 0.000172673, 0.0001677412, 0.000113554, 8.083438e-05, 
    6.756397e-05, 5.484123e-05, 3.493025e-05, 2.178456e-05, 1.467924e-05,
  3.142635e-06, 4.084324e-06, 5.265096e-06, 5.869922e-06, 6.192954e-06, 
    1.955332e-05, 2.929769e-05, 2.638966e-05, 2.247435e-05, 1.084831e-05, 
    2.100001e-06, 8.375109e-07, 1.212927e-06, 1.660135e-06, 4.080379e-06,
  3.215111e-06, 2.63172e-06, 2.619789e-06, 2.873217e-06, 3.668442e-06, 
    4.810827e-06, 7.137346e-06, 1.212167e-05, 8.79967e-06, 5.219661e-06, 
    5.27873e-07, 2.436037e-07, 1.291405e-07, 1.723232e-06, 4.872552e-07,
  3.911585e-06, 2.571393e-06, 2.025544e-06, 1.86485e-06, 1.591541e-06, 
    1.844825e-06, 2.188458e-06, 2.706259e-06, 2.906895e-06, 3.133451e-06, 
    9.923607e-07, 4.309678e-07, 1.586625e-07, 1.186419e-06, 2.076112e-07,
  4.068236e-06, 3.892393e-06, 2.837025e-06, 2.074926e-06, 2.287053e-06, 
    1.655538e-06, 9.939688e-07, 2.083872e-06, 1.386724e-06, 8.024094e-07, 
    9.092567e-07, 4.311754e-07, 1.921723e-07, 7.135977e-08, 4.089639e-08,
  4.854714e-06, 4.686781e-06, 4.478329e-06, 3.363265e-06, 3.235521e-06, 
    2.837381e-06, 1.59162e-06, 1.528801e-06, 1.576689e-06, 9.940416e-07, 
    7.907234e-07, 4.7512e-07, 3.622388e-07, 1.789095e-07, 1.406463e-08,
  4.602746e-06, 3.975896e-06, 3.366713e-06, 3.645016e-06, 3.392351e-06, 
    2.97536e-06, 2.714637e-06, 1.674005e-06, 1.030846e-06, 5.848142e-07, 
    1.668032e-07, 1.515247e-07, 1.623736e-08, 6.18102e-08, 5.28491e-08,
  5.015017e-06, 4.314334e-06, 3.879602e-06, 3.518616e-06, 3.346374e-06, 
    2.300498e-06, 1.814817e-06, 1.575121e-06, 1.566949e-06, 1.205531e-06, 
    6.55754e-07, 2.748192e-07, 1.116859e-07, 1.40939e-07, 1.673951e-06,
  4.282536e-06, 3.409521e-06, 3.903422e-06, 3.040758e-06, 2.912846e-06, 
    1.721609e-06, 1.420111e-06, 1.679515e-06, 1.483845e-06, 2.401677e-06, 
    8.244391e-07, 1.13529e-06, 9.337914e-07, 9.303975e-07, 1.208289e-06,
  5.264995e-06, 3.518102e-06, 1.856319e-06, 3.954432e-06, 2.793249e-06, 
    1.807796e-06, 1.635157e-06, 1.887337e-06, 2.391735e-06, 2.534832e-06, 
    2.115029e-06, 2.589562e-07, 2.099225e-06, 2.633181e-06, 4.702841e-06,
  8.14129e-07, 1.137343e-06, 3.37926e-06, 1.289913e-05, 5.544711e-05, 
    0.000176524, 0.0003310281, 0.0004166446, 0.000308799, 0.0001414815, 
    4.875374e-05, 2.060564e-05, 9.31222e-06, 5.620698e-06, 6.204568e-06,
  8.777685e-07, 1.146814e-06, 9.25419e-07, 3.244863e-06, 1.833953e-05, 
    7.998695e-05, 0.0001996684, 0.000299798, 0.0003058547, 0.0001853874, 
    7.068148e-05, 2.569175e-05, 9.495418e-06, 5.810967e-06, 6.217569e-06,
  1.626803e-06, 1.790686e-06, 2.0086e-06, 2.457705e-06, 4.735472e-06, 
    2.133163e-05, 6.451941e-05, 0.0001458862, 0.0002091007, 0.0001798052, 
    9.082047e-05, 3.284652e-05, 1.523554e-05, 1.037259e-05, 9.107719e-06,
  2.447707e-06, 2.569048e-06, 2.125356e-06, 1.597615e-06, 2.151944e-06, 
    3.364338e-06, 1.850818e-05, 5.523748e-05, 0.0001059023, 0.000119344, 
    8.39837e-05, 4.38475e-05, 2.14753e-05, 1.419257e-05, 1.121945e-05,
  2.708178e-06, 1.756637e-06, 1.059587e-06, 1.304234e-06, 2.093361e-06, 
    1.058571e-06, 1.069915e-06, 8.145952e-06, 3.412529e-05, 5.998062e-05, 
    6.555849e-05, 4.303183e-05, 1.981954e-05, 1.189209e-05, 9.387425e-06,
  2.474771e-06, 1.99122e-06, 1.200199e-06, 1.283129e-06, 1.580687e-06, 
    1.441704e-06, 8.095533e-07, 1.332866e-06, 4.317225e-06, 1.599257e-05, 
    3.079209e-05, 2.788654e-05, 1.40965e-05, 6.419472e-06, 4.893771e-06,
  3.897581e-06, 3.075229e-06, 1.892247e-06, 1.218647e-06, 8.81118e-07, 
    7.907958e-07, 8.360693e-07, 5.069822e-07, 7.341056e-07, 1.603217e-06, 
    7.792156e-06, 1.374977e-05, 1.146107e-05, 5.344975e-06, 3.268669e-06,
  4.701174e-06, 3.335242e-06, 2.004685e-06, 1.178433e-06, 1.100135e-06, 
    3.658655e-07, 1.231712e-06, 2.549808e-07, 1.931846e-07, 2.850211e-07, 
    2.568064e-07, 1.882815e-07, 1.618971e-06, 4.69235e-06, 6.081718e-06,
  5.064996e-06, 3.9346e-06, 2.387311e-06, 2.016197e-06, 2.179381e-06, 
    1.572909e-06, 1.669397e-06, 1.803342e-06, 1.967955e-06, 2.29603e-06, 
    1.609549e-06, 1.164494e-06, 4.989059e-07, 1.088258e-06, 7.474459e-06,
  5.695629e-06, 4.793463e-06, 3.372636e-06, 1.908238e-06, 2.104748e-06, 
    2.082782e-06, 1.097837e-06, 2.654774e-06, 5.262336e-06, 4.360955e-06, 
    2.481903e-06, 2.568718e-06, 5.183472e-06, 6.065917e-06, 6.771477e-06,
  1.301139e-06, 1.139128e-06, 1.105324e-06, 1.31152e-06, 4.227725e-08, 
    2.589393e-07, 1.178425e-06, 5.821654e-06, 6.300522e-06, 1.389296e-05, 
    1.153667e-05, 9.28669e-06, 8.081381e-06, 7.15936e-06, 8.403824e-06,
  3.041693e-06, 8.283237e-07, 1.905033e-06, 1.598158e-06, 3.341297e-07, 
    9.581716e-08, 3.013742e-06, 1.14141e-05, 1.826568e-05, 9.26339e-06, 
    3.233761e-06, 5.006046e-06, 5.88162e-06, 7.335733e-06, 1.535472e-05,
  2.326999e-06, 1.101187e-06, 1.464414e-06, 2.758973e-06, 3.214472e-06, 
    1.728771e-06, 1.296313e-05, 2.512644e-05, 4.87723e-05, 4.231504e-05, 
    8.432929e-06, 3.564641e-06, 4.740996e-06, 1.844697e-05, 2.36539e-05,
  1.648706e-06, 2.619132e-06, 9.930358e-07, 1.049697e-06, 1.799004e-06, 
    8.639987e-06, 2.334415e-05, 2.604408e-05, 4.406729e-05, 7.18247e-05, 
    4.311428e-05, 9.946468e-06, 1.100227e-05, 2.072901e-05, 2.040864e-05,
  1.56183e-06, 1.084278e-06, 8.569701e-07, 5.362144e-07, 6.616419e-07, 
    3.297023e-07, 4.159816e-06, 8.731844e-06, 2.817372e-05, 0.0001076521, 
    0.0001275941, 4.698642e-05, 1.654688e-05, 1.030867e-05, 1.260643e-05,
  2.476086e-06, 1.287959e-06, 1.068742e-06, 5.212059e-07, 5.463126e-07, 
    7.551946e-07, 5.782402e-07, 6.356215e-06, 4.13797e-05, 0.0001784676, 
    0.0002250899, 0.0001004913, 2.592733e-05, 1.169356e-05, 1.50309e-05,
  2.182763e-06, 2.311552e-06, 2.140984e-06, 1.243903e-06, 2.602563e-06, 
    2.111509e-06, 8.75232e-06, 2.054875e-05, 7.424705e-05, 0.0002204324, 
    0.0002710415, 0.0001541777, 5.079097e-05, 2.186686e-05, 2.038408e-05,
  5.051452e-06, 2.585778e-06, 5.257441e-06, 1.787349e-06, 1.917926e-06, 
    2.619405e-06, 1.904733e-05, 4.981293e-05, 0.0001039314, 0.0001843612, 
    0.0002280892, 0.0001514107, 6.146434e-05, 2.707184e-05, 2.170658e-05,
  6.46762e-06, 3.56068e-06, 2.947854e-06, 2.815161e-06, 2.11795e-06, 
    3.653094e-06, 8.129802e-06, 4.438464e-05, 9.909236e-05, 0.0001575373, 
    0.0001741225, 0.0001002988, 3.579048e-05, 1.639644e-05, 3.009543e-05,
  2.924787e-06, 3.109714e-06, 3.795913e-06, 3.670305e-06, 2.994452e-06, 
    6.785494e-06, 4.21114e-06, 1.568957e-05, 5.621775e-05, 0.0001158605, 
    0.0001280669, 7.546106e-05, 3.286076e-05, 2.572637e-05, 3.29131e-05,
  1.336813e-06, 8.715846e-07, 2.604096e-07, 9.742404e-07, 9.171661e-08, 
    1.439319e-07, 1.784609e-06, 1.200102e-05, 1.892041e-05, 1.078393e-05, 
    8.984642e-06, 9.070588e-06, 9.790396e-06, 1.203242e-05, 3.436734e-05,
  2.470378e-06, 1.717105e-06, 5.772532e-07, 1.244906e-06, 1.719258e-07, 
    3.621737e-07, 1.25667e-06, 7.974087e-06, 1.829079e-05, 1.608486e-05, 
    9.200653e-06, 9.950973e-06, 8.736293e-06, 1.127515e-05, 0.0001297733,
  2.716991e-06, 1.462657e-06, 9.35197e-07, 1.705614e-06, 2.745729e-07, 
    8.444089e-07, 2.423842e-06, 7.085297e-06, 1.42671e-05, 1.930417e-05, 
    1.295509e-05, 9.573847e-06, 7.288246e-06, 3.630307e-05, 0.0002249947,
  3.02386e-06, 3.28066e-06, 3.536743e-06, 2.126513e-06, 1.371586e-06, 
    1.201926e-06, 3.142279e-06, 8.480049e-06, 1.275099e-05, 1.782976e-05, 
    1.490867e-05, 1.231819e-05, 1.939413e-05, 0.0001441898, 0.0002724302,
  2.792262e-06, 2.910906e-06, 1.031809e-06, 2.550423e-06, 1.545213e-06, 
    9.47654e-07, 3.569335e-06, 1.058963e-05, 1.191006e-05, 1.594087e-05, 
    1.890929e-05, 2.341635e-05, 8.120008e-05, 0.0002049093, 0.0002344454,
  3.704188e-06, 2.635354e-06, 2.06011e-06, 2.738629e-06, 8.798782e-07, 
    4.939339e-07, 3.139125e-06, 9.083355e-06, 1.472963e-05, 1.649743e-05, 
    2.858119e-05, 5.473247e-05, 0.0001447191, 0.0001794835, 9.479815e-05,
  3.578928e-06, 1.908798e-06, 3.722493e-06, 2.309593e-06, 1.824491e-06, 
    2.335272e-07, 4.073712e-06, 1.078163e-05, 1.824219e-05, 3.195188e-05, 
    5.124075e-05, 0.0001112085, 0.0001279737, 8.365248e-05, 4.603174e-05,
  2.148627e-06, 1.413282e-06, 3.983668e-06, 2.848393e-06, 1.738905e-06, 
    2.626413e-06, 1.111739e-05, 2.015155e-05, 3.176915e-05, 4.941793e-05, 
    0.0001028676, 0.0001332192, 9.330759e-05, 4.709461e-05, 5.33749e-05,
  2.044055e-06, 1.225506e-06, 2.457542e-06, 3.98108e-06, 3.110245e-06, 
    2.118825e-06, 1.018436e-05, 2.465888e-05, 4.684542e-05, 9.455522e-05, 
    0.0001179097, 0.0001048377, 6.865554e-05, 5.402719e-05, 2.878559e-05,
  3.407488e-06, 3.52066e-06, 3.565723e-06, 7.149124e-06, 4.193437e-06, 
    7.522697e-06, 1.209939e-05, 4.252984e-05, 9.566132e-05, 0.0001194062, 
    0.0001039419, 7.560366e-05, 5.985152e-05, 3.00947e-05, 1.562389e-05,
  4.932751e-06, 5.356095e-06, 7.050798e-06, 7.400702e-06, 9.631927e-06, 
    1.543592e-05, 1.592352e-05, 1.154099e-05, 8.459259e-06, 9.56359e-06, 
    7.416357e-06, 4.600296e-06, 2.503515e-06, 2.660371e-06, 3.130765e-06,
  5.078013e-06, 7.60762e-06, 8.063977e-06, 8.941843e-06, 1.059762e-05, 
    1.674233e-05, 1.536546e-05, 1.239947e-05, 8.550832e-06, 7.291081e-06, 
    4.132209e-06, 2.727699e-06, 2.329794e-06, 2.234447e-06, 4.078444e-06,
  7.644109e-06, 7.569374e-06, 6.708917e-06, 8.604869e-06, 1.148622e-05, 
    1.865478e-05, 1.63695e-05, 1.021838e-05, 7.417724e-06, 5.344658e-06, 
    5.979578e-06, 3.998181e-06, 4.168392e-06, 4.577838e-06, 5.614511e-06,
  1.068871e-05, 9.968435e-06, 8.251061e-06, 1.0867e-05, 1.531615e-05, 
    1.983856e-05, 1.807461e-05, 1.143526e-05, 5.823978e-06, 7.422956e-06, 
    6.034597e-06, 5.318515e-06, 6.212378e-06, 5.876279e-06, 6.329307e-06,
  1.493381e-05, 1.413041e-05, 1.306357e-05, 1.296025e-05, 1.816317e-05, 
    1.841239e-05, 1.362201e-05, 8.886002e-06, 6.331137e-06, 6.93789e-06, 
    6.486851e-06, 5.587073e-06, 5.224991e-06, 3.910413e-06, 4.572439e-06,
  1.965426e-05, 1.693237e-05, 1.416282e-05, 1.279371e-05, 1.484702e-05, 
    1.543072e-05, 1.29847e-05, 7.428955e-06, 7.425027e-06, 8.404851e-06, 
    6.307137e-06, 3.124204e-06, 3.548153e-06, 3.782768e-06, 3.916481e-06,
  2.50659e-05, 2.162715e-05, 1.680163e-05, 1.22395e-05, 1.286488e-05, 
    1.201254e-05, 9.908052e-06, 8.519974e-06, 1.297207e-05, 1.067227e-05, 
    4.364314e-06, 3.025732e-06, 3.597205e-06, 3.540446e-06, 3.575679e-06,
  2.880427e-05, 2.302106e-05, 1.488929e-05, 1.019296e-05, 1.239107e-05, 
    1.096419e-05, 1.097912e-05, 1.663636e-05, 2.185723e-05, 1.255512e-05, 
    4.799356e-06, 3.459245e-06, 2.60406e-06, 3.125995e-06, 5.016161e-06,
  3.097488e-05, 2.247655e-05, 1.542766e-05, 1.173902e-05, 1.106371e-05, 
    1.676519e-05, 2.217793e-05, 2.668494e-05, 2.068134e-05, 9.082823e-06, 
    4.493847e-06, 3.585586e-06, 2.658488e-06, 4.076769e-06, 5.20754e-06,
  3.578899e-05, 2.268568e-05, 2.085316e-05, 2.360883e-05, 2.660431e-05, 
    3.358733e-05, 3.8501e-05, 3.198432e-05, 1.537062e-05, 5.474118e-06, 
    3.650016e-06, 2.834608e-06, 2.197139e-06, 8.294611e-07, 1.195617e-06,
  5.397183e-06, 4.912785e-06, 4.031062e-06, 5.357857e-06, 8.929952e-06, 
    6.871896e-06, 7.174854e-06, 7.343935e-06, 6.409868e-06, 6.212642e-06, 
    5.048547e-06, 4.012961e-06, 5.504124e-06, 9.692625e-06, 1.383936e-05,
  5.294374e-06, 4.336501e-06, 3.977595e-06, 9.535672e-06, 9.714549e-06, 
    8.455399e-06, 7.905953e-06, 7.879449e-06, 7.41135e-06, 6.032348e-06, 
    5.77482e-06, 4.86373e-06, 4.674534e-06, 4.864608e-06, 9.454165e-06,
  3.901808e-06, 5.572741e-06, 5.569929e-06, 8.598478e-06, 1.01272e-05, 
    7.066928e-06, 6.060787e-06, 8.864807e-06, 6.203653e-06, 5.312513e-06, 
    7.077374e-06, 4.356688e-06, 3.824355e-06, 3.628047e-06, 5.292967e-06,
  4.82559e-06, 6.208754e-06, 6.577061e-06, 5.731958e-06, 6.50534e-06, 
    6.632185e-06, 5.675836e-06, 5.976487e-06, 8.017936e-06, 8.506182e-06, 
    6.824803e-06, 4.074614e-06, 2.184322e-06, 2.963242e-06, 3.735556e-06,
  3.914332e-06, 3.067005e-06, 4.274447e-06, 3.982398e-06, 4.242026e-06, 
    4.078659e-06, 5.179067e-06, 4.422096e-06, 7.211509e-06, 8.000563e-06, 
    8.586258e-06, 8.148412e-06, 5.995295e-06, 3.312898e-06, 3.657572e-06,
  3.843347e-06, 3.289049e-06, 4.323099e-06, 3.488836e-06, 3.333413e-06, 
    4.364553e-06, 5.412425e-06, 5.461401e-06, 4.04186e-06, 6.635742e-06, 
    6.785522e-06, 7.823286e-06, 7.317152e-06, 7.588607e-06, 4.129163e-06,
  5.50616e-06, 6.591405e-06, 5.057056e-06, 6.122294e-06, 5.11448e-06, 
    5.105408e-06, 5.480908e-06, 6.143449e-06, 4.799278e-06, 4.652525e-06, 
    5.824738e-06, 6.531147e-06, 4.62041e-06, 4.007697e-06, 5.666145e-06,
  6.495744e-06, 6.243776e-06, 6.228244e-06, 7.582955e-06, 6.504701e-06, 
    8.294465e-06, 8.151737e-06, 7.800603e-06, 6.462521e-06, 5.757201e-06, 
    5.312344e-06, 4.523589e-06, 3.661228e-06, 5.723187e-06, 5.797177e-06,
  6.078788e-06, 6.823094e-06, 8.16285e-06, 9.214776e-06, 1.028356e-05, 
    1.016372e-05, 1.016432e-05, 7.568841e-06, 7.751612e-06, 9.141615e-06, 
    8.106192e-06, 7.44267e-06, 6.634973e-06, 8.089057e-06, 7.5076e-06,
  7.235495e-06, 8.788765e-06, 9.259148e-06, 1.163662e-05, 1.166326e-05, 
    1.180599e-05, 1.02039e-05, 1.020102e-05, 9.811612e-06, 1.080431e-05, 
    1.00256e-05, 8.049138e-06, 8.545075e-06, 8.37147e-06, 8.942753e-06,
  6.277444e-06, 4.479393e-06, 4.149152e-06, 3.621337e-06, 3.345631e-06, 
    4.255173e-06, 1.007205e-05, 9.112038e-06, 6.35732e-06, 5.071292e-06, 
    4.544816e-06, 5.989966e-06, 6.917442e-06, 5.494191e-06, 4.427735e-06,
  7.381715e-06, 5.392723e-06, 4.114717e-06, 5.776874e-06, 3.358069e-06, 
    4.372761e-06, 7.113338e-06, 8.63323e-06, 6.739488e-06, 7.414895e-06, 
    2.693091e-06, 4.592107e-06, 5.858922e-06, 7.950175e-06, 7.067658e-06,
  7.93724e-06, 6.960901e-06, 7.676857e-06, 2.120074e-06, 1.208833e-06, 
    1.732412e-06, 2.021483e-06, 5.384522e-06, 7.238546e-06, 4.968254e-06, 
    2.969004e-06, 3.093739e-06, 3.919685e-06, 6.523014e-06, 6.374348e-06,
  8.716429e-06, 7.933347e-06, 6.482469e-06, 5.493035e-06, 3.586635e-06, 
    2.123634e-06, 1.511635e-06, 3.633706e-06, 2.190483e-06, 6.527856e-06, 
    5.488405e-06, 1.358952e-06, 3.470086e-06, 7.187041e-06, 5.527305e-06,
  6.269517e-06, 6.487353e-06, 4.509758e-06, 6.016236e-06, 5.834923e-06, 
    4.840354e-06, 2.764961e-06, 3.334349e-06, 5.288547e-06, 5.490031e-06, 
    2.828297e-06, 3.175451e-06, 4.767312e-06, 5.72374e-06, 7.242991e-06,
  6.103585e-06, 5.916999e-06, 6.287269e-06, 5.677739e-06, 4.965809e-06, 
    3.14025e-06, 4.786432e-06, 2.034385e-06, 2.22397e-06, 4.739948e-06, 
    2.203407e-06, 2.11553e-06, 5.900159e-06, 6.230982e-06, 1.129931e-05,
  5.57767e-06, 7.025623e-06, 5.961108e-06, 4.559082e-06, 4.490701e-06, 
    4.378055e-06, 4.459768e-06, 3.514025e-06, 2.381063e-06, 2.071606e-06, 
    3.493885e-06, 2.132596e-06, 4.063143e-06, 9.933214e-06, 1.290417e-05,
  4.71691e-06, 4.523393e-06, 3.945644e-06, 3.668545e-06, 2.871021e-06, 
    3.549106e-06, 3.820001e-06, 4.978622e-06, 3.693021e-06, 2.890438e-06, 
    3.590752e-06, 1.903723e-06, 5.374127e-06, 1.030902e-05, 1.871245e-05,
  4.027152e-06, 2.92165e-06, 2.697495e-06, 2.643181e-06, 1.916301e-06, 
    2.663239e-06, 2.607135e-06, 4.147885e-06, 4.548383e-06, 4.224802e-06, 
    3.622383e-06, 3.295008e-06, 7.62809e-06, 1.295653e-05, 1.637305e-05,
  3.715319e-06, 2.63417e-06, 2.68064e-06, 2.273985e-06, 2.360846e-06, 
    2.390687e-06, 2.203437e-06, 2.484979e-06, 4.004684e-06, 5.029171e-06, 
    4.25048e-06, 5.003851e-06, 1.178257e-05, 1.272563e-05, 1.682589e-05,
  3.126151e-06, 1.790514e-06, 4.770513e-06, 2.325812e-06, 2.393514e-06, 
    2.830807e-06, 4.577464e-06, 6.753207e-06, 6.768473e-06, 8.819693e-06, 
    4.68816e-06, 2.300202e-06, 6.689223e-07, 2.820793e-06, 7.379384e-06,
  2.119411e-06, 1.211104e-06, 1.711505e-06, 4.39196e-06, 1.272351e-06, 
    1.778654e-06, 4.10201e-06, 5.652843e-06, 7.36044e-06, 6.8631e-06, 
    4.533411e-06, 1.114908e-06, 8.581123e-07, 2.917707e-06, 9.627121e-06,
  3.332297e-06, 1.810386e-06, 1.750119e-06, 3.227914e-06, 3.517886e-06, 
    2.521416e-06, 3.223802e-06, 3.209584e-06, 4.293994e-06, 2.796551e-06, 
    3.752381e-06, 2.996948e-06, 3.978556e-07, 2.479409e-06, 8.12759e-06,
  4.491837e-06, 2.602496e-06, 2.528133e-06, 1.687716e-06, 2.905388e-06, 
    1.22387e-06, 1.289641e-06, 4.74825e-06, 2.303315e-06, 2.07731e-06, 
    1.571725e-06, 2.391325e-06, 2.594046e-06, 4.699217e-06, 1.874603e-05,
  5.649004e-06, 8.261787e-06, 2.685216e-06, 2.472293e-06, 3.051512e-06, 
    1.867182e-06, 1.318761e-07, 1.698297e-06, 4.180131e-06, 4.097773e-06, 
    1.542292e-06, 2.878438e-06, 4.212268e-06, 1.032405e-05, 4.831175e-05,
  4.492536e-06, 7.595436e-06, 5.046623e-06, 2.244935e-06, 2.632288e-06, 
    1.704724e-06, 8.719787e-07, 1.449994e-06, 3.659729e-06, 2.202955e-06, 
    1.271341e-06, 3.235465e-06, 5.632629e-06, 2.380404e-05, 8.20642e-05,
  5.128805e-06, 8.090575e-06, 4.916404e-06, 2.230468e-06, 1.601855e-06, 
    4.570901e-06, 2.045152e-07, 8.490886e-07, 3.713823e-06, 1.13303e-06, 
    2.051856e-06, 5.641153e-06, 1.242016e-05, 2.550529e-05, 8.711204e-05,
  4.583392e-06, 4.065676e-06, 4.627642e-06, 2.419873e-06, 1.903692e-06, 
    1.937765e-06, 3.081524e-07, 1.787406e-06, 1.028833e-06, 1.313445e-06, 
    3.874997e-06, 7.400025e-06, 1.412379e-05, 2.780363e-05, 6.946986e-05,
  5.02186e-06, 3.717749e-06, 3.78236e-06, 1.510579e-06, 5.965375e-06, 
    2.63748e-06, 2.635545e-06, 1.479398e-06, 1.961073e-07, 1.585968e-06, 
    3.758333e-06, 7.150031e-06, 1.575754e-05, 2.546789e-05, 4.441644e-05,
  3.30834e-06, 3.286257e-06, 4.060163e-06, 3.197119e-06, 5.674342e-06, 
    5.798255e-06, 2.011867e-06, 7.423723e-07, 2.178426e-07, 2.535745e-06, 
    6.762657e-06, 7.832582e-06, 1.168086e-05, 1.83101e-05, 2.807333e-05,
  2.849006e-06, 1.835946e-06, 4.751822e-06, 2.447384e-06, 3.537008e-06, 
    3.076037e-06, 4.185954e-06, 3.823122e-06, 1.475093e-06, 3.112192e-06, 
    1.163865e-05, 1.772733e-05, 1.923911e-05, 1.8146e-05, 2.125359e-05,
  4.182927e-06, 5.675977e-06, 5.239897e-06, 5.311453e-06, 3.90839e-06, 
    2.017856e-06, 1.129563e-06, 3.172401e-06, 2.158351e-06, 3.973839e-06, 
    8.560005e-06, 1.426914e-05, 1.827824e-05, 2.038278e-05, 2.72042e-05,
  3.850688e-06, 4.671223e-06, 3.258943e-06, 3.370054e-06, 6.041745e-06, 
    2.644789e-06, 2.554782e-06, 1.671638e-06, 2.694278e-06, 4.639102e-06, 
    6.877096e-06, 9.435591e-06, 1.474229e-05, 2.015345e-05, 2.69274e-05,
  5.380193e-06, 2.8774e-06, 4.099964e-06, 4.645184e-06, 5.571377e-06, 
    3.768311e-06, 3.920162e-06, 3.925787e-06, 2.159148e-06, 4.55338e-06, 
    7.065829e-06, 8.627037e-06, 1.504063e-05, 2.057517e-05, 2.74988e-05,
  4.565594e-06, 3.386815e-06, 4.537437e-06, 4.629459e-06, 4.469007e-06, 
    4.521517e-06, 2.766892e-06, 3.453026e-06, 2.022787e-06, 4.660888e-06, 
    6.650319e-06, 8.897965e-06, 1.564257e-05, 2.413346e-05, 3.214718e-05,
  6.190326e-06, 4.047091e-06, 3.109417e-06, 5.086304e-06, 6.391391e-06, 
    6.864818e-06, 3.342098e-06, 3.194894e-06, 1.687666e-06, 4.667672e-06, 
    4.867226e-06, 8.612073e-06, 1.580717e-05, 2.571321e-05, 3.686187e-05,
  4.436195e-06, 3.586854e-06, 6.728587e-06, 7.055386e-06, 9.209145e-06, 
    6.714627e-06, 3.137504e-06, 7.306521e-07, 1.829263e-06, 2.23877e-06, 
    4.119514e-06, 7.917509e-06, 1.797752e-05, 3.06898e-05, 4.828957e-05,
  4.501324e-06, 6.481631e-06, 7.705075e-06, 6.059658e-06, 9.694784e-06, 
    6.326884e-06, 2.923236e-06, 2.22224e-06, 3.541764e-07, 1.33909e-06, 
    4.467128e-06, 9.996239e-06, 2.099058e-05, 3.764874e-05, 6.356509e-05,
  4.850163e-06, 6.20923e-06, 8.206264e-06, 8.964392e-06, 1.075149e-05, 
    5.852587e-06, 2.635527e-06, 1.547453e-06, 1.20077e-07, 7.732284e-07, 
    3.816213e-06, 1.355722e-05, 2.228992e-05, 4.082466e-05, 7.9825e-05,
  4.764051e-06, 6.648581e-06, 9.698349e-06, 7.886964e-06, 1.20094e-05, 
    6.693802e-06, 1.918634e-06, 8.334784e-07, 1.538056e-08, 5.947294e-07, 
    4.923489e-06, 1.481724e-05, 2.504072e-05, 5.213098e-05, 9.695601e-05,
  1.867191e-06, 2.372631e-06, 2.348356e-06, 2.204858e-06, 1.658866e-06, 
    1.299163e-06, 2.028099e-07, 2.832177e-06, 2.085194e-05, 7.060624e-05, 
    0.0001011392, 0.0002026467, 0.0002197794, 6.764618e-05, 5.668566e-06,
  1.965924e-06, 2.618973e-06, 1.900842e-06, 1.481724e-06, 7.041614e-07, 
    1.928377e-07, 5.024923e-08, 7.703094e-06, 6.921624e-05, 0.0001016779, 
    8.667591e-05, 0.0001312411, 0.0001300169, 2.791455e-05, 1.769378e-05,
  1.83394e-06, 2.516513e-06, 2.313569e-06, 2.173223e-06, 3.838746e-07, 
    2.163318e-08, 1.505789e-06, 2.735451e-05, 0.0001024742, 9.144595e-05, 
    2.735052e-05, 2.972143e-05, 4.624832e-05, 1.816197e-05, 2.308984e-05,
  1.708094e-06, 1.816756e-06, 2.181549e-06, 1.774878e-06, 2.161424e-07, 
    8.062928e-08, 8.553922e-06, 6.319873e-05, 9.235308e-05, 3.679071e-05, 
    2.758378e-06, 1.013034e-05, 1.957721e-05, 1.470187e-05, 2.28008e-05,
  1.634166e-06, 2.77907e-06, 1.709214e-06, 1.014879e-06, 4.744945e-07, 
    8.572136e-07, 2.509158e-05, 6.724603e-05, 4.994435e-05, 1.35554e-05, 
    4.340342e-06, 7.220643e-06, 9.059853e-06, 9.401061e-06, 8.443372e-06,
  2.731663e-06, 2.719147e-06, 3.491527e-06, 1.254124e-06, 3.224056e-07, 
    3.628672e-06, 3.384128e-05, 4.682425e-05, 2.75e-05, 1.120099e-05, 
    6.052488e-06, 7.064566e-06, 5.467947e-06, 2.582002e-06, 1.617381e-06,
  3.833663e-06, 3.177462e-06, 2.859589e-06, 1.074325e-06, 2.182303e-07, 
    6.284156e-06, 2.939687e-05, 2.899138e-05, 1.847387e-05, 1.178707e-05, 
    7.671393e-06, 6.433005e-06, 4.887176e-06, 3.505484e-06, 3.138155e-06,
  4.408728e-06, 3.869396e-06, 2.926452e-06, 6.913785e-07, 4.76109e-07, 
    9.468431e-06, 2.305316e-05, 1.837975e-05, 1.496375e-05, 1.278451e-05, 
    8.53837e-06, 6.541447e-06, 5.48006e-06, 3.966607e-06, 3.334087e-06,
  3.100759e-06, 3.366159e-06, 2.001083e-06, 8.841861e-07, 1.144865e-06, 
    1.09724e-05, 2.04106e-05, 1.244148e-05, 1.610557e-05, 1.659063e-05, 
    1.083484e-05, 7.489265e-06, 5.505721e-06, 3.428177e-06, 2.208585e-06,
  4.314174e-06, 2.334621e-06, 1.915306e-06, 1.019106e-06, 1.398287e-06, 
    1.119621e-05, 1.73736e-05, 1.066774e-05, 1.531207e-05, 1.78037e-05, 
    1.287169e-05, 7.23588e-06, 3.998293e-06, 1.886329e-06, 4.228079e-06,
  2.708383e-06, 2.3263e-06, 3.586605e-06, 4.587504e-06, 4.792908e-06, 
    4.873194e-06, 3.792688e-06, 4.894745e-06, 3.8255e-06, 3.15958e-06, 
    6.208024e-07, 1.085104e-05, 0.0001179111, 0.000356948, 0.0003985082,
  2.592415e-06, 3.884506e-06, 2.866483e-06, 2.856677e-06, 2.590842e-06, 
    3.536406e-06, 3.320686e-06, 4.157755e-06, 1.659905e-06, 1.786443e-06, 
    3.089817e-06, 5.598697e-05, 0.0001979083, 0.0004176081, 0.0003964804,
  2.137473e-06, 2.654335e-06, 2.779421e-06, 2.216401e-06, 2.334302e-06, 
    2.374227e-06, 2.683843e-06, 1.63042e-06, 9.465925e-07, 7.92346e-06, 
    2.878181e-05, 0.000101713, 0.0002256569, 0.0003172551, 0.0003323689,
  2.166599e-06, 2.755112e-06, 2.529483e-06, 1.808091e-06, 8.833453e-07, 
    1.346198e-06, 2.501559e-06, 4.83044e-06, 1.340642e-05, 3.500134e-05, 
    4.784652e-05, 0.0001158844, 0.0002174457, 0.0002390638, 0.0003288128,
  2.291949e-06, 2.42955e-06, 2.067126e-06, 1.264467e-06, 6.449566e-07, 
    2.251112e-06, 1.222309e-05, 1.497163e-05, 2.501549e-05, 5.148953e-05, 
    7.314288e-05, 0.0001310142, 0.0001863566, 0.0002025935, 0.0003304123,
  2.229616e-06, 2.00121e-06, 1.193669e-06, 6.048525e-07, 1.172839e-06, 
    9.152341e-06, 2.280752e-05, 1.736883e-05, 3.403731e-05, 5.033414e-05, 
    6.148216e-05, 0.0001149374, 0.0001537389, 0.0001725457, 0.0003057341,
  1.385831e-06, 3.457845e-06, 1.701028e-06, 1.534242e-06, 1.016519e-06, 
    1.752087e-05, 2.551903e-05, 2.508664e-05, 2.453758e-05, 3.356662e-05, 
    5.75377e-05, 9.824238e-05, 0.0001268016, 0.0001387644, 0.0002470277,
  1.081722e-06, 2.84034e-06, 1.21396e-06, 1.249814e-06, 3.054878e-06, 
    2.043559e-05, 3.210022e-05, 2.399591e-05, 2.060911e-05, 3.069455e-05, 
    5.900471e-05, 9.464595e-05, 0.0001109428, 0.0001155785, 0.0002030497,
  4.480527e-06, 2.753903e-06, 1.256831e-06, 5.515903e-07, 7.425426e-06, 
    2.607179e-05, 2.103493e-05, 2.098691e-05, 1.704182e-05, 2.111801e-05, 
    4.31377e-05, 7.803223e-05, 8.229194e-05, 9.829232e-05, 0.0001727749,
  3.738551e-06, 1.276761e-06, 7.533874e-07, 1.66256e-06, 1.410822e-05, 
    3.01765e-05, 1.941999e-05, 1.288543e-05, 6.721195e-06, 1.037296e-05, 
    2.299691e-05, 5.201868e-05, 6.178694e-05, 8.990587e-05, 0.0001395773,
  6.830382e-05, 9.570626e-05, 9.19364e-05, 2.278592e-05, 8.058489e-07, 
    8.272722e-07, 1.546019e-06, 2.399017e-06, 7.50335e-07, 1.345406e-05, 
    3.642172e-05, 6.542735e-05, 6.406641e-05, 3.710245e-05, 8.114842e-06,
  5.033768e-05, 9.504068e-05, 0.0001163304, 9.510687e-05, 2.805663e-06, 
    1.104842e-06, 1.133435e-06, 1.100416e-06, 1.820711e-06, 2.535953e-05, 
    6.638156e-05, 0.0001728662, 0.0001155732, 7.345498e-05, 3.083841e-05,
  2.084745e-05, 7.520935e-05, 0.0001194797, 0.0001242393, 6.491613e-05, 
    2.662439e-06, 1.273138e-06, 3.611818e-07, 2.647965e-07, 2.232096e-05, 
    6.034732e-05, 0.0001107924, 0.0001190484, 0.0001030406, 5.591054e-05,
  7.746262e-06, 5.032555e-05, 0.0001061245, 0.0001200051, 0.0001199415, 
    6.246646e-06, 1.995366e-07, 5.469709e-07, 9.558603e-08, 1.756118e-05, 
    5.163056e-05, 0.0001004433, 0.0001151757, 0.000124336, 8.770089e-05,
  2.621174e-06, 2.776567e-05, 7.811013e-05, 0.0001059095, 0.0001375601, 
    8.731354e-05, 1.863031e-07, 3.80121e-07, 3.017096e-08, 1.480588e-05, 
    4.589702e-05, 9.564021e-05, 0.000119458, 0.0001449849, 0.0001195442,
  2.320097e-06, 1.24172e-05, 4.260514e-05, 7.295628e-05, 0.0001269664, 
    0.0001364577, 2.076597e-06, 2.262944e-07, 2.022117e-07, 9.633538e-06, 
    3.97785e-05, 9.548135e-05, 0.0001259159, 0.0001707502, 0.0001544536,
  2.362513e-06, 2.234157e-06, 1.124595e-05, 2.762759e-05, 8.433302e-05, 
    0.000153081, 6.23975e-05, 6.537952e-07, 2.253028e-07, 3.622817e-06, 
    3.059035e-05, 9.405217e-05, 0.0001356531, 0.0001881054, 0.0001824914,
  2.482917e-06, 3.122911e-06, 3.098965e-06, 4.561076e-06, 2.986822e-05, 
    0.0001371511, 0.0001365236, 3.456597e-06, 3.797691e-07, 9.543224e-07, 
    2.346586e-05, 9.266637e-05, 0.0001453568, 0.0002044458, 0.0001829152,
  4.579042e-06, 4.21391e-06, 2.751576e-06, 2.044514e-06, 3.028787e-06, 
    0.0001066983, 0.000154362, 1.492944e-05, 5.945907e-07, 5.103876e-07, 
    1.787096e-05, 8.759086e-05, 0.0001450491, 0.0002105929, 0.0001828881,
  5.5218e-06, 5.31326e-06, 4.261129e-06, 9.581634e-07, 1.866488e-06, 
    6.458742e-05, 0.0001704581, 8.294026e-05, 2.555063e-06, 1.659234e-06, 
    1.50156e-05, 7.936193e-05, 0.0001350859, 0.0002119248, 0.000190417,
  3.490453e-05, 2.808589e-05, 1.377489e-05, 1.662585e-07, 4.326758e-07, 
    1.173836e-05, 5.821109e-05, 7.809672e-05, 4.086164e-05, 4.417353e-06, 
    2.598619e-06, 1.51098e-06, 2.021291e-06, 2.139482e-06, 4.233477e-06,
  3.314891e-05, 3.644521e-05, 3.247407e-05, 1.40112e-05, 5.86593e-07, 
    8.894875e-06, 5.155016e-05, 5.596244e-05, 8.445792e-06, 3.241888e-06, 
    2.658812e-06, 8.615645e-07, 2.113559e-06, 2.389349e-06, 3.251474e-06,
  2.588578e-05, 4.230079e-05, 4.125997e-05, 3.596692e-05, 7.463177e-06, 
    2.172161e-06, 2.413849e-05, 2.24743e-05, 5.598518e-06, 3.632457e-06, 
    3.912188e-06, 1.039582e-06, 2.677276e-06, 2.308228e-06, 4.674937e-06,
  1.041702e-05, 3.26175e-05, 5.158425e-05, 4.583557e-05, 3.748823e-05, 
    2.741606e-06, 1.67582e-05, 1.100669e-05, 3.779078e-06, 3.864015e-06, 
    5.909972e-06, 1.578052e-06, 3.493504e-06, 3.315875e-06, 6.332009e-06,
  6.28853e-06, 2.216011e-05, 6.297773e-05, 5.140822e-05, 6.583422e-05, 
    2.234842e-05, 6.028389e-06, 1.135218e-05, 2.056615e-06, 5.765984e-06, 
    8.447199e-06, 3.121474e-06, 4.412854e-06, 5.354006e-06, 7.672538e-06,
  7.136746e-06, 1.699298e-05, 6.499349e-05, 5.964808e-05, 8.663539e-05, 
    6.477466e-05, 1.686802e-06, 7.254667e-06, 3.015656e-06, 9.398158e-06, 
    9.236756e-06, 4.546595e-06, 3.854136e-06, 6.88648e-06, 1.003738e-05,
  7.807925e-06, 1.053176e-05, 6.374725e-05, 7.925733e-05, 9.303019e-05, 
    0.0001167551, 1.896091e-05, 8.27751e-06, 2.790475e-06, 9.400431e-06, 
    1.056833e-05, 6.569275e-06, 4.942637e-06, 8.353302e-06, 1.288867e-05,
  8.573498e-06, 1.039909e-05, 6.123788e-05, 0.0001032505, 9.786487e-05, 
    0.0001490337, 7.570886e-05, 2.63818e-06, 3.505713e-06, 1.053051e-05, 
    1.029042e-05, 7.498384e-06, 6.46955e-06, 8.891087e-06, 1.89414e-05,
  1.021855e-05, 1.067783e-05, 5.298042e-05, 0.0001232923, 0.0001060041, 
    0.0001661998, 0.0001459784, 3.499629e-06, 2.567477e-06, 9.094958e-06, 
    1.008391e-05, 1.099765e-05, 8.761413e-06, 1.074601e-05, 1.550505e-05,
  6.112118e-06, 7.109099e-06, 3.80806e-05, 0.000135041, 0.0001248386, 
    0.0001717938, 0.0001862486, 1.739691e-05, 1.703627e-06, 8.443394e-06, 
    1.035598e-05, 1.351373e-05, 7.496678e-06, 1.361139e-05, 1.285819e-05,
  1.729597e-05, 1.722599e-05, 8.792878e-06, 3.816387e-06, 3.230352e-06, 
    4.049488e-06, 2.61591e-06, 3.289888e-06, 1.327915e-06, 1.898988e-06, 
    9.589425e-07, 2.227454e-06, 1.575983e-06, 8.30656e-07, 5.346948e-07,
  1.422e-05, 2.051956e-05, 2.556033e-05, 3.221087e-06, 3.309608e-06, 
    4.104497e-06, 3.982105e-06, 1.812625e-06, 8.081046e-07, 1.077295e-06, 
    1.315143e-06, 1.355082e-06, 7.191397e-07, 2.646239e-07, 1.577436e-07,
  2.170048e-05, 2.428554e-05, 4.851962e-05, 3.446745e-06, 1.308767e-06, 
    5.840967e-06, 5.107124e-06, 1.121034e-06, 8.193396e-07, 6.983057e-07, 
    1.500462e-06, 1.509588e-06, 5.118883e-07, 2.772572e-07, 6.408554e-07,
  3.179619e-05, 3.017298e-05, 8.001606e-05, 4.504864e-06, 1.352842e-06, 
    3.29892e-06, 4.284335e-06, 6.552921e-07, 1.020228e-06, 9.54172e-07, 
    1.505782e-06, 1.140198e-06, 5.401897e-07, 4.508633e-07, 5.875282e-07,
  5.269513e-05, 4.253335e-05, 0.0001163171, 9.424308e-06, 1.110936e-06, 
    2.898316e-06, 3.323551e-06, 8.308481e-07, 1.254831e-06, 1.852305e-06, 
    1.330007e-06, 1.300023e-06, 9.635971e-07, 7.65779e-07, 9.261823e-07,
  6.721242e-05, 5.576501e-05, 0.0001505197, 4.026291e-05, 2.402263e-07, 
    1.822854e-06, 2.675518e-06, 9.207611e-07, 1.450574e-06, 1.756493e-06, 
    1.544406e-06, 1.125747e-06, 1.117627e-06, 1.653559e-06, 1.588031e-06,
  9.715088e-05, 6.014438e-05, 0.0001772839, 7.696029e-05, 5.508098e-07, 
    1.961461e-06, 2.186882e-06, 5.165149e-07, 1.674665e-06, 1.192636e-06, 
    1.720398e-06, 1.46947e-06, 1.674636e-06, 1.826643e-06, 1.423149e-06,
  0.0001238286, 6.417729e-05, 0.0002001776, 0.0001107858, 2.033443e-07, 
    1.44487e-06, 1.842171e-06, 5.949237e-07, 2.11472e-06, 1.998571e-06, 
    2.564985e-06, 1.259805e-06, 1.335609e-06, 1.167673e-06, 1.539382e-06,
  0.0001431384, 6.712737e-05, 0.0002102759, 0.0001533992, 3.639544e-07, 
    1.479568e-06, 1.836512e-06, 6.97981e-07, 2.570266e-06, 1.570238e-06, 
    2.433718e-06, 1.447041e-06, 3.359259e-06, 3.278006e-06, 3.358019e-06,
  0.0001631348, 7.354475e-05, 0.0002156686, 0.0001932679, 6.947433e-07, 
    1.721037e-06, 1.830555e-06, 8.648165e-07, 3.338235e-06, 2.656676e-06, 
    5.326316e-06, 3.808866e-06, 4.328605e-06, 6.450968e-06, 6.42e-06,
  4.161744e-05, 5.518761e-05, 2.557884e-05, 5.843226e-06, 1.18392e-05, 
    1.756462e-05, 1.277732e-05, 9.897975e-06, 1.065318e-05, 1.525602e-05, 
    1.65691e-05, 1.475213e-05, 1.309859e-05, 1.219503e-05, 1.584805e-05,
  3.6597e-05, 4.400067e-05, 6.739084e-06, 5.263477e-06, 1.094016e-05, 
    1.20609e-05, 9.02389e-06, 9.258646e-06, 9.531472e-06, 1.096795e-05, 
    1.022555e-05, 1.014379e-05, 1.094177e-05, 1.194498e-05, 9.378216e-06,
  1.169443e-05, 1.030022e-05, 7.350266e-06, 5.239673e-06, 7.169186e-06, 
    7.891518e-06, 7.857759e-06, 9.028339e-06, 8.710418e-06, 1.003916e-05, 
    5.872978e-06, 8.644808e-06, 7.941173e-06, 6.813632e-06, 4.582e-06,
  1.336431e-06, 4.596946e-06, 4.826192e-06, 4.916279e-06, 5.958307e-06, 
    5.309306e-06, 7.829722e-06, 8.120806e-06, 8.044462e-06, 6.049459e-06, 
    6.347413e-06, 7.503119e-06, 4.679765e-06, 4.122757e-06, 5.753364e-06,
  2.306745e-06, 3.409788e-06, 3.536784e-06, 3.050239e-06, 4.270499e-06, 
    4.744054e-06, 6.374536e-06, 7.730946e-06, 7.844981e-06, 5.721591e-06, 
    6.68746e-06, 4.980823e-06, 4.05073e-06, 3.989828e-06, 4.914251e-06,
  1.639876e-06, 3.389137e-06, 3.635194e-06, 2.879983e-06, 2.709931e-06, 
    2.631199e-06, 6.011689e-06, 6.576683e-06, 5.502533e-06, 5.681656e-06, 
    7.395535e-06, 5.573246e-06, 4.639153e-06, 4.591946e-06, 5.014651e-06,
  1.2559e-06, 3.023561e-06, 3.385126e-06, 1.604741e-06, 1.56317e-06, 
    4.248561e-06, 5.536347e-06, 3.940287e-06, 5.406206e-06, 6.488171e-06, 
    6.626451e-06, 4.71568e-06, 5.91933e-06, 5.36762e-06, 6.187362e-06,
  6.375916e-07, 8.825581e-07, 1.110782e-06, 6.03306e-07, 1.578191e-06, 
    4.761969e-06, 4.853694e-06, 4.769104e-06, 6.202301e-06, 5.404989e-06, 
    5.047911e-06, 4.935368e-06, 7.090332e-06, 6.348127e-06, 3.348085e-06,
  6.464542e-07, 3.760638e-07, 7.294494e-07, 3.444707e-07, 2.103255e-06, 
    4.182127e-06, 3.499816e-06, 4.697426e-06, 5.532596e-06, 4.241968e-06, 
    5.290873e-06, 5.032965e-06, 4.987919e-06, 4.985493e-06, 4.077887e-06,
  3.276815e-07, 2.780043e-07, 4.969769e-07, 2.509639e-07, 2.655756e-06, 
    4.165758e-06, 2.961066e-06, 3.434739e-06, 4.257576e-06, 5.07591e-06, 
    4.589898e-06, 5.364679e-06, 5.006283e-06, 3.428082e-06, 3.827658e-06,
  0.0006443481, 0.000793707, 0.0007128783, 0.0004097166, 0.0002012593, 
    0.0001103464, 7.331451e-05, 4.846687e-05, 3.094519e-05, 2.32176e-05, 
    2.278721e-05, 1.661247e-05, 1.286371e-05, 1.186472e-05, 1.155766e-05,
  0.0005105612, 0.0006132656, 0.000566155, 0.0003467082, 0.0001143127, 
    3.320803e-05, 1.921753e-05, 1.453734e-05, 1.28833e-05, 1.536259e-05, 
    1.394958e-05, 1.229728e-05, 1.005867e-05, 1.274513e-05, 1.300255e-05,
  0.0002784021, 0.0003520618, 0.0003755586, 0.00020062, 3.32878e-05, 
    1.154349e-05, 1.18147e-05, 1.291489e-05, 1.023204e-05, 1.014592e-05, 
    1.035926e-05, 1.175231e-05, 5.518153e-06, 6.407975e-06, 8.153549e-06,
  9.735522e-05, 0.0001329337, 0.0001726496, 7.376781e-05, 1.080289e-05, 
    9.035317e-06, 1.012214e-05, 9.029042e-06, 9.487228e-06, 8.455205e-06, 
    8.096998e-06, 1.014821e-05, 6.361485e-06, 3.119272e-06, 2.829821e-06,
  1.691661e-05, 1.761537e-05, 3.438234e-05, 9.007948e-06, 9.80031e-06, 
    9.010892e-06, 9.758208e-06, 8.658815e-06, 9.502057e-06, 8.5232e-06, 
    5.353002e-06, 4.351547e-06, 8.229128e-06, 5.585276e-06, 7.64788e-06,
  7.980594e-06, 1.121006e-05, 5.348374e-06, 9.471631e-06, 6.756221e-06, 
    9.552489e-06, 9.739705e-06, 7.387181e-06, 7.183795e-06, 6.856051e-06, 
    7.448312e-06, 5.99417e-06, 4.652378e-06, 3.234397e-06, 3.607343e-06,
  4.76732e-06, 6.745257e-06, 6.244836e-06, 7.026279e-06, 7.685192e-06, 
    4.725371e-06, 5.584367e-06, 6.976918e-06, 6.533971e-06, 6.352222e-06, 
    5.325718e-06, 4.17095e-06, 6.925888e-06, 3.297152e-06, 7.070661e-06,
  6.390569e-06, 4.78546e-06, 8.623972e-06, 6.309797e-06, 7.088441e-06, 
    4.789722e-06, 4.704097e-06, 4.180109e-06, 7.973194e-06, 6.394601e-06, 
    3.420572e-06, 3.430843e-06, 4.928211e-06, 8.034136e-06, 6.619559e-06,
  4.094544e-06, 6.867871e-06, 9.290985e-06, 5.855404e-06, 6.790852e-06, 
    5.457341e-06, 4.194492e-06, 4.115191e-06, 6.270444e-06, 6.623643e-06, 
    3.533844e-06, 3.974553e-06, 5.255265e-06, 9.299257e-06, 6.814593e-06,
  6.217896e-06, 2.218519e-06, 2.776943e-06, 3.110926e-06, 5.409062e-06, 
    3.856358e-06, 4.761321e-06, 3.889427e-06, 4.107421e-06, 3.108038e-06, 
    3.756676e-06, 3.024634e-06, 5.419506e-06, 5.919196e-06, 6.332255e-06,
  5.481419e-05, 6.348783e-05, 5.600892e-05, 5.902079e-05, 9.690595e-05, 
    0.0001885016, 0.00032511, 0.0004508739, 0.0004723943, 0.0003002587, 
    0.000121745, 6.801986e-05, 2.083399e-05, 9.750197e-06, 1.68095e-05,
  0.0001142708, 0.0001371715, 0.0001317625, 0.0001457304, 0.0001832696, 
    0.000252907, 0.0003162645, 0.000380571, 0.0003360766, 0.0002025867, 
    5.110593e-05, 4.119544e-05, 2.010639e-05, 1.10277e-05, 1.908573e-05,
  0.0002210132, 0.000233615, 0.0002223517, 0.0002096556, 0.000195604, 
    0.0002202173, 0.0002455108, 0.0002721117, 0.0002466654, 0.0001409644, 
    2.700348e-05, 3.576479e-05, 1.317817e-05, 9.692781e-06, 2.003649e-05,
  0.0002857725, 0.000295245, 0.0002828671, 0.000252348, 0.000213183, 
    0.0002101822, 0.0002217625, 0.000246101, 0.0002199262, 0.0001003476, 
    2.165326e-05, 1.892648e-05, 7.219172e-06, 1.062533e-05, 1.777622e-05,
  0.0002664791, 0.0003234206, 0.0003355222, 0.0003028198, 0.0002499196, 
    0.0002398077, 0.0002274941, 0.0002056735, 0.0001853877, 8.16307e-05, 
    2.493373e-05, 1.11295e-05, 7.221869e-06, 1.515463e-05, 1.798902e-05,
  0.0002355153, 0.0003052659, 0.0003457938, 0.0003186232, 0.0002886093, 
    0.0002548867, 0.0002150507, 0.0001748684, 0.0001501435, 8.672618e-05, 
    1.918781e-05, 8.47465e-06, 9.971505e-06, 1.472337e-05, 1.689708e-05,
  0.0002121762, 0.0003008253, 0.0003374515, 0.0003353647, 0.0002903373, 
    0.0002519748, 0.0001987936, 0.0001313232, 0.0001071879, 8.031235e-05, 
    1.577117e-05, 8.006871e-06, 1.176298e-05, 1.457809e-05, 1.448167e-05,
  0.0001860012, 0.0002898812, 0.00032467, 0.000302671, 0.0002542468, 
    0.000210758, 0.0001444664, 7.375002e-05, 8.017757e-05, 6.559888e-05, 
    9.634191e-06, 1.092832e-05, 1.105759e-05, 9.983502e-06, 1.252271e-05,
  0.0001903751, 0.0003044603, 0.0003127582, 0.0002545522, 0.0001902702, 
    0.0001490085, 9.481019e-05, 4.076075e-05, 5.272769e-05, 3.794844e-05, 
    9.449736e-06, 1.122425e-05, 9.100228e-06, 9.680605e-06, 1.259408e-05,
  0.0001951868, 0.000296297, 0.00025661, 0.0001749497, 0.0001224441, 
    9.204235e-05, 5.091614e-05, 1.869908e-05, 3.028371e-05, 1.923494e-05, 
    1.110803e-05, 6.474582e-06, 9.065118e-06, 9.018416e-06, 9.457141e-06,
  1.875947e-05, 2.223551e-05, 2.682882e-05, 2.468869e-05, 2.277707e-05, 
    2.12555e-05, 2.752258e-05, 3.169955e-05, 1.919397e-05, 1.37378e-05, 
    1.215871e-05, 9.563845e-06, 1.104583e-05, 9.345031e-06, 8.799156e-06,
  1.931774e-05, 3.069162e-05, 3.716525e-05, 2.94354e-05, 2.419969e-05, 
    2.260398e-05, 3.505774e-05, 4.419552e-05, 2.611596e-05, 1.752244e-05, 
    1.258089e-05, 9.721257e-06, 1.20297e-05, 1.07901e-05, 7.742255e-06,
  2.554539e-05, 3.117495e-05, 3.875387e-05, 3.184988e-05, 2.771819e-05, 
    2.829602e-05, 5.521551e-05, 7.031209e-05, 3.367347e-05, 1.900511e-05, 
    1.251844e-05, 1.144478e-05, 1.264149e-05, 1.101133e-05, 1.186557e-05,
  2.74376e-05, 3.504783e-05, 3.753086e-05, 3.590197e-05, 3.25918e-05, 
    3.800075e-05, 0.0001000282, 0.0001095757, 4.804262e-05, 2.441231e-05, 
    1.350849e-05, 1.154109e-05, 1.34489e-05, 1.25018e-05, 1.196653e-05,
  4.879201e-05, 3.897757e-05, 4.004336e-05, 4.052196e-05, 4.098277e-05, 
    8.44672e-05, 0.0001910389, 0.0001620662, 6.533477e-05, 2.736399e-05, 
    1.447095e-05, 1.240858e-05, 1.417549e-05, 1.366195e-05, 1.179571e-05,
  6.587903e-05, 4.688805e-05, 4.045358e-05, 4.185368e-05, 4.884424e-05, 
    0.0001411438, 0.0002825788, 0.0002841947, 8.84368e-05, 2.287991e-05, 
    1.512088e-05, 1.366683e-05, 1.276762e-05, 1.206718e-05, 9.92011e-06,
  7.518732e-05, 5.774149e-05, 3.873561e-05, 2.9341e-05, 5.891258e-05, 
    0.0001700696, 0.000334975, 0.000423524, 0.0001442122, 2.437867e-05, 
    1.581544e-05, 1.11044e-05, 1.358411e-05, 1.279256e-05, 1.026053e-05,
  9.802145e-05, 7.905011e-05, 3.260968e-05, 1.797754e-05, 7.20615e-05, 
    0.0002160713, 0.0004298414, 0.0004906585, 0.0002183504, 2.192358e-05, 
    1.70957e-05, 1.277257e-05, 1.389222e-05, 1.155033e-05, 7.942591e-06,
  0.000140334, 0.0001086512, 3.569076e-05, 2.498396e-05, 0.0001120864, 
    0.0002610818, 0.0004723386, 0.0005316262, 0.0002705397, 2.023425e-05, 
    1.615539e-05, 1.575332e-05, 1.338509e-05, 9.162794e-06, 8.126417e-06,
  0.0002087949, 0.0001684373, 7.565915e-05, 5.447843e-05, 0.0001656391, 
    0.0003003434, 0.0004258975, 0.0005030713, 0.0002802488, 9.609105e-06, 
    1.598889e-05, 1.532055e-05, 1.045347e-05, 8.785311e-06, 7.371731e-06,
  7.459284e-06, 7.066368e-06, 6.274522e-06, 5.461911e-06, 4.782132e-06, 
    3.851271e-06, 4.107243e-06, 4.837649e-06, 5.680705e-06, 4.766571e-06, 
    4.585652e-06, 4.346737e-06, 5.297878e-06, 5.256129e-06, 5.05203e-06,
  9.356266e-06, 8.548345e-06, 6.491018e-06, 6.240967e-06, 3.934795e-06, 
    4.828134e-06, 5.674272e-06, 5.521515e-06, 5.856196e-06, 4.893433e-06, 
    4.978768e-06, 4.480498e-06, 4.517929e-06, 5.187385e-06, 3.872066e-06,
  1.066611e-05, 9.463713e-06, 1.017977e-05, 5.811457e-06, 6.104465e-06, 
    6.946814e-06, 5.876207e-06, 6.538603e-06, 5.960398e-06, 6.213245e-06, 
    4.961568e-06, 5.11417e-06, 6.261728e-06, 6.346853e-06, 7.298147e-06,
  1.419349e-05, 1.482669e-05, 1.183401e-05, 6.640875e-06, 9.445018e-06, 
    8.58222e-06, 6.879602e-06, 6.920127e-06, 6.352765e-06, 6.287351e-06, 
    6.332545e-06, 6.831397e-06, 7.419905e-06, 7.375359e-06, 1.1124e-05,
  1.880907e-05, 1.94983e-05, 1.563306e-05, 1.196698e-05, 1.184227e-05, 
    1.031164e-05, 8.598066e-06, 7.138351e-06, 7.667393e-06, 7.319202e-06, 
    8.469722e-06, 6.610472e-06, 8.366919e-06, 8.982114e-06, 1.035205e-05,
  2.501457e-05, 1.872326e-05, 2.029914e-05, 1.731587e-05, 1.500433e-05, 
    1.26364e-05, 9.269788e-06, 8.269493e-06, 8.289971e-06, 7.78004e-06, 
    8.742639e-06, 8.293458e-06, 9.18254e-06, 8.916198e-06, 8.994237e-06,
  2.788836e-05, 2.798965e-05, 2.807851e-05, 2.808596e-05, 2.13991e-05, 
    1.689161e-05, 1.027471e-05, 8.847658e-06, 1.011267e-05, 9.969906e-06, 
    8.326689e-06, 7.788007e-06, 8.530998e-06, 9.285677e-06, 9.624321e-06,
  2.788593e-05, 2.30456e-05, 3.555896e-05, 4.960669e-05, 4.036842e-05, 
    2.685242e-05, 1.491855e-05, 9.865382e-06, 1.160077e-05, 1.060695e-05, 
    8.084568e-06, 7.792122e-06, 8.820401e-06, 1.158117e-05, 9.630374e-06,
  2.780523e-05, 3.330708e-05, 4.744934e-05, 5.604027e-05, 4.876099e-05, 
    4.188779e-05, 2.372883e-05, 1.340309e-05, 1.191046e-05, 1.221832e-05, 
    8.351081e-06, 7.226962e-06, 9.836315e-06, 1.023889e-05, 1.022005e-05,
  2.619589e-05, 3.76091e-05, 3.835049e-05, 3.296368e-05, 2.443333e-05, 
    2.792194e-05, 2.70612e-05, 1.578526e-05, 1.340909e-05, 1.266816e-05, 
    1.124669e-05, 9.657077e-06, 7.499652e-06, 1.09338e-05, 1.15141e-05,
  6.642932e-07, 1.564648e-06, 2.272617e-06, 1.802541e-06, 1.700595e-06, 
    1.759244e-06, 2.821063e-06, 1.873147e-06, 2.537714e-06, 5.028633e-06, 
    7.590948e-06, 8.168511e-06, 1.070548e-05, 1.133336e-05, 1.077261e-05,
  2.502571e-06, 1.425377e-06, 1.489046e-06, 1.262092e-06, 1.523713e-06, 
    2.525974e-06, 2.362966e-06, 2.644761e-06, 2.303992e-06, 2.46239e-06, 
    4.604181e-06, 4.605407e-06, 3.642872e-06, 5.114564e-06, 5.678625e-06,
  2.279346e-06, 1.259621e-06, 1.672822e-06, 2.150537e-06, 3.309045e-06, 
    4.35643e-06, 5.025098e-06, 4.11775e-06, 4.537156e-06, 5.971442e-06, 
    6.823389e-06, 6.0366e-06, 7.176288e-06, 7.340797e-06, 7.630601e-06,
  3.05507e-06, 3.488732e-06, 3.94277e-06, 3.90444e-06, 4.196514e-06, 
    4.397054e-06, 5.823915e-06, 5.031631e-06, 5.141368e-06, 8.858128e-06, 
    7.653979e-06, 8.29415e-06, 8.579457e-06, 9.036237e-06, 8.534952e-06,
  3.188557e-06, 4.560872e-06, 3.654301e-06, 2.826692e-06, 2.45417e-06, 
    2.814003e-06, 2.861287e-06, 2.547642e-06, 2.40474e-06, 2.23301e-06, 
    2.787402e-06, 4.470584e-06, 3.729957e-06, 3.067042e-06, 3.751564e-06,
  3.631304e-06, 3.917269e-06, 2.990857e-06, 2.970279e-06, 2.578442e-06, 
    2.409959e-06, 2.521771e-06, 2.034529e-06, 1.858132e-06, 1.474326e-06, 
    2.457913e-07, 2.019722e-07, 7.628598e-08, 5.37199e-07, 2.510729e-07,
  4.683973e-06, 4.098974e-06, 2.99461e-06, 3.174674e-06, 2.983924e-06, 
    3.338453e-06, 3.175259e-06, 2.457511e-06, 2.42785e-06, 1.374071e-06, 
    8.897634e-07, 6.677928e-07, 8.508547e-08, 1.37594e-07, 2.505199e-06,
  4.175998e-06, 4.506751e-06, 3.790024e-06, 3.503989e-06, 3.83155e-06, 
    3.848555e-06, 3.570819e-06, 3.864508e-06, 3.663788e-06, 3.785487e-06, 
    3.574511e-06, 3.557484e-06, 1.608691e-06, 1.024015e-06, 2.710097e-06,
  5.741852e-06, 5.303917e-06, 4.495741e-06, 4.475471e-06, 5.625152e-06, 
    6.186814e-06, 4.74378e-06, 5.172373e-06, 4.138079e-06, 4.78114e-06, 
    4.724489e-06, 4.913313e-06, 4.880511e-06, 3.24859e-06, 2.088105e-06,
  5.856925e-06, 5.343218e-06, 6.092607e-06, 5.325493e-06, 7.629539e-06, 
    6.878479e-06, 6.374918e-06, 5.116082e-06, 6.632541e-06, 6.59947e-06, 
    5.687571e-06, 5.842002e-06, 7.273011e-06, 4.289285e-06, 4.377127e-06,
  5.190433e-06, 4.728389e-06, 7.435914e-06, 3.744189e-05, 0.0001025064, 
    0.000178496, 0.0002626211, 0.0003407295, 0.0004272766, 0.0004485227, 
    0.0005414434, 0.0005596883, 0.000434211, 0.0002418165, 7.411464e-05,
  5.534949e-06, 6.16745e-06, 5.509169e-06, 8.376136e-06, 2.900035e-05, 
    6.195171e-05, 0.0001167844, 0.0001753126, 0.0002242265, 0.0002639368, 
    0.0003575434, 0.0004299711, 0.0004033001, 0.0002558787, 0.0001224299,
  5.667093e-06, 6.193143e-06, 7.361713e-06, 7.284405e-06, 7.648628e-06, 
    1.978799e-05, 4.796227e-05, 7.915907e-05, 0.0001131488, 0.0001255741, 
    0.0001736001, 0.0002949345, 0.0003396851, 0.0002666522, 0.0001741786,
  5.994221e-06, 6.082319e-06, 7.351894e-06, 7.813234e-06, 8.258293e-06, 
    1.001162e-05, 1.583005e-05, 3.337174e-05, 5.414417e-05, 5.707786e-05, 
    6.511519e-05, 0.0001187409, 0.0001977246, 0.00022383, 0.0002035707,
  3.398928e-06, 3.205025e-06, 3.47931e-06, 3.910336e-06, 5.174603e-06, 
    7.459615e-06, 6.81277e-06, 1.05938e-05, 1.735011e-05, 2.051611e-05, 
    2.44289e-05, 3.643192e-05, 7.62735e-05, 0.0001341508, 0.0001679792,
  2.37442e-06, 2.226612e-06, 1.696752e-06, 2.088751e-06, 1.60378e-06, 
    1.999775e-06, 2.216713e-06, 2.998838e-06, 5.574349e-06, 7.590944e-06, 
    8.214422e-06, 1.153415e-05, 1.987864e-05, 4.883654e-05, 7.830722e-05,
  1.723791e-06, 2.218093e-06, 2.559023e-06, 2.283057e-06, 2.137897e-06, 
    1.759361e-06, 1.750906e-06, 6.763948e-07, 1.436179e-06, 4.685135e-06, 
    3.387188e-06, 4.519872e-06, 7.234655e-06, 8.086798e-06, 1.650807e-05,
  2.597529e-06, 1.917773e-06, 2.52601e-06, 2.77327e-06, 2.61497e-06, 
    3.131401e-06, 2.733939e-06, 1.301716e-06, 4.749615e-06, 3.778481e-06, 
    2.073941e-06, 1.464877e-06, 3.191142e-06, 3.244091e-06, 4.900255e-06,
  1.609292e-06, 2.540964e-06, 1.57921e-06, 3.24467e-06, 3.452928e-06, 
    4.878854e-06, 4.889911e-06, 4.731313e-06, 4.22021e-06, 3.016864e-06, 
    2.419967e-06, 3.298331e-06, 1.899488e-06, 1.984689e-06, 4.422811e-06,
  3.706929e-06, 4.003868e-06, 7.068283e-07, 1.660887e-06, 3.811352e-06, 
    6.661488e-06, 6.011024e-06, 2.619799e-06, 2.478434e-06, 2.354393e-06, 
    3.233697e-06, 3.334454e-06, 1.66601e-06, 3.576223e-06, 4.047294e-06,
  0.0006515467, 0.001108036, 0.001432085, 0.001366027, 0.0008586898, 
    0.0004135679, 0.0001784799, 5.739002e-05, 1.118653e-05, 8.301799e-06, 
    1.948533e-05, 2.745628e-05, 2.993376e-05, 3.00876e-05, 2.803392e-05,
  0.0007341559, 0.001176839, 0.001461928, 0.001240386, 0.000691277, 
    0.0003268745, 0.00014773, 5.872795e-05, 2.234732e-05, 1.065109e-05, 
    1.555527e-05, 2.978412e-05, 3.374488e-05, 3.016331e-05, 2.068929e-05,
  0.0006978182, 0.001036606, 0.001230445, 0.0009789587, 0.0004046882, 
    0.0002025275, 0.0001177352, 7.488943e-05, 4.384374e-05, 1.824476e-05, 
    1.651288e-05, 2.834946e-05, 4.962105e-05, 4.999385e-05, 3.732217e-05,
  0.0005098064, 0.0007493497, 0.0009340747, 0.0007444972, 0.0002697331, 
    0.0001373971, 0.0001131042, 9.010825e-05, 6.755397e-05, 4.796494e-05, 
    3.279656e-05, 4.387115e-05, 8.28202e-05, 0.0001063629, 9.440701e-05,
  0.0001968326, 0.0003914445, 0.0005090645, 0.000450184, 0.0002160653, 
    0.0001110476, 0.0001140557, 0.0001137301, 9.077758e-05, 7.128455e-05, 
    6.412633e-05, 6.547941e-05, 0.0001215512, 0.0001919391, 0.0002133336,
  3.130972e-05, 8.634781e-05, 0.0001637261, 0.0001798506, 0.0001284123, 
    9.192144e-05, 9.166094e-05, 0.0001035435, 0.0001011589, 8.559554e-05, 
    6.293827e-05, 5.125204e-05, 8.629109e-05, 0.0002019531, 0.0002938778,
  8.978657e-06, 1.513335e-05, 2.650501e-05, 5.337702e-05, 5.65342e-05, 
    5.885066e-05, 6.052273e-05, 8.043624e-05, 0.0001001468, 8.173056e-05, 
    5.931551e-05, 4.055722e-05, 4.354087e-05, 0.000111717, 0.0002417831,
  5.384915e-06, 5.187392e-06, 6.800654e-06, 9.84241e-06, 2.446737e-05, 
    4.073733e-05, 4.628297e-05, 6.180199e-05, 9.365076e-05, 9.13511e-05, 
    6.80151e-05, 4.320439e-05, 3.740585e-05, 6.45192e-05, 0.0001494707,
  5.478882e-06, 5.824593e-06, 4.848654e-06, 6.143965e-06, 6.647809e-06, 
    1.395862e-05, 2.31101e-05, 3.88677e-05, 6.216639e-05, 7.512189e-05, 
    6.450756e-05, 4.533099e-05, 3.124181e-05, 4.38561e-05, 9.293265e-05,
  4.902348e-06, 6.236412e-06, 6.322422e-06, 5.462685e-06, 3.886823e-06, 
    3.795443e-06, 8.195428e-06, 1.597296e-05, 2.936989e-05, 3.862047e-05, 
    3.646667e-05, 2.904336e-05, 2.005523e-05, 1.962137e-05, 3.487962e-05,
  0.0004015615, 0.0005753497, 0.0003881392, 3.99197e-05, 9.999652e-06, 
    7.577856e-06, 1.022601e-05, 2.319604e-05, 2.44129e-05, 2.045408e-05, 
    1.814617e-05, 1.141575e-05, 9.742424e-06, 1.039066e-05, 8.161021e-06,
  0.0007803364, 0.0008740277, 0.0003365577, 1.457907e-05, 7.502017e-06, 
    9.814586e-06, 1.401763e-05, 2.029049e-05, 1.878331e-05, 1.726332e-05, 
    1.232568e-05, 8.028101e-06, 9.113562e-06, 5.31388e-06, 6.909865e-06,
  0.001126096, 0.0009846311, 0.0002202503, 9.715402e-06, 5.088569e-06, 
    7.999503e-06, 9.533146e-06, 1.085169e-05, 1.189661e-05, 1.255041e-05, 
    1.393648e-05, 1.274105e-05, 8.838776e-06, 7.371223e-06, 7.242917e-06,
  0.001259908, 0.0007974147, 0.0002653474, 4.423039e-05, 5.71076e-06, 
    6.187888e-06, 9.088439e-06, 8.284967e-06, 9.999721e-06, 1.006904e-05, 
    8.693242e-06, 8.74237e-06, 1.143835e-05, 1.054535e-05, 8.018582e-06,
  0.001108726, 0.0006715572, 0.0004076706, 0.0001718994, 2.123516e-05, 
    8.176052e-06, 1.075142e-05, 1.098559e-05, 1.163954e-05, 9.656452e-06, 
    6.832393e-06, 8.213548e-06, 1.381325e-05, 1.269153e-05, 9.203853e-06,
  0.001015334, 0.0007258446, 0.0005018737, 0.0002767317, 8.256883e-05, 
    1.418211e-05, 1.107498e-05, 1.36946e-05, 1.495175e-05, 1.051031e-05, 
    9.712063e-06, 1.04435e-05, 1.359642e-05, 1.433101e-05, 9.774451e-06,
  0.0008653229, 0.0006655825, 0.0004733789, 0.0003042954, 0.0001317452, 
    2.49333e-05, 9.615793e-06, 2.05345e-05, 2.850886e-05, 2.362226e-05, 
    1.516606e-05, 1.159527e-05, 1.114032e-05, 1.111158e-05, 8.662616e-06,
  0.0005877372, 0.0005089361, 0.0003797806, 0.0002732423, 0.0001562619, 
    6.072005e-05, 1.557683e-05, 2.578158e-05, 4.734427e-05, 4.449187e-05, 
    3.204698e-05, 2.042747e-05, 1.144988e-05, 1.067838e-05, 1.211921e-05,
  0.0003332559, 0.0002939325, 0.0002427939, 0.000215361, 0.0001846471, 
    0.0001150707, 4.637261e-05, 4.343129e-05, 8.232135e-05, 0.0001026764, 
    7.998562e-05, 4.950495e-05, 2.931925e-05, 1.874319e-05, 1.264159e-05,
  0.0001735566, 0.0002084062, 0.0002074895, 0.0001991272, 0.0002142969, 
    0.0001887019, 9.800593e-05, 4.806265e-05, 7.898806e-05, 0.0001361101, 
    0.0001413291, 0.000102026, 6.112616e-05, 2.832116e-05, 1.207431e-05,
  1.143671e-05, 1.302141e-05, 1.312695e-05, 1.503866e-05, 1.588471e-05, 
    1.568733e-05, 1.566765e-05, 1.286729e-05, 1.136802e-05, 1.323239e-05, 
    1.677019e-05, 1.68675e-05, 1.808698e-05, 1.730391e-05, 1.7122e-05,
  5.87833e-06, 7.668561e-06, 9.605184e-06, 1.530029e-05, 1.721379e-05, 
    1.4791e-05, 1.340783e-05, 1.49436e-05, 1.414057e-05, 1.309617e-05, 
    7.812939e-06, 8.557479e-06, 1.531828e-05, 2.09795e-05, 1.777682e-05,
  7.678975e-06, 1.01837e-05, 1.02864e-05, 1.114004e-05, 1.367396e-05, 
    1.236374e-05, 1.600346e-05, 1.248146e-05, 1.209067e-05, 5.614706e-06, 
    9.889756e-06, 1.433745e-05, 1.404805e-05, 1.557879e-05, 1.539843e-05,
  1.02035e-05, 6.130098e-06, 1.016595e-05, 1.147999e-05, 1.153683e-05, 
    1.061359e-05, 9.349867e-06, 1.289651e-05, 1.068747e-05, 8.943894e-06, 
    4.22574e-06, 6.324507e-06, 1.110874e-05, 1.223213e-05, 1.309235e-05,
  1.273947e-05, 6.980671e-06, 7.330797e-06, 1.04259e-05, 1.018352e-05, 
    1.134798e-05, 1.071305e-05, 9.777737e-06, 7.724744e-06, 8.391983e-06, 
    4.077566e-06, 2.505812e-06, 9.620476e-06, 1.208958e-05, 1.119514e-05,
  1.654953e-05, 7.606273e-06, 7.889688e-06, 1.127698e-05, 1.326705e-05, 
    1.228561e-05, 1.178886e-05, 1.214526e-05, 9.790327e-06, 7.397958e-06, 
    6.413869e-06, 3.998111e-06, 6.324105e-06, 1.108289e-05, 1.324697e-05,
  3.728298e-05, 1.254097e-05, 5.832024e-06, 9.721662e-06, 1.236765e-05, 
    1.322021e-05, 1.417396e-05, 1.183158e-05, 1.134262e-05, 9.536309e-06, 
    7.636379e-06, 2.763963e-06, 9.749631e-06, 1.248251e-05, 1.554692e-05,
  6.363972e-05, 2.186279e-05, 7.98322e-06, 5.240184e-06, 1.222983e-05, 
    1.421767e-05, 1.353667e-05, 1.16184e-05, 1.054921e-05, 9.307208e-06, 
    9.653958e-06, 4.366938e-06, 1.011719e-05, 1.066221e-05, 1.914343e-05,
  9.76306e-05, 3.759809e-05, 1.55471e-05, 1.102095e-05, 1.04161e-05, 
    1.123659e-05, 9.820874e-06, 1.14712e-05, 1.141683e-05, 1.027921e-05, 
    7.429603e-06, 7.519667e-06, 9.766764e-06, 9.380075e-06, 1.803708e-05,
  0.0001235153, 5.32106e-05, 3.003318e-05, 1.616697e-05, 1.253679e-05, 
    1.106706e-05, 1.122389e-05, 1.076855e-05, 1.192552e-05, 1.071879e-05, 
    9.226241e-06, 6.429688e-06, 1.31661e-05, 1.041629e-05, 1.496258e-05,
  1.600116e-05, 1.834655e-05, 1.537496e-05, 1.753646e-05, 1.405347e-05, 
    1.296376e-05, 5.746234e-06, 4.310798e-06, 3.845529e-06, 4.59842e-06, 
    1.78599e-06, 2.898013e-06, 3.406904e-06, 3.750061e-06, 5.524146e-06,
  8.087763e-06, 1.747835e-05, 1.793673e-05, 1.782198e-05, 1.798469e-05, 
    1.516532e-05, 9.411679e-06, 7.545096e-06, 4.224776e-06, 3.313607e-06, 
    3.232344e-06, 2.333476e-06, 7.564793e-06, 4.992966e-06, 5.934946e-06,
  1.524294e-05, 1.370739e-05, 1.500945e-05, 1.689851e-05, 1.825085e-05, 
    1.499677e-05, 1.068316e-05, 5.31865e-06, 6.209075e-06, 4.703994e-06, 
    4.138219e-06, 3.113491e-06, 4.901623e-06, 5.480159e-06, 5.939949e-06,
  1.587595e-05, 1.740571e-05, 1.808972e-05, 1.516259e-05, 1.802983e-05, 
    1.447822e-05, 9.654706e-06, 5.221931e-06, 6.172826e-06, 6.656294e-06, 
    5.956318e-06, 4.448138e-06, 5.400991e-06, 7.263307e-06, 8.566388e-06,
  1.851002e-05, 1.919948e-05, 2.033553e-05, 1.478554e-05, 1.812328e-05, 
    1.324536e-05, 8.544336e-06, 4.053798e-06, 3.475178e-06, 3.724499e-06, 
    5.029072e-06, 4.830059e-06, 6.432739e-06, 7.632892e-06, 9.077165e-06,
  2.010597e-05, 1.71986e-05, 2.120494e-05, 1.722096e-05, 1.363998e-05, 
    1.371761e-05, 9.257945e-06, 6.869097e-06, 4.478978e-06, 3.340712e-06, 
    4.169911e-06, 5.749334e-06, 6.710487e-06, 1.023721e-05, 1.082627e-05,
  2.09361e-05, 1.96088e-05, 2.017722e-05, 2.046202e-05, 1.622235e-05, 
    1.438999e-05, 1.132442e-05, 1.113991e-05, 7.138273e-06, 4.244476e-06, 
    4.416397e-06, 7.989645e-06, 1.049525e-05, 1.109845e-05, 1.314767e-05,
  1.777379e-05, 2.02042e-05, 2.143291e-05, 2.067984e-05, 2.012971e-05, 
    1.237027e-05, 1.095747e-05, 1.013056e-05, 9.76934e-06, 5.360035e-06, 
    3.789593e-06, 9.832003e-06, 1.238669e-05, 1.501527e-05, 1.404948e-05,
  1.728003e-05, 1.799575e-05, 1.949609e-05, 2.140242e-05, 2.07713e-05, 
    1.470726e-05, 1.049454e-05, 1.34498e-05, 1.09893e-05, 7.436748e-06, 
    4.494267e-06, 8.601464e-06, 1.659315e-05, 2.079146e-05, 2.107663e-05,
  1.704865e-05, 1.827037e-05, 2.002345e-05, 1.796324e-05, 1.857315e-05, 
    1.713597e-05, 1.202128e-05, 1.053171e-05, 1.219696e-05, 1.024967e-05, 
    5.097877e-06, 9.125318e-06, 1.960417e-05, 2.832867e-05, 2.804412e-05,
  6.86929e-06, 4.678698e-06, 3.143594e-06, 3.286321e-07, 1.104168e-06, 
    1.363827e-06, 1.061372e-06, 1.021021e-06, 1.179722e-06, 8.432356e-07, 
    1.370504e-06, 9.100509e-07, 2.182526e-06, 1.138871e-06, 2.194549e-06,
  6.633926e-06, 3.652505e-06, 2.072012e-06, 1.356406e-06, 8.970786e-07, 
    7.743064e-07, 1.111254e-06, 1.135438e-06, 1.07263e-06, 1.174665e-06, 
    9.532247e-07, 8.997978e-07, 2.180229e-06, 2.237623e-06, 3.270764e-06,
  5.541879e-06, 3.783543e-06, 2.153707e-06, 1.012602e-06, 1.321348e-06, 
    9.015819e-07, 8.698578e-07, 9.439498e-07, 1.13717e-06, 1.538506e-06, 
    8.503902e-07, 1.091372e-06, 1.997669e-06, 4.124235e-06, 4.683349e-06,
  4.073082e-06, 2.213502e-06, 2.096086e-06, 7.091474e-07, 7.944467e-07, 
    1.266506e-06, 8.074271e-07, 1.204541e-06, 1.515921e-06, 1.872784e-06, 
    2.190633e-06, 2.339435e-06, 4.37696e-06, 5.086634e-06, 4.822346e-06,
  5.546548e-06, 3.626176e-06, 1.865594e-06, 4.629158e-07, 9.99158e-07, 
    1.545366e-06, 1.108264e-06, 1.383271e-06, 1.851693e-06, 2.133267e-06, 
    2.390453e-06, 3.129061e-06, 4.669464e-06, 5.69618e-06, 5.144557e-06,
  9.532385e-06, 4.8623e-06, 2.267576e-06, 1.313679e-06, 1.165892e-06, 
    1.470569e-06, 1.429286e-06, 1.606922e-06, 2.263513e-06, 2.268351e-06, 
    2.76251e-06, 3.624759e-06, 4.581083e-06, 5.322761e-06, 4.870714e-06,
  8.461532e-06, 8.761162e-06, 3.506271e-06, 1.07957e-06, 1.091673e-06, 
    1.408863e-06, 1.529274e-06, 1.649849e-06, 2.316647e-06, 2.159697e-06, 
    2.665286e-06, 4.743014e-06, 4.670424e-06, 4.929968e-06, 5.183671e-06,
  5.568667e-06, 5.024166e-06, 1.969737e-06, 9.383112e-07, 1.372339e-06, 
    1.463369e-06, 1.510269e-06, 1.947973e-06, 2.571725e-06, 2.870328e-06, 
    2.827343e-06, 4.64552e-06, 6.60502e-06, 5.392093e-06, 6.652817e-06,
  9.513066e-06, 2.784119e-06, 1.442576e-06, 1.295989e-06, 1.307514e-06, 
    1.827593e-06, 1.711036e-06, 2.563173e-06, 2.555219e-06, 3.214437e-06, 
    4.043087e-06, 6.226342e-06, 7.843133e-06, 7.583933e-06, 8.150668e-06,
  9.331348e-06, 3.940876e-06, 2.420203e-06, 1.051334e-06, 1.602409e-06, 
    1.822065e-06, 2.018697e-06, 3.49045e-06, 3.520833e-06, 3.416406e-06, 
    5.577318e-06, 8.785372e-06, 1.056039e-05, 1.066605e-05, 1.145375e-05,
  3.228713e-06, 3.704394e-06, 2.337868e-06, 3.48176e-06, 1.907264e-06, 
    2.043034e-06, 1.257211e-06, 1.781708e-07, 9.815288e-07, 5.368134e-07, 
    8.42619e-07, 2.108118e-06, 4.089251e-06, 7.533373e-06, 8.050347e-06,
  5.653028e-06, 3.08798e-06, 3.437537e-06, 2.353444e-06, 5.723676e-07, 
    1.243537e-06, 1.061049e-06, 1.454049e-06, 1.098165e-06, 1.121408e-06, 
    1.250751e-06, 3.129222e-06, 5.941816e-06, 1.013524e-05, 1.179276e-05,
  2.709751e-06, 2.195952e-06, 1.265956e-06, 1.450881e-06, 1.040498e-06, 
    6.098983e-07, 1.674104e-06, 1.12185e-06, 1.564704e-06, 1.905099e-06, 
    3.441936e-06, 4.884413e-06, 9.051115e-06, 1.148471e-05, 1.157909e-05,
  1.441072e-06, 7.355658e-07, 5.322702e-07, 7.595654e-07, 7.973302e-07, 
    1.077987e-06, 1.721647e-06, 1.417229e-06, 1.581034e-06, 3.207284e-06, 
    3.937414e-06, 7.208858e-06, 1.092433e-05, 1.161589e-05, 9.568682e-06,
  2.17374e-07, 1.762512e-07, 2.278084e-07, 1.943341e-06, 1.521037e-06, 
    5.074023e-07, 1.30544e-06, 1.435192e-06, 2.448727e-06, 2.929578e-06, 
    6.684426e-06, 8.234018e-06, 8.540256e-06, 8.010828e-06, 7.523241e-06,
  4.500192e-08, 3.752513e-08, 3.161373e-07, 2.310909e-06, 1.07962e-06, 
    1.142206e-06, 1.426111e-06, 1.464524e-06, 4.868068e-06, 6.179322e-06, 
    6.679132e-06, 7.186723e-06, 7.18939e-06, 6.613062e-06, 6.44019e-06,
  4.311767e-08, 2.953914e-07, 1.334247e-06, 2.123941e-06, 1.174517e-06, 
    1.370827e-06, 1.377007e-06, 3.985021e-06, 4.124554e-06, 4.927706e-06, 
    6.352989e-06, 8.2487e-06, 8.487179e-06, 1.015935e-05, 8.057713e-06,
  2.132933e-07, 1.973269e-07, 5.683956e-07, 2.680614e-06, 4.793026e-07, 
    6.058254e-07, 2.651595e-06, 2.254803e-06, 3.894533e-06, 5.563259e-06, 
    6.98689e-06, 8.216872e-06, 9.013726e-06, 9.837911e-06, 1.097187e-05,
  2.573738e-07, 2.465406e-07, 1.650642e-06, 9.456745e-07, 4.483301e-07, 
    2.47066e-06, 2.161782e-06, 2.591815e-06, 4.097256e-06, 4.828153e-06, 
    6.733592e-06, 7.223559e-06, 9.993773e-06, 8.408309e-06, 7.750328e-06,
  1.541762e-06, 2.17059e-06, 1.085118e-06, 1.036847e-06, 1.980747e-06, 
    2.118677e-06, 2.009395e-06, 3.028562e-06, 4.943333e-06, 8.166088e-06, 
    5.923207e-06, 8.038672e-06, 6.880569e-06, 6.439354e-06, 5.418827e-06,
  6.061619e-05, 3.740932e-05, 6.510576e-05, 0.000125473, 0.0002039761, 
    0.0004109469, 0.0007290174, 0.000818332, 0.000784833, 0.0002514227, 
    1.028956e-06, 6.884417e-06, 3.226455e-06, 4.242456e-06, 7.719754e-06,
  7.984032e-05, 6.352131e-05, 6.593578e-05, 0.000151207, 0.0002779947, 
    0.0004773628, 0.0006150241, 0.0006111567, 0.0005657301, 8.798606e-05, 
    5.403937e-07, 3.827705e-06, 3.480287e-06, 6.853888e-06, 8.751124e-06,
  9.652579e-05, 9.167456e-05, 6.930497e-05, 0.0001718039, 0.0003043727, 
    0.0004243412, 0.0004163572, 0.0003913011, 0.0003572039, 1.061207e-05, 
    1.081444e-06, 2.988391e-06, 5.429572e-06, 9.594285e-06, 7.833979e-06,
  8.704576e-05, 0.000121772, 0.0001106001, 0.000176206, 0.0002840561, 
    0.0003193301, 0.0002773107, 0.0002266726, 0.0001400665, 1.075048e-06, 
    1.775248e-06, 2.884326e-06, 8.563556e-06, 7.677269e-06, 5.692651e-06,
  6.964667e-05, 0.0001495205, 0.0001619379, 0.0001712261, 0.0002150605, 
    0.0001880568, 0.0001605672, 0.0001266507, 2.13465e-05, 1.737082e-06, 
    1.439643e-06, 7.236556e-06, 8.712947e-06, 7.323425e-06, 4.052924e-06,
  5.790089e-05, 0.0001674389, 0.0002081156, 0.0001546988, 0.0001099317, 
    8.787353e-05, 7.952e-05, 4.032117e-05, 1.693663e-06, 2.227729e-06, 
    4.113827e-06, 8.25685e-06, 8.480663e-06, 7.262813e-06, 5.508985e-06,
  4.380276e-05, 0.0001786253, 0.0002357324, 0.0001374348, 4.128592e-05, 
    3.438701e-05, 4.26976e-05, 3.849574e-06, 2.797732e-06, 3.173604e-06, 
    7.701148e-06, 1.178462e-05, 7.735522e-06, 5.221775e-06, 8.559024e-06,
  3.776018e-05, 0.0001806981, 0.0002366639, 0.0001286372, 2.180256e-05, 
    1.479727e-05, 2.051323e-05, 3.747386e-06, 2.793202e-06, 5.237772e-06, 
    9.360403e-06, 9.057776e-06, 5.825864e-06, 1.818892e-06, 7.512022e-06,
  3.283556e-05, 0.0001655711, 0.0002079731, 0.0001099369, 2.20232e-05, 
    9.759348e-06, 5.832946e-06, 3.069547e-06, 5.009003e-06, 7.810663e-06, 
    7.422934e-07, 3.962322e-06, 1.349743e-06, 2.489496e-06, 4.943806e-06,
  2.765979e-05, 0.0001343529, 0.0001620804, 9.221e-05, 2.314446e-05, 
    8.241826e-06, 2.974966e-06, 3.783813e-06, 5.117548e-06, 2.594312e-06, 
    5.416341e-07, 3.21709e-06, 1.509818e-06, 3.387971e-06, 7.984881e-06,
  2.329523e-05, 2.637843e-05, 2.389476e-05, 8.727879e-06, 0.0001467715, 
    0.000573792, 0.0007115916, 0.0001850276, 1.813204e-05, 5.78751e-06, 
    7.6672e-06, 9.415148e-06, 9.058974e-06, 1.001319e-05, 1.078411e-05,
  2.333694e-05, 3.020555e-05, 1.782229e-05, 8.215867e-06, 4.478282e-05, 
    0.0005216873, 0.00106814, 0.0006992017, 4.381681e-05, 3.041649e-06, 
    7.002548e-06, 7.568082e-06, 6.273754e-06, 8.042321e-06, 9.267518e-06,
  2.74274e-05, 2.994868e-05, 1.732222e-05, 5.988732e-06, 1.669197e-05, 
    0.0003520919, 0.0008590165, 0.0009390182, 0.0001365468, 9.46365e-06, 
    5.767259e-06, 6.424812e-06, 5.092997e-06, 6.85685e-06, 6.894858e-06,
  2.6167e-05, 3.33975e-05, 2.284245e-05, 9.676319e-06, 4.159219e-05, 
    0.0001963581, 0.0005612068, 0.0006536505, 0.0002418477, 2.889121e-06, 
    3.615739e-06, 3.957792e-06, 4.368238e-06, 5.557834e-06, 8.927252e-06,
  3.788986e-05, 3.292351e-05, 2.91435e-05, 3.043181e-05, 9.81357e-05, 
    0.0002158015, 0.0003190109, 0.0004090093, 0.0002159076, 4.016578e-06, 
    3.521665e-06, 2.380096e-06, 3.783653e-06, 5.393113e-06, 8.620729e-06,
  0.0001081697, 3.378347e-05, 3.678044e-05, 6.008345e-05, 0.0001631363, 
    0.0002526061, 0.0002770355, 0.0003137979, 0.0001876635, 3.219171e-06, 
    1.813742e-06, 7.431192e-07, 2.1714e-06, 4.983383e-06, 6.402561e-06,
  0.0002265986, 6.423357e-05, 4.638225e-05, 8.985669e-05, 0.0001985496, 
    0.0002499937, 0.0002494727, 0.0002742861, 0.0001299729, 9.780327e-08, 
    1.39279e-06, 1.130142e-06, 3.54324e-06, 6.789594e-06, 3.153827e-06,
  0.0003220272, 0.0002037555, 6.088497e-05, 9.709565e-05, 0.0001984169, 
    0.0002165033, 0.0002093645, 0.0001770454, 5.082611e-05, 1.810646e-07, 
    1.455254e-06, 9.791929e-07, 4.352485e-06, 6.161859e-06, 3.211994e-06,
  0.0003430014, 0.000334226, 0.0001243489, 0.0001045113, 0.0001795165, 
    0.0001831542, 0.0001674842, 9.311811e-05, 2.079646e-05, 7.664963e-07, 
    1.627132e-06, 2.044415e-06, 4.089944e-06, 5.647729e-06, 2.458351e-06,
  0.0002803895, 0.0004470474, 0.000229311, 0.0001103524, 0.0001620949, 
    0.0001681997, 0.0001415312, 6.110687e-05, 4.520376e-06, 1.859569e-06, 
    2.321409e-06, 2.316174e-06, 6.791214e-06, 4.228262e-06, 2.442238e-06,
  1.175139e-05, 3.691151e-06, 1.192251e-05, 2.40934e-05, 2.5975e-05, 
    4.103653e-05, 1.732338e-05, 8.218995e-06, 3.995734e-06, 5.026162e-06, 
    7.323665e-06, 5.807469e-06, 5.772661e-06, 5.435209e-06, 5.211684e-06,
  5.655333e-05, 1.242758e-05, 9.329158e-06, 2.121704e-05, 2.001946e-05, 
    3.134135e-05, 3.186165e-05, 1.134923e-05, 3.090622e-06, 5.749638e-06, 
    5.798755e-06, 5.501789e-06, 3.62187e-06, 4.103034e-06, 3.811952e-06,
  6.690462e-05, 5.780132e-05, 5.626852e-05, 7.615921e-05, 1.410859e-05, 
    2.209664e-05, 3.510041e-05, 1.424757e-05, 2.222112e-06, 3.793911e-06, 
    5.537982e-06, 4.983045e-06, 3.825311e-06, 4.416143e-06, 3.502703e-06,
  1.432046e-05, 5.163501e-05, 0.0001498168, 0.0001658874, 1.983516e-05, 
    1.890062e-05, 3.125309e-05, 1.511574e-05, 2.882924e-06, 2.910818e-06, 
    4.875233e-06, 4.282541e-06, 3.618538e-06, 3.498356e-06, 2.363524e-06,
  2.554332e-05, 4.988749e-05, 0.000157983, 0.0001328325, 2.876977e-05, 
    2.525601e-05, 2.632966e-05, 1.080665e-05, 2.208554e-06, 2.022356e-06, 
    5.290941e-06, 3.521121e-06, 3.515109e-06, 4.101182e-06, 3.126371e-06,
  0.0001682298, 1.138894e-05, 4.500948e-05, 4.818099e-05, 4.050085e-05, 
    3.371257e-05, 3.074959e-05, 1.734419e-05, 3.016408e-05, 2.949547e-06, 
    5.21077e-06, 2.276214e-06, 3.058688e-06, 2.849264e-06, 2.921363e-06,
  0.0005411984, 4.274567e-05, 2.271147e-05, 4.843434e-05, 4.585278e-05, 
    4.418515e-05, 5.355353e-05, 7.495579e-05, 0.000136147, 2.523256e-06, 
    4.328392e-06, 2.203556e-06, 2.166539e-06, 3.292126e-06, 2.676634e-06,
  0.0008171785, 0.0002148162, 1.80137e-05, 7.705954e-05, 6.277215e-05, 
    5.832952e-05, 9.55531e-05, 0.0002073373, 0.0002204092, 2.208355e-06, 
    3.276079e-06, 3.015104e-06, 4.014778e-06, 4.586247e-06, 3.635882e-06,
  0.0009070293, 0.0003485329, 3.736148e-05, 6.876532e-05, 5.515093e-05, 
    6.850654e-05, 0.0001401062, 0.0002896256, 0.0001818729, 2.06348e-06, 
    2.651072e-06, 2.441127e-06, 3.354949e-06, 4.592476e-06, 4.085224e-06,
  0.0008795607, 0.0004341718, 8.555614e-05, 3.444052e-05, 3.804379e-05, 
    6.539211e-05, 0.0001811052, 0.0003048638, 0.0001007797, 2.495555e-06, 
    3.799463e-06, 2.696945e-06, 3.765009e-06, 3.935198e-06, 4.593855e-06,
  5.188867e-05, 7.806895e-05, 8.707902e-05, 0.0001143957, 0.0001784143, 
    0.0002613964, 0.0001375909, 1.117263e-05, 6.380991e-06, 5.957336e-06, 
    6.307413e-06, 6.647437e-06, 7.300875e-06, 5.82126e-06, 5.797958e-06,
  4.078884e-05, 4.169451e-05, 5.823108e-05, 0.0001164881, 0.0001952116, 
    0.0002951314, 0.0001494289, 1.172927e-05, 6.635241e-06, 5.036821e-06, 
    6.310826e-06, 6.564471e-06, 6.781857e-06, 6.538158e-06, 5.261403e-06,
  1.986549e-05, 2.454085e-05, 3.886993e-05, 0.000117233, 0.0001735018, 
    0.0002382332, 0.0001091619, 5.242763e-06, 6.776349e-06, 5.548964e-06, 
    5.750602e-06, 8.183802e-06, 7.0181e-06, 6.974214e-06, 5.55339e-06,
  7.892367e-06, 1.520523e-05, 3.066226e-05, 0.0001473963, 0.0001327898, 
    0.000178585, 7.978113e-05, 5.907594e-06, 6.392916e-06, 6.920834e-06, 
    6.25767e-06, 8.218011e-06, 5.701031e-06, 5.578715e-06, 4.094687e-06,
  8.330358e-06, 7.785511e-06, 7.874642e-05, 0.0001131683, 8.059031e-05, 
    0.0001149968, 3.807252e-05, 4.797644e-06, 6.882064e-06, 7.122202e-06, 
    7.375288e-06, 6.107131e-06, 4.403105e-06, 5.216834e-06, 4.950423e-06,
  6.939407e-06, 1.058529e-05, 3.877561e-05, 6.484356e-05, 1.841983e-05, 
    2.619923e-05, 6.667925e-06, 5.656299e-06, 7.313579e-06, 8.157983e-06, 
    7.070583e-06, 6.420535e-06, 5.70379e-06, 2.767175e-06, 5.532232e-06,
  8.375826e-06, 1.290617e-05, 2.869872e-05, 5.009282e-05, 7.697026e-06, 
    6.381938e-06, 6.117386e-06, 9.190763e-06, 6.321566e-06, 8.340897e-06, 
    7.406114e-06, 5.648227e-06, 4.59511e-06, 3.355279e-06, 2.151708e-06,
  8.419826e-06, 7.02649e-06, 2.410877e-05, 3.233479e-05, 4.781959e-06, 
    5.672562e-06, 3.37117e-06, 2.030733e-06, 4.550424e-06, 5.870869e-06, 
    9.473469e-06, 5.137406e-06, 4.185798e-06, 1.815739e-06, 1.38202e-06,
  1.186344e-05, 7.134695e-06, 1.313079e-05, 1.439696e-05, 4.945196e-06, 
    3.805791e-06, 4.066756e-06, 1.250402e-06, 3.154875e-06, 5.163259e-06, 
    6.802784e-06, 4.644812e-06, 2.636947e-06, 2.437182e-06, 2.227642e-06,
  1.080931e-05, 6.437925e-06, 6.935456e-06, 6.330379e-06, 3.868021e-06, 
    2.973861e-06, 3.322401e-06, 1.270794e-06, 1.443545e-06, 2.369869e-06, 
    2.01479e-06, 9.669059e-07, 1.347853e-07, 2.128044e-06, 4.083944e-06,
  3.4875e-05, 1.721124e-05, 1.810773e-05, 3.490087e-05, 8.384966e-05, 
    0.0002448643, 0.0004565692, 0.0003394695, 0.000104888, 7.009469e-05, 
    4.957561e-05, 2.53601e-05, 1.243007e-05, 1.289282e-05, 9.683386e-06,
  8.720182e-06, 7.114585e-06, 8.991424e-06, 1.362903e-05, 3.166029e-05, 
    0.0001374742, 0.0003792144, 0.0003551851, 8.316657e-05, 4.833417e-05, 
    3.994603e-05, 2.475958e-05, 1.607966e-05, 1.232206e-05, 9.926894e-06,
  6.770512e-06, 6.806168e-06, 9.624539e-06, 9.520092e-06, 1.042014e-05, 
    1.610178e-05, 0.0001235572, 0.0001022872, 1.663801e-05, 1.599374e-05, 
    2.269922e-05, 1.959587e-05, 1.182529e-05, 7.706081e-06, 6.276454e-06,
  7.886882e-06, 1.252919e-05, 1.076869e-05, 7.941061e-06, 7.624045e-06, 
    1.163725e-05, 6.262363e-05, 2.443454e-05, 1.095649e-05, 1.010045e-05, 
    8.887165e-06, 8.277423e-06, 6.279271e-06, 5.373854e-06, 3.958797e-06,
  9.286708e-06, 8.433709e-06, 1.135868e-05, 9.110078e-06, 6.67079e-06, 
    3.277027e-05, 6.80174e-05, 2.625179e-05, 6.163915e-06, 7.847801e-06, 
    6.935349e-06, 5.930368e-06, 6.436574e-06, 4.440224e-06, 3.935355e-06,
  7.935377e-06, 1.173469e-05, 1.404098e-05, 1.573978e-05, 8.364996e-06, 
    2.214669e-05, 2.01944e-05, 6.335572e-06, 4.569312e-06, 6.593111e-06, 
    5.983163e-06, 5.523315e-06, 3.860123e-06, 3.549355e-06, 3.398354e-06,
  8.939352e-06, 8.487109e-06, 1.032021e-05, 1.547783e-05, 1.896826e-05, 
    9.195807e-06, 8.046823e-06, 7.819272e-06, 3.48514e-06, 8.774118e-06, 
    6.556346e-06, 5.129435e-06, 5.888013e-06, 5.476427e-06, 5.386539e-06,
  4.820854e-06, 6.260171e-06, 9.27566e-06, 5.208527e-06, 7.522675e-06, 
    7.700598e-06, 4.554094e-06, 6.819806e-06, 7.814182e-06, 1.484668e-05, 
    9.80914e-06, 7.022798e-06, 6.713368e-06, 4.040347e-06, 2.444362e-06,
  1.532318e-06, 1.130714e-05, 7.334916e-06, 4.174193e-06, 2.704172e-06, 
    6.142151e-07, 2.060089e-06, 1.341025e-06, 3.831534e-06, 4.79113e-06, 
    5.579691e-06, 8.256682e-06, 6.909086e-06, 4.94622e-06, 2.621051e-06,
  1.265888e-05, 5.1279e-06, 3.369337e-06, 4.248217e-06, 2.40024e-06, 
    2.002223e-06, 1.190258e-06, 1.924928e-06, 3.886924e-06, 5.543754e-06, 
    7.750625e-06, 1.121383e-05, 5.370522e-06, 3.964874e-06, 3.27604e-06,
  1.382802e-05, 1.236901e-05, 8.366193e-06, 7.87834e-06, 5.681739e-06, 
    1.142938e-05, 4.039694e-05, 6.435122e-05, 6.64579e-05, 4.610397e-05, 
    4.249185e-05, 4.869119e-05, 5.785904e-05, 6.285181e-05, 7.774575e-05,
  8.555197e-06, 8.236195e-06, 5.349275e-06, 7.057274e-06, 6.86999e-06, 
    5.961584e-06, 6.665349e-06, 3.191081e-05, 4.483375e-05, 3.938395e-05, 
    3.736456e-05, 4.384031e-05, 5.165859e-05, 6.413225e-05, 7.640828e-05,
  4.053928e-06, 4.404036e-06, 6.218506e-06, 5.459728e-06, 6.356355e-06, 
    3.502132e-06, 4.377388e-06, 3.582388e-06, 1.800287e-05, 2.496766e-05, 
    3.027269e-05, 3.808559e-05, 4.699449e-05, 5.337487e-05, 6.196883e-05,
  7.044378e-06, 7.319228e-06, 5.9911e-06, 3.393452e-06, 3.456856e-06, 
    3.212896e-06, 3.834027e-06, 2.853007e-06, 3.661926e-06, 7.301888e-06, 
    1.756168e-05, 2.929733e-05, 3.831906e-05, 4.43744e-05, 5.508477e-05,
  6.820991e-06, 8.542271e-06, 7.563744e-06, 4.273364e-06, 4.352755e-06, 
    2.590315e-06, 1.677556e-06, 2.90502e-06, 3.889207e-06, 2.675911e-06, 
    5.324209e-06, 1.930993e-05, 3.782039e-05, 4.191672e-05, 5.054734e-05,
  1.013262e-05, 8.388368e-06, 1.11537e-05, 6.979493e-06, 5.324431e-06, 
    4.347104e-06, 2.394003e-06, 2.723948e-06, 3.718204e-06, 3.058178e-06, 
    3.232259e-06, 1.026329e-05, 3.033343e-05, 4.349561e-05, 5.109488e-05,
  1.665131e-05, 1.685979e-05, 1.233434e-05, 9.782471e-06, 6.954013e-06, 
    4.90108e-06, 4.831954e-06, 5.367386e-06, 4.561612e-06, 3.753732e-06, 
    3.16004e-06, 4.133881e-06, 2.068374e-05, 3.861948e-05, 5.115966e-05,
  3.801677e-05, 2.704975e-05, 2.241317e-05, 1.586197e-05, 8.66911e-06, 
    5.978717e-06, 9.232399e-06, 1.147507e-05, 9.940966e-06, 6.912742e-06, 
    6.286625e-06, 3.85615e-06, 6.000546e-06, 2.514166e-05, 4.233161e-05,
  0.000177534, 8.50397e-05, 2.441574e-05, 2.857481e-05, 2.048155e-05, 
    9.467726e-06, 6.345399e-06, 1.260599e-05, 1.29497e-05, 1.037119e-05, 
    1.128096e-05, 8.223131e-06, 3.51167e-06, 2.728955e-06, 1.991496e-05,
  0.0004188569, 0.0001992183, 3.950471e-05, 2.666295e-05, 3.423851e-05, 
    1.716946e-05, 6.503231e-06, 1.263973e-05, 1.405459e-05, 1.516418e-05, 
    1.454025e-05, 1.196011e-05, 7.168907e-06, 6.786016e-06, 4.552948e-06,
  2.238051e-05, 3.952968e-05, 6.744535e-05, 0.0001138854, 0.0002116585, 
    0.0002288053, 8.086555e-05, 3.374216e-05, 1.849589e-05, 1.324883e-05, 
    8.174258e-06, 2.863236e-05, 3.088579e-05, 1.743011e-05, 1.068475e-05,
  1.583445e-05, 3.019879e-05, 6.74148e-05, 0.0001225313, 0.0002582933, 
    0.0002804811, 0.0001521578, 7.771566e-05, 4.503673e-05, 2.757523e-05, 
    1.706287e-05, 1.92917e-05, 1.913649e-05, 1.381503e-05, 1.17473e-05,
  4.159671e-06, 1.208849e-05, 5.594302e-05, 0.0001286958, 0.0003052539, 
    0.0002896156, 0.0001562988, 0.0001115631, 8.295447e-05, 5.001149e-05, 
    2.714755e-05, 1.440887e-05, 1.000333e-05, 1.033454e-05, 1.148361e-05,
  4.66355e-06, 1.75146e-05, 6.70808e-05, 0.000148492, 0.0003006853, 
    0.0002675581, 0.0001228522, 9.961784e-05, 9.540995e-05, 7.292101e-05, 
    4.385184e-05, 1.790537e-05, 9.68836e-06, 1.029537e-05, 1.490018e-05,
  8.575169e-06, 3.359815e-05, 9.408556e-05, 0.0001657294, 0.0002836569, 
    0.0002392259, 9.792742e-05, 8.997736e-05, 9.410638e-05, 7.980634e-05, 
    5.362722e-05, 3.325686e-05, 1.541396e-05, 1.23381e-05, 1.567193e-05,
  1.320406e-05, 5.243837e-05, 0.0001023542, 0.0001799536, 0.0002499995, 
    0.0002131267, 8.651579e-05, 8.628717e-05, 9.794814e-05, 8.042022e-05, 
    6.456506e-05, 4.846886e-05, 3.337922e-05, 1.79977e-05, 1.663902e-05,
  3.745324e-05, 7.616987e-05, 0.0001029855, 0.0001655258, 0.0002126847, 
    0.0001867034, 8.381482e-05, 8.926367e-05, 0.000101977, 9.022582e-05, 
    7.079197e-05, 6.002088e-05, 5.47588e-05, 3.147677e-05, 2.179706e-05,
  7.082289e-05, 9.397927e-05, 0.0001079037, 0.0001567464, 0.0001825406, 
    0.0001503638, 8.351389e-05, 9.605273e-05, 0.0001088646, 9.645796e-05, 
    7.490171e-05, 6.519913e-05, 7.4737e-05, 6.076949e-05, 4.141374e-05,
  5.995797e-05, 9.225502e-05, 0.0001232429, 0.0001494135, 0.000150471, 
    0.0001177276, 8.236966e-05, 9.876761e-05, 0.0001094395, 9.233574e-05, 
    7.554371e-05, 6.669819e-05, 7.772486e-05, 8.491453e-05, 6.683331e-05,
  1.613426e-05, 6.101284e-05, 0.000105572, 0.0001234821, 0.0001104632, 
    9.216123e-05, 9.053572e-05, 0.0001102065, 0.0001085643, 8.610157e-05, 
    6.354538e-05, 6.590785e-05, 7.345112e-05, 8.274538e-05, 8.611353e-05,
  1.4299e-05, 2.462305e-05, 3.598149e-05, 3.838256e-05, 1.35954e-05, 
    1.266771e-05, 8.643312e-06, 1.599267e-05, 7.903963e-06, 1.246713e-05, 
    8.339428e-06, 7.049023e-06, 4.899558e-06, 4.48775e-06, 6.255391e-06,
  2.577146e-05, 3.545755e-05, 4.546741e-05, 6.225159e-05, 4.065031e-05, 
    1.672558e-05, 1.3887e-05, 1.197572e-05, 1.340041e-05, 1.089473e-05, 
    1.817851e-05, 5.536543e-06, 5.319901e-06, 5.966729e-06, 6.044168e-06,
  3.299478e-05, 4.625417e-05, 5.771983e-05, 8.103702e-05, 6.297058e-05, 
    2.450599e-05, 1.374705e-05, 8.516831e-06, 9.701194e-06, 7.415802e-06, 
    5.947919e-06, 4.815405e-06, 6.134627e-06, 7.139807e-06, 7.449421e-06,
  3.590695e-05, 4.876876e-05, 6.376421e-05, 8.853739e-05, 8.888853e-05, 
    3.361274e-05, 9.190448e-06, 7.633845e-06, 5.589394e-06, 3.88435e-06, 
    5.313283e-06, 5.695907e-06, 6.730169e-06, 8.776175e-06, 8.685374e-06,
  3.911804e-05, 5.118356e-05, 6.167191e-05, 9.799281e-05, 0.0001088467, 
    4.20429e-05, 6.850071e-06, 6.949593e-06, 4.460878e-06, 3.978673e-06, 
    6.426457e-06, 5.048287e-06, 6.977657e-06, 5.63499e-06, 7.497392e-06,
  4.616957e-05, 5.54994e-05, 7.108803e-05, 0.0001072491, 0.0001301941, 
    6.240995e-05, 9.63154e-06, 5.826103e-06, 4.831847e-06, 3.411506e-06, 
    4.321167e-06, 4.91529e-06, 6.875458e-06, 5.273663e-06, 5.517252e-06,
  5.189123e-05, 6.001658e-05, 7.64478e-05, 0.0001456858, 0.0001661217, 
    9.070225e-05, 1.396092e-05, 5.453655e-06, 6.290789e-06, 4.065198e-06, 
    5.236217e-06, 5.600522e-06, 4.677976e-06, 4.63829e-06, 4.273461e-06,
  6.765557e-05, 7.133884e-05, 8.032729e-05, 0.0002199522, 0.0002206147, 
    0.0001212474, 1.153695e-05, 4.459136e-06, 6.74266e-06, 4.810487e-06, 
    4.183718e-06, 5.712887e-06, 5.021976e-06, 4.003791e-06, 4.297948e-06,
  8.949402e-05, 9.727755e-05, 0.0001347727, 0.0003002534, 0.0002764162, 
    0.0001514642, 7.673638e-06, 5.096445e-06, 7.916324e-06, 6.338229e-06, 
    5.000769e-06, 4.846128e-06, 5.459969e-06, 4.001232e-06, 3.256201e-06,
  0.0001020935, 0.0001509268, 0.000233802, 0.0003649025, 0.0003275612, 
    0.0001642328, 6.212964e-06, 6.003954e-06, 8.542289e-06, 7.639709e-06, 
    4.906523e-06, 6.051415e-06, 7.953663e-06, 4.594712e-06, 3.518469e-06,
  3.612816e-06, 8.682323e-07, 4.714305e-07, 1.112646e-06, 4.716977e-07, 
    1.51218e-06, 1.562441e-06, 1.984297e-06, 2.478143e-06, 1.447129e-06, 
    3.469758e-06, 7.795476e-06, 7.273213e-06, 7.751412e-06, 1.010791e-05,
  3.201508e-06, 2.858134e-06, 2.356544e-06, 8.520452e-07, 7.416119e-07, 
    2.039099e-06, 2.331153e-06, 2.450341e-06, 2.247307e-06, 1.813674e-06, 
    4.4683e-06, 5.792123e-06, 5.016726e-06, 6.078238e-06, 8.366615e-06,
  3.824184e-06, 3.358252e-06, 2.301973e-06, 1.407486e-06, 2.706295e-07, 
    1.639202e-06, 3.534283e-06, 2.667573e-06, 2.896696e-06, 3.486442e-06, 
    6.298105e-06, 6.627772e-06, 5.778724e-06, 9.847513e-06, 1.596355e-05,
  1.887436e-06, 2.743627e-06, 1.483397e-06, 1.869755e-06, 1.40957e-06, 
    1.758025e-06, 3.740676e-06, 3.91367e-06, 4.031906e-06, 5.8036e-06, 
    6.78137e-06, 6.940524e-06, 8.218643e-06, 9.830464e-06, 1.486413e-05,
  3.036141e-06, 5.679284e-06, 1.923675e-06, 3.802631e-06, 8.962096e-07, 
    4.060632e-06, 3.462123e-06, 4.352909e-06, 4.3287e-06, 5.881439e-06, 
    7.44326e-06, 6.364291e-06, 7.75019e-06, 1.229658e-05, 1.041632e-05,
  6.730621e-06, 7.448676e-06, 3.860958e-06, 3.50107e-06, 2.399573e-06, 
    1.452495e-06, 3.745705e-06, 5.371639e-06, 6.083616e-06, 7.091033e-06, 
    6.813956e-06, 5.897147e-06, 1.273421e-05, 7.30367e-06, 6.93501e-06,
  6.520738e-06, 5.226591e-06, 4.313925e-06, 3.649554e-06, 1.200976e-06, 
    9.85473e-07, 4.068846e-06, 5.04349e-06, 6.313896e-06, 8.404973e-06, 
    5.820538e-06, 8.007938e-06, 7.583834e-06, 4.571929e-06, 3.285074e-06,
  2.842938e-06, 4.817127e-06, 5.261822e-06, 2.243022e-06, 1.231986e-06, 
    1.757221e-06, 6.564681e-06, 5.884494e-06, 6.437625e-06, 7.734724e-06, 
    5.213388e-06, 5.053708e-06, 6.839107e-06, 4.442298e-06, 2.875918e-06,
  4.879413e-06, 4.455949e-06, 4.585931e-06, 3.940105e-06, 3.736477e-06, 
    3.505646e-06, 6.078657e-06, 7.498027e-06, 7.270449e-06, 7.572183e-06, 
    8.077309e-06, 4.117393e-06, 5.057486e-06, 3.01716e-06, 1.767434e-06,
  3.636759e-06, 4.232108e-06, 3.432286e-06, 1.698298e-06, 9.963109e-07, 
    3.880756e-06, 4.928881e-06, 6.106574e-06, 8.815068e-06, 7.855057e-06, 
    7.389358e-06, 5.66437e-06, 3.002498e-06, 2.88083e-06, 3.242673e-06,
  8.929136e-06, 1.469001e-05, 1.783233e-05, 1.4683e-05, 9.365344e-06, 
    6.425469e-06, 4.166746e-06, 4.05042e-06, 6.857954e-06, 7.168221e-06, 
    8.356321e-06, 1.000684e-05, 1.007969e-05, 5.479802e-06, 9.182595e-06,
  8.721144e-06, 1.105473e-05, 9.76749e-06, 8.439391e-06, 7.725589e-06, 
    5.543741e-06, 3.430079e-06, 2.946174e-06, 7.730086e-06, 7.391576e-06, 
    8.305091e-06, 7.430536e-06, 7.682769e-06, 6.096309e-06, 1.041769e-05,
  9.607009e-06, 9.133903e-06, 6.083686e-06, 5.479593e-06, 6.823843e-06, 
    5.215041e-06, 3.030279e-06, 4.331528e-06, 6.724349e-06, 7.571524e-06, 
    8.449354e-06, 5.623389e-06, 7.028926e-06, 6.881418e-06, 6.816821e-06,
  7.572391e-06, 6.072849e-06, 5.471787e-06, 4.263839e-06, 4.320882e-06, 
    3.609716e-06, 5.429605e-06, 4.861162e-06, 5.627123e-06, 4.878682e-06, 
    1.050499e-05, 9.092266e-06, 5.813078e-06, 3.056784e-06, 7.328988e-06,
  6.628356e-06, 5.462904e-06, 3.981319e-06, 4.777693e-06, 3.105877e-06, 
    3.322814e-06, 4.10617e-06, 4.345356e-06, 4.700379e-06, 3.920842e-06, 
    6.741458e-06, 9.063836e-06, 2.578765e-06, 2.399724e-06, 2.647358e-06,
  6.057376e-06, 4.197313e-06, 1.601235e-06, 2.328699e-06, 3.393554e-06, 
    2.900322e-06, 3.35284e-06, 3.617682e-06, 2.474152e-06, 6.020499e-06, 
    6.371406e-06, 4.337753e-06, 4.827112e-06, 1.577571e-06, 6.296429e-07,
  4.788059e-06, 2.341993e-06, 3.581091e-06, 2.562515e-06, 1.947089e-06, 
    1.525883e-06, 2.156508e-06, 2.707079e-06, 2.242856e-06, 3.742957e-06, 
    2.458158e-06, 3.025918e-06, 2.046223e-06, 3.195206e-06, 9.914352e-07,
  2.807343e-06, 2.148206e-06, 3.020064e-06, 1.985033e-06, 1.741541e-06, 
    3.073798e-06, 1.981691e-06, 2.18567e-06, 2.367727e-06, 2.030708e-06, 
    1.777902e-07, 9.411428e-07, 3.504269e-06, 2.785596e-06, 7.539833e-07,
  1.077121e-06, 1.362468e-06, 1.888346e-06, 2.329963e-06, 2.021668e-06, 
    4.71432e-06, 4.492953e-06, 2.935516e-06, 1.643162e-06, 1.990579e-06, 
    2.330563e-06, 8.906246e-07, 2.065039e-06, 2.272686e-06, 8.169466e-07,
  2.355629e-06, 1.364719e-06, 1.520762e-06, 1.641947e-06, 3.65165e-06, 
    5.493664e-06, 3.228243e-06, 2.509187e-06, 1.072612e-06, 5.322004e-06, 
    3.496385e-06, 3.942979e-06, 3.011556e-06, 1.17897e-06, 4.811619e-07,
  0.0002793806, 0.000216931, 0.0001725806, 0.0001011204, 3.025469e-05, 
    1.463363e-05, 1.460608e-05, 1.315085e-05, 1.346558e-05, 9.502747e-06, 
    1.419573e-05, 1.358078e-05, 3.015095e-05, 3.160854e-05, 2.518645e-05,
  0.0002616494, 0.000202302, 0.0001719139, 8.718274e-05, 2.698902e-05, 
    1.638442e-05, 1.468624e-05, 1.401147e-05, 1.234062e-05, 1.425641e-05, 
    1.790329e-05, 2.115863e-05, 2.540769e-05, 3.833183e-05, 4.241118e-05,
  0.0002216075, 0.0001719589, 0.0001096601, 5.867532e-05, 2.184528e-05, 
    1.658017e-05, 1.599299e-05, 1.390565e-05, 1.37553e-05, 1.190559e-05, 
    1.613616e-05, 2.117383e-05, 3.588082e-05, 3.609502e-05, 3.523493e-05,
  0.0002341247, 0.0001407582, 8.613718e-05, 4.197927e-05, 1.966786e-05, 
    1.883766e-05, 1.613381e-05, 1.339568e-05, 1.967062e-05, 1.944051e-05, 
    1.750294e-05, 2.198594e-05, 3.041122e-05, 4.69816e-05, 5.019653e-05,
  0.0002241854, 0.0001178256, 7.094524e-05, 3.474257e-05, 2.420745e-05, 
    1.889989e-05, 1.778384e-05, 1.862233e-05, 2.879033e-05, 2.142744e-05, 
    2.050958e-05, 2.813561e-05, 4.794343e-05, 5.080634e-05, 4.908415e-05,
  0.0002162783, 0.0001057627, 5.333691e-05, 3.450827e-05, 2.384221e-05, 
    1.749603e-05, 1.522018e-05, 2.301809e-05, 2.381796e-05, 2.362702e-05, 
    2.339601e-05, 3.052699e-05, 6.715261e-05, 4.875585e-05, 5.509932e-05,
  0.0002054891, 9.582244e-05, 3.957972e-05, 3.888408e-05, 2.594057e-05, 
    1.597906e-05, 1.897929e-05, 2.52924e-05, 2.61153e-05, 2.007214e-05, 
    2.741378e-05, 5.328135e-05, 3.808274e-05, 4.77813e-05, 5.718929e-05,
  0.0001988764, 9.481666e-05, 4.980004e-05, 3.523393e-05, 2.515638e-05, 
    1.908192e-05, 2.213823e-05, 2.265736e-05, 3.060044e-05, 3.336142e-05, 
    2.795723e-05, 7.504794e-05, 4.725001e-05, 5.689035e-05, 8.086428e-05,
  0.0001713495, 8.691507e-05, 5.172929e-05, 3.911234e-05, 2.292708e-05, 
    2.167415e-05, 2.496637e-05, 2.337365e-05, 3.267375e-05, 2.307551e-05, 
    2.847859e-05, 4.095133e-05, 6.318332e-05, 7.583008e-05, 8.883636e-05,
  0.000149935, 8.036318e-05, 5.674156e-05, 3.109899e-05, 2.461587e-05, 
    1.762114e-05, 1.794919e-05, 2.328676e-05, 2.845435e-05, 4.3299e-05, 
    4.020739e-05, 5.647274e-05, 8.569154e-05, 8.773094e-05, 0.0001046503,
  3.020485e-06, 2.285172e-06, 1.420956e-06, 1.705822e-07, 2.667046e-08, 
    3.676771e-08, 1.427435e-07, 2.504893e-07, 5.862867e-07, 1.02275e-06, 
    3.055447e-07, 2.381117e-07, 1.553975e-07, 6.056692e-08, 1.404137e-07,
  5.396853e-06, 3.030221e-06, 6.054353e-07, 5.831912e-08, 6.427089e-08, 
    1.59595e-07, 2.770416e-07, 3.38097e-07, 4.868722e-07, 1.955814e-07, 
    8.657451e-08, 1.024922e-07, 1.411277e-07, 4.518794e-07, 8.474604e-07,
  9.137295e-06, 2.880503e-06, 5.28607e-07, 9.694868e-08, 1.754272e-07, 
    2.084717e-07, 4.387222e-08, 9.282762e-08, 2.161938e-07, 1.739921e-07, 
    1.625992e-07, 2.436287e-07, 4.976652e-07, 1.881401e-06, 4.050961e-06,
  9.700873e-06, 4.825655e-06, 4.21291e-07, 7.299207e-08, 1.015439e-07, 
    8.324887e-08, 6.647834e-08, 9.177064e-08, 2.128582e-07, 1.197603e-07, 
    3.704778e-07, 4.870028e-07, 1.678524e-06, 2.969301e-06, 3.637704e-06,
  9.479992e-06, 6.438766e-06, 9.131813e-07, 3.683e-08, 5.018456e-08, 
    6.509065e-08, 8.930687e-08, 1.109241e-08, 6.780467e-08, 2.33999e-07, 
    8.904731e-07, 1.786613e-06, 2.756119e-06, 5.143247e-06, 3.134125e-06,
  1.337506e-05, 7.42413e-06, 1.110776e-07, 6.945394e-09, 9.201252e-09, 
    6.470371e-08, 5.281187e-08, 7.323576e-09, 9.99357e-08, 5.44959e-07, 
    1.698038e-06, 2.548379e-06, 2.710726e-06, 2.892359e-06, 3.134004e-06,
  1.963826e-05, 1.23449e-05, 4.335375e-07, 2.001954e-09, 4.053818e-09, 
    8.186717e-09, 4.037874e-09, 6.631499e-08, 1.677202e-07, 9.182356e-07, 
    1.914631e-06, 2.747432e-06, 1.507947e-06, 3.829515e-06, 3.809325e-06,
  2.356745e-05, 8.699652e-06, 1.856106e-07, 4.192036e-09, 2.523655e-09, 
    3.767294e-10, 1.778388e-08, 7.771136e-08, 4.621471e-07, 9.978824e-07, 
    1.863302e-06, 2.574183e-06, 2.544341e-06, 2.174112e-06, 2.597857e-06,
  3.132191e-05, 1.202541e-05, 9.192288e-06, 3.526604e-09, 3.668256e-09, 
    5.238604e-08, 2.090584e-08, 3.205402e-07, 1.000952e-06, 1.883184e-06, 
    1.988163e-06, 1.958036e-06, 1.949234e-06, 2.345575e-06, 2.285175e-06,
  2.859751e-05, 1.563477e-05, 4.07388e-06, 1.930182e-09, 7.921037e-08, 
    1.686394e-07, 3.822801e-07, 6.925093e-07, 1.422615e-06, 1.148503e-06, 
    1.543824e-06, 1.939182e-06, 2.239753e-06, 3.332221e-06, 4.582775e-06,
  7.526157e-06, 5.950816e-06, 1.770164e-06, 7.948156e-08, 4.852561e-08, 
    1.48911e-07, 3.596075e-08, 3.327677e-07, 1.788916e-06, 2.919743e-06, 
    3.693408e-06, 3.911921e-06, 3.046807e-06, 2.196348e-06, 2.884889e-06,
  5.169472e-07, 8.345567e-08, 6.096408e-08, 3.565896e-09, 4.713296e-08, 
    4.83242e-08, 3.420201e-07, 6.995501e-07, 2.353834e-06, 2.420196e-06, 
    3.078115e-06, 2.263573e-06, 3.810555e-06, 3.35687e-06, 3.847768e-06,
  3.631205e-08, 7.954124e-09, 2.289752e-09, 8.669032e-09, 4.089695e-08, 
    1.135378e-07, 2.500808e-06, 2.468634e-06, 3.138551e-06, 3.48989e-06, 
    2.030823e-06, 4.665486e-06, 4.053237e-06, 3.848435e-06, 3.652511e-06,
  2.36969e-09, 7.908608e-09, 3.241911e-08, 1.555749e-08, 1.019947e-07, 
    1.624309e-06, 1.848754e-06, 1.783006e-06, 4.07902e-06, 1.806393e-06, 
    3.364327e-06, 3.466591e-06, 4.641834e-06, 4.012521e-06, 4.86201e-06,
  2.651693e-09, 8.880999e-08, 1.884495e-07, 7.230403e-08, 2.770528e-07, 
    1.742979e-06, 3.133233e-06, 1.697922e-06, 2.114987e-06, 3.694772e-06, 
    3.991157e-06, 4.146611e-06, 4.122841e-06, 5.226846e-06, 8.889277e-06,
  6.089021e-08, 4.401876e-07, 3.066782e-07, 4.944099e-07, 1.676644e-06, 
    2.260452e-06, 2.282371e-06, 2.862733e-06, 2.911062e-06, 3.207846e-06, 
    3.025605e-06, 3.694125e-06, 3.112978e-06, 4.159586e-06, 1.060142e-05,
  1.853141e-08, 1.575452e-07, 2.50632e-07, 1.138941e-06, 1.655442e-06, 
    3.155463e-06, 5.554028e-06, 2.386375e-06, 4.307522e-06, 3.09542e-06, 
    3.805376e-06, 4.651685e-06, 6.245611e-06, 8.081336e-06, 1.137019e-05,
  6.116311e-08, 2.936984e-07, 1.728283e-06, 3.055667e-06, 3.217587e-06, 
    2.94488e-06, 2.28439e-06, 2.744119e-06, 4.592593e-06, 4.65775e-06, 
    5.094488e-06, 3.724464e-06, 7.903147e-06, 8.876492e-06, 8.364565e-06,
  1.845543e-07, 1.348243e-06, 3.0226e-06, 3.84395e-06, 4.357146e-06, 
    4.362699e-06, 3.485054e-06, 3.769307e-06, 4.854683e-06, 7.937277e-06, 
    6.31843e-06, 4.899315e-06, 5.397673e-06, 5.860613e-06, 5.524694e-06,
  1.464548e-06, 3.007715e-06, 4.375654e-06, 5.431791e-06, 6.057329e-06, 
    6.254273e-06, 3.557832e-06, 3.034857e-06, 5.498438e-06, 6.291666e-06, 
    3.373916e-06, 4.135826e-06, 5.131839e-06, 5.815642e-06, 4.938436e-06,
  0.0001879227, 0.0004250692, 0.0007606511, 0.0007235756, 0.0002703401, 
    8.182201e-06, 4.295786e-06, 2.897267e-06, 3.034739e-06, 6.36768e-06, 
    7.380968e-06, 6.384991e-06, 5.798541e-06, 3.723568e-06, 4.841994e-06,
  0.0001470016, 0.0003735845, 0.0006926416, 0.0007405134, 0.0003106031, 
    1.167706e-05, 3.47774e-06, 3.495265e-06, 2.614281e-06, 3.786373e-06, 
    3.836788e-06, 3.708367e-06, 4.656812e-06, 5.875333e-06, 4.992838e-06,
  0.0001209628, 0.0003548569, 0.0006142655, 0.0006446177, 0.0002465771, 
    1.140817e-05, 4.142865e-06, 3.503802e-06, 3.014185e-06, 4.193484e-06, 
    5.348094e-06, 3.354969e-06, 5.432081e-06, 5.584692e-06, 5.092073e-06,
  8.407039e-05, 0.0003387966, 0.000552003, 0.0005279945, 0.0001897707, 
    1.5349e-05, 3.768422e-06, 4.657173e-06, 6.008855e-06, 4.549961e-06, 
    4.221613e-06, 2.758266e-06, 5.277911e-06, 5.316586e-06, 5.084925e-06,
  7.317311e-05, 0.0002812065, 0.0004131375, 0.0003460985, 0.0001130335, 
    1.397342e-05, 5.001843e-06, 4.131188e-06, 3.408969e-06, 2.729255e-06, 
    2.190564e-06, 3.826229e-06, 4.408368e-06, 4.372645e-06, 7.509492e-06,
  6.497723e-05, 0.0002178228, 0.0002857491, 0.0001857636, 4.788293e-05, 
    6.13426e-06, 2.519428e-06, 2.605648e-06, 4.660328e-06, 3.745801e-06, 
    7.812411e-06, 8.960632e-06, 5.224391e-06, 4.865439e-06, 6.964389e-06,
  6.028646e-05, 0.0001326784, 0.0001274544, 7.337228e-05, 1.196617e-05, 
    2.331745e-06, 2.322944e-06, 2.328641e-06, 4.079702e-06, 4.143426e-06, 
    4.854715e-06, 8.043902e-06, 8.025277e-06, 9.085443e-06, 8.266008e-06,
  2.816804e-05, 4.022611e-05, 2.631627e-05, 7.694717e-06, 5.082421e-06, 
    2.456562e-06, 2.524218e-06, 3.434921e-06, 5.636159e-06, 6.486725e-06, 
    6.880546e-06, 1.105149e-05, 1.087277e-05, 9.596673e-06, 1.188665e-05,
  5.068791e-06, 5.917759e-06, 3.32043e-06, 2.960435e-06, 4.75212e-06, 
    4.112866e-06, 3.412169e-06, 5.387454e-06, 7.982037e-06, 6.720225e-06, 
    9.489858e-06, 7.060094e-06, 7.787638e-06, 7.674847e-06, 1.274141e-05,
  3.252822e-06, 3.281607e-06, 3.686522e-06, 2.632967e-06, 4.944241e-06, 
    5.50168e-06, 3.518964e-06, 5.464574e-06, 5.203256e-06, 1.279687e-05, 
    9.718894e-06, 1.098384e-05, 7.083333e-06, 1.041895e-05, 1.051545e-05,
  1.323472e-05, 5.921467e-06, 2.114866e-05, 1.597131e-05, 6.443264e-06, 
    4.923374e-06, 4.803876e-06, 4.074246e-06, 3.39606e-06, 3.436882e-06, 
    5.513451e-06, 5.175645e-06, 2.541087e-06, 2.029796e-06, 3.679753e-06,
  1.979786e-05, 5.373839e-05, 9.764246e-05, 5.281934e-05, 1.034867e-05, 
    5.76254e-06, 3.103038e-06, 2.947589e-06, 3.412903e-06, 3.854131e-06, 
    4.497836e-06, 3.259552e-06, 3.187982e-06, 1.886548e-06, 1.359358e-06,
  3.5042e-05, 0.000173705, 0.0002482501, 0.0001405323, 1.226505e-05, 
    5.51009e-06, 4.821429e-06, 3.623683e-06, 5.223505e-06, 4.407116e-06, 
    6.244241e-06, 5.73239e-06, 2.876818e-06, 2.961271e-06, 4.665539e-06,
  4.906364e-05, 0.0003187617, 0.0004472871, 0.0002424533, 1.993808e-05, 
    5.264267e-06, 2.930421e-06, 4.269863e-06, 5.05938e-06, 4.892095e-06, 
    5.484692e-06, 6.352589e-06, 4.695185e-06, 8.429846e-06, 7.157135e-06,
  7.682318e-05, 0.0005025491, 0.0006893643, 0.0002951788, 2.032123e-05, 
    4.796542e-06, 3.142838e-06, 5.024923e-06, 5.490665e-06, 4.397346e-06, 
    6.387795e-06, 8.387751e-06, 7.809433e-06, 9.432498e-06, 1.095677e-05,
  0.0002767423, 0.0007556276, 0.0008989692, 0.0002861475, 2.121425e-05, 
    5.031489e-06, 3.852033e-06, 5.038275e-06, 5.285518e-06, 6.596275e-06, 
    4.251585e-06, 7.747677e-06, 6.906139e-06, 8.394886e-06, 7.34566e-06,
  0.000508938, 0.0009618512, 0.0008649635, 0.0002101549, 1.961941e-05, 
    5.76266e-06, 3.710919e-06, 5.609298e-06, 5.456963e-06, 6.18009e-06, 
    7.983642e-06, 9.157301e-06, 7.833044e-06, 7.96894e-06, 5.932984e-06,
  0.0007154686, 0.001061552, 0.0007182508, 0.0001066041, 1.334973e-05, 
    2.949325e-06, 3.936126e-06, 5.108473e-06, 5.38618e-06, 6.223909e-06, 
    5.396456e-06, 1.135169e-05, 1.070938e-05, 6.694552e-06, 4.873149e-06,
  0.0008671237, 0.0009760448, 0.0004307121, 3.936512e-05, 4.786664e-06, 
    3.582385e-06, 6.012958e-06, 7.398167e-06, 6.09964e-06, 7.103515e-06, 
    9.7688e-06, 9.653462e-06, 5.367114e-06, 6.22606e-06, 8.280087e-06,
  0.0008930493, 0.0007006621, 0.0001491174, 2.025305e-05, 3.891358e-06, 
    5.106284e-06, 5.912795e-06, 5.059143e-06, 6.052644e-06, 7.53699e-06, 
    9.498514e-06, 9.618037e-06, 8.126143e-06, 9.463422e-06, 8.496986e-06,
  6.000157e-06, 5.020523e-06, 6.886794e-06, 6.483046e-06, 5.853655e-06, 
    3.480311e-06, 5.254947e-06, 3.134914e-06, 3.843444e-06, 4.641217e-06, 
    2.779454e-06, 4.166791e-06, 5.560161e-06, 8.003942e-06, 8.751155e-06,
  1.284828e-06, 3.266174e-06, 6.523261e-06, 5.049314e-06, 5.041262e-06, 
    4.354751e-06, 3.452405e-06, 3.530026e-06, 2.623847e-06, 4.235738e-06, 
    6.883158e-06, 1.035592e-05, 1.304208e-05, 1.511952e-05, 1.054658e-05,
  2.015051e-06, 5.151807e-06, 5.155797e-06, 3.487015e-06, 3.473186e-06, 
    4.363273e-06, 3.200302e-06, 3.876699e-06, 4.112788e-06, 7.16099e-06, 
    8.665505e-06, 7.351565e-06, 6.648166e-06, 4.557521e-06, 3.217137e-06,
  6.017252e-06, 4.827887e-06, 3.733918e-06, 4.153361e-06, 3.918683e-06, 
    4.433116e-06, 4.507611e-06, 4.818647e-06, 7.655555e-06, 7.491071e-06, 
    5.264781e-06, 2.602916e-06, 3.918668e-06, 1.748578e-06, 2.183898e-07,
  6.152287e-06, 4.48004e-06, 2.981532e-06, 1.955981e-06, 3.719276e-06, 
    5.160917e-06, 6.109347e-06, 7.900783e-06, 4.568401e-06, 6.487972e-06, 
    5.39858e-06, 3.143429e-06, 3.689703e-06, 4.076595e-07, 4.525252e-07,
  5.14703e-06, 2.873644e-06, 3.225668e-06, 4.327709e-06, 5.961998e-06, 
    5.891472e-06, 7.381922e-06, 5.341821e-06, 2.127008e-06, 7.201333e-06, 
    7.870194e-06, 7.686634e-06, 5.353721e-06, 1.418039e-06, 1.624057e-06,
  4.596528e-06, 3.545687e-06, 4.428216e-06, 4.682101e-06, 5.262222e-06, 
    4.937011e-06, 8.713609e-06, 3.502266e-06, 9.744908e-06, 8.557507e-06, 
    1.070939e-05, 9.470993e-06, 6.558401e-06, 4.218297e-06, 7.597859e-07,
  4.260032e-06, 3.609076e-06, 4.008823e-06, 3.835331e-06, 5.470766e-06, 
    5.062095e-06, 5.693495e-06, 6.439177e-06, 7.815349e-06, 1.118526e-05, 
    1.170143e-05, 8.949525e-06, 6.282109e-06, 4.487536e-06, 1.456697e-06,
  4.903884e-06, 5.094515e-06, 4.968222e-06, 4.921761e-06, 6.052844e-06, 
    8.715525e-06, 6.357134e-06, 8.458948e-06, 1.010225e-05, 9.513638e-06, 
    8.760018e-06, 8.272086e-06, 7.931623e-06, 6.871255e-06, 4.160199e-06,
  5.017933e-06, 5.83476e-06, 6.069613e-06, 5.533831e-06, 6.120113e-06, 
    4.259983e-06, 4.985208e-06, 6.474045e-06, 7.968481e-06, 7.357276e-06, 
    8.517754e-06, 6.779621e-06, 5.948331e-06, 5.291606e-06, 2.503082e-06,
  9.413567e-06, 8.160534e-06, 7.56737e-06, 3.816133e-06, 4.050326e-06, 
    3.456332e-06, 2.555204e-06, 2.97914e-06, 3.69435e-06, 5.071694e-06, 
    5.473758e-06, 4.854621e-06, 5.106773e-06, 5.67032e-06, 5.906868e-06,
  5.203347e-06, 5.533206e-06, 6.498707e-06, 4.703501e-06, 6.123699e-06, 
    4.301106e-06, 3.164148e-06, 3.803658e-06, 5.097469e-06, 4.489482e-06, 
    6.403095e-06, 6.542547e-06, 7.324639e-06, 8.354646e-06, 7.359245e-06,
  5.251093e-06, 6.387883e-06, 6.670477e-06, 7.642771e-06, 4.868614e-06, 
    3.515393e-06, 6.126107e-06, 7.282201e-06, 8.250036e-06, 7.828348e-06, 
    6.805431e-06, 1.033466e-05, 7.606747e-06, 8.21821e-06, 7.147927e-06,
  4.9064e-06, 7.397039e-06, 1.021975e-05, 9.153739e-06, 6.407062e-06, 
    5.200032e-06, 4.943356e-06, 4.869679e-06, 4.615171e-06, 5.416759e-06, 
    6.328223e-06, 7.260071e-06, 3.574949e-06, 4.897709e-06, 1.988752e-06,
  5.369909e-06, 5.74152e-06, 2.386766e-06, 2.56856e-06, 2.101761e-06, 
    1.622186e-06, 3.211847e-06, 3.998124e-06, 7.350985e-06, 7.288148e-06, 
    7.893251e-06, 9.948263e-06, 1.004787e-05, 8.043769e-06, 5.033563e-06,
  4.195297e-06, 2.504469e-06, 2.507326e-06, 4.127956e-06, 3.530984e-06, 
    3.795336e-06, 4.753288e-06, 8.469926e-06, 8.534989e-06, 9.126138e-06, 
    1.079754e-05, 1.151738e-05, 1.191559e-05, 1.11801e-05, 7.813657e-06,
  3.807347e-06, 4.060359e-06, 5.990165e-06, 7.481076e-06, 8.434896e-06, 
    8.93796e-06, 1.172537e-05, 1.045351e-05, 1.001058e-05, 9.164462e-06, 
    8.136495e-06, 1.20186e-05, 1.36984e-05, 1.303361e-05, 7.028745e-06,
  4.501886e-06, 5.845505e-06, 8.353875e-06, 1.081274e-05, 1.228517e-05, 
    1.094178e-05, 1.022148e-05, 7.803024e-06, 7.779479e-06, 7.228426e-06, 
    5.818406e-06, 8.001271e-06, 6.982284e-06, 9.181714e-06, 4.59712e-06,
  7.118333e-06, 8.088715e-06, 9.941617e-06, 1.171633e-05, 1.35485e-05, 
    8.844737e-06, 9.307087e-06, 8.407276e-06, 7.949448e-06, 6.748975e-06, 
    3.191213e-06, 3.075757e-06, 5.711749e-06, 7.866137e-06, 5.512566e-06,
  7.171236e-06, 7.725101e-06, 9.159281e-06, 1.030254e-05, 1.167286e-05, 
    1.040551e-05, 9.359115e-06, 8.298563e-06, 6.403735e-06, 6.096102e-06, 
    4.251914e-06, 4.304698e-06, 5.382939e-06, 1.029873e-05, 9.419248e-06,
  4.013817e-06, 2.600068e-06, 6.677133e-06, 2.46768e-06, 2.101697e-06, 
    1.658035e-06, 1.37043e-06, 2.224048e-06, 1.486663e-05, 8.188879e-05, 
    0.0001802034, 0.0004511219, 0.0007763086, 0.0009509656, 0.0008473029,
  3.952012e-06, 4.843013e-06, 4.343433e-06, 3.71018e-06, 2.610309e-06, 
    1.976369e-06, 1.880099e-06, 2.860402e-06, 4.587007e-06, 1.932542e-05, 
    0.0001140338, 0.0002255573, 0.0003950548, 0.0005358215, 0.0005036068,
  5.384201e-06, 6.132912e-06, 5.604357e-06, 4.719589e-06, 5.45705e-06, 
    4.152653e-06, 3.807264e-06, 2.049007e-06, 3.86401e-06, 5.002455e-06, 
    2.285114e-05, 7.764853e-05, 0.0001527783, 0.0002271452, 0.0002394164,
  5.962361e-06, 4.881333e-06, 4.982728e-06, 5.236161e-06, 6.299235e-06, 
    5.203444e-06, 4.39096e-06, 9.405406e-07, 3.823389e-06, 4.067561e-06, 
    5.576835e-06, 1.018008e-05, 2.974308e-05, 7.918709e-05, 7.993021e-05,
  4.874189e-06, 4.325383e-06, 3.797513e-06, 7.333905e-06, 7.336111e-06, 
    9.713875e-06, 5.942394e-06, 4.26792e-06, 6.593473e-06, 3.89993e-06, 
    3.182312e-06, 3.790286e-06, 3.695538e-06, 8.927097e-06, 1.306579e-05,
  1.122432e-05, 7.188875e-06, 6.602331e-06, 7.835053e-06, 8.397511e-06, 
    8.275084e-06, 7.167032e-06, 7.509494e-06, 6.906767e-06, 6.030033e-06, 
    7.59248e-06, 6.525545e-06, 5.121234e-06, 3.174671e-06, 6.296435e-06,
  9.419775e-06, 1.332967e-05, 1.052164e-05, 1.386805e-05, 1.246396e-05, 
    1.424586e-05, 1.0608e-05, 9.774199e-06, 9.305769e-06, 1.02133e-05, 
    9.045043e-06, 7.983949e-06, 5.199492e-06, 5.705255e-06, 7.191126e-06,
  6.742659e-06, 1.166404e-05, 1.571252e-05, 1.486587e-05, 1.579093e-05, 
    1.362416e-05, 7.004723e-06, 5.966896e-06, 7.295094e-06, 1.038066e-05, 
    7.26707e-06, 8.855414e-06, 8.102021e-06, 1.054507e-05, 7.850838e-06,
  7.963009e-06, 9.273245e-06, 1.269353e-05, 1.356668e-05, 1.646525e-05, 
    1.136429e-05, 9.344964e-06, 1.078864e-05, 1.220888e-05, 1.27493e-05, 
    1.153002e-05, 1.034476e-05, 1.101492e-05, 1.202848e-05, 1.063342e-05,
  5.533044e-06, 5.223229e-06, 8.008497e-06, 1.130368e-05, 1.231084e-05, 
    1.012759e-05, 9.731374e-06, 9.473921e-06, 1.109834e-05, 1.392772e-05, 
    1.376936e-05, 1.344775e-05, 1.466045e-05, 1.288015e-05, 1.273088e-05,
  6.84042e-06, 5.404711e-06, 6.890822e-06, 3.42828e-05, 5.597761e-05, 
    4.366077e-05, 3.222298e-05, 2.785537e-05, 3.048973e-05, 4.634889e-05, 
    0.0001721111, 0.0003595866, 0.0005057629, 0.0006146142, 0.0006026216,
  3.09721e-06, 5.248605e-06, 4.344841e-06, 1.64164e-05, 4.178358e-05, 
    3.734301e-05, 2.723332e-05, 2.234084e-05, 2.765315e-05, 4.502248e-05, 
    0.0001280299, 0.0004489646, 0.0007386165, 0.0009234432, 0.0009228538,
  8.569689e-07, 3.244009e-06, 4.241399e-06, 6.2628e-06, 2.616759e-05, 
    3.330549e-05, 2.463389e-05, 1.969485e-05, 2.29363e-05, 4.013711e-05, 
    9.012531e-05, 0.0004556347, 0.0008655833, 0.001112222, 0.001026071,
  7.66231e-07, 1.382023e-06, 3.434445e-06, 4.796178e-06, 1.522735e-05, 
    2.598749e-05, 2.457963e-05, 1.825985e-05, 1.794338e-05, 3.027802e-05, 
    5.944621e-05, 0.0003633926, 0.0007750868, 0.001026824, 0.001138745,
  7.852236e-07, 1.487286e-06, 2.020669e-06, 4.409213e-06, 1.04787e-05, 
    2.03729e-05, 2.453281e-05, 2.219006e-05, 1.794146e-05, 2.332086e-05, 
    4.61554e-05, 0.0002734947, 0.0006499239, 0.001024889, 0.001104786,
  1.928346e-06, 2.476942e-06, 1.266847e-06, 1.950523e-06, 6.437727e-06, 
    1.551426e-05, 2.317751e-05, 2.430734e-05, 2.215182e-05, 2.261382e-05, 
    3.927341e-05, 0.0002164187, 0.0005390017, 0.0009473178, 0.001125054,
  4.2584e-06, 3.360574e-06, 7.292186e-07, 9.654897e-07, 2.226796e-06, 
    1.031434e-05, 1.774546e-05, 2.400226e-05, 2.237794e-05, 2.343798e-05, 
    3.039616e-05, 0.0001522958, 0.0004275384, 0.0008184313, 0.001099927,
  5.698482e-06, 4.546144e-06, 3.638803e-06, 1.754943e-06, 1.022776e-06, 
    4.229956e-06, 1.415341e-05, 2.201956e-05, 2.397373e-05, 2.163531e-05, 
    2.789824e-05, 8.97205e-05, 0.0003142878, 0.0006946531, 0.001043343,
  9.75345e-06, 6.197007e-06, 4.727677e-06, 2.457724e-06, 1.707831e-06, 
    3.394101e-06, 1.003643e-05, 1.8593e-05, 2.421823e-05, 2.44554e-05, 
    2.749621e-05, 6.759361e-05, 0.0002391496, 0.0005987203, 0.0009906336,
  1.114514e-05, 1.080032e-05, 6.025106e-06, 3.916106e-06, 5.12622e-06, 
    5.681827e-06, 5.371792e-06, 1.325397e-05, 2.190941e-05, 2.554932e-05, 
    2.77194e-05, 5.797611e-05, 0.0002043276, 0.0005317237, 0.0009434046,
  0.0002940624, 0.0003611919, 0.0001611289, 5.988691e-05, 7.516304e-06, 
    5.243022e-06, 1.17691e-06, 2.532882e-06, 4.512973e-06, 4.089383e-06, 
    3.597502e-06, 3.342654e-06, 4.980697e-06, 6.403436e-06, 1.246195e-05,
  0.0003327023, 0.0004132438, 0.0001835661, 8.224096e-05, 1.958739e-05, 
    6.200312e-06, 4.125278e-06, 3.855961e-06, 7.479065e-06, 4.519535e-06, 
    5.077545e-06, 3.965794e-06, 5.484194e-06, 7.184653e-06, 1.030566e-05,
  0.0003194067, 0.0004164703, 0.0001758471, 9.652148e-05, 3.383022e-05, 
    8.322977e-06, 6.147212e-06, 5.087563e-06, 5.028582e-06, 2.922357e-06, 
    5.479491e-06, 4.962836e-06, 4.970175e-06, 7.491311e-06, 1.28676e-05,
  0.0003145419, 0.0003991371, 0.0001892954, 0.0001010259, 4.704341e-05, 
    1.420681e-05, 6.09452e-06, 4.268249e-06, 4.487664e-06, 5.632699e-06, 
    6.462138e-06, 5.960565e-06, 7.687793e-06, 9.737601e-06, 1.402606e-05,
  0.0002774342, 0.0003535332, 0.0001958376, 0.0001050401, 5.603048e-05, 
    2.409377e-05, 6.753008e-06, 4.114318e-06, 4.105566e-06, 7.846807e-06, 
    4.917223e-06, 6.422123e-06, 8.287025e-06, 1.030382e-05, 1.522035e-05,
  0.0002437209, 0.000310174, 0.0002088256, 0.0001149684, 6.453036e-05, 
    3.461465e-05, 1.392815e-05, 5.345789e-06, 5.374921e-06, 3.9377e-06, 
    5.770067e-06, 5.093257e-06, 7.470609e-06, 1.073544e-05, 1.356756e-05,
  0.0002594862, 0.000293335, 0.000219286, 0.0001191918, 6.379143e-05, 
    4.041823e-05, 2.271798e-05, 1.131373e-05, 5.754565e-06, 3.894627e-06, 
    4.976394e-06, 7.053003e-06, 9.962543e-06, 1.042138e-05, 1.618727e-05,
  0.0002835169, 0.0002999378, 0.0002199701, 0.0001297465, 7.085806e-05, 
    4.443952e-05, 3.03038e-05, 1.81498e-05, 8.201397e-06, 4.893852e-06, 
    5.013613e-06, 6.221529e-06, 9.281634e-06, 1.028724e-05, 1.1445e-05,
  0.0002842853, 0.0002811977, 0.0002167572, 0.000128582, 7.451876e-05, 
    4.866607e-05, 3.634615e-05, 2.405804e-05, 1.584833e-05, 5.477636e-06, 
    3.653744e-06, 7.239988e-06, 9.351918e-06, 9.424743e-06, 1.120095e-05,
  0.0002177636, 0.0002559507, 0.0002050494, 0.0001215203, 7.431836e-05, 
    4.733876e-05, 4.289712e-05, 3.158718e-05, 2.060752e-05, 1.399337e-05, 
    5.361888e-06, 7.71308e-06, 9.425066e-06, 8.099425e-06, 7.979374e-06,
  0.0005584733, 0.000289372, 6.452717e-05, 9.659904e-06, 8.477988e-06, 
    9.283867e-06, 1.255542e-05, 8.834363e-06, 8.411092e-06, 9.850134e-06, 
    1.07479e-05, 8.400979e-06, 7.595589e-06, 8.262272e-06, 5.937697e-06,
  0.000559205, 0.0002780331, 4.296682e-05, 7.604221e-06, 7.525154e-06, 
    8.507703e-06, 7.061183e-06, 8.451792e-06, 5.294823e-06, 7.425581e-06, 
    6.755909e-06, 7.911709e-06, 5.906586e-06, 6.340762e-06, 6.412713e-06,
  0.0005150727, 0.0002476704, 2.337178e-05, 7.825783e-06, 5.810797e-06, 
    7.968853e-06, 9.395562e-06, 7.969302e-06, 3.95476e-06, 4.271961e-06, 
    8.53709e-06, 6.637372e-06, 5.804781e-06, 5.837562e-06, 6.059967e-06,
  0.000463993, 0.0002213677, 1.579088e-05, 7.2222e-06, 5.221222e-06, 
    6.800568e-06, 5.557668e-06, 3.171447e-06, 4.009628e-06, 5.387737e-06, 
    7.78965e-06, 5.336006e-06, 6.160886e-06, 7.013755e-06, 6.060245e-06,
  0.0004148889, 0.0001935399, 1.362286e-05, 7.380316e-06, 5.04423e-06, 
    5.707502e-06, 6.031068e-06, 4.345933e-06, 4.093578e-06, 6.710623e-06, 
    5.607349e-06, 4.144606e-06, 4.448715e-06, 5.218861e-06, 4.859893e-06,
  0.0003766766, 0.0001507814, 1.100246e-05, 5.832921e-06, 4.868851e-06, 
    5.723337e-06, 5.307634e-06, 2.320437e-06, 3.502904e-06, 6.028483e-06, 
    5.678587e-06, 4.441629e-06, 3.109503e-06, 3.164602e-06, 5.672318e-06,
  0.0003339564, 0.0001272791, 8.560804e-06, 4.867708e-06, 4.515573e-06, 
    5.014544e-06, 4.249807e-06, 2.30097e-06, 3.361149e-06, 6.849712e-06, 
    4.703486e-06, 3.993623e-06, 4.230785e-06, 4.803101e-06, 4.357997e-06,
  0.0003151941, 0.0001024582, 6.944147e-06, 3.182397e-06, 3.925415e-06, 
    5.168992e-06, 3.035688e-06, 2.996448e-06, 4.036278e-06, 5.683628e-06, 
    5.210172e-06, 4.543577e-06, 4.226433e-06, 4.688437e-06, 3.417621e-06,
  0.0003180222, 9.596221e-05, 7.297184e-06, 2.789771e-06, 5.035279e-06, 
    4.834387e-06, 3.019419e-06, 2.484951e-06, 3.504819e-06, 5.575483e-06, 
    5.174369e-06, 3.787795e-06, 3.702027e-06, 4.088198e-06, 4.585349e-06,
  0.000364358, 0.0001058155, 8.685782e-06, 2.854804e-06, 4.569045e-06, 
    4.93505e-06, 2.720207e-06, 2.35878e-06, 4.620982e-06, 4.84649e-06, 
    4.257396e-06, 3.415177e-06, 4.580849e-06, 3.174022e-06, 3.804083e-06,
  5.873789e-06, 7.959516e-06, 8.828485e-06, 9.348259e-06, 1.019887e-05, 
    8.790347e-06, 7.814354e-06, 8.430748e-06, 6.818256e-06, 5.746582e-06, 
    5.744134e-06, 4.931203e-06, 7.25886e-06, 7.466328e-06, 3.227927e-06,
  6.069199e-06, 7.685186e-06, 7.824645e-06, 8.406293e-06, 9.436695e-06, 
    9.279433e-06, 8.823714e-06, 8.410342e-06, 5.476609e-06, 3.550596e-06, 
    4.856609e-06, 5.406382e-06, 9.18886e-06, 8.167623e-06, 2.512496e-06,
  9.235856e-06, 6.994653e-06, 7.716741e-06, 9.154115e-06, 1.161187e-05, 
    9.901216e-06, 9.445444e-06, 4.640085e-06, 4.043397e-06, 4.81522e-06, 
    4.953703e-06, 6.549474e-06, 8.588308e-06, 2.88845e-06, 2.786239e-06,
  1.057033e-05, 6.92013e-06, 8.777974e-06, 9.837562e-06, 9.23868e-06, 
    8.685539e-06, 7.783996e-06, 4.062211e-06, 3.709102e-06, 4.289242e-06, 
    5.778199e-06, 8.031792e-06, 7.174016e-06, 3.284187e-06, 3.870803e-06,
  1.247238e-05, 7.733483e-06, 8.252381e-06, 8.18938e-06, 9.350631e-06, 
    9.978843e-06, 5.604039e-06, 3.258165e-06, 4.454056e-06, 5.070897e-06, 
    7.139697e-06, 9.29319e-06, 5.836615e-06, 5.025185e-06, 8.103417e-06,
  1.232923e-05, 6.818168e-06, 7.753336e-06, 8.687787e-06, 9.890319e-06, 
    7.356992e-06, 5.685794e-06, 3.74127e-06, 5.407706e-06, 5.476434e-06, 
    7.830085e-06, 9.010927e-06, 3.03824e-06, 6.78071e-06, 1.072329e-05,
  7.600734e-06, 5.898687e-06, 6.921033e-06, 8.918295e-06, 9.95469e-06, 
    5.079688e-06, 5.010934e-06, 4.011814e-06, 5.446124e-06, 6.508923e-06, 
    9.105698e-06, 7.399968e-06, 3.077022e-06, 4.883432e-06, 6.671637e-06,
  9.407953e-06, 6.022386e-06, 9.595633e-06, 1.09869e-05, 7.487373e-06, 
    5.403156e-06, 3.76136e-06, 4.399068e-06, 6.196231e-06, 6.94325e-06, 
    8.535045e-06, 8.970564e-06, 4.946321e-06, 4.173075e-06, 5.664805e-06,
  3.900147e-06, 2.486336e-06, 3.808967e-06, 6.992004e-06, 5.389541e-06, 
    4.630846e-06, 3.951226e-06, 5.638236e-06, 5.536566e-06, 4.454619e-06, 
    7.344364e-06, 6.777798e-06, 5.13637e-06, 3.474978e-06, 2.321336e-06,
  3.173026e-06, 1.50261e-06, 5.51312e-06, 4.317154e-06, 4.651825e-06, 
    4.8893e-06, 4.635253e-06, 4.825417e-06, 6.521303e-06, 5.069854e-06, 
    4.49007e-06, 5.713474e-06, 5.883904e-06, 7.314265e-06, 4.05125e-06,
  1.307153e-05, 1.042264e-05, 1.111832e-05, 9.839193e-06, 7.764296e-06, 
    8.402799e-06, 6.555433e-06, 6.527368e-06, 6.894451e-06, 1.245845e-05, 
    1.641865e-05, 1.672913e-05, 1.066903e-05, 7.897747e-06, 9.125235e-06,
  1.079952e-05, 8.609391e-06, 1.201796e-05, 7.842305e-06, 8.989752e-06, 
    9.324103e-06, 7.25725e-06, 7.38372e-06, 8.94294e-06, 1.328933e-05, 
    1.39175e-05, 1.23172e-05, 5.929752e-06, 8.366895e-06, 7.902897e-06,
  8.715717e-06, 9.695132e-06, 9.668364e-06, 1.016036e-05, 1.042626e-05, 
    1.06158e-05, 9.993004e-06, 9.494403e-06, 1.360636e-05, 1.203284e-05, 
    1.148233e-05, 8.131064e-06, 6.286346e-06, 3.187753e-06, 5.322009e-06,
  9.967767e-06, 9.931662e-06, 1.316178e-05, 9.512662e-06, 8.977137e-06, 
    9.915911e-06, 9.456032e-06, 1.011035e-05, 1.326483e-05, 1.163894e-05, 
    8.712076e-06, 8.420363e-06, 8.877331e-06, 5.941903e-06, 3.692716e-06,
  1.041548e-05, 1.149453e-05, 1.335799e-05, 1.029395e-05, 9.884729e-06, 
    1.051831e-05, 9.025631e-06, 1.016045e-05, 1.504094e-05, 1.163576e-05, 
    1.047374e-05, 9.23612e-06, 7.555712e-06, 7.417181e-06, 6.091484e-06,
  1.222791e-05, 1.133611e-05, 1.21293e-05, 1.071336e-05, 8.36678e-06, 
    1.033043e-05, 9.849196e-06, 1.512782e-05, 1.529131e-05, 9.702578e-06, 
    1.001983e-05, 1.079387e-05, 5.501485e-06, 6.442931e-06, 7.549035e-06,
  1.345137e-05, 9.712712e-06, 1.372724e-05, 1.208822e-05, 1.254201e-05, 
    1.656556e-05, 1.520787e-05, 1.569327e-05, 1.207894e-05, 1.061514e-05, 
    1.216581e-05, 1.093806e-05, 7.334037e-06, 6.732794e-06, 7.568935e-06,
  8.639194e-06, 1.171661e-05, 1.429277e-05, 1.420246e-05, 1.585109e-05, 
    1.072794e-05, 1.257019e-05, 1.410831e-05, 1.212056e-05, 1.323288e-05, 
    1.325886e-05, 1.088253e-05, 8.348004e-06, 8.290225e-06, 5.766148e-06,
  6.802087e-06, 8.902956e-06, 1.507245e-05, 1.422855e-05, 1.112267e-05, 
    1.183177e-05, 1.204021e-05, 1.266324e-05, 1.350322e-05, 1.717991e-05, 
    1.148528e-05, 1.039128e-05, 8.3789e-06, 5.388628e-06, 5.382542e-06,
  5.124666e-06, 8.401789e-06, 1.047032e-05, 1.112854e-05, 7.483502e-06, 
    1.009401e-05, 1.177258e-05, 1.28186e-05, 1.328252e-05, 1.183771e-05, 
    9.754702e-06, 8.3248e-06, 1.01883e-05, 6.633963e-06, 7.058141e-06,
  1.586266e-05, 1.198938e-05, 9.92108e-06, 8.590341e-06, 9.093752e-06, 
    6.05128e-06, 5.13228e-06, 4.356938e-06, 3.999057e-06, 3.804423e-06, 
    3.245705e-06, 3.377153e-06, 6.183433e-06, 6.170761e-06, 9.709625e-06,
  1.577659e-05, 1.399736e-05, 1.090693e-05, 8.638121e-06, 6.612877e-06, 
    6.025001e-06, 4.807787e-06, 5.149958e-06, 4.940267e-06, 3.789303e-06, 
    3.27266e-06, 2.226278e-06, 5.772954e-06, 7.594148e-06, 7.327681e-06,
  1.715692e-05, 1.465936e-05, 1.123705e-05, 8.260941e-06, 7.675959e-06, 
    6.353661e-06, 6.859577e-06, 6.440816e-06, 6.424709e-06, 5.30641e-06, 
    6.240522e-06, 2.280762e-06, 3.204322e-06, 8.606188e-06, 8.169841e-06,
  1.795608e-05, 1.302119e-05, 1.207684e-05, 9.527957e-06, 1.017743e-05, 
    1.061648e-05, 1.240073e-05, 1.300674e-05, 1.074962e-05, 9.131756e-06, 
    5.604709e-06, 2.53351e-06, 3.263332e-06, 6.830541e-06, 1.031483e-05,
  2.018031e-05, 1.606807e-05, 1.574504e-05, 1.411891e-05, 1.37805e-05, 
    1.532472e-05, 1.033795e-05, 1.140333e-05, 1.003624e-05, 1.233337e-05, 
    1.136161e-05, 4.719117e-06, 4.261125e-06, 6.251153e-06, 1.077608e-05,
  2.594302e-05, 2.320701e-05, 2.353553e-05, 2.08934e-05, 2.001974e-05, 
    1.509083e-05, 9.27724e-06, 6.695961e-06, 1.064654e-05, 1.098934e-05, 
    1.373754e-05, 8.813361e-06, 5.777319e-06, 7.710806e-06, 7.721377e-06,
  3.441206e-05, 3.453354e-05, 3.037569e-05, 3.003616e-05, 2.170708e-05, 
    1.183906e-05, 5.537514e-06, 6.113737e-06, 3.684062e-06, 1.107368e-05, 
    1.166786e-05, 1.146118e-05, 1.593234e-05, 6.478337e-06, 8.336317e-06,
  2.894676e-05, 2.922589e-05, 2.106381e-05, 2.088725e-05, 1.795197e-05, 
    1.123929e-05, 4.016913e-06, 3.526503e-06, 3.824014e-06, 5.098264e-06, 
    7.879427e-06, 7.345758e-06, 1.196617e-05, 8.156414e-06, 9.273404e-06,
  2.215275e-05, 2.117123e-05, 2.280578e-05, 1.729528e-05, 1.473419e-05, 
    1.00955e-05, 4.511735e-06, 2.394098e-06, 2.538496e-06, 2.068691e-06, 
    3.612185e-06, 5.939352e-06, 7.944093e-06, 9.374068e-06, 6.917126e-06,
  2.460397e-05, 2.180471e-05, 1.590415e-05, 1.433138e-05, 1.234357e-05, 
    8.029613e-06, 3.116689e-06, 2.678915e-06, 1.788569e-06, 1.6616e-06, 
    2.480723e-06, 3.921902e-06, 5.236794e-06, 8.157912e-06, 5.836548e-06,
  5.223184e-06, 4.083242e-06, 4.322143e-06, 4.417975e-06, 4.098783e-06, 
    4.319207e-06, 4.246963e-06, 7.29329e-06, 5.40478e-06, 1.091661e-05, 
    7.067482e-06, 6.891102e-06, 2.575328e-05, 7.364369e-05, 0.000108601,
  4.500057e-06, 3.725997e-06, 4.119597e-06, 3.841202e-06, 4.075705e-06, 
    4.460603e-06, 5.282219e-06, 5.146574e-06, 8.779737e-06, 6.964508e-06, 
    8.16463e-06, 9.208647e-06, 3.74849e-05, 8.851473e-05, 0.0001199216,
  6.297948e-06, 3.283775e-06, 4.328628e-06, 3.976907e-06, 4.919706e-06, 
    3.567298e-06, 5.184308e-06, 4.550071e-06, 9.430247e-06, 9.712437e-06, 
    7.962022e-06, 8.525308e-06, 3.638191e-05, 9.357063e-05, 0.0001208325,
  6.668752e-06, 5.987885e-06, 3.123075e-06, 5.079435e-06, 4.905199e-06, 
    2.799109e-06, 4.88229e-06, 8.449836e-06, 5.76703e-06, 7.911088e-06, 
    8.690949e-06, 9.132898e-06, 2.946266e-05, 9.505149e-05, 0.0001194583,
  5.949486e-06, 6.753005e-06, 4.109553e-06, 3.734895e-06, 3.926643e-06, 
    3.384746e-06, 5.254927e-06, 1.055892e-05, 7.767328e-06, 7.260234e-06, 
    6.760994e-06, 8.951502e-06, 3.414313e-05, 9.403193e-05, 0.0001098184,
  6.103551e-06, 5.621093e-06, 3.540686e-06, 3.455589e-06, 5.171679e-06, 
    4.636609e-06, 5.113296e-06, 1.011568e-05, 8.156664e-06, 8.446359e-06, 
    7.260838e-06, 7.460755e-06, 4.051358e-05, 8.439447e-05, 9.581301e-05,
  6.112278e-06, 5.749443e-06, 5.293532e-06, 4.856976e-06, 3.512118e-06, 
    4.018522e-06, 8.636401e-06, 1.10549e-05, 1.041798e-05, 9.720654e-06, 
    8.701923e-06, 8.379856e-06, 3.98256e-05, 8.455918e-05, 7.943641e-05,
  7.680215e-06, 5.861691e-06, 5.933687e-06, 4.844741e-06, 4.165545e-06, 
    4.927675e-06, 7.530657e-06, 8.663945e-06, 1.029176e-05, 1.178743e-05, 
    9.463742e-06, 9.026e-06, 5.315136e-05, 8.020613e-05, 5.881874e-05,
  1.268787e-05, 6.673552e-06, 5.991833e-06, 6.088953e-06, 4.997425e-06, 
    8.240509e-06, 9.210991e-06, 7.038377e-06, 9.477597e-06, 1.011049e-05, 
    9.973128e-06, 9.654796e-06, 5.035411e-05, 7.016954e-05, 5.001292e-05,
  3.124064e-05, 8.139214e-06, 7.958834e-06, 7.180532e-06, 4.625719e-06, 
    5.918867e-06, 9.244017e-06, 8.275778e-06, 9.172331e-06, 1.032087e-05, 
    8.543569e-06, 7.967214e-06, 4.413835e-05, 5.271069e-05, 4.529058e-05,
  8.794183e-06, 8.548735e-06, 9.904294e-06, 2.00988e-05, 2.162303e-05, 
    2.441174e-05, 2.687463e-05, 2.69949e-05, 2.847279e-05, 3.529825e-05, 
    4.660955e-05, 5.724869e-05, 5.499265e-05, 2.499951e-05, 6.24624e-06,
  7.353474e-06, 6.96497e-06, 9.825876e-06, 1.711652e-05, 2.271622e-05, 
    2.607001e-05, 2.707839e-05, 2.796121e-05, 3.72364e-05, 4.603964e-05, 
    5.623745e-05, 6.614187e-05, 5.690372e-05, 1.976792e-05, 6.806252e-06,
  9.951905e-06, 7.616085e-06, 1.13056e-05, 1.763977e-05, 2.176557e-05, 
    2.595859e-05, 2.90461e-05, 3.073505e-05, 4.090299e-05, 5.055395e-05, 
    5.64373e-05, 6.455459e-05, 5.864885e-05, 1.847544e-05, 7.821863e-06,
  7.589183e-06, 1.020837e-05, 1.128684e-05, 2.015478e-05, 2.336394e-05, 
    2.746869e-05, 3.004854e-05, 3.865383e-05, 5.240416e-05, 5.452511e-05, 
    5.691724e-05, 6.132155e-05, 6.145089e-05, 1.618552e-05, 8.150848e-06,
  7.312187e-06, 7.829236e-06, 1.172614e-05, 2.043279e-05, 2.379003e-05, 
    2.62633e-05, 3.139181e-05, 4.63559e-05, 6.26976e-05, 6.101899e-05, 
    6.062309e-05, 6.680026e-05, 5.794293e-05, 1.726914e-05, 1.066898e-05,
  5.80618e-06, 7.330128e-06, 1.222251e-05, 2.25496e-05, 2.465378e-05, 
    2.826129e-05, 3.468535e-05, 5.212087e-05, 7.615705e-05, 6.7833e-05, 
    5.841305e-05, 6.598388e-05, 5.642437e-05, 1.716986e-05, 1.301643e-05,
  6.107914e-06, 8.3592e-06, 9.000759e-06, 2.023556e-05, 3.639365e-05, 
    3.274889e-05, 4.923438e-05, 6.224665e-05, 7.155937e-05, 7.158524e-05, 
    5.981891e-05, 6.222757e-05, 4.951038e-05, 2.046055e-05, 1.717848e-05,
  5.841288e-06, 8.264305e-06, 8.430367e-06, 1.788249e-05, 2.651084e-05, 
    4.087379e-05, 4.48609e-05, 7.042157e-05, 7.573152e-05, 7.295578e-05, 
    5.776958e-05, 6.121592e-05, 4.449057e-05, 2.117265e-05, 2.040565e-05,
  4.692215e-06, 6.922263e-06, 7.277658e-06, 2.098979e-05, 3.420704e-05, 
    3.532441e-05, 5.336006e-05, 6.174722e-05, 7.558538e-05, 8.314048e-05, 
    5.212897e-05, 5.602529e-05, 4.517091e-05, 2.604657e-05, 2.499281e-05,
  4.310726e-06, 6.378119e-06, 7.064802e-06, 1.179145e-05, 3.268755e-05, 
    3.856646e-05, 5.336763e-05, 7.285573e-05, 7.69222e-05, 7.077738e-05, 
    5.48417e-05, 5.555333e-05, 4.554485e-05, 2.338194e-05, 3.439687e-05,
  1.831606e-05, 9.626469e-06, 4.757712e-06, 3.208252e-06, 3.98754e-06, 
    3.912432e-06, 4.122551e-06, 3.520528e-06, 3.189916e-06, 4.392985e-06, 
    3.844315e-06, 3.089979e-06, 2.005857e-06, 1.86767e-06, 6.222657e-06,
  9.678299e-06, 7.600979e-06, 5.684704e-06, 3.151794e-06, 2.503211e-06, 
    3.153814e-06, 2.927982e-06, 2.906895e-06, 2.670501e-06, 3.650898e-06, 
    3.959794e-06, 3.156177e-06, 2.542754e-06, 3.344426e-06, 7.271171e-06,
  1.562357e-05, 8.997908e-06, 8.117141e-06, 3.09744e-06, 2.653675e-06, 
    4.247483e-06, 3.774637e-06, 2.379903e-06, 2.67149e-06, 3.840539e-06, 
    2.831973e-06, 3.014029e-06, 2.929825e-06, 4.259258e-06, 7.247439e-06,
  1.817665e-05, 1.622582e-05, 9.89314e-06, 4.549538e-06, 2.935996e-06, 
    3.728381e-06, 2.83482e-06, 2.701092e-06, 2.758846e-06, 2.637136e-06, 
    2.390099e-06, 2.637107e-06, 3.332256e-06, 4.668125e-06, 7.013311e-06,
  1.880243e-05, 9.234457e-06, 1.040873e-05, 4.338373e-06, 2.538364e-06, 
    3.080557e-06, 2.585228e-06, 3.067271e-06, 2.273012e-06, 2.485215e-06, 
    2.535878e-06, 2.73684e-06, 3.686155e-06, 5.897899e-06, 7.41526e-06,
  1.342536e-05, 1.43961e-05, 1.177991e-05, 5.427575e-06, 3.294594e-06, 
    2.985488e-06, 3.359077e-06, 2.884032e-06, 3.297929e-06, 2.178751e-06, 
    3.089758e-06, 3.548136e-06, 4.415101e-06, 5.751776e-06, 8.022714e-06,
  2.209953e-05, 1.459352e-05, 1.471674e-05, 5.944838e-06, 3.064684e-06, 
    2.391058e-06, 2.753388e-06, 3.268884e-06, 3.012062e-06, 2.352833e-06, 
    2.820667e-06, 3.800622e-06, 4.574405e-06, 5.772642e-06, 7.345175e-06,
  1.806094e-05, 1.133669e-05, 1.353286e-05, 9.954952e-06, 2.933687e-06, 
    3.426195e-06, 2.739289e-06, 3.631053e-06, 2.444846e-06, 2.570194e-06, 
    3.094887e-06, 4.337754e-06, 5.391891e-06, 5.802795e-06, 7.123856e-06,
  2.135077e-05, 1.426366e-05, 1.72132e-05, 9.554977e-06, 3.132923e-06, 
    3.035669e-06, 3.096432e-06, 3.948629e-06, 3.142446e-06, 3.571991e-06, 
    4.127604e-06, 5.101083e-06, 5.843525e-06, 6.579188e-06, 7.377535e-06,
  1.729669e-05, 1.026344e-05, 1.193418e-05, 2.204025e-05, 3.521882e-06, 
    2.295586e-06, 2.843962e-06, 4.367502e-06, 3.764654e-06, 3.124608e-06, 
    4.054536e-06, 4.843513e-06, 5.744977e-06, 5.577886e-06, 6.841437e-06,
  2.282682e-06, 4.919714e-06, 7.191878e-06, 8.927073e-06, 9.628832e-06, 
    6.811193e-06, 4.747331e-06, 7.054204e-06, 4.081898e-06, 2.62295e-06, 
    1.020833e-06, 1.018028e-06, 4.196559e-06, 1.003822e-05, 8.219537e-06,
  4.271997e-06, 5.706041e-06, 7.219796e-06, 8.886071e-06, 5.922104e-06, 
    5.74005e-06, 5.007914e-06, 5.637608e-06, 3.139657e-06, 2.665066e-06, 
    1.02932e-06, 1.654009e-06, 4.217778e-06, 5.690079e-06, 2.687463e-06,
  3.816049e-06, 5.92229e-06, 7.564776e-06, 5.933784e-06, 6.429472e-06, 
    5.124586e-06, 5.166008e-06, 3.115872e-06, 1.964603e-06, 8.411682e-07, 
    1.936023e-06, 6.268038e-06, 6.79699e-06, 5.659586e-06, 2.672663e-06,
  6.431318e-06, 8.446822e-06, 5.402914e-06, 4.147467e-06, 2.649186e-06, 
    2.307048e-06, 3.328299e-06, 2.083854e-06, 1.347162e-06, 1.130839e-06, 
    1.966659e-06, 5.655968e-06, 7.269424e-06, 3.470185e-06, 2.177874e-06,
  7.918289e-06, 6.099109e-06, 3.815429e-06, 3.315195e-06, 1.842995e-06, 
    2.070801e-06, 1.782472e-06, 1.281524e-06, 1.690424e-06, 1.391425e-06, 
    2.086381e-06, 2.831139e-06, 2.945784e-06, 2.156555e-06, 1.580012e-06,
  5.205381e-06, 4.40708e-06, 2.514478e-06, 2.278705e-06, 2.350936e-06, 
    1.499912e-06, 1.326912e-06, 2.696713e-06, 2.079577e-06, 2.354332e-06, 
    2.603063e-06, 2.700842e-06, 2.474727e-06, 1.106619e-06, 1.624136e-06,
  4.156257e-06, 2.549651e-06, 2.262953e-06, 2.960143e-06, 2.435175e-06, 
    1.188269e-06, 2.359151e-06, 1.614313e-06, 2.308998e-06, 3.127828e-06, 
    3.286705e-06, 3.445098e-06, 3.306752e-06, 2.325004e-06, 2.508432e-06,
  4.372189e-06, 2.509e-06, 2.398125e-06, 2.885954e-06, 1.93994e-06, 
    1.566486e-06, 1.759466e-06, 2.234587e-06, 3.049455e-06, 4.124088e-06, 
    3.536858e-06, 2.569202e-06, 3.05618e-06, 2.810646e-06, 2.481518e-06,
  3.980677e-06, 1.960544e-06, 2.371798e-06, 2.255739e-06, 1.730562e-06, 
    1.929214e-06, 1.153898e-06, 2.302551e-06, 3.204676e-06, 2.479061e-06, 
    2.415262e-06, 2.321117e-06, 2.874878e-06, 3.654393e-06, 3.516875e-06,
  2.178098e-06, 1.14754e-06, 1.140489e-06, 1.03392e-06, 1.70258e-06, 
    2.278583e-06, 2.183779e-06, 2.198249e-06, 2.426883e-06, 3.336262e-06, 
    1.96776e-06, 2.479218e-06, 3.737564e-06, 4.172846e-06, 3.695835e-06,
  1.544946e-05, 1.157456e-05, 1.025661e-05, 1.23445e-05, 5.339028e-06, 
    6.43768e-06, 7.632595e-06, 6.008725e-06, 5.65316e-06, 3.74252e-06, 
    5.862179e-06, 7.335539e-06, 6.443653e-06, 3.481412e-06, 4.165905e-06,
  9.280794e-06, 1.258969e-05, 1.385164e-05, 6.845406e-06, 6.121531e-06, 
    7.895575e-06, 5.164435e-06, 2.824304e-06, 4.435535e-06, 4.083615e-06, 
    5.035106e-06, 4.459827e-06, 3.522444e-06, 2.714405e-06, 2.51387e-06,
  1.476666e-05, 1.19789e-05, 7.980874e-06, 4.620356e-06, 6.136254e-06, 
    3.618204e-06, 4.725401e-06, 3.228378e-06, 2.983822e-06, 4.042933e-06, 
    4.809215e-06, 2.394721e-06, 2.518565e-06, 1.893179e-06, 1.296745e-06,
  9.496104e-06, 7.468308e-06, 4.10853e-06, 4.181457e-06, 4.160356e-06, 
    1.550187e-06, 3.523493e-06, 4.401204e-06, 4.586897e-06, 3.236078e-06, 
    3.345464e-06, 3.439256e-06, 1.891848e-06, 4.638412e-07, 3.878059e-07,
  7.339733e-06, 6.393541e-06, 3.546159e-06, 4.053072e-06, 3.486435e-06, 
    3.287055e-06, 3.247752e-06, 5.021147e-06, 3.745736e-06, 2.41981e-06, 
    9.280161e-07, 8.291629e-07, 1.619071e-06, 1.928813e-06, 1.878541e-06,
  7.099618e-06, 3.767077e-06, 3.389742e-06, 2.849491e-06, 3.537384e-06, 
    3.406084e-06, 3.341934e-06, 3.466329e-06, 2.342021e-06, 2.105947e-06, 
    1.875992e-06, 2.45105e-06, 3.800964e-06, 2.411299e-06, 2.884453e-06,
  3.908137e-06, 4.193461e-06, 3.426093e-06, 2.571056e-06, 3.868193e-06, 
    2.40689e-06, 2.337778e-06, 2.482198e-06, 3.19544e-06, 3.222938e-06, 
    3.114161e-06, 2.947789e-06, 3.373167e-06, 3.76102e-06, 4.10261e-06,
  3.860109e-06, 3.823592e-06, 2.743496e-06, 3.153317e-06, 1.954985e-06, 
    2.554509e-06, 2.251795e-06, 3.613053e-06, 4.140335e-06, 3.716022e-06, 
    3.047608e-06, 3.635482e-06, 3.14683e-06, 4.065484e-06, 3.761035e-06,
  2.978757e-06, 4.682037e-06, 2.775943e-06, 2.027286e-06, 3.11726e-06, 
    2.760733e-06, 2.669845e-06, 3.517878e-06, 3.764647e-06, 4.344795e-06, 
    3.993746e-06, 4.359641e-06, 3.852335e-06, 4.141904e-06, 7.400129e-06,
  4.621366e-06, 3.671594e-06, 3.203802e-06, 4.338404e-06, 2.8473e-06, 
    3.525038e-06, 2.930909e-06, 2.145543e-06, 5.394795e-06, 5.535483e-06, 
    6.170166e-06, 4.404656e-06, 3.813467e-06, 3.636931e-06, 4.322373e-06,
  0.0007083581, 0.0001909735, 2.409785e-05, 2.102794e-05, 1.146756e-05, 
    6.487877e-06, 5.846115e-06, 1.583746e-05, 1.107647e-05, 1.646408e-05, 
    1.837585e-05, 1.528321e-05, 1.242518e-05, 1.150062e-05, 1.004431e-05,
  0.0004404121, 7.469432e-05, 1.328729e-05, 1.250182e-05, 1.189704e-05, 
    8.562397e-06, 1.425421e-05, 1.741185e-05, 9.485215e-06, 1.153471e-05, 
    1.191544e-05, 1.049813e-05, 8.736925e-06, 1.060082e-05, 1.103282e-05,
  0.0001284566, 1.903496e-05, 1.059545e-05, 7.559179e-06, 5.222744e-06, 
    1.334616e-05, 1.081539e-05, 1.48128e-05, 7.131816e-06, 6.277188e-06, 
    8.686613e-06, 7.752985e-06, 6.808499e-06, 8.803555e-06, 1.02157e-05,
  2.77126e-05, 1.234451e-05, 7.297282e-06, 4.891874e-06, 6.528355e-06, 
    9.776707e-06, 1.119717e-05, 6.190435e-06, 5.217375e-06, 8.068366e-06, 
    8.676759e-06, 5.893389e-06, 8.773264e-06, 9.92359e-06, 1.067077e-05,
  8.893507e-06, 7.171791e-06, 3.440936e-06, 3.292297e-06, 6.626979e-06, 
    5.615015e-06, 5.530288e-06, 2.362672e-06, 3.785283e-06, 5.028604e-06, 
    7.037272e-06, 5.012347e-06, 8.854667e-06, 1.400672e-05, 1.440519e-05,
  5.350503e-06, 5.995595e-06, 1.922513e-06, 2.913159e-06, 3.5643e-06, 
    5.227473e-06, 5.274939e-06, 3.268774e-06, 7.419478e-06, 6.951808e-06, 
    7.708525e-06, 8.498624e-06, 1.140141e-05, 9.482033e-06, 1.366438e-05,
  4.779229e-06, 3.165187e-06, 1.351363e-06, 3.622768e-06, 3.674607e-06, 
    2.658934e-06, 4.843463e-06, 5.188889e-06, 9.236424e-06, 9.853028e-06, 
    1.160487e-05, 1.017951e-05, 6.325839e-06, 6.760777e-06, 8.959544e-06,
  1.645706e-06, 2.293892e-06, 2.426911e-06, 3.739472e-06, 3.040298e-06, 
    3.675256e-06, 3.901469e-06, 8.758098e-06, 1.108996e-05, 1.09099e-05, 
    1.105176e-05, 1.10466e-05, 8.533621e-06, 7.492832e-06, 4.184568e-06,
  3.077276e-06, 2.68232e-06, 1.414929e-06, 3.019353e-06, 4.776178e-06, 
    5.25597e-06, 7.228462e-06, 8.521902e-06, 1.226538e-05, 1.28487e-05, 
    7.778155e-06, 9.208818e-06, 5.120567e-06, 3.890187e-06, 3.538253e-06,
  1.587196e-06, 2.778086e-06, 4.707141e-06, 5.811567e-06, 7.83125e-06, 
    8.969349e-06, 9.898729e-06, 1.365525e-05, 1.272316e-05, 1.198318e-05, 
    1.027907e-05, 6.84349e-06, 3.644115e-06, 4.455028e-06, 1.361205e-05,
  0.0004076023, 0.0001103388, 3.970963e-05, 1.766716e-05, 2.564909e-06, 
    3.703084e-06, 4.333762e-06, 7.352128e-06, 6.770069e-06, 7.255312e-06, 
    6.94583e-06, 7.432351e-06, 1.229011e-05, 2.922288e-05, 1.583451e-05,
  0.0008297606, 0.0004819505, 0.0002077828, 3.804322e-05, 3.686238e-06, 
    3.176004e-06, 5.480646e-06, 7.984757e-06, 8.911237e-06, 7.056638e-06, 
    6.284214e-06, 7.023607e-06, 1.386463e-05, 2.745371e-05, 1.382198e-05,
  0.0009853321, 0.0007781625, 0.0005364515, 0.0001552208, 5.503079e-06, 
    3.233545e-06, 6.704498e-06, 7.227966e-06, 8.125903e-06, 7.159028e-06, 
    5.863074e-06, 8.74299e-06, 1.49317e-05, 2.342135e-05, 1.495047e-05,
  0.0008950953, 0.0008297953, 0.0007337934, 0.0004023315, 3.868193e-05, 
    3.399191e-06, 8.636157e-06, 7.726881e-06, 7.00612e-06, 5.676022e-06, 
    9.908709e-06, 1.278424e-05, 1.520098e-05, 2.433126e-05, 1.492172e-05,
  0.000662382, 0.0006880578, 0.000724206, 0.0005536584, 0.0001803871, 
    3.327755e-06, 8.718991e-06, 5.089876e-06, 6.534588e-06, 8.505e-06, 
    9.868429e-06, 1.223069e-05, 1.671916e-05, 2.552222e-05, 1.509723e-05,
  0.0004018963, 0.0004560518, 0.0006511721, 0.0006089342, 0.000310126, 
    3.780597e-06, 6.783589e-06, 6.495806e-06, 5.991572e-06, 6.946284e-06, 
    8.339995e-06, 9.832432e-06, 1.724893e-05, 2.644483e-05, 1.58331e-05,
  0.0002178331, 0.0003180883, 0.0005481345, 0.0006162026, 0.0003445728, 
    3.956054e-06, 6.67244e-06, 5.607319e-06, 6.393603e-06, 6.652379e-06, 
    9.097357e-06, 1.027437e-05, 1.585707e-05, 2.304534e-05, 1.54584e-05,
  0.0001361703, 0.0002574193, 0.0004754736, 0.0005645401, 0.0003240997, 
    3.418039e-06, 2.962735e-06, 2.934822e-06, 5.432475e-06, 7.351502e-06, 
    9.710318e-06, 1.01269e-05, 1.015331e-05, 1.865939e-05, 1.387915e-05,
  0.0001288222, 0.0002329853, 0.0003853581, 0.0004547873, 0.0002657567, 
    2.094459e-06, 1.719097e-06, 2.472141e-06, 5.71511e-06, 7.18301e-06, 
    7.497914e-06, 6.992576e-06, 9.861679e-06, 2.399465e-05, 1.820056e-05,
  0.0001226919, 0.0001797081, 0.0002573141, 0.0003073843, 0.0001773624, 
    2.27461e-06, 4.054329e-06, 4.74269e-06, 4.332465e-06, 5.163214e-06, 
    8.413203e-06, 1.239018e-05, 2.80181e-05, 6.576854e-05, 5.058491e-05,
  1.059014e-05, 8.185177e-06, 7.580225e-06, 8.688388e-06, 1.577031e-05, 
    1.696829e-05, 1.619405e-05, 1.767673e-05, 1.514339e-05, 1.394335e-05, 
    1.040916e-05, 7.169864e-06, 4.845248e-06, 5.533634e-06, 5.201407e-06,
  8.877895e-06, 6.81578e-06, 8.111747e-06, 7.432267e-06, 1.080457e-05, 
    1.331273e-05, 1.28986e-05, 1.280445e-05, 1.220897e-05, 1.110998e-05, 
    6.474256e-06, 4.822726e-06, 3.966681e-06, 4.510201e-06, 6.118749e-06,
  1.014411e-05, 7.993316e-06, 7.753541e-06, 8.955091e-06, 1.162582e-05, 
    1.343693e-05, 1.475304e-05, 1.186381e-05, 1.03586e-05, 1.061591e-05, 
    6.681961e-06, 4.697376e-06, 4.493864e-06, 3.078638e-06, 3.088011e-06,
  1.058177e-05, 8.498439e-06, 6.819926e-06, 7.460805e-06, 9.075616e-06, 
    1.099735e-05, 1.323846e-05, 1.159026e-05, 9.078338e-06, 7.68775e-06, 
    7.672033e-06, 4.749179e-06, 2.699636e-06, 1.79595e-06, 1.777214e-06,
  6.119246e-05, 1.985912e-05, 1.102469e-05, 8.116435e-06, 8.999216e-06, 
    8.181843e-06, 1.361106e-05, 1.185507e-05, 1.071182e-05, 8.099186e-06, 
    8.480614e-06, 2.869857e-06, 1.884902e-06, 1.680459e-06, 7.263133e-07,
  0.0001541757, 5.26579e-05, 3.134485e-05, 9.697595e-06, 5.794844e-06, 
    7.46988e-06, 1.253082e-05, 1.206371e-05, 1.133866e-05, 1.198012e-05, 
    7.40261e-06, 2.267282e-06, 1.256432e-06, 6.959595e-07, 5.383766e-07,
  0.0002484269, 0.0001149031, 6.915989e-05, 2.288561e-05, 8.042187e-06, 
    6.797899e-06, 1.698803e-05, 1.085177e-05, 1.284547e-05, 9.636115e-06, 
    5.207355e-06, 2.214789e-06, 3.098707e-07, 3.046221e-07, 3.46221e-08,
  0.0003100692, 0.0001729076, 0.0001226161, 5.146555e-05, 5.690126e-06, 
    5.178407e-06, 9.505982e-06, 4.966664e-06, 7.148892e-06, 1.029466e-05, 
    4.12595e-06, 1.184819e-06, 5.608862e-07, 3.530995e-07, 5.282445e-07,
  0.0003358186, 0.0002310625, 0.0002057185, 0.0001061252, 1.189709e-05, 
    3.827578e-06, 7.884682e-06, 7.284391e-06, 9.956255e-06, 3.774964e-06, 
    2.086788e-06, 6.327409e-07, 2.687568e-07, 7.385293e-07, 2.584411e-06,
  0.0003879038, 0.0003308832, 0.0003193189, 0.0001785839, 3.413125e-05, 
    4.7024e-06, 6.735035e-06, 8.686568e-06, 6.660808e-06, 4.378399e-06, 
    2.705477e-06, 4.264062e-07, 1.142877e-06, 2.85878e-06, 1.636584e-06,
  8.230715e-06, 7.851639e-06, 7.393401e-06, 7.73864e-06, 9.618012e-06, 
    7.903797e-06, 7.741621e-06, 3.966645e-06, 1.012644e-06, 9.617033e-07, 
    1.725336e-06, 2.617751e-06, 3.066313e-06, 5.412719e-06, 5.651765e-06,
  6.654485e-06, 5.151559e-06, 4.263647e-06, 3.739186e-06, 4.265218e-06, 
    5.8384e-06, 1.251379e-06, 1.036907e-06, 2.571611e-06, 2.64725e-06, 
    2.259808e-06, 3.581725e-06, 4.840531e-06, 5.21131e-06, 7.089562e-06,
  5.978155e-06, 5.11031e-06, 3.565165e-06, 2.121238e-06, 4.100549e-06, 
    3.629225e-06, 7.917374e-07, 1.747673e-06, 2.200285e-06, 1.764667e-06, 
    2.426992e-06, 1.348103e-06, 1.501502e-06, 1.416185e-06, 1.554652e-06,
  6.074976e-06, 5.878157e-06, 2.395877e-06, 2.163788e-06, 2.070872e-06, 
    2.603089e-06, 5.884146e-06, 4.894839e-06, 3.276119e-06, 2.54868e-06, 
    2.456136e-06, 2.404755e-06, 2.448407e-06, 3.548155e-06, 3.802479e-06,
  6.039885e-06, 3.776972e-06, 3.852341e-06, 2.963336e-06, 3.203482e-06, 
    2.832809e-06, 4.545722e-06, 6.616263e-06, 7.897247e-06, 7.002722e-06, 
    4.020785e-06, 4.630054e-06, 2.952051e-06, 3.694636e-06, 3.914244e-06,
  7.169964e-06, 5.331406e-06, 5.334583e-06, 3.731293e-06, 3.802358e-06, 
    8.162984e-06, 9.611172e-06, 8.81682e-06, 8.994476e-06, 9.525515e-06, 
    6.389816e-06, 5.408229e-06, 4.889692e-06, 5.655419e-06, 3.386182e-06,
  9.205341e-06, 1.062448e-05, 8.18574e-06, 9.839515e-06, 1.090217e-05, 
    1.217038e-05, 1.175385e-05, 1.239756e-05, 1.306487e-05, 1.049596e-05, 
    9.553075e-06, 9.13165e-06, 7.616316e-06, 5.70501e-06, 5.974603e-06,
  1.284141e-05, 1.18283e-05, 1.486476e-05, 1.203218e-05, 1.005064e-05, 
    1.418347e-05, 1.201361e-05, 1.429e-05, 1.659879e-05, 1.693729e-05, 
    1.537678e-05, 1.340788e-05, 1.321479e-05, 1.327408e-05, 9.518974e-06,
  1.27e-05, 1.325336e-05, 1.705365e-05, 1.610507e-05, 1.44451e-05, 
    1.316467e-05, 1.586595e-05, 1.821898e-05, 2.154692e-05, 2.424827e-05, 
    2.162476e-05, 1.893496e-05, 1.988648e-05, 1.559712e-05, 1.480427e-05,
  9.601145e-06, 1.399697e-05, 1.748686e-05, 1.768125e-05, 1.608653e-05, 
    1.905237e-05, 2.264828e-05, 2.19718e-05, 2.539734e-05, 2.940134e-05, 
    2.676857e-05, 2.776249e-05, 2.505896e-05, 2.464828e-05, 1.969173e-05,
  1.93743e-06, 1.790077e-06, 1.81875e-06, 4.017773e-06, 1.81503e-06, 
    5.275356e-06, 4.789695e-06, 3.398159e-06, 3.59555e-06, 1.956498e-06, 
    1.613197e-06, 6.256447e-07, 6.094431e-07, 6.719191e-07, 7.23431e-07,
  8.256325e-07, 2.108983e-06, 2.320903e-06, 2.290195e-06, 3.400786e-06, 
    3.258739e-06, 6.390581e-07, 4.197721e-07, 7.538277e-07, 1.099782e-06, 
    5.15503e-07, 4.505889e-07, 1.875407e-07, 1.016494e-07, 1.737011e-07,
  4.94342e-07, 8.623561e-07, 4.897542e-07, 3.432809e-07, 4.58276e-07, 
    1.668342e-07, 5.302708e-07, 6.86743e-07, 8.626512e-07, 1.214944e-06, 
    1.27862e-06, 1.488309e-06, 1.043314e-06, 9.364082e-07, 6.181594e-07,
  4.452637e-07, 4.236828e-07, 2.050795e-07, 2.145128e-07, 2.6565e-07, 
    2.344678e-07, 7.013851e-07, 1.502738e-06, 1.832931e-06, 2.5414e-06, 
    3.278728e-06, 3.256988e-06, 3.40125e-06, 2.855835e-06, 1.818124e-06,
  6.874785e-07, 2.826781e-07, 1.514653e-07, 2.028601e-07, 6.591712e-07, 
    1.131145e-06, 1.846665e-06, 2.28939e-06, 4.092815e-06, 4.49969e-06, 
    3.741885e-06, 3.824648e-06, 5.334736e-06, 4.536654e-06, 3.743804e-06,
  4.025907e-07, 2.981878e-07, 5.073614e-08, 5.706599e-07, 1.99632e-06, 
    1.793416e-06, 3.538692e-06, 5.382105e-06, 5.623386e-06, 4.984141e-06, 
    3.840486e-06, 5.20119e-06, 6.17349e-06, 8.498376e-06, 8.791512e-06,
  8.120977e-07, 5.77774e-07, 9.141188e-08, 4.529038e-07, 3.038169e-06, 
    4.647516e-06, 7.115628e-06, 6.291477e-06, 8.782631e-06, 8.158648e-06, 
    9.837231e-06, 8.848519e-06, 1.056024e-05, 1.088824e-05, 1.194584e-05,
  1.339182e-06, 1.076364e-06, 7.324008e-07, 9.222758e-07, 3.348084e-06, 
    5.065742e-06, 6.845572e-06, 8.428537e-06, 9.418256e-06, 1.251674e-05, 
    1.400675e-05, 1.540552e-05, 1.546531e-05, 1.347525e-05, 1.356167e-05,
  2.325555e-06, 1.393244e-06, 1.324351e-06, 2.828384e-06, 4.902049e-06, 
    7.08616e-06, 8.660234e-06, 9.474856e-06, 1.077442e-05, 1.334702e-05, 
    1.522607e-05, 1.441664e-05, 1.532384e-05, 1.6061e-05, 1.481394e-05,
  3.318443e-06, 1.578604e-06, 3.651643e-06, 6.125841e-06, 6.05458e-06, 
    7.111163e-06, 9.506236e-06, 1.187434e-05, 1.363891e-05, 1.778749e-05, 
    1.526054e-05, 1.782874e-05, 1.572442e-05, 1.568092e-05, 1.348664e-05,
  2.23664e-06, 4.120317e-06, 2.043255e-06, 2.39045e-06, 1.285694e-06, 
    1.602163e-06, 1.089292e-06, 1.500625e-07, 1.768751e-07, 9.228949e-08, 
    1.512409e-07, 1.333738e-06, 1.349487e-06, 1.807551e-06, 9.250314e-07,
  4.221889e-06, 7.73642e-06, 5.574406e-06, 3.359377e-06, 3.099558e-06, 
    2.805018e-06, 2.592333e-06, 2.075048e-06, 4.865715e-07, 1.183752e-06, 
    1.415193e-06, 3.233616e-07, 1.210857e-06, 2.133468e-06, 2.635324e-06,
  1.053438e-05, 9.391052e-06, 7.608051e-06, 7.321873e-06, 5.456876e-06, 
    6.865279e-06, 5.669534e-06, 4.479082e-06, 5.376866e-06, 4.327867e-06, 
    2.831098e-06, 3.353265e-06, 1.774254e-06, 2.054848e-06, 1.321528e-06,
  1.923347e-05, 1.531548e-05, 1.185278e-05, 9.95071e-06, 8.997437e-06, 
    9.599893e-06, 9.342518e-06, 7.513233e-06, 6.963201e-06, 5.075473e-06, 
    5.18233e-06, 4.465099e-06, 3.132443e-06, 2.348494e-06, 1.109464e-06,
  2.595281e-05, 1.960166e-05, 1.808695e-05, 1.963683e-05, 1.259487e-05, 
    1.100856e-05, 9.653241e-06, 8.124084e-06, 6.514305e-06, 5.295765e-06, 
    4.744256e-06, 3.244545e-06, 2.384745e-06, 1.882601e-06, 1.685532e-06,
  3.256636e-05, 3.098785e-05, 2.687987e-05, 2.480461e-05, 2.38326e-05, 
    1.334683e-05, 1.24384e-05, 8.648066e-06, 7.429409e-06, 5.171784e-06, 
    3.978144e-06, 3.15372e-06, 2.70307e-06, 3.194039e-06, 2.694165e-06,
  4.518973e-05, 4.411886e-05, 3.621034e-05, 3.948732e-05, 2.64612e-05, 
    2.865859e-05, 1.484886e-05, 9.847624e-06, 9.240136e-06, 7.016046e-06, 
    4.701998e-06, 5.009786e-06, 3.400324e-06, 3.351278e-06, 2.736567e-06,
  6.560612e-05, 6.818154e-05, 4.91291e-05, 4.608914e-05, 4.383435e-05, 
    3.699137e-05, 2.465641e-05, 2.049707e-05, 1.242035e-05, 9.54389e-06, 
    6.467913e-06, 5.18039e-06, 5.001069e-06, 4.285871e-06, 3.497754e-06,
  7.586996e-05, 8.420464e-05, 7.434619e-05, 6.270249e-05, 6.134907e-05, 
    4.632549e-05, 3.796536e-05, 2.935893e-05, 2.884019e-05, 2.043794e-05, 
    1.086986e-05, 7.302997e-06, 6.147086e-06, 4.059019e-06, 3.168883e-06,
  0.0001156108, 8.929698e-05, 8.999148e-05, 8.658683e-05, 7.36096e-05, 
    7.132539e-05, 5.196531e-05, 4.407873e-05, 4.289576e-05, 3.215106e-05, 
    2.215327e-05, 1.473717e-05, 7.977193e-06, 5.313047e-06, 3.578622e-06,
  8.490856e-08, 1.782639e-07, 2.281614e-08, 7.395727e-08, 1.81464e-07, 
    1.527552e-06, 4.983079e-06, 7.326818e-06, 1.035809e-05, 3.310243e-05, 
    5.924145e-05, 8.849792e-05, 0.0001322512, 0.0001800198, 0.000266398,
  6.631745e-07, 7.587146e-07, 4.740432e-08, 3.263601e-08, 3.873099e-08, 
    1.357789e-07, 1.407871e-06, 2.715932e-06, 4.281939e-06, 1.413783e-05, 
    2.581154e-05, 3.336798e-05, 5.278847e-05, 9.466276e-05, 0.0001335484,
  4.427662e-07, 1.13637e-07, 4.67361e-08, 4.36536e-08, 5.225457e-08, 
    3.205318e-08, 9.534544e-08, 3.851721e-07, 3.5467e-06, 3.689323e-06, 
    7.406249e-06, 1.499329e-05, 2.136798e-05, 3.936179e-05, 6.262676e-05,
  3.329462e-06, 1.176845e-06, 8.31188e-07, 4.663105e-08, 6.592803e-08, 
    6.581853e-07, 1.274521e-07, 1.431306e-07, 1.206367e-07, 1.005008e-07, 
    2.680578e-06, 4.739381e-06, 7.726638e-06, 1.390439e-05, 1.805671e-05,
  6.249892e-06, 6.279141e-06, 1.65956e-06, 1.425077e-06, 2.257912e-06, 
    1.700815e-07, 7.555868e-07, 1.780917e-07, 3.346065e-07, 1.443011e-07, 
    1.195694e-07, 1.665473e-06, 2.60617e-06, 3.90759e-06, 6.148637e-06,
  1.105457e-05, 1.254258e-05, 6.624632e-06, 4.485406e-06, 3.064534e-06, 
    2.522669e-06, 9.408092e-07, 7.45796e-07, 6.08031e-07, 2.502929e-07, 
    1.066217e-08, 2.934746e-09, 5.967598e-08, 2.620925e-07, 4.094395e-07,
  1.546717e-05, 1.857688e-05, 1.441377e-05, 1.004233e-05, 9.04465e-06, 
    5.184782e-06, 4.086976e-06, 1.909839e-06, 1.314523e-06, 2.513683e-07, 
    7.605559e-07, 9.60602e-09, 1.552388e-08, 1.740679e-08, 3.910559e-08,
  2.079844e-05, 2.179701e-05, 1.849254e-05, 1.494668e-05, 1.321842e-05, 
    1.12889e-05, 6.532176e-06, 4.469768e-06, 3.04715e-06, 1.670053e-06, 
    1.225814e-06, 3.386225e-07, 4.947313e-07, 7.506918e-08, 1.590774e-08,
  2.596535e-05, 2.812159e-05, 2.386514e-05, 2.158328e-05, 1.784165e-05, 
    1.726945e-05, 1.046958e-05, 9.638095e-06, 4.778473e-06, 2.35263e-06, 
    3.018753e-06, 1.257418e-06, 9.372494e-07, 9.246626e-07, 2.421828e-07,
  3.172652e-05, 3.409886e-05, 3.126674e-05, 2.733667e-05, 2.139174e-05, 
    1.720436e-05, 1.357297e-05, 1.811556e-05, 8.347799e-06, 6.747467e-06, 
    5.335872e-06, 2.758768e-06, 2.224175e-06, 1.924257e-06, 1.65757e-06,
  4.880695e-06, 1.973993e-05, 5.58605e-05, 0.000105618, 0.000138937, 
    0.0001537672, 0.0001683319, 0.0001684698, 0.0001612604, 0.0001561059, 
    0.0001451305, 0.0001328764, 0.0001300863, 0.0001430543, 0.0001651588,
  2.958514e-06, 5.507943e-06, 1.533434e-05, 4.817309e-05, 9.370343e-05, 
    0.0001230987, 0.0001390241, 0.0001509767, 0.000158793, 0.0001589181, 
    0.0001587484, 0.0001532083, 0.000142573, 0.0001386661, 0.0001459128,
  1.895311e-06, 3.039812e-06, 2.838427e-06, 8.245333e-06, 2.448436e-05, 
    5.926691e-05, 9.814218e-05, 0.0001234101, 0.000142905, 0.000165127, 
    0.0001754919, 0.0001969989, 0.000194482, 0.0002044288, 0.0001872564,
  5.349562e-06, 3.468498e-06, 2.846554e-06, 3.301583e-06, 2.308318e-06, 
    4.547855e-06, 1.565869e-05, 3.633056e-05, 6.571531e-05, 9.87515e-05, 
    0.0001284664, 0.0001559391, 0.0001778655, 0.0001994499, 0.0002213083,
  7.360822e-06, 6.662553e-06, 6.410443e-06, 3.100304e-06, 4.659029e-06, 
    5.100513e-06, 4.125126e-06, 4.059043e-06, 7.616719e-06, 1.765438e-05, 
    3.64087e-05, 5.984592e-05, 9.004075e-05, 0.0001223646, 0.0001385782,
  8.865306e-06, 8.428717e-06, 6.866603e-06, 5.335986e-06, 4.221156e-06, 
    4.923315e-06, 4.772428e-06, 4.695489e-06, 4.001799e-06, 4.989715e-06, 
    4.237693e-06, 1.003596e-05, 2.090567e-05, 3.980183e-05, 5.534875e-05,
  1.083264e-05, 1.023385e-05, 8.903438e-06, 7.175032e-06, 4.88e-06, 
    5.023789e-06, 4.107515e-06, 5.132465e-06, 5.554713e-06, 4.423893e-06, 
    3.789235e-06, 1.346488e-06, 4.372318e-06, 7.156955e-06, 1.186745e-05,
  1.353642e-05, 1.12129e-05, 1.077423e-05, 8.062295e-06, 6.517972e-06, 
    5.183304e-06, 4.810042e-06, 4.750993e-06, 5.284379e-06, 4.931102e-06, 
    5.104763e-06, 5.316972e-06, 3.996949e-06, 3.096767e-06, 3.614167e-06,
  1.810988e-05, 1.625537e-05, 1.401999e-05, 1.078098e-05, 8.100824e-06, 
    5.964389e-06, 4.256412e-06, 4.928062e-06, 5.331205e-06, 5.066096e-06, 
    4.53423e-06, 5.024735e-06, 5.630054e-06, 4.881019e-06, 3.550496e-06,
  1.960459e-05, 1.986802e-05, 1.800436e-05, 1.472807e-05, 1.151777e-05, 
    7.497536e-06, 5.849452e-06, 5.490835e-06, 4.26626e-06, 4.712971e-06, 
    5.595176e-06, 3.105411e-06, 4.872519e-06, 6.290064e-06, 6.269732e-06,
  0.0003859893, 0.0003529299, 0.0002823983, 0.0001936218, 0.0001040425, 
    5.275485e-05, 2.962898e-05, 1.676591e-05, 1.937847e-05, 1.826931e-05, 
    1.515575e-05, 1.481211e-05, 2.497185e-05, 2.135588e-05, 1.318761e-05,
  0.0003753502, 0.0004045195, 0.0003719371, 0.0003224884, 0.0002319667, 
    0.0001564037, 0.0001017003, 6.736418e-05, 4.442213e-05, 3.991314e-05, 
    2.560343e-05, 1.90906e-05, 1.957087e-05, 2.950422e-05, 3.606286e-05,
  0.0003094438, 0.00032334, 0.0003278744, 0.0003295788, 0.0003079008, 
    0.0002722937, 0.0002360331, 0.0002076559, 0.0001694085, 0.0001094443, 
    6.259971e-05, 3.474395e-05, 2.343082e-05, 2.136384e-05, 3.877472e-05,
  0.0002061462, 0.0002256636, 0.0002468977, 0.0002477437, 0.00024101, 
    0.0002643622, 0.0002814972, 0.000284643, 0.0002881444, 0.0002485171, 
    0.0001849543, 0.000104748, 5.952606e-05, 4.24257e-05, 3.906778e-05,
  0.0001692886, 0.0001822087, 0.0001967199, 0.0001818566, 0.0001590527, 
    0.0001722468, 0.0002081155, 0.0002663476, 0.0002988276, 0.0002964184, 
    0.0002727982, 0.0002274765, 0.0001697488, 0.0001050783, 7.676845e-05,
  0.0001420278, 0.0001600851, 0.0001728745, 0.0001616699, 0.0001303987, 
    0.0001103007, 0.0001247399, 0.0001792704, 0.0002256659, 0.0002429184, 
    0.0002478759, 0.0002202649, 0.0002074206, 0.0001937123, 0.000162069,
  0.0001166919, 0.0001179067, 0.0001082756, 0.0001127952, 0.0001023978, 
    8.838905e-05, 9.732772e-05, 0.0001389913, 0.0001747311, 0.0001760758, 
    0.0001609398, 0.0001355084, 0.0001276117, 0.0001484445, 0.0001695124,
  5.232654e-05, 5.550817e-05, 5.148867e-05, 5.400372e-05, 5.008537e-05, 
    4.246195e-05, 4.800044e-05, 7.486809e-05, 0.0001201869, 0.0001458654, 
    0.000136234, 0.0001075926, 8.936244e-05, 7.639472e-05, 8.250874e-05,
  9.033008e-06, 1.152599e-05, 1.048477e-05, 1.283442e-05, 1.153053e-05, 
    8.42018e-06, 1.129874e-05, 2.059156e-05, 5.64647e-05, 9.122652e-05, 
    9.443611e-05, 7.762128e-05, 5.980951e-05, 5.184385e-05, 4.560731e-05,
  4.221865e-06, 5.891628e-06, 4.309899e-06, 3.43398e-06, 5.890996e-06, 
    5.845491e-06, 4.365052e-06, 6.28927e-06, 1.53925e-05, 3.911207e-05, 
    5.207902e-05, 4.478593e-05, 3.369416e-05, 2.733504e-05, 2.255985e-05,
  3.896904e-05, 5.032365e-05, 7.373425e-06, 1.4398e-05, 4.878772e-05, 
    4.374217e-05, 5.122571e-05, 3.873718e-05, 5.798728e-05, 6.819054e-05, 
    4.581437e-05, 1.858986e-05, 1.569685e-05, 2.207878e-05, 1.00732e-05,
  3.511335e-05, 1.081127e-05, 1.342871e-05, 2.300788e-05, 5.577306e-05, 
    0.0001244494, 4.119963e-05, 2.125559e-05, 8.727538e-05, 2.936375e-05, 
    4.695552e-05, 1.233576e-05, 2.328352e-05, 1.109137e-05, 1.005952e-05,
  3.83726e-05, 1.915021e-05, 1.153163e-05, 1.473681e-05, 3.662912e-05, 
    0.0001279406, 2.710153e-05, 1.888602e-05, 3.059159e-05, 2.535339e-05, 
    1.253857e-05, 1.955275e-05, 1.672816e-05, 1.688998e-05, 8.312941e-06,
  1.707767e-05, 1.480354e-05, 1.569913e-05, 1.580118e-05, 3.037068e-05, 
    3.713535e-05, 2.335892e-05, 2.024233e-05, 1.711979e-05, 6.636534e-06, 
    1.425911e-05, 1.931437e-05, 2.089969e-05, 2.039967e-05, 1.762556e-05,
  2.772944e-05, 2.652195e-05, 2.014981e-05, 1.715913e-05, 2.123064e-05, 
    2.607358e-05, 1.839555e-05, 2.745449e-05, 7.508448e-06, 1.124274e-05, 
    1.661279e-05, 2.086472e-05, 1.805065e-05, 1.823001e-05, 2.355894e-05,
  5.28232e-05, 4.198274e-05, 3.715435e-05, 3.221156e-05, 2.997826e-05, 
    2.348997e-05, 1.964894e-05, 1.229497e-05, 1.174225e-05, 1.431084e-05, 
    1.93148e-05, 2.135994e-05, 2.117604e-05, 2.639067e-05, 2.612311e-05,
  8.404681e-05, 7.207046e-05, 7.208464e-05, 6.605949e-05, 6.029183e-05, 
    4.959658e-05, 3.238465e-05, 1.940105e-05, 1.574804e-05, 1.383041e-05, 
    1.409281e-05, 1.672587e-05, 2.352442e-05, 2.341632e-05, 1.977698e-05,
  9.54408e-05, 9.795731e-05, 0.0001022009, 9.830183e-05, 9.562029e-05, 
    7.63958e-05, 5.723658e-05, 3.849016e-05, 3.209608e-05, 2.364845e-05, 
    1.873549e-05, 1.623918e-05, 1.984414e-05, 1.632181e-05, 1.366215e-05,
  8.582265e-05, 9.335668e-05, 9.8497e-05, 0.0001042447, 9.209261e-05, 
    7.095671e-05, 5.383139e-05, 4.550294e-05, 5.026233e-05, 5.230548e-05, 
    4.471339e-05, 3.024865e-05, 2.62622e-05, 2.260014e-05, 1.942585e-05,
  6.494114e-05, 7.733431e-05, 8.104569e-05, 9.042312e-05, 8.358958e-05, 
    6.41993e-05, 4.617463e-05, 4.110279e-05, 5.331231e-05, 7.278602e-05, 
    7.352134e-05, 5.038063e-05, 4.093794e-05, 4.150683e-05, 3.770377e-05,
  2.743469e-05, 2.024028e-05, 2.044612e-05, 1.41272e-05, 1.279249e-05, 
    1.066615e-05, 2.81082e-06, 3.154421e-06, 2.75098e-06, 9.125996e-06, 
    1.328394e-05, 2.056301e-05, 2.936917e-05, 1.619894e-05, 1.406679e-05,
  1.773843e-05, 3.701801e-05, 2.87554e-05, 1.307205e-05, 1.564147e-05, 
    8.688166e-06, 5.803954e-06, 5.055399e-06, 5.360858e-06, 2.934188e-06, 
    1.388874e-06, 3.676236e-06, 1.718764e-06, 6.967432e-06, 1.358426e-05,
  1.42339e-05, 3.024522e-05, 3.901607e-05, 3.529747e-05, 2.652201e-05, 
    3.242841e-05, 8.427835e-06, 7.171655e-06, 1.396273e-05, 6.769929e-06, 
    2.866833e-06, 2.470244e-06, 1.857972e-06, 2.845159e-06, 7.030624e-06,
  2.906312e-05, 3.529639e-05, 3.98439e-05, 1.657367e-05, 2.212403e-05, 
    2.746106e-05, 1.518989e-05, 9.62065e-06, 1.774985e-05, 1.096624e-05, 
    6.999552e-06, 4.848167e-06, 3.772481e-06, 2.857243e-06, 3.368767e-06,
  3.348281e-05, 2.888174e-05, 1.947551e-05, 1.739819e-05, 2.968772e-05, 
    2.243078e-05, 2.408205e-05, 1.475375e-05, 1.405788e-05, 8.887778e-06, 
    1.071556e-05, 7.635773e-06, 3.902184e-06, 4.214766e-06, 3.538327e-06,
  2.36414e-05, 1.723991e-05, 3.118738e-05, 2.358543e-05, 3.983084e-05, 
    2.754106e-05, 2.964445e-05, 1.594988e-05, 1.019635e-05, 1.535917e-05, 
    9.463269e-06, 6.108658e-06, 5.17561e-06, 5.651133e-06, 3.70494e-06,
  9.474797e-06, 1.481731e-05, 3.31646e-05, 2.802007e-05, 4.48129e-05, 
    2.779638e-05, 1.332826e-05, 8.750926e-06, 1.569747e-05, 2.061485e-05, 
    1.31399e-05, 8.459744e-06, 1.042562e-05, 8.626292e-06, 8.287365e-06,
  9.518911e-06, 1.431198e-05, 2.983056e-05, 4.031045e-05, 3.22823e-05, 
    3.716775e-05, 1.183391e-05, 1.267571e-05, 2.017933e-05, 1.704143e-05, 
    1.64848e-05, 1.453801e-05, 9.676882e-06, 1.137853e-05, 2.018829e-05,
  8.894693e-06, 4.206925e-06, 1.582369e-05, 2.663031e-05, 3.770446e-05, 
    3.522108e-05, 9.931065e-06, 1.461449e-05, 1.066526e-05, 1.52972e-05, 
    1.799078e-05, 1.484026e-05, 1.581571e-05, 2.819026e-05, 4.444407e-05,
  8.381279e-06, 4.51197e-06, 8.081233e-06, 2.167722e-05, 1.728032e-05, 
    1.751992e-05, 8.438473e-06, 8.282981e-06, 1.244515e-05, 1.278982e-05, 
    1.037368e-05, 1.270368e-05, 1.732502e-05, 3.329029e-05, 4.855458e-05,
  1.374609e-05, 1.685746e-05, 2.460935e-05, 4.557015e-05, 4.474304e-05, 
    5.75506e-05, 7.524778e-05, 7.822586e-05, 7.627043e-05, 6.808005e-05, 
    5.230953e-05, 4.435002e-05, 3.892314e-05, 2.15146e-05, 1.114247e-05,
  7.400718e-06, 1.185775e-05, 2.160532e-05, 3.834197e-05, 2.679421e-05, 
    4.780171e-05, 4.731588e-05, 8.022665e-05, 7.293295e-05, 6.022379e-05, 
    6.774555e-05, 4.997114e-05, 4.695249e-05, 4.453991e-05, 1.676119e-05,
  1.11143e-06, 1.59111e-05, 1.283974e-05, 3.980062e-05, 3.816608e-05, 
    4.27289e-05, 4.476506e-05, 7.346481e-05, 7.608339e-05, 5.674873e-05, 
    4.072786e-05, 7.074102e-05, 4.594361e-05, 3.962896e-05, 3.734676e-05,
  3.929629e-07, 6.386127e-07, 7.45569e-06, 2.582704e-05, 2.655661e-05, 
    4.091233e-05, 4.550891e-05, 5.236109e-05, 6.87158e-05, 5.596537e-05, 
    5.578197e-05, 4.824511e-05, 5.566669e-05, 4.903944e-05, 3.257496e-05,
  9.633231e-07, 1.141798e-06, 3.186505e-06, 1.206389e-05, 3.233911e-05, 
    1.818179e-05, 2.846804e-05, 4.351025e-05, 5.531314e-05, 5.526789e-05, 
    5.182358e-05, 4.860886e-05, 6.836693e-05, 9.042983e-05, 8.179465e-05,
  2.178532e-06, 1.854617e-06, 2.249245e-06, 7.84058e-06, 1.284168e-05, 
    7.176201e-06, 1.83787e-05, 3.25877e-05, 4.588356e-05, 4.309238e-05, 
    3.705516e-05, 4.814981e-05, 8.748528e-05, 0.000118223, 9.167054e-05,
  5.560581e-06, 1.863339e-06, 4.493484e-06, 3.635162e-06, 2.513532e-06, 
    3.022609e-06, 7.672358e-06, 1.230346e-05, 7.67059e-06, 2.824194e-05, 
    2.554062e-05, 3.958665e-05, 7.569363e-05, 8.022352e-05, 5.893963e-05,
  9.227862e-06, 4.458981e-06, 4.340102e-06, 6.907487e-06, 3.866129e-06, 
    1.905266e-06, 3.462368e-06, 4.167915e-06, 1.141376e-05, 1.381627e-05, 
    1.034288e-05, 1.129071e-05, 3.104305e-05, 3.952841e-05, 6.27082e-05,
  1.270946e-05, 1.287694e-05, 7.411429e-06, 8.710514e-06, 1.164244e-05, 
    3.749598e-06, 3.452906e-06, 2.221911e-06, 2.967837e-06, 2.24971e-06, 
    2.791854e-06, 1.334774e-06, 3.848507e-06, 7.319924e-06, 1.233124e-05,
  1.761873e-05, 1.505915e-05, 7.031056e-06, 1.176484e-05, 1.681334e-05, 
    1.368997e-05, 2.859638e-06, 3.325893e-06, 2.420698e-06, 3.952374e-06, 
    3.517438e-06, 3.236827e-06, 1.186743e-06, 1.552686e-06, 2.26095e-06,
  7.335533e-05, 4.89765e-05, 7.162388e-05, 5.343244e-05, 3.336707e-05, 
    1.789401e-05, 1.91433e-05, 3.78783e-05, 9.76405e-05, 0.0001000674, 
    4.247779e-05, 3.32084e-05, 2.401243e-05, 1.979496e-05, 1.661839e-05,
  8.036374e-05, 7.752936e-05, 6.135398e-05, 5.538061e-05, 5.467203e-05, 
    3.106973e-05, 2.644607e-05, 5.288987e-05, 7.663217e-05, 4.231848e-05, 
    3.384772e-05, 2.657611e-05, 2.711537e-05, 1.804032e-05, 1.44586e-05,
  5.643312e-05, 6.215467e-05, 6.691477e-05, 5.133976e-05, 4.907938e-05, 
    3.509086e-05, 2.437018e-05, 3.944398e-05, 3.844052e-05, 2.594265e-05, 
    2.923489e-05, 3.249191e-05, 3.265079e-05, 3.932881e-05, 4.867338e-05,
  8.283454e-05, 8.129347e-05, 0.0001007983, 8.221131e-05, 4.750955e-05, 
    4.265597e-05, 3.019774e-05, 3.786712e-05, 2.728551e-05, 2.002306e-05, 
    2.314784e-05, 4.000002e-05, 6.189938e-05, 8.990549e-05, 8.620699e-05,
  3.349513e-05, 0.0001144478, 0.0001486658, 8.314253e-05, 7.556753e-05, 
    5.576609e-05, 5.782116e-05, 2.763666e-05, 2.02345e-05, 1.735995e-05, 
    3.100914e-05, 4.648452e-05, 5.796953e-05, 8.118746e-05, 7.157299e-05,
  1.420969e-05, 4.501216e-05, 8.020641e-05, 0.0001219066, 8.625212e-05, 
    5.653231e-05, 8.36886e-05, 3.760895e-05, 3.177411e-05, 3.791431e-05, 
    3.314256e-05, 3.331694e-05, 5.273108e-05, 4.771957e-05, 4.813749e-05,
  2.750423e-06, 6.970575e-06, 8.424891e-05, 7.407197e-05, 0.0001222774, 
    5.871228e-05, 5.197727e-05, 6.822632e-05, 4.997651e-05, 5.106574e-05, 
    4.755956e-05, 3.860011e-05, 5.124702e-05, 4.589544e-05, 5.197392e-05,
  1.209886e-06, 1.275824e-06, 6.22478e-06, 9.217792e-05, 0.0001292338, 
    5.633019e-05, 8.721445e-05, 0.0001057733, 5.100515e-05, 3.653466e-05, 
    4.402694e-05, 6.086686e-05, 5.256855e-05, 5.91281e-05, 5.166447e-05,
  1.063095e-06, 1.713619e-07, 1.2723e-06, 2.115191e-05, 6.862987e-05, 
    4.07575e-05, 4.107722e-05, 8.407036e-05, 7.717531e-05, 1.464667e-05, 
    1.608215e-05, 3.36102e-05, 4.275535e-05, 7.236206e-05, 5.661231e-05,
  6.335432e-07, 2.287515e-07, 1.545199e-06, 9.760241e-07, 2.04891e-05, 
    2.897679e-05, 5.130918e-05, 5.847854e-05, 9.563098e-05, 1.25843e-05, 
    4.500198e-06, 9.450267e-06, 3.225968e-05, 3.659913e-05, 4.906839e-05,
  4.466659e-07, 1.140975e-06, 2.335857e-06, 2.795139e-06, 5.671096e-06, 
    1.374525e-05, 8.573385e-06, 4.216837e-06, 6.84991e-06, 1.840224e-05, 
    1.253853e-05, 1.651002e-05, 2.01745e-05, 2.732172e-05, 3.241625e-05,
  3.395989e-07, 7.693926e-07, 1.981675e-06, 3.234783e-06, 6.393396e-06, 
    1.935486e-05, 1.96305e-05, 4.907678e-06, 2.941193e-06, 4.056368e-06, 
    7.703574e-06, 1.133034e-05, 8.996078e-06, 8.7563e-06, 1.39012e-05,
  1.466431e-05, 6.520073e-07, 1.217099e-06, 3.281399e-06, 6.341108e-06, 
    2.028355e-05, 5.178606e-05, 1.224047e-05, 5.195148e-06, 6.81137e-06, 
    6.96566e-06, 4.592989e-06, 3.694702e-06, 2.049984e-06, 1.01623e-06,
  3.460794e-05, 2.286912e-05, 2.446429e-06, 3.713851e-06, 6.508702e-06, 
    2.205004e-05, 4.876412e-05, 2.616071e-05, 1.341559e-05, 1.028332e-05, 
    1.002686e-05, 9.929932e-06, 8.118761e-06, 6.127005e-06, 3.305047e-06,
  0.0001173381, 3.686639e-05, 1.384285e-05, 1.921997e-06, 7.437957e-06, 
    1.929531e-05, 4.183598e-05, 4.106776e-05, 2.911985e-05, 1.5827e-05, 
    2.026975e-05, 1.660125e-05, 1.304333e-05, 9.604281e-06, 6.923352e-06,
  5.8894e-05, 8.428919e-05, 3.886843e-05, 6.508236e-06, 5.464039e-06, 
    1.750889e-05, 3.707907e-05, 4.151912e-05, 2.667643e-05, 2.899566e-05, 
    2.676429e-05, 1.944097e-05, 1.503444e-05, 6.978234e-06, 5.416015e-06,
  5.018827e-05, 0.0001074257, 0.0001152739, 3.144493e-05, 5.864809e-06, 
    1.449145e-05, 3.348388e-05, 4.794537e-05, 4.61827e-05, 2.944249e-05, 
    1.970113e-05, 2.409576e-05, 1.31104e-05, 5.496442e-06, 4.131961e-06,
  3.180089e-05, 4.219842e-05, 0.0001150699, 0.0001214171, 3.235245e-05, 
    1.509156e-05, 3.148358e-05, 6.141829e-05, 5.810654e-05, 2.968817e-05, 
    2.296253e-05, 2.664551e-05, 1.868577e-05, 1.623872e-05, 7.784002e-06,
  2.055163e-05, 4.290462e-05, 0.0001406131, 0.0002175397, 0.0001263932, 
    3.249512e-05, 3.083271e-05, 4.914376e-05, 4.624264e-05, 3.384396e-05, 
    2.515063e-05, 4.79651e-05, 3.817416e-05, 2.175226e-05, 1.958214e-05,
  1.330092e-05, 2.553653e-05, 8.972572e-05, 0.0001624064, 0.0002311298, 
    0.0001081175, 3.043146e-05, 3.473297e-05, 4.958287e-05, 4.716337e-05, 
    4.931984e-05, 4.607588e-05, 3.728793e-05, 3.821562e-05, 2.842106e-05,
  7.403976e-09, 2.082123e-07, 1.43126e-06, 2.350068e-06, 3.05703e-06, 
    5.836628e-06, 7.463695e-06, 7.715538e-06, 4.176077e-06, 3.392691e-06, 
    4.171016e-06, 5.316379e-06, 6.288578e-06, 9.54826e-06, 1.504317e-05,
  4.093139e-12, 1.195267e-07, 2.794382e-07, 1.447274e-07, 6.115289e-07, 
    5.058749e-07, 6.190861e-07, 3.40298e-06, 3.672108e-06, 2.293224e-06, 
    4.722792e-06, 6.761109e-06, 8.304874e-06, 1.155365e-05, 1.533245e-05,
  2.791748e-11, 1.364611e-07, 2.832455e-07, 3.419351e-07, 1.935861e-07, 
    6.18931e-08, 7.56282e-08, 1.71557e-06, 2.00326e-06, 1.70006e-06, 
    3.062653e-06, 5.047884e-06, 7.37977e-06, 1.077367e-05, 9.991447e-06,
  2.292977e-12, 1.766114e-07, 3.587393e-07, 4.94705e-07, 3.183315e-07, 
    2.986338e-08, 5.017833e-08, 4.588935e-07, 2.724423e-06, 3.921388e-06, 
    2.492044e-06, 3.995363e-06, 6.332884e-06, 5.907428e-06, 2.342048e-06,
  3.63255e-09, 1.388563e-07, 3.768165e-07, 4.586261e-07, 4.352155e-07, 
    3.752662e-07, 3.719112e-07, 3.068358e-07, 8.402014e-07, 4.226998e-06, 
    1.692922e-06, 1.911459e-06, 3.828259e-06, 4.977738e-06, 2.763056e-06,
  2.13893e-08, 2.5073e-07, 6.653332e-07, 4.532154e-07, 4.506392e-07, 
    4.594996e-07, 1.091332e-06, 1.843812e-06, 3.340315e-06, 4.756907e-06, 
    7.949544e-06, 2.58362e-06, 2.601577e-06, 1.966544e-06, 2.789612e-06,
  1.522342e-07, 5.673995e-07, 1.076774e-06, 1.426814e-06, 7.740336e-07, 
    6.790698e-07, 7.787206e-07, 1.285132e-06, 2.687213e-06, 2.708534e-06, 
    3.253953e-06, 1.86992e-06, 2.734301e-06, 2.161138e-06, 4.123006e-06,
  4.777061e-07, 1.122725e-06, 1.884121e-06, 2.109857e-06, 8.33823e-07, 
    1.223291e-06, 1.088842e-06, 2.633438e-06, 4.777151e-06, 4.432225e-06, 
    3.954834e-06, 3.31539e-06, 3.748547e-06, 3.674056e-06, 5.232395e-06,
  2.479865e-06, 1.611612e-06, 2.557055e-06, 2.225375e-06, 1.999085e-06, 
    2.051571e-06, 2.580114e-06, 3.208804e-06, 5.569872e-06, 4.009772e-06, 
    4.29848e-06, 3.55518e-06, 3.590844e-06, 4.769089e-06, 6.338974e-06,
  9.073937e-06, 3.187464e-06, 3.231686e-06, 4.601535e-06, 4.10043e-06, 
    4.584248e-06, 4.644258e-06, 6.049684e-06, 9.334401e-06, 6.42951e-06, 
    6.342711e-06, 4.939399e-06, 4.626696e-06, 6.691406e-06, 9.623518e-06,
  1.035704e-06, 2.607185e-07, 9.568687e-09, 2.675139e-08, 2.223541e-07, 
    3.442843e-06, 4.419884e-06, 6.001966e-06, 1.591495e-05, 5.097065e-05, 
    9.223197e-05, 0.0001103005, 0.0001642714, 0.000220765, 0.000290463,
  4.643737e-07, 1.721389e-07, 2.176661e-07, 8.133288e-09, 1.76825e-06, 
    1.18536e-06, 5.229687e-06, 5.54468e-06, 2.218202e-05, 7.402566e-05, 
    0.0001287556, 0.0001601248, 0.0002196795, 0.0003098952, 0.0003244037,
  5.007956e-08, 4.146565e-08, 2.165058e-07, 1.000775e-07, 5.844702e-07, 
    2.837133e-06, 5.140987e-06, 6.654189e-06, 2.494696e-05, 8.932983e-05, 
    0.0001572319, 0.0002028147, 0.0002768883, 0.0003323062, 0.0002738139,
  1.262722e-07, 7.186461e-09, 8.740047e-08, 2.14486e-07, 6.695143e-07, 
    1.277442e-06, 6.154905e-06, 6.40302e-06, 2.076076e-05, 8.64777e-05, 
    0.0001688654, 0.0002268386, 0.0002833764, 0.0002745996, 0.0001981969,
  2.443722e-07, 2.41849e-07, 6.082082e-08, 3.147913e-07, 1.13448e-06, 
    2.248996e-06, 4.39212e-06, 4.718231e-06, 7.939634e-06, 9.087526e-05, 
    0.0001917298, 0.0002440994, 0.0002592728, 0.000212352, 0.0001430867,
  3.11545e-07, 6.515364e-07, 3.61529e-07, 3.088387e-07, 8.031839e-07, 
    3.620386e-06, 6.194852e-06, 5.454805e-06, 3.585185e-06, 6.239025e-05, 
    0.0002041123, 0.0002484501, 0.0002307774, 0.0001711141, 0.0001110335,
  4.098699e-07, 7.311941e-07, 1.143078e-06, 1.049301e-06, 1.367015e-06, 
    4.620778e-06, 8.584324e-06, 5.43347e-06, 3.12594e-06, 4.474103e-05, 
    0.0001916005, 0.0002312575, 0.0001802762, 0.0001313553, 9.261496e-05,
  9.158788e-07, 2.032566e-06, 1.585188e-06, 1.744607e-06, 2.030259e-06, 
    3.554641e-06, 5.085617e-06, 3.921915e-06, 6.482439e-06, 3.55133e-05, 
    0.0001727404, 0.0001949659, 0.0001489706, 0.0001023094, 7.388826e-05,
  1.74157e-06, 2.895165e-06, 4.246826e-06, 3.513485e-06, 3.963619e-06, 
    3.995011e-06, 5.381061e-06, 4.38217e-06, 4.653565e-06, 3.71727e-05, 
    0.0001462759, 0.0001617093, 0.0001301677, 8.70518e-05, 6.635884e-05,
  3.066138e-06, 3.823597e-06, 4.416343e-06, 4.577166e-06, 4.357787e-06, 
    4.38257e-06, 3.418515e-06, 3.547145e-06, 2.608687e-06, 3.333556e-05, 
    0.0001189067, 0.0001359428, 0.000112562, 8.292154e-05, 6.465852e-05,
  4.642339e-06, 5.537298e-06, 1.181464e-05, 2.496159e-05, 2.132902e-05, 
    1.38311e-05, 1.226639e-05, 1.989487e-05, 2.147683e-05, 7.067729e-06, 
    1.957787e-08, 1.67459e-08, 1.220221e-07, 2.48931e-07, 4.084329e-07,
  5.321581e-06, 4.692834e-06, 9.114428e-06, 2.173958e-05, 2.39243e-05, 
    1.898481e-05, 1.661727e-05, 2.976437e-05, 3.43573e-05, 9.836911e-06, 
    4.237658e-07, 6.876144e-08, 6.858619e-08, 2.210529e-07, 1.439738e-06,
  8.423863e-06, 5.942307e-06, 7.454773e-06, 2.19735e-05, 3.108713e-05, 
    2.4627e-05, 2.709854e-05, 4.090749e-05, 4.951549e-05, 1.758752e-05, 
    1.057248e-06, 2.719303e-07, 2.812901e-07, 3.605009e-07, 1.742871e-06,
  1.2904e-05, 7.569244e-06, 5.024724e-06, 2.086278e-05, 3.428263e-05, 
    3.178215e-05, 3.434921e-05, 5.591494e-05, 6.793814e-05, 3.413303e-05, 
    3.158765e-06, 3.386781e-07, 4.51143e-07, 9.438265e-07, 7.426684e-07,
  1.113422e-05, 1.126303e-05, 1.046917e-05, 2.726698e-05, 4.531537e-05, 
    5.310855e-05, 5.573005e-05, 7.244027e-05, 9.60821e-05, 5.823186e-05, 
    9.343205e-06, 5.024959e-07, 9.780883e-07, 1.365702e-06, 1.181414e-06,
  1.156147e-05, 1.49418e-05, 1.608573e-05, 1.776131e-05, 4.698827e-05, 
    6.918092e-05, 6.966489e-05, 9.121582e-05, 0.0001173575, 9.030577e-05, 
    2.867019e-05, 2.137599e-06, 1.283093e-06, 1.501704e-06, 1.966585e-06,
  8.841474e-06, 1.139612e-05, 1.997767e-05, 2.414934e-05, 4.584874e-05, 
    7.169862e-05, 9.013853e-05, 0.0001122244, 0.0001208165, 0.0001257351, 
    5.147918e-05, 4.349568e-06, 1.48836e-06, 1.538396e-06, 1.281967e-06,
  7.344215e-06, 9.79653e-06, 1.521978e-05, 3.980624e-05, 3.751971e-05, 
    7.32687e-05, 9.786055e-05, 0.0001164815, 0.0001389161, 0.0001400932, 
    6.526184e-05, 9.149244e-06, 2.276862e-06, 2.341307e-06, 1.904789e-06,
  8.428492e-06, 8.777416e-06, 9.805967e-06, 1.825084e-05, 3.037944e-05, 
    7.544634e-05, 0.0001112784, 0.0001302703, 0.0001260871, 0.0001363749, 
    7.129752e-05, 1.470582e-05, 3.276335e-06, 3.767914e-06, 2.258665e-06,
  7.377389e-06, 8.70999e-06, 8.102873e-06, 1.399302e-05, 2.497481e-05, 
    7.07656e-05, 0.0001187912, 0.0001333177, 0.0001183238, 0.0001199828, 
    6.227969e-05, 1.299066e-05, 4.478358e-06, 3.571863e-06, 2.991335e-06,
  3.671053e-06, 1.459041e-06, 6.762655e-08, 1.089897e-07, 3.18553e-07, 
    6.132572e-07, 1.497616e-06, 2.640332e-06, 4.699362e-06, 5.21288e-06, 
    3.997276e-06, 4.552539e-06, 2.739225e-06, 9.079671e-06, 4.080737e-05,
  2.45992e-06, 4.048707e-07, 6.303075e-09, 2.593121e-09, 4.586341e-08, 
    3.796262e-07, 7.234762e-07, 1.851895e-06, 3.209114e-06, 5.385542e-06, 
    2.201202e-06, 4.437188e-06, 7.464671e-06, 1.310369e-05, 4.883358e-05,
  3.232875e-06, 3.113819e-07, 2.691222e-08, 6.09779e-09, 2.480839e-09, 
    5.556043e-08, 3.167524e-07, 6.04775e-07, 2.17192e-06, 5.518508e-06, 
    2.761948e-06, 2.952196e-06, 5.752764e-06, 9.365088e-06, 4.213918e-05,
  5.409524e-06, 1.782489e-06, 4.846242e-08, 4.71209e-08, 1.721217e-08, 
    1.70263e-08, 1.789477e-07, 5.621104e-07, 1.272305e-06, 4.933242e-06, 
    2.907303e-06, 4.475811e-06, 5.875232e-06, 7.792339e-06, 3.537354e-05,
  6.381978e-06, 3.616318e-06, 2.421997e-07, 1.841645e-08, 7.556261e-09, 
    1.12122e-07, 2.03469e-07, 7.940947e-07, 9.17574e-07, 3.993915e-06, 
    3.950089e-06, 5.332233e-06, 6.397794e-06, 8.06708e-06, 3.954687e-05,
  7.953189e-06, 4.260115e-06, 9.291041e-07, 1.566529e-08, 2.276681e-08, 
    7.909566e-08, 6.211088e-08, 3.703648e-07, 9.132402e-07, 2.781e-06, 
    5.603951e-06, 5.968918e-06, 7.478954e-06, 1.094766e-05, 3.744041e-05,
  6.571017e-06, 5.497632e-06, 2.386572e-06, 2.043166e-07, 2.969931e-07, 
    2.977696e-07, 2.546677e-07, 9.709354e-07, 1.361414e-06, 2.427979e-06, 
    2.328456e-06, 3.944624e-06, 9.234695e-06, 1.085925e-05, 3.271818e-05,
  8.568008e-06, 6.349567e-06, 4.604962e-06, 7.165838e-07, 3.363738e-07, 
    3.371281e-07, 1.03276e-06, 3.265227e-06, 1.601342e-06, 2.852237e-06, 
    2.94425e-06, 3.060662e-06, 1.003002e-05, 1.486691e-05, 2.645278e-05,
  8.415394e-06, 6.161567e-06, 4.691415e-06, 1.938709e-06, 2.221974e-07, 
    3.29758e-07, 9.509637e-07, 2.04004e-06, 4.37021e-06, 5.687243e-06, 
    5.669776e-06, 5.659419e-06, 9.208427e-06, 1.416731e-05, 2.490806e-05,
  7.061879e-06, 9.410363e-06, 6.448955e-06, 1.597772e-06, 1.132043e-07, 
    1.355622e-07, 5.186843e-07, 2.807157e-06, 4.231415e-06, 6.763739e-06, 
    6.731174e-06, 6.987561e-06, 7.077459e-06, 1.205528e-05, 2.324228e-05,
  9.37926e-06, 1.231521e-05, 1.60308e-05, 1.4408e-05, 1.570554e-05, 
    1.11087e-05, 3.52871e-06, 3.743178e-06, 8.452276e-05, 0.0001398252, 
    0.0001401137, 8.674037e-05, 9.368065e-05, 8.247922e-05, 5.594359e-05,
  9.275616e-06, 7.418624e-06, 1.292711e-05, 1.100317e-05, 1.301036e-05, 
    1.214574e-05, 4.981273e-06, 1.788055e-06, 6.002261e-05, 0.0001375674, 
    0.0001613267, 0.0001095542, 0.0001144912, 9.65301e-05, 8.178211e-05,
  1.236125e-05, 1.197744e-05, 1.242732e-05, 1.021816e-05, 1.077072e-05, 
    7.010879e-06, 5.505316e-06, 3.446761e-06, 2.33052e-05, 0.0001185392, 
    0.0001376894, 0.0001201783, 0.0001164014, 0.0001107077, 9.818255e-05,
  1.060119e-05, 1.224107e-05, 1.871866e-05, 9.806876e-06, 8.026835e-06, 
    4.104143e-06, 3.416386e-06, 2.936029e-06, 9.95341e-06, 9.492863e-05, 
    9.547373e-05, 0.0001180455, 0.0001193436, 0.0001200116, 9.791167e-05,
  8.266823e-06, 1.043297e-05, 1.425781e-05, 1.474021e-05, 7.467222e-06, 
    4.690788e-06, 2.352094e-06, 3.268776e-06, 1.057485e-05, 6.379925e-05, 
    7.267938e-05, 0.000125319, 0.0001344834, 0.0001375477, 0.0001075301,
  7.244798e-06, 1.17516e-05, 9.435672e-06, 1.271087e-05, 8.745635e-06, 
    3.671362e-06, 1.579341e-06, 2.620061e-06, 1.542846e-05, 4.287011e-05, 
    7.12093e-05, 0.0001498928, 0.000152622, 0.0001518589, 0.0001208963,
  8.383801e-06, 9.623376e-06, 9.147942e-06, 1.004176e-05, 6.477534e-06, 
    3.316286e-06, 9.889751e-07, 1.755555e-06, 2.558912e-05, 2.522287e-05, 
    7.30248e-05, 0.0001701157, 0.0001631046, 0.0001543007, 0.0001369849,
  6.249974e-06, 8.914267e-06, 1.022334e-05, 1.00267e-05, 3.933731e-06, 
    2.417853e-06, 1.244106e-06, 1.760367e-06, 2.937521e-05, 1.449949e-05, 
    7.028751e-05, 0.0001823006, 0.0001648256, 0.0001588975, 0.0001448498,
  5.048325e-06, 1.03166e-05, 9.425848e-06, 6.164783e-06, 5.935148e-06, 
    2.703954e-06, 9.744552e-07, 2.034422e-06, 2.708141e-05, 1.374816e-05, 
    7.776756e-05, 0.000184325, 0.0001587126, 0.0001624869, 0.000136358,
  5.418127e-06, 7.914762e-06, 6.111945e-06, 5.853678e-06, 3.106831e-06, 
    1.733776e-06, 1.445145e-06, 2.164297e-06, 2.03524e-05, 1.642908e-05, 
    8.479192e-05, 0.0001790334, 0.0001482391, 0.0001630291, 0.0001138949,
  2.165175e-05, 3.073052e-05, 4.79664e-05, 4.689578e-05, 4.473272e-05, 
    6.040691e-05, 9.153794e-05, 0.0001250783, 0.0001268247, 8.539426e-05, 
    2.335605e-05, 1.261496e-05, 1.493811e-05, 1.187479e-05, 1.093406e-05,
  1.723375e-05, 4.820915e-05, 8.257201e-05, 7.771021e-05, 7.034821e-05, 
    9.037514e-05, 0.0001473432, 0.0002107247, 0.0002065972, 0.0001229138, 
    2.897787e-05, 2.030311e-05, 2.237458e-05, 1.658333e-05, 1.84915e-05,
  1.005876e-05, 4.259733e-05, 9.373188e-05, 8.87748e-05, 7.474793e-05, 
    9.773811e-05, 0.0001683344, 0.0002548777, 0.0002564693, 0.0001792898, 
    4.403768e-05, 2.161048e-05, 1.959061e-05, 1.641716e-05, 1.711111e-05,
  8.457956e-06, 2.531564e-05, 8.293055e-05, 8.647321e-05, 6.542095e-05, 
    9.133498e-05, 0.0001628652, 0.0002588205, 0.0002423323, 0.0001862367, 
    5.287684e-05, 1.50769e-05, 1.591356e-05, 1.645555e-05, 1.471024e-05,
  7.924158e-06, 1.266741e-05, 6.581019e-05, 8.845093e-05, 6.736413e-05, 
    9.426006e-05, 0.0001771975, 0.0002673044, 0.0002307158, 0.0001935703, 
    6.116621e-05, 1.427884e-05, 1.659538e-05, 1.689846e-05, 1.313111e-05,
  7.525301e-06, 6.975115e-06, 4.169735e-05, 8.982593e-05, 7.837301e-05, 
    9.950018e-05, 0.0001757131, 0.0002672973, 0.0002347338, 0.0001711721, 
    6.3871e-05, 1.666357e-05, 1.61572e-05, 1.695402e-05, 1.563369e-05,
  7.938401e-06, 3.362997e-06, 1.957063e-05, 7.789724e-05, 8.391707e-05, 
    0.0001039085, 0.0001755493, 0.0002637016, 0.000237652, 0.0001787524, 
    6.760917e-05, 2.023166e-05, 1.554547e-05, 1.861976e-05, 1.731144e-05,
  5.411043e-06, 3.261313e-06, 5.588323e-06, 5.477228e-05, 8.094685e-05, 
    0.0001064627, 0.0001698604, 0.0002596779, 0.0002338021, 0.0001786856, 
    8.865796e-05, 2.486481e-05, 1.802125e-05, 1.978642e-05, 1.769879e-05,
  6.026616e-06, 4.686427e-06, 1.557299e-06, 3.370736e-05, 7.513316e-05, 
    0.0001012528, 0.0001656417, 0.0002487015, 0.0002250133, 0.0001741614, 
    0.0001063594, 3.672498e-05, 1.481283e-05, 1.717717e-05, 1.901234e-05,
  6.041838e-06, 4.66875e-06, 1.263477e-06, 1.028872e-05, 5.855596e-05, 
    0.0001006184, 0.0001576444, 0.0002502695, 0.0002310688, 0.0001766179, 
    0.0001505083, 5.168692e-05, 1.717376e-05, 1.861433e-05, 2.372307e-05,
  4.150071e-05, 1.518593e-05, 4.394974e-06, 2.75754e-06, 3.528967e-06, 
    5.60752e-06, 8.683921e-06, 1.270974e-05, 1.679829e-05, 1.626989e-05, 
    1.745789e-05, 1.670096e-05, 1.842483e-05, 1.78499e-05, 1.945726e-05,
  5.832634e-05, 3.130375e-05, 7.109292e-06, 3.471101e-06, 3.943596e-06, 
    8.10349e-06, 1.220086e-05, 1.754007e-05, 1.863087e-05, 1.872543e-05, 
    1.790351e-05, 1.853753e-05, 2.314792e-05, 1.889618e-05, 1.979537e-05,
  5.824455e-05, 3.724615e-05, 1.044142e-05, 3.668898e-06, 4.444109e-06, 
    1.017699e-05, 1.82964e-05, 2.093876e-05, 2.215387e-05, 2.031384e-05, 
    1.98735e-05, 2.458578e-05, 2.511845e-05, 2.519283e-05, 2.240298e-05,
  5.818822e-05, 4.826915e-05, 1.898884e-05, 4.27058e-06, 6.762914e-06, 
    1.478622e-05, 2.230744e-05, 2.307693e-05, 2.450125e-05, 2.525561e-05, 
    2.713667e-05, 2.875658e-05, 2.950411e-05, 3.209138e-05, 3.017202e-05,
  5.884085e-05, 6.256602e-05, 3.465161e-05, 6.533528e-06, 9.473404e-06, 
    2.11781e-05, 2.693954e-05, 2.925747e-05, 3.03104e-05, 3.193074e-05, 
    3.270413e-05, 3.368759e-05, 3.502635e-05, 3.34123e-05, 2.693261e-05,
  5.903442e-05, 6.639049e-05, 5.431185e-05, 1.454847e-05, 1.071215e-05, 
    2.354552e-05, 3.082966e-05, 3.433712e-05, 4.125205e-05, 4.118799e-05, 
    3.585281e-05, 3.576938e-05, 3.788024e-05, 3.490409e-05, 2.997451e-05,
  6.51264e-05, 6.771107e-05, 7.332253e-05, 2.893458e-05, 1.861911e-05, 
    4.075255e-05, 4.948298e-05, 4.076622e-05, 4.709178e-05, 5.33423e-05, 
    4.105394e-05, 4.120554e-05, 3.819175e-05, 3.405483e-05, 3.881241e-05,
  6.57664e-05, 6.531797e-05, 8.26892e-05, 4.926527e-05, 4.349135e-05, 
    6.309985e-05, 5.339634e-05, 4.690448e-05, 6.585438e-05, 4.456264e-05, 
    4.140957e-05, 3.765662e-05, 4.175207e-05, 4.763143e-05, 6.117109e-05,
  7.213819e-05, 6.396595e-05, 8.237264e-05, 6.928143e-05, 5.187114e-05, 
    5.422794e-05, 5.71059e-05, 4.204802e-05, 3.878362e-05, 3.999026e-05, 
    3.562577e-05, 4.087469e-05, 4.950841e-05, 5.420383e-05, 7.594099e-05,
  8.096298e-05, 6.847823e-05, 8.252605e-05, 8.494951e-05, 5.11516e-05, 
    5.227994e-05, 3.457134e-05, 4.522129e-05, 3.591794e-05, 4.245909e-05, 
    4.535604e-05, 4.93792e-05, 8.136567e-05, 7.941315e-05, 7.678394e-05,
  3.178748e-05, 2.93202e-05, 2.349694e-05, 2.168569e-05, 2.530281e-05, 
    2.510854e-05, 2.212552e-05, 2.087019e-05, 2.449361e-05, 2.045373e-05, 
    2.074549e-05, 1.913291e-05, 1.989387e-05, 1.811722e-05, 1.574143e-05,
  3.126207e-05, 2.699696e-05, 2.398144e-05, 2.483266e-05, 2.563526e-05, 
    2.312527e-05, 1.717336e-05, 1.797017e-05, 1.875581e-05, 1.817808e-05, 
    2.164316e-05, 2.328776e-05, 2.176795e-05, 1.957692e-05, 1.933232e-05,
  3.005601e-05, 2.683289e-05, 2.568656e-05, 2.555653e-05, 2.700466e-05, 
    2.324001e-05, 1.434273e-05, 1.251444e-05, 1.497755e-05, 1.693946e-05, 
    1.7683e-05, 1.869754e-05, 1.992197e-05, 1.984899e-05, 1.925402e-05,
  2.770943e-05, 2.906471e-05, 2.894257e-05, 2.794886e-05, 2.77046e-05, 
    2.09478e-05, 1.346309e-05, 1.21552e-05, 1.505253e-05, 1.693564e-05, 
    1.435343e-05, 1.514784e-05, 1.72801e-05, 1.746073e-05, 1.788562e-05,
  3.137668e-05, 3.185778e-05, 2.907124e-05, 3.32526e-05, 2.980849e-05, 
    2.146741e-05, 1.325273e-05, 1.299408e-05, 1.75934e-05, 1.838507e-05, 
    1.692225e-05, 1.532785e-05, 1.535898e-05, 1.630785e-05, 1.59386e-05,
  3.109469e-05, 2.982406e-05, 3.734684e-05, 4.368227e-05, 4.340364e-05, 
    2.492355e-05, 1.398876e-05, 1.874402e-05, 2.738631e-05, 2.646835e-05, 
    2.533581e-05, 2.358951e-05, 1.856676e-05, 1.491686e-05, 1.468667e-05,
  3.451339e-05, 3.579089e-05, 4.504024e-05, 5.379833e-05, 4.71627e-05, 
    2.969482e-05, 2.316114e-05, 2.991381e-05, 4.648188e-05, 4.629966e-05, 
    3.924095e-05, 2.976796e-05, 2.460667e-05, 2.120635e-05, 1.928031e-05,
  6.182721e-05, 6.483769e-05, 7.03043e-05, 8.464542e-05, 4.997352e-05, 
    3.808876e-05, 3.610825e-05, 4.598415e-05, 5.479365e-05, 8.067032e-05, 
    7.124546e-05, 5.684948e-05, 4.324583e-05, 3.547634e-05, 2.730138e-05,
  7.160185e-05, 6.610175e-05, 6.682678e-05, 8.484171e-05, 5.961327e-05, 
    5.118045e-05, 4.983908e-05, 5.966904e-05, 7.124902e-05, 9.893807e-05, 
    8.412622e-05, 0.0001003276, 7.756746e-05, 5.905776e-05, 4.298422e-05,
  6.490637e-05, 5.35476e-05, 8.225915e-05, 6.872472e-05, 6.25506e-05, 
    5.533345e-05, 5.701701e-05, 6.558203e-05, 7.478796e-05, 8.806957e-05, 
    0.0001076322, 9.747846e-05, 9.535206e-05, 8.612004e-05, 7.018731e-05,
  2.181952e-05, 2.137341e-05, 2.052469e-05, 1.80361e-05, 2.080871e-05, 
    1.895621e-05, 1.260656e-05, 1.000152e-05, 8.376944e-06, 6.748379e-06, 
    5.457724e-06, 6.531447e-06, 5.191498e-06, 5.603012e-06, 5.296889e-06,
  2.414776e-05, 2.534042e-05, 2.314001e-05, 2.426298e-05, 2.545541e-05, 
    2.321272e-05, 1.633625e-05, 1.624662e-05, 1.478138e-05, 1.180439e-05, 
    9.005859e-06, 6.428875e-06, 4.607527e-06, 4.887176e-06, 6.028824e-06,
  2.923189e-05, 3.057469e-05, 3.138e-05, 2.527604e-05, 2.464061e-05, 
    2.638663e-05, 2.464793e-05, 2.195843e-05, 2.002031e-05, 1.794183e-05, 
    1.366644e-05, 7.478703e-06, 5.275951e-06, 5.074221e-06, 3.321393e-06,
  4.817204e-05, 3.524071e-05, 3.898088e-05, 3.369122e-05, 3.280755e-05, 
    3.323792e-05, 2.904275e-05, 2.439259e-05, 2.723389e-05, 2.307023e-05, 
    1.927841e-05, 1.433319e-05, 8.385056e-06, 6.390541e-06, 3.810229e-06,
  7.074977e-05, 6.393301e-05, 4.557384e-05, 4.297236e-05, 5.144705e-05, 
    3.784195e-05, 3.604491e-05, 3.647788e-05, 3.364061e-05, 2.801057e-05, 
    2.67772e-05, 2.308953e-05, 1.552981e-05, 1.009719e-05, 5.180158e-06,
  7.674879e-05, 5.49073e-05, 8.355058e-05, 6.833947e-05, 5.318504e-05, 
    7.149364e-05, 5.290228e-05, 4.478228e-05, 3.591998e-05, 2.384433e-05, 
    3.541241e-05, 3.071676e-05, 3.010809e-05, 1.783383e-05, 1.174052e-05,
  9.722784e-05, 6.630766e-05, 8.866756e-05, 0.0001081717, 0.0001037768, 
    6.219301e-05, 5.550894e-05, 4.898082e-05, 4.228992e-05, 3.048144e-05, 
    3.300067e-05, 3.725146e-05, 2.803739e-05, 2.092051e-05, 2.161883e-05,
  0.0001311091, 0.0001092743, 9.225307e-05, 9.999495e-05, 8.522861e-05, 
    7.944406e-05, 8.403589e-05, 7.891243e-05, 4.851982e-05, 3.560756e-05, 
    3.019728e-05, 2.919824e-05, 3.148345e-05, 3.273034e-05, 2.165155e-05,
  0.0001056043, 9.500547e-05, 0.0001144716, 0.0001085354, 0.0001028553, 
    9.754035e-05, 0.0001034701, 7.937771e-05, 6.196766e-05, 4.185181e-05, 
    3.363165e-05, 3.106082e-05, 2.899627e-05, 2.817982e-05, 2.723818e-05,
  0.0001208632, 0.0001481671, 0.0001330863, 0.0001289692, 0.0001324003, 
    9.025668e-05, 0.0001066897, 7.870339e-05, 8.857693e-05, 4.290036e-05, 
    3.732552e-05, 3.123479e-05, 2.850038e-05, 2.621235e-05, 1.953703e-05,
  2.512224e-05, 2.674962e-05, 2.417747e-05, 1.987222e-05, 1.929117e-05, 
    1.982619e-05, 1.716458e-05, 1.680194e-05, 1.983235e-05, 1.791406e-05, 
    1.558071e-05, 1.677205e-05, 1.578515e-05, 1.313174e-05, 1.166133e-05,
  1.960754e-05, 2.540655e-05, 2.253186e-05, 2.557334e-05, 2.676677e-05, 
    2.850684e-05, 2.32154e-05, 2.076291e-05, 2.244477e-05, 2.309711e-05, 
    2.013758e-05, 1.682742e-05, 1.266306e-05, 1.25619e-05, 1.049364e-05,
  1.292971e-05, 1.651077e-05, 1.849729e-05, 1.935075e-05, 2.366855e-05, 
    3.013645e-05, 2.970698e-05, 2.896518e-05, 3.180647e-05, 2.966302e-05, 
    2.616168e-05, 2.227556e-05, 1.895613e-05, 1.764848e-05, 1.126919e-05,
  1.007033e-05, 1.219319e-05, 1.201974e-05, 1.01255e-05, 1.292477e-05, 
    1.867839e-05, 2.00032e-05, 2.497797e-05, 3.277495e-05, 3.744534e-05, 
    3.237195e-05, 3.469063e-05, 2.808762e-05, 2.760005e-05, 1.453748e-05,
  8.731286e-06, 9.930488e-06, 9.678475e-06, 9.32129e-06, 8.346677e-06, 
    8.943969e-06, 1.260704e-05, 1.212314e-05, 1.725327e-05, 2.24344e-05, 
    3.038095e-05, 3.808186e-05, 4.458868e-05, 2.615203e-05, 2.752723e-05,
  7.15377e-06, 8.242495e-06, 8.059246e-06, 8.279801e-06, 7.842026e-06, 
    6.572172e-06, 7.46901e-06, 7.652901e-06, 1.083632e-05, 1.220688e-05, 
    1.357216e-05, 1.262918e-05, 1.978646e-05, 2.602062e-05, 3.806741e-05,
  6.075894e-06, 8.460261e-06, 9.339315e-06, 6.77818e-06, 8.297022e-06, 
    6.960638e-06, 5.90775e-06, 7.363439e-06, 7.517428e-06, 9.023511e-06, 
    5.941415e-06, 1.015966e-05, 8.040135e-06, 1.930754e-05, 1.984316e-05,
  8.969624e-06, 9.51063e-06, 1.080571e-05, 7.936331e-06, 9.559699e-06, 
    9.125454e-06, 5.200615e-06, 5.754582e-06, 7.04895e-06, 8.098429e-06, 
    6.438964e-06, 9.347167e-06, 8.270048e-06, 9.182957e-06, 1.054122e-05,
  1.216057e-05, 1.114218e-05, 1.159425e-05, 1.230625e-05, 1.221036e-05, 
    1.25745e-05, 6.936203e-06, 6.725392e-06, 6.904619e-06, 7.867277e-06, 
    6.642013e-06, 6.922265e-06, 1.091917e-05, 1.145728e-05, 1.005526e-05,
  1.662587e-05, 1.56386e-05, 1.566268e-05, 1.442264e-05, 1.382701e-05, 
    1.481351e-05, 1.11708e-05, 9.811151e-06, 1.006437e-05, 8.542709e-06, 
    6.118618e-06, 6.927494e-06, 3.816808e-06, 5.167345e-06, 5.113699e-06,
  1.838634e-05, 1.655042e-05, 1.637367e-05, 1.625984e-05, 1.622242e-05, 
    1.813726e-05, 1.130642e-05, 8.767583e-06, 1.05502e-05, 1.205532e-05, 
    1.132297e-05, 1.03851e-05, 7.575711e-06, 6.383889e-06, 4.419725e-06,
  2.003543e-05, 1.663602e-05, 1.632179e-05, 1.385596e-05, 1.692802e-05, 
    1.743539e-05, 1.125014e-05, 1.081238e-05, 1.239819e-05, 1.327895e-05, 
    1.265505e-05, 1.101241e-05, 9.250498e-06, 6.115737e-06, 5.463042e-06,
  1.487028e-05, 1.861673e-05, 1.704893e-05, 1.721549e-05, 1.771873e-05, 
    1.540049e-05, 1.22249e-05, 1.211045e-05, 1.163568e-05, 1.332859e-05, 
    1.088988e-05, 8.902789e-06, 7.229715e-06, 8.698971e-06, 8.408096e-06,
  1.434859e-05, 1.59867e-05, 1.940743e-05, 1.841193e-05, 1.783897e-05, 
    1.495342e-05, 1.303353e-05, 1.050011e-05, 1.138024e-05, 1.352869e-05, 
    1.13404e-05, 9.133794e-06, 9.076086e-06, 1.059707e-05, 8.990377e-06,
  1.472802e-05, 1.860803e-05, 1.901001e-05, 1.955074e-05, 1.572598e-05, 
    1.529923e-05, 1.377293e-05, 1.074495e-05, 1.285582e-05, 1.36898e-05, 
    1.024878e-05, 8.709994e-06, 1.036937e-05, 7.554011e-06, 7.317253e-06,
  1.747772e-05, 2.24707e-05, 2.055486e-05, 1.914684e-05, 1.887353e-05, 
    1.869567e-05, 1.391345e-05, 1.268293e-05, 1.35213e-05, 1.325031e-05, 
    1.169306e-05, 6.270567e-06, 7.160952e-06, 4.467674e-06, 8.142993e-06,
  2.013957e-05, 2.145142e-05, 2.358443e-05, 2.477553e-05, 2.422986e-05, 
    1.706538e-05, 1.609077e-05, 1.560072e-05, 1.423662e-05, 1.109871e-05, 
    7.055981e-06, 7.950278e-06, 7.433542e-06, 7.058491e-06, 6.175955e-06,
  2.176645e-05, 2.290091e-05, 2.180475e-05, 2.129678e-05, 2.748574e-05, 
    2.622792e-05, 2.322772e-05, 2.273903e-05, 2.061153e-05, 1.577591e-05, 
    1.079106e-05, 8.683195e-06, 8.750316e-06, 5.823202e-06, 5.75063e-06,
  2.940429e-05, 2.27742e-05, 2.134855e-05, 2.252742e-05, 2.45932e-05, 
    2.271989e-05, 1.955373e-05, 2.309297e-05, 2.85046e-05, 2.895726e-05, 
    2.08451e-05, 1.702086e-05, 1.007406e-05, 8.314651e-06, 6.298061e-06,
  3.074503e-05, 3.063252e-05, 2.771003e-05, 2.365059e-05, 2.505533e-05, 
    2.644416e-05, 2.046252e-05, 1.768896e-05, 2.267162e-05, 2.536227e-05, 
    3.10444e-05, 2.657855e-05, 2.003687e-05, 1.845143e-05, 1.060949e-05,
  6.848734e-06, 5.0569e-06, 5.352788e-06, 5.708363e-06, 6.32928e-06, 
    5.728826e-06, 4.96246e-06, 5.818033e-06, 7.701471e-06, 7.82286e-06, 
    2.974131e-06, 2.848181e-06, 6.461781e-06, 1.073897e-05, 8.274288e-06,
  9.156002e-06, 7.216384e-06, 7.28069e-06, 6.573754e-06, 7.107879e-06, 
    9.239133e-06, 7.538963e-06, 6.789049e-06, 8.089008e-06, 8.211989e-06, 
    4.886056e-06, 1.947615e-06, 4.774386e-06, 7.642003e-06, 1.016512e-05,
  1.152294e-05, 9.79252e-06, 9.453518e-06, 8.11159e-06, 1.052774e-05, 
    1.341638e-05, 1.099877e-05, 8.965941e-06, 8.341399e-06, 8.109392e-06, 
    4.619891e-06, 2.498213e-06, 6.362852e-06, 7.972523e-06, 7.328898e-06,
  1.288978e-05, 1.065289e-05, 1.074881e-05, 9.798669e-06, 1.039475e-05, 
    1.142203e-05, 8.076158e-06, 8.137934e-06, 9.526265e-06, 8.573904e-06, 
    7.660732e-06, 2.696875e-06, 4.61604e-06, 7.143592e-06, 8.901783e-06,
  1.292488e-05, 1.271419e-05, 1.099277e-05, 8.368354e-06, 1.102619e-05, 
    7.658963e-06, 6.892281e-06, 7.137515e-06, 7.778483e-06, 9.780386e-06, 
    8.007492e-06, 2.854283e-06, 3.668319e-06, 6.624131e-06, 6.538516e-06,
  1.460226e-05, 1.201242e-05, 1.170129e-05, 1.11661e-05, 9.441119e-06, 
    8.276295e-06, 5.688639e-06, 7.535983e-06, 8.541077e-06, 6.209365e-06, 
    2.655184e-06, 2.862984e-06, 5.335999e-06, 8.689164e-06, 4.798041e-06,
  1.350894e-05, 1.116131e-05, 1.128474e-05, 1.084778e-05, 1.107362e-05, 
    9.424794e-06, 6.281247e-06, 7.931343e-06, 8.25098e-06, 7.069878e-06, 
    4.315717e-06, 3.154251e-06, 5.113959e-06, 8.939611e-06, 6.731219e-06,
  1.14664e-05, 9.616895e-06, 1.027363e-05, 1.113801e-05, 1.251344e-05, 
    9.431171e-06, 6.793364e-06, 6.929486e-06, 8.243022e-06, 7.27515e-06, 
    6.035018e-06, 4.549939e-06, 6.928119e-06, 6.903972e-06, 4.49968e-06,
  1.296246e-05, 1.000665e-05, 1.103537e-05, 1.156904e-05, 1.172048e-05, 
    1.177685e-05, 8.023344e-06, 6.186166e-06, 6.653949e-06, 7.514475e-06, 
    5.279948e-06, 4.625045e-06, 4.762748e-06, 5.676085e-06, 4.25101e-06,
  1.144571e-05, 1.249034e-05, 1.07722e-05, 1.07316e-05, 1.217345e-05, 
    1.169069e-05, 1.10108e-05, 7.208304e-06, 7.153726e-06, 7.203347e-06, 
    3.987121e-06, 4.383074e-06, 4.845351e-06, 4.776963e-06, 6.574155e-06,
  9.511091e-06, 8.345382e-06, 7.223845e-06, 8.792345e-06, 7.958261e-06, 
    6.242321e-06, 5.585569e-06, 4.140464e-06, 3.120851e-06, 1.289597e-05, 
    1.034118e-05, 9.500518e-06, 1.030401e-05, 9.765739e-06, 7.897953e-06,
  1.035192e-05, 9.246291e-06, 8.093877e-06, 8.528243e-06, 7.041473e-06, 
    5.877301e-06, 5.441621e-06, 7.410708e-06, 9.181305e-06, 1.170807e-05, 
    8.891828e-06, 7.595165e-06, 8.440737e-06, 1.037313e-05, 1.050366e-05,
  1.385303e-05, 1.282766e-05, 6.486869e-06, 7.436959e-06, 7.263625e-06, 
    8.138648e-06, 9.597828e-06, 9.915309e-06, 9.486524e-06, 8.742907e-06, 
    7.365074e-06, 7.784133e-06, 8.516475e-06, 1.099613e-05, 1.405651e-05,
  1.888592e-05, 1.035252e-05, 8.435543e-06, 6.929286e-06, 7.977636e-06, 
    7.827299e-06, 4.187324e-06, 6.16435e-06, 7.755926e-06, 5.050196e-06, 
    4.929124e-06, 6.917435e-06, 1.054088e-05, 8.57592e-06, 1.670831e-05,
  1.321242e-05, 9.900406e-06, 6.819592e-06, 6.692039e-06, 7.257383e-06, 
    6.167478e-06, 5.677225e-06, 7.147254e-06, 6.014574e-06, 4.483589e-06, 
    3.980866e-06, 6.560847e-06, 8.265642e-06, 1.121336e-05, 1.233118e-05,
  8.407848e-06, 5.805591e-06, 5.443915e-06, 8.236353e-06, 8.538663e-06, 
    7.281896e-06, 5.48658e-06, 6.113153e-06, 3.638744e-06, 3.063989e-06, 
    5.452676e-06, 6.837446e-06, 7.028666e-06, 9.140079e-06, 1.579245e-05,
  8.788712e-06, 4.045834e-06, 4.012195e-06, 8.808371e-06, 1.009869e-05, 
    6.209792e-06, 3.193278e-06, 4.586693e-06, 3.716912e-06, 3.663509e-06, 
    3.327148e-06, 5.210817e-06, 8.207006e-06, 9.416863e-06, 8.438014e-06,
  5.265742e-06, 5.200201e-06, 6.957611e-06, 8.660178e-06, 7.072527e-06, 
    5.915537e-06, 3.502545e-06, 4.259809e-06, 7.345754e-06, 5.329235e-06, 
    3.984959e-06, 5.831543e-06, 9.228515e-06, 1.003585e-05, 6.935755e-06,
  7.141559e-06, 7.054894e-06, 7.788749e-06, 9.677473e-06, 7.075937e-06, 
    5.609133e-06, 4.994624e-06, 5.880683e-06, 7.572007e-06, 4.177804e-06, 
    2.61206e-06, 3.523154e-06, 8.487775e-06, 8.894814e-06, 5.991156e-06,
  1.03893e-05, 6.39926e-06, 7.503613e-06, 7.685048e-06, 5.285243e-06, 
    5.228824e-06, 4.933363e-06, 7.832829e-06, 7.775108e-06, 6.532061e-06, 
    6.583569e-06, 3.97741e-06, 3.411756e-06, 4.765253e-06, 5.085276e-06,
  6.215293e-06, 7.407049e-06, 9.552692e-06, 1.014858e-05, 1.016865e-05, 
    1.044918e-05, 1.229359e-05, 1.593859e-05, 1.233832e-05, 1.208314e-05, 
    9.618179e-06, 8.31696e-06, 7.777655e-06, 7.424635e-06, 5.809414e-06,
  9.613002e-06, 1.038732e-05, 1.003144e-05, 1.035735e-05, 1.275947e-05, 
    1.312589e-05, 1.632613e-05, 1.493978e-05, 1.558221e-05, 1.828745e-05, 
    1.216886e-05, 1.132204e-05, 1.186747e-05, 1.205059e-05, 9.042812e-06,
  1.31297e-05, 1.2211e-05, 1.106038e-05, 1.364267e-05, 1.625006e-05, 
    1.46665e-05, 1.749973e-05, 1.853732e-05, 1.740932e-05, 1.740612e-05, 
    1.657772e-05, 1.224063e-05, 1.242817e-05, 1.404932e-05, 1.517149e-05,
  1.389224e-05, 1.162572e-05, 1.506973e-05, 1.705915e-05, 1.695982e-05, 
    1.396168e-05, 1.784085e-05, 1.834505e-05, 1.441583e-05, 1.696551e-05, 
    1.318843e-05, 9.441838e-06, 1.115455e-05, 1.267352e-05, 9.560204e-06,
  1.209819e-05, 1.422525e-05, 1.660542e-05, 1.641593e-05, 1.656836e-05, 
    1.591449e-05, 1.690926e-05, 1.80894e-05, 1.840829e-05, 1.207748e-05, 
    7.269574e-06, 8.624598e-06, 1.362909e-05, 7.56344e-06, 5.366247e-06,
  7.848793e-06, 1.600895e-05, 1.336834e-05, 1.341814e-05, 1.27945e-05, 
    1.342277e-05, 1.399445e-05, 1.411391e-05, 1.568468e-05, 1.145785e-05, 
    6.95079e-06, 1.355767e-05, 8.903048e-06, 6.162273e-06, 3.96114e-06,
  8.131854e-06, 1.153011e-05, 1.194703e-05, 1.022738e-05, 1.229046e-05, 
    1.172383e-05, 9.321771e-06, 1.303265e-05, 1.251947e-05, 1.132003e-05, 
    8.279851e-06, 7.999734e-06, 4.896936e-06, 3.763223e-06, 4.797808e-06,
  9.188447e-06, 1.105434e-05, 1.449468e-05, 1.158974e-05, 1.037114e-05, 
    1.223073e-05, 9.109872e-06, 1.051471e-05, 1.225697e-05, 1.272949e-05, 
    1.030351e-05, 1.136055e-05, 7.514785e-06, 8.358809e-06, 4.572324e-06,
  1.23372e-05, 1.33626e-05, 1.546748e-05, 1.315697e-05, 1.260223e-05, 
    1.303175e-05, 1.049849e-05, 1.239705e-05, 1.545576e-05, 1.404318e-05, 
    8.572873e-06, 9.693425e-06, 1.165201e-05, 1.366612e-05, 1.600858e-05,
  1.483547e-05, 1.716219e-05, 1.366371e-05, 1.089961e-05, 1.04695e-05, 
    9.397603e-06, 1.106117e-05, 1.316577e-05, 1.179574e-05, 9.537262e-06, 
    8.858739e-06, 8.876171e-06, 8.954355e-06, 1.137632e-05, 1.237245e-05,
  1.079944e-05, 1.064172e-05, 1.030564e-05, 1.33419e-05, 1.482878e-05, 
    1.364235e-05, 1.121702e-05, 9.714047e-06, 1.257722e-05, 1.912535e-05, 
    1.961959e-05, 1.457164e-05, 7.643986e-06, 7.789193e-06, 4.837767e-06,
  1.06952e-05, 1.203705e-05, 1.36912e-05, 1.337512e-05, 1.428432e-05, 
    1.345339e-05, 9.213642e-06, 8.909898e-06, 1.09058e-05, 1.414711e-05, 
    1.646071e-05, 1.053096e-05, 9.54168e-06, 7.460452e-06, 8.828369e-06,
  7.839218e-06, 1.017637e-05, 1.177056e-05, 1.309434e-05, 1.42255e-05, 
    1.190544e-05, 1.302457e-05, 9.286602e-06, 1.033616e-05, 1.076228e-05, 
    1.290356e-05, 1.472512e-05, 1.171809e-05, 1.269971e-05, 1.49011e-05,
  7.185284e-06, 7.407354e-06, 9.544687e-06, 1.096348e-05, 1.242565e-05, 
    1.296655e-05, 9.666464e-06, 9.236577e-06, 1.037617e-05, 8.327013e-06, 
    8.213514e-06, 1.039086e-05, 1.571683e-05, 2.072238e-05, 2.17537e-05,
  6.835779e-06, 4.824936e-06, 7.22309e-06, 8.239586e-06, 8.547699e-06, 
    9.763308e-06, 1.173826e-05, 1.183765e-05, 1.365795e-05, 1.134383e-05, 
    8.364622e-06, 9.01829e-06, 1.246714e-05, 1.409014e-05, 1.382366e-05,
  4.379665e-06, 4.940511e-06, 4.418032e-06, 6.27992e-06, 4.982073e-06, 
    4.085071e-06, 8.697519e-06, 1.165063e-05, 1.819241e-05, 1.536555e-05, 
    8.290079e-06, 6.139694e-06, 1.009294e-05, 1.262188e-05, 8.602283e-06,
  3.523222e-06, 7.535366e-06, 4.659406e-06, 4.732708e-06, 5.457915e-06, 
    5.093692e-06, 8.675278e-06, 1.014384e-05, 1.429002e-05, 1.134396e-05, 
    1.052483e-05, 8.198946e-06, 9.489711e-06, 9.254859e-06, 8.592937e-06,
  2.595172e-06, 6.140743e-06, 3.847224e-06, 3.938907e-06, 3.164922e-06, 
    3.555566e-06, 4.985364e-06, 9.281027e-06, 7.396958e-06, 1.052195e-05, 
    1.165971e-05, 9.164059e-06, 3.332291e-06, 6.366187e-06, 8.849001e-06,
  3.444715e-06, 2.730258e-06, 3.193275e-06, 6.535468e-06, 5.403712e-06, 
    3.71895e-06, 6.621774e-06, 6.902578e-06, 6.910784e-06, 6.926639e-06, 
    1.275229e-05, 1.22602e-05, 4.414257e-06, 6.259016e-06, 6.84368e-06,
  1.687466e-06, 1.245559e-06, 2.179362e-06, 3.615668e-06, 6.576615e-06, 
    7.871392e-06, 7.619046e-06, 9.186882e-06, 6.522783e-06, 6.487578e-06, 
    6.587095e-06, 7.681797e-06, 6.549647e-06, 6.760331e-06, 8.974418e-06,
  9.257927e-07, 1.107121e-06, 1.744787e-06, 2.937141e-06, 6.9526e-06, 
    3.907333e-06, 2.803539e-06, 3.259521e-06, 5.143484e-06, 6.458943e-06, 
    7.369963e-06, 1.110809e-05, 8.32082e-06, 9.818569e-06, 5.491187e-06,
  7.774613e-07, 1.228851e-06, 3.826255e-06, 2.553877e-06, 2.54246e-06, 
    5.560676e-06, 4.822727e-06, 5.673819e-06, 5.065142e-06, 7.149904e-06, 
    9.327779e-06, 1.014431e-05, 8.78532e-06, 1.129907e-05, 6.55438e-06,
  4.806969e-07, 3.049232e-07, 1.466935e-06, 1.406786e-06, 1.835704e-06, 
    4.128578e-06, 4.751009e-06, 4.101761e-06, 5.386805e-06, 6.92069e-06, 
    7.224769e-06, 8.360721e-06, 9.207522e-06, 1.027613e-05, 5.754463e-06,
  7.013071e-07, 2.052489e-07, 7.436172e-07, 2.59183e-06, 3.341628e-06, 
    3.9812e-06, 2.961404e-06, 3.622514e-06, 4.867894e-06, 5.694189e-06, 
    6.80428e-06, 9.176792e-06, 8.905362e-06, 6.911594e-06, 6.26587e-06,
  5.421758e-07, 8.160253e-07, 1.568987e-06, 4.47713e-06, 6.028436e-06, 
    9.855251e-06, 3.384479e-06, 2.584037e-06, 4.686222e-06, 6.738551e-06, 
    6.018609e-06, 6.636335e-06, 7.727166e-06, 6.349776e-06, 4.087871e-06,
  1.191748e-06, 2.464677e-06, 4.604327e-06, 9.847082e-06, 7.733121e-06, 
    8.140121e-06, 9.020567e-06, 5.265336e-06, 5.845e-06, 7.621004e-06, 
    7.163939e-06, 6.954034e-06, 3.630099e-06, 6.59236e-06, 3.789458e-06,
  5.964277e-06, 3.585298e-06, 6.026683e-06, 6.93592e-06, 5.289387e-06, 
    6.220925e-06, 4.813824e-06, 3.754618e-06, 3.645663e-06, 8.797771e-06, 
    8.775459e-06, 5.93914e-06, 4.355947e-06, 6.633888e-06, 4.85559e-06,
  4.641677e-06, 3.454395e-06, 2.438234e-06, 4.922453e-06, 6.378667e-06, 
    5.457974e-06, 4.262971e-06, 1.626001e-06, 4.696212e-06, 7.956657e-06, 
    9.825314e-06, 5.58467e-06, 2.572787e-06, 7.605212e-06, 6.265635e-06,
  1.263841e-06, 6.974781e-07, 1.533923e-07, 3.795363e-06, 7.813752e-06, 
    7.4862e-06, 9.294231e-06, 7.90452e-06, 4.115309e-06, 6.505711e-06, 
    8.951817e-06, 2.380439e-06, 4.749503e-06, 7.373813e-06, 5.108748e-06,
  3.271308e-07, 9.534484e-08, 2.283582e-09, 8.46084e-07, 7.710794e-06, 
    1.003612e-05, 1.07535e-05, 5.144943e-06, 4.62753e-06, 7.336749e-06, 
    5.976901e-06, 5.161083e-06, 4.906793e-06, 8.227924e-06, 4.531118e-06,
  0.0001513461, 0.0001800286, 0.0002022414, 0.0002402669, 0.0002697068, 
    0.000255654, 0.0002040752, 0.0001450608, 5.925721e-05, 1.312782e-05, 
    5.895962e-06, 4.472664e-06, 2.712257e-06, 4.784695e-06, 4.393996e-06,
  0.0001076665, 0.0001557154, 0.0001915468, 0.0002019243, 0.0001963576, 
    0.0002061196, 0.0001722917, 0.0001436611, 8.166715e-05, 2.615674e-05, 
    6.823405e-06, 4.415369e-06, 4.733254e-06, 4.092368e-06, 5.407687e-06,
  9.929827e-05, 0.0001341411, 0.0001635224, 0.0001686615, 0.0001403816, 
    0.0001209311, 0.0001102327, 0.0001003655, 8.560805e-05, 3.490709e-05, 
    9.107974e-06, 3.485615e-06, 4.319149e-06, 1.97593e-06, 2.601084e-06,
  9.52086e-05, 0.0001231706, 0.0001453663, 0.000147242, 0.0001292193, 
    8.407189e-05, 4.527923e-05, 6.570682e-05, 7.022832e-05, 3.688674e-05, 
    1.16479e-05, 2.874648e-06, 2.78494e-06, 4.999787e-07, 5.147819e-07,
  7.602488e-05, 0.0001125264, 0.0001369795, 0.000130243, 0.0001157529, 
    8.28035e-05, 2.393064e-05, 1.966262e-05, 4.805221e-05, 3.10312e-05, 
    9.447809e-06, 2.380465e-06, 2.709916e-06, 1.835533e-06, 1.174656e-08,
  2.727949e-05, 5.635238e-05, 8.098713e-05, 9.20322e-05, 9.950531e-05, 
    6.316407e-05, 2.338542e-05, 1.228372e-05, 2.590913e-05, 2.250618e-05, 
    6.792908e-06, 1.700964e-06, 1.603834e-06, 6.675096e-07, 2.655332e-08,
  2.963013e-06, 4.473822e-06, 1.872019e-05, 3.828178e-05, 4.033603e-05, 
    2.942539e-05, 1.666549e-05, 2.144922e-05, 1.474937e-05, 9.74673e-06, 
    5.080934e-06, 1.376757e-06, 1.214585e-06, 2.943128e-07, 6.282907e-08,
  5.959477e-06, 5.539279e-06, 4.402403e-06, 1.080828e-05, 1.157899e-05, 
    1.094404e-05, 9.172183e-06, 9.320658e-06, 1.613668e-05, 6.546464e-06, 
    5.270636e-06, 3.554098e-07, 6.677649e-07, 1.808909e-06, 1.819612e-06,
  5.663117e-06, 5.19476e-06, 3.085151e-06, 3.099117e-06, 4.760113e-06, 
    4.03258e-06, 3.411079e-06, 3.114208e-06, 5.849879e-06, 1.345409e-05, 
    6.64438e-06, 2.22605e-06, 3.879878e-07, 2.570139e-06, 5.369789e-06,
  3.694154e-06, 3.23484e-06, 6.28005e-07, 9.807598e-07, 3.604355e-06, 
    4.592845e-06, 5.991066e-06, 3.907845e-06, 4.156322e-06, 9.103367e-06, 
    9.424908e-06, 1.96937e-06, 1.226057e-06, 4.860065e-06, 7.599561e-06,
  0.0001290491, 0.0001459284, 0.0001581836, 0.0001295601, 7.04508e-05, 
    5.294478e-05, 7.560822e-05, 0.0001173787, 0.0001173443, 5.724247e-05, 
    4.261057e-05, 4.158137e-05, 3.105477e-05, 2.521588e-05, 2.226731e-05,
  0.0001225396, 0.0001737457, 0.0002046528, 0.0001524219, 7.947975e-05, 
    6.693646e-05, 6.485289e-05, 9.523845e-05, 0.0001588336, 0.0001367362, 
    6.456781e-05, 5.122312e-05, 4.487224e-05, 3.522358e-05, 1.243257e-05,
  0.000104222, 0.0001782385, 0.0002135832, 0.000148787, 9.171035e-05, 
    7.679734e-05, 7.570571e-05, 8.491504e-05, 0.0001387134, 0.0001960089, 
    0.0001755548, 0.0001076389, 8.171076e-05, 5.449234e-05, 2.547208e-05,
  8.781654e-05, 0.0001619496, 0.0002019284, 0.0001363506, 9.45536e-05, 
    9.240284e-05, 9.682884e-05, 9.643942e-05, 0.0001385942, 0.000235544, 
    0.0002365123, 0.0001833519, 0.0001255788, 7.15487e-05, 3.510262e-05,
  9.39789e-05, 0.0001463912, 0.0001858701, 0.0001251597, 9.345214e-05, 
    0.0001028115, 0.0001279191, 0.0001277701, 0.0001370224, 0.0001975071, 
    0.0002219372, 0.0001991392, 0.0001534302, 0.000103272, 4.591758e-05,
  0.0001832714, 0.0001977147, 0.0002123316, 0.0001463572, 0.0001197761, 
    0.0001308308, 0.0001529557, 0.0001415456, 0.0001424943, 0.0001438058, 
    0.0001707136, 0.0001654631, 0.0001336554, 9.689845e-05, 6.315444e-05,
  0.0002099142, 0.0002340746, 0.000249281, 0.0002126628, 0.0001656273, 
    0.0001658281, 0.0001643162, 0.0001507708, 0.0001572258, 0.0001460894, 
    0.0001408735, 0.0001378171, 0.0001119038, 7.573953e-05, 5.855701e-05,
  0.0001468807, 0.0001300835, 0.0001751536, 0.0001842238, 0.0001684184, 
    0.0001622111, 0.0001487558, 0.0001457629, 0.0001511258, 0.0001851303, 
    0.0001838173, 0.0001429841, 0.0001114939, 6.566844e-05, 4.645803e-05,
  0.0001369754, 6.047825e-05, 6.557895e-05, 9.913442e-05, 0.0001286435, 
    0.0001351406, 0.0001266456, 0.0001286177, 0.0001441726, 0.0002029435, 
    0.0002389767, 0.0001849701, 0.0001268894, 7.016723e-05, 3.572049e-05,
  0.0001618598, 6.289468e-05, 2.968803e-05, 4.323968e-05, 7.418393e-05, 
    0.0001014962, 0.0001092358, 0.0001134254, 0.0001391285, 0.0001996301, 
    0.0002494545, 0.0002039268, 0.000141347, 7.639654e-05, 3.009467e-05,
  9.838655e-05, 6.704631e-05, 3.836977e-05, 2.683537e-05, 1.973456e-05, 
    2.431613e-05, 2.615882e-05, 3.854158e-05, 3.554114e-05, 3.702759e-05, 
    2.8729e-05, 2.122433e-05, 1.315001e-05, 1.257793e-05, 9.977947e-06,
  6.1996e-05, 3.519071e-05, 3.250869e-05, 1.978576e-05, 2.370745e-05, 
    3.072431e-05, 3.415417e-05, 3.831733e-05, 4.922331e-05, 4.068993e-05, 
    2.791349e-05, 2.452405e-05, 1.381905e-05, 1.19859e-05, 8.228677e-06,
  6.794349e-05, 3.140982e-05, 3.29026e-05, 2.275142e-05, 2.954946e-05, 
    3.544131e-05, 4.347703e-05, 6.368297e-05, 7.835463e-05, 6.291514e-05, 
    4.136032e-05, 2.152158e-05, 1.267402e-05, 9.94545e-06, 6.933252e-06,
  9.817532e-05, 3.740454e-05, 2.332221e-05, 3.00018e-05, 4.137387e-05, 
    4.80848e-05, 6.526502e-05, 8.968718e-05, 0.0001136478, 0.0001075725, 
    6.871361e-05, 2.981875e-05, 1.347953e-05, 1.000736e-05, 8.820898e-06,
  0.0001433278, 5.38996e-05, 2.960107e-05, 3.53269e-05, 4.953857e-05, 
    5.901094e-05, 8.265166e-05, 0.0001256924, 0.0001627419, 0.0001544696, 
    0.0001085361, 5.012181e-05, 1.892895e-05, 9.96977e-06, 6.292974e-06,
  0.000190963, 9.290347e-05, 3.412426e-05, 4.07542e-05, 4.170309e-05, 
    6.480448e-05, 9.61286e-05, 0.0001520392, 0.0001876815, 0.000158232, 
    0.0001062746, 5.295761e-05, 2.384513e-05, 1.037354e-05, 6.491821e-06,
  0.000235131, 0.0001609929, 7.284861e-05, 4.635433e-05, 3.461871e-05, 
    5.573922e-05, 9.741703e-05, 0.0001597532, 0.000173989, 0.0001138355, 
    6.111427e-05, 3.873562e-05, 2.047053e-05, 1.141755e-05, 6.95664e-06,
  0.0002046387, 0.0002215119, 0.0001605968, 8.097294e-05, 3.830194e-05, 
    5.48297e-05, 9.358882e-05, 0.0001464112, 0.0001403516, 8.121914e-05, 
    3.845834e-05, 2.297052e-05, 1.265205e-05, 9.745482e-06, 5.971486e-06,
  0.0001993839, 0.0002015847, 0.0002169795, 0.0001288066, 5.494592e-05, 
    4.744377e-05, 8.648662e-05, 0.0001384825, 0.0001063688, 9.132392e-05, 
    9.544604e-05, 4.033328e-05, 8.92824e-06, 1.023104e-05, 9.922249e-06,
  0.0002455737, 0.0001613521, 0.0002187621, 0.0001567684, 6.141183e-05, 
    4.322049e-05, 7.096625e-05, 0.0001181052, 9.075179e-05, 0.0001402207, 
    0.0001916179, 8.275941e-05, 1.487161e-05, 1.57831e-05, 1.064015e-05,
  6.281794e-06, 5.879104e-06, 5.678919e-06, 4.70838e-06, 6.112848e-06, 
    5.186796e-06, 5.562541e-06, 6.592081e-06, 7.1192e-06, 6.576829e-06, 
    7.67146e-06, 8.288822e-06, 8.40241e-06, 9.332874e-06, 9.062166e-06,
  6.790701e-06, 6.873092e-06, 6.449754e-06, 5.993612e-06, 6.281882e-06, 
    7.253476e-06, 6.447067e-06, 7.79432e-06, 8.984946e-06, 8.695067e-06, 
    7.764609e-06, 8.522651e-06, 1.058374e-05, 1.101834e-05, 1.045766e-05,
  8.006527e-06, 6.427091e-06, 6.492309e-06, 7.089813e-06, 6.552716e-06, 
    8.153434e-06, 7.283682e-06, 7.274632e-06, 1.086641e-05, 9.87597e-06, 
    7.84794e-06, 9.113101e-06, 9.922918e-06, 1.076704e-05, 1.082521e-05,
  7.233547e-06, 7.944787e-06, 8.364397e-06, 7.399571e-06, 8.986708e-06, 
    9.577591e-06, 7.922806e-06, 9.015608e-06, 1.050799e-05, 1.205066e-05, 
    1.040309e-05, 1.070937e-05, 1.018286e-05, 1.002094e-05, 1.087192e-05,
  1.012092e-05, 8.940941e-06, 1.101373e-05, 1.029914e-05, 9.590856e-06, 
    9.390109e-06, 1.145163e-05, 1.172319e-05, 1.203526e-05, 1.285758e-05, 
    1.255552e-05, 1.186954e-05, 1.077776e-05, 1.098137e-05, 1.414068e-05,
  1.18039e-05, 1.073267e-05, 1.195648e-05, 1.068035e-05, 1.252712e-05, 
    1.187156e-05, 1.133944e-05, 1.49654e-05, 1.536295e-05, 1.514582e-05, 
    1.444544e-05, 1.329443e-05, 1.369312e-05, 1.394535e-05, 1.545611e-05,
  1.167564e-05, 1.336094e-05, 1.269072e-05, 1.647665e-05, 1.588399e-05, 
    1.539604e-05, 1.306695e-05, 1.546573e-05, 1.749837e-05, 2.139721e-05, 
    1.891443e-05, 1.585455e-05, 1.56363e-05, 2.058973e-05, 1.671388e-05,
  1.166524e-05, 1.376376e-05, 1.400292e-05, 1.471902e-05, 1.732805e-05, 
    1.719575e-05, 1.858072e-05, 1.739567e-05, 1.818343e-05, 1.990093e-05, 
    2.258115e-05, 1.997124e-05, 2.279604e-05, 2.218771e-05, 1.630847e-05,
  1.25802e-05, 1.101974e-05, 1.381297e-05, 1.877191e-05, 1.986683e-05, 
    2.259771e-05, 1.72492e-05, 2.224073e-05, 1.903054e-05, 2.778154e-05, 
    2.956121e-05, 2.385167e-05, 2.319494e-05, 2.977756e-05, 1.988487e-05,
  1.178929e-05, 1.335327e-05, 1.436007e-05, 2.101126e-05, 2.091586e-05, 
    2.963853e-05, 2.806435e-05, 2.776922e-05, 3.231833e-05, 3.744337e-05, 
    4.38906e-05, 4.833504e-05, 3.362403e-05, 4.149842e-05, 3.171812e-05,
  9.802917e-06, 9.291658e-06, 9.94269e-06, 8.746189e-06, 9.486838e-06, 
    6.933178e-06, 5.293814e-06, 5.555893e-06, 7.113676e-06, 6.789878e-06, 
    5.972734e-06, 4.498419e-06, 3.858614e-06, 4.705833e-06, 3.633091e-06,
  9.963814e-06, 8.611148e-06, 7.936632e-06, 8.028767e-06, 7.856219e-06, 
    7.328575e-06, 4.377654e-06, 6.301312e-06, 1.006688e-05, 6.358979e-06, 
    6.73306e-06, 6.563019e-06, 6.64654e-06, 5.370564e-06, 5.138834e-06,
  9.280717e-06, 8.658029e-06, 7.708615e-06, 7.599875e-06, 8.754042e-06, 
    9.157267e-06, 8.45916e-06, 7.869312e-06, 9.379065e-06, 9.500943e-06, 
    9.295673e-06, 8.481475e-06, 7.320411e-06, 8.068137e-06, 6.306649e-06,
  9.100049e-06, 8.070058e-06, 8.710344e-06, 8.282851e-06, 9.843652e-06, 
    1.333137e-05, 1.050818e-05, 1.279402e-05, 1.46825e-05, 1.315506e-05, 
    1.252515e-05, 1.275512e-05, 1.529131e-05, 1.377798e-05, 1.715568e-05,
  1.163069e-05, 1.100193e-05, 1.025059e-05, 1.089129e-05, 1.137186e-05, 
    1.100259e-05, 1.243622e-05, 1.443321e-05, 1.936979e-05, 2.072741e-05, 
    2.083223e-05, 2.232646e-05, 2.383382e-05, 2.307353e-05, 2.546942e-05,
  1.512599e-05, 1.408682e-05, 1.184087e-05, 1.004086e-05, 1.241374e-05, 
    1.290347e-05, 1.046506e-05, 1.238871e-05, 1.494737e-05, 1.799705e-05, 
    1.677265e-05, 1.71885e-05, 1.565386e-05, 2.324775e-05, 1.056126e-05,
  1.499683e-05, 1.338627e-05, 1.281165e-05, 1.311538e-05, 1.210207e-05, 
    1.030261e-05, 8.664735e-06, 9.373402e-06, 1.320286e-05, 1.30779e-05, 
    8.318257e-06, 1.005692e-05, 9.745992e-06, 1.225734e-05, 6.808395e-06,
  1.521059e-05, 1.244283e-05, 1.212508e-05, 1.177782e-05, 1.222835e-05, 
    9.551516e-06, 8.575003e-06, 9.283559e-06, 1.017623e-05, 8.858029e-06, 
    6.876016e-06, 7.565306e-06, 6.75469e-06, 5.138519e-06, 5.724361e-06,
  1.55019e-05, 1.547886e-05, 1.487863e-05, 1.353276e-05, 1.192276e-05, 
    9.930545e-06, 9.524344e-06, 7.239442e-06, 7.424146e-06, 9.730153e-06, 
    6.802238e-06, 6.23902e-06, 5.057536e-06, 4.399868e-06, 3.067838e-06,
  1.856521e-05, 1.799259e-05, 1.695759e-05, 1.504808e-05, 1.267636e-05, 
    1.246767e-05, 1.03265e-05, 7.842406e-06, 7.449249e-06, 7.355182e-06, 
    6.374843e-06, 6.830566e-06, 3.873481e-06, 2.643851e-06, 1.533711e-06,
  7.431626e-06, 7.631022e-06, 1.097362e-05, 1.247328e-05, 1.595229e-05, 
    3.262111e-05, 9.113988e-05, 0.000160966, 0.0001852222, 0.0001609238, 
    0.0001385029, 0.0001171562, 0.0001196198, 0.0001271289, 0.0001354965,
  6.004781e-06, 7.312442e-06, 1.00045e-05, 1.430816e-05, 2.097449e-05, 
    3.430384e-05, 6.939828e-05, 0.0001225131, 0.0001711072, 0.0001595586, 
    0.0001210992, 8.704953e-05, 6.997627e-05, 6.788799e-05, 7.199506e-05,
  3.321376e-06, 5.164703e-06, 9.686665e-06, 1.172913e-05, 1.286484e-05, 
    2.669813e-05, 6.367079e-05, 0.0001050232, 0.00013364, 0.000137486, 
    0.0001222361, 0.0001002489, 7.375646e-05, 6.713984e-05, 6.32253e-05,
  4.465424e-06, 6.54084e-06, 8.979651e-06, 1.10848e-05, 9.491259e-06, 
    1.49389e-05, 3.263198e-05, 6.833823e-05, 8.879205e-05, 0.0001013324, 
    0.0001027423, 9.60531e-05, 8.158276e-05, 7.497422e-05, 7.242766e-05,
  5.415281e-06, 7.232314e-06, 7.124931e-06, 9.943344e-06, 1.052969e-05, 
    1.123904e-05, 1.472466e-05, 2.315888e-05, 5.055732e-05, 6.97068e-05, 
    7.865143e-05, 8.336606e-05, 8.513586e-05, 8.060255e-05, 8.479617e-05,
  3.521646e-06, 4.825066e-06, 6.720717e-06, 8.961181e-06, 8.513577e-06, 
    1.014867e-05, 1.246704e-05, 1.180497e-05, 1.973298e-05, 3.153154e-05, 
    4.753321e-05, 6.212785e-05, 7.131731e-05, 7.964612e-05, 8.772156e-05,
  2.57081e-06, 2.214938e-06, 3.136397e-06, 6.181087e-06, 9.650994e-06, 
    5.339189e-06, 6.959664e-06, 9.656035e-06, 9.064582e-06, 1.034915e-05, 
    1.443478e-05, 2.639691e-05, 4.930165e-05, 6.13567e-05, 7.50422e-05,
  6.198441e-07, 1.497825e-06, 1.831217e-06, 3.556033e-06, 6.266806e-06, 
    5.619198e-06, 4.056214e-06, 5.753644e-06, 6.734329e-06, 5.355298e-06, 
    5.263475e-06, 6.278115e-06, 1.39053e-05, 2.923741e-05, 4.648527e-05,
  1.213233e-06, 1.45128e-06, 1.101612e-06, 1.56158e-06, 2.590888e-06, 
    3.883558e-06, 3.336955e-06, 2.47712e-06, 3.884061e-06, 4.877324e-06, 
    2.567702e-06, 1.58874e-06, 2.455705e-06, 7.458957e-06, 1.25732e-05,
  4.055554e-06, 3.336682e-06, 2.507973e-06, 4.794834e-06, 2.246624e-06, 
    2.221559e-06, 3.007322e-06, 2.793078e-06, 2.794591e-06, 3.754474e-06, 
    3.685766e-06, 1.256315e-06, 1.514358e-06, 2.486764e-06, 2.674112e-06,
  1.025747e-05, 3.373729e-05, 0.0001456996, 0.0003213999, 0.0004345768, 
    0.0003182783, 0.000167935, 7.695427e-05, 2.871109e-05, 3.372921e-05, 
    6.705186e-05, 0.0001156889, 0.0001541507, 0.0001546549, 0.000124756,
  3.065623e-05, 5.230451e-05, 0.0002325913, 0.0004869926, 0.0005255315, 
    0.0003166741, 0.0002020888, 0.0001315269, 6.449225e-05, 2.951265e-05, 
    5.323753e-05, 0.000101709, 0.0001761846, 0.0001309327, 8.101609e-05,
  4.518736e-05, 8.909811e-05, 0.0003487291, 0.00065669, 0.0006341779, 
    0.0003658008, 0.0002259181, 0.0001689805, 0.0001036457, 5.645029e-05, 
    5.325584e-05, 9.612164e-05, 0.0001380829, 8.069498e-05, 5.26518e-05,
  5.853389e-05, 0.0001287799, 0.0004756801, 0.0007499175, 0.0006317442, 
    0.000383068, 0.000269088, 0.0001976699, 0.000133325, 8.156127e-05, 
    6.119499e-05, 9.889741e-05, 9.368684e-05, 4.406292e-05, 3.720392e-05,
  8.225963e-05, 0.0002591567, 0.0005685121, 0.0007198215, 0.0004802133, 
    0.0003262133, 0.0002691789, 0.0002162735, 0.0001541489, 9.780088e-05, 
    7.488234e-05, 8.953425e-05, 6.366039e-05, 3.461908e-05, 4.737191e-05,
  0.0001510963, 0.0003375873, 0.0005587475, 0.0005856282, 0.0003696806, 
    0.0002777997, 0.000238034, 0.0001985661, 0.0001678895, 0.0001241667, 
    9.131264e-05, 7.797503e-05, 5.093627e-05, 4.285618e-05, 8.663921e-05,
  0.0001584307, 0.0002914032, 0.0004446099, 0.0004328574, 0.0002829924, 
    0.0002221669, 0.0001930219, 0.0001692173, 0.0001569703, 0.0001392264, 
    0.0001163159, 9.768492e-05, 6.960328e-05, 7.339974e-05, 0.0001497751,
  7.548363e-05, 0.0001626348, 0.0002610054, 0.0002773394, 0.0002110441, 
    0.0001615675, 0.0001512911, 0.0001408749, 0.0001384604, 0.0001354007, 
    0.0001311002, 0.0001207769, 0.0001094274, 0.0001226942, 0.0002240774,
  1.858731e-05, 4.847804e-05, 0.000110268, 0.0001382353, 0.0001336001, 
    0.0001309329, 0.0001174401, 0.0001103778, 0.000117087, 0.0001237338, 
    0.0001316243, 0.0001293737, 0.0001294513, 0.000164, 0.0003005764,
  7.487777e-06, 1.556317e-05, 2.879919e-05, 4.025918e-05, 6.68977e-05, 
    9.048658e-05, 9.826552e-05, 9.904835e-05, 9.64756e-05, 0.0001078304, 
    0.0001279693, 0.0001318465, 0.0001306367, 0.0001752949, 0.0003379182,
  0.0003579546, 0.0001469968, 9.889053e-05, 0.0002035554, 0.0003921092, 
    0.0003364728, 0.0002140604, 0.0001626068, 0.0001528038, 0.0001140555, 
    7.946569e-05, 3.158104e-05, 1.263758e-05, 7.206617e-06, 5.987694e-06,
  0.0004000124, 0.0002094172, 9.861556e-05, 0.0001753306, 0.0004151046, 
    0.0003603506, 0.000186181, 0.0001103988, 0.0001055647, 8.192773e-05, 
    6.105482e-05, 2.926322e-05, 1.282549e-05, 8.527694e-06, 7.560018e-06,
  0.000482776, 0.000398845, 0.0002152913, 0.000207282, 0.0003623326, 
    0.0003234356, 0.0001278626, 6.504424e-05, 6.421214e-05, 5.621586e-05, 
    4.625183e-05, 2.637898e-05, 1.436186e-05, 1.031758e-05, 9.093525e-06,
  0.0005084344, 0.0005391451, 0.0004720558, 0.0003442672, 0.0003692679, 
    0.0002806326, 6.876561e-05, 3.465076e-05, 3.939835e-05, 4.473012e-05, 
    3.577287e-05, 2.956938e-05, 1.721575e-05, 9.844417e-06, 9.236584e-06,
  0.0004623064, 0.000561801, 0.0006872141, 0.0006110992, 0.0004656584, 
    0.0002951118, 3.500253e-05, 2.635208e-05, 3.457569e-05, 3.42067e-05, 
    3.404298e-05, 3.10751e-05, 1.504926e-05, 9.274956e-06, 8.796682e-06,
  0.0003171775, 0.0004903522, 0.000780726, 0.0008198259, 0.0005285495, 
    0.0003048075, 1.953067e-05, 1.876844e-05, 3.31418e-05, 3.083907e-05, 
    3.247533e-05, 3.016552e-05, 1.274469e-05, 7.840183e-06, 8.658833e-06,
  0.000195419, 0.0003905733, 0.0007764194, 0.0008724572, 0.0005107973, 
    0.0002941024, 1.759069e-05, 1.763085e-05, 3.452212e-05, 2.998781e-05, 
    2.777064e-05, 1.847694e-05, 9.944607e-06, 9.555428e-06, 8.448358e-06,
  0.0001178159, 0.0003275016, 0.0007553016, 0.0008553177, 0.0004873854, 
    0.000290251, 3.384533e-05, 1.700086e-05, 2.891983e-05, 2.995572e-05, 
    1.77031e-05, 9.210606e-06, 9.617565e-06, 1.130678e-05, 1.082103e-05,
  8.682322e-05, 0.0002124405, 0.0006289329, 0.0007843029, 0.0004599223, 
    0.0002937917, 7.467117e-05, 1.948173e-05, 1.86868e-05, 2.757444e-05, 
    1.23742e-05, 6.529249e-06, 8.482636e-06, 1.198327e-05, 9.50904e-06,
  4.776526e-05, 0.0001397828, 0.0004749656, 0.0006898918, 0.0004513356, 
    0.0003093244, 0.0001462332, 2.627016e-05, 1.111283e-05, 2.425022e-05, 
    1.431419e-05, 7.675229e-06, 1.016556e-05, 1.057682e-05, 1.046764e-05,
  3.701934e-05, 2.154978e-05, 1.351902e-05, 9.077009e-06, 1.297608e-05, 
    1.156761e-05, 9.35783e-06, 6.095466e-06, 7.151863e-06, 6.169924e-06, 
    6.626149e-06, 6.678282e-06, 5.6215e-06, 7.720304e-06, 1.103431e-05,
  9.904161e-05, 4.453738e-05, 1.752042e-05, 1.043525e-05, 1.204708e-05, 
    1.086612e-05, 9.135711e-06, 7.49442e-06, 6.9741e-06, 6.132724e-06, 
    6.296488e-06, 4.899701e-06, 3.871737e-06, 5.850865e-06, 9.50204e-06,
  0.0001910616, 0.0001362253, 4.700447e-05, 1.294426e-05, 1.178006e-05, 
    1.2184e-05, 1.083563e-05, 8.152091e-06, 6.393621e-06, 4.622324e-06, 
    4.684613e-06, 4.378533e-06, 2.286719e-06, 2.740005e-06, 7.843561e-06,
  0.0001967013, 0.0002599632, 0.0001431275, 1.363878e-05, 1.189264e-05, 
    1.268353e-05, 9.38525e-06, 9.550375e-06, 7.918113e-06, 4.672718e-06, 
    3.366318e-06, 3.426122e-06, 2.146387e-06, 1.848829e-06, 4.855399e-06,
  0.0001633306, 0.0004319387, 0.0002729137, 3.723789e-05, 1.654046e-05, 
    1.16351e-05, 8.798343e-06, 8.906679e-06, 8.482893e-06, 4.782388e-06, 
    2.575346e-06, 2.051232e-06, 1.974361e-06, 1.862073e-06, 3.172022e-06,
  0.0002212734, 0.0005743693, 0.0004464326, 9.840278e-05, 1.211231e-05, 
    1.249289e-05, 7.924795e-06, 8.570551e-06, 7.918215e-06, 5.67644e-06, 
    2.781971e-06, 1.64064e-06, 1.809754e-06, 1.617074e-06, 1.880335e-06,
  0.0002331392, 0.000605514, 0.0006798127, 0.000224455, 1.492371e-05, 
    1.377267e-05, 1.080599e-05, 9.52205e-06, 8.798379e-06, 4.692609e-06, 
    2.125192e-06, 2.112472e-06, 1.652277e-06, 7.829626e-07, 1.030031e-06,
  0.0002098092, 0.0005232657, 0.0008301024, 0.0003689666, 4.747372e-05, 
    9.444464e-06, 1.301204e-05, 8.060249e-06, 7.447812e-06, 4.627808e-06, 
    4.2303e-06, 2.311612e-06, 1.203237e-06, 1.838223e-06, 1.338785e-06,
  0.0001937057, 0.0004626338, 0.000808911, 0.0006318099, 0.0001244983, 
    4.759181e-06, 1.29916e-05, 8.320735e-06, 5.881163e-06, 5.148357e-06, 
    1.864289e-06, 1.767749e-06, 1.654195e-06, 1.162305e-06, 1.572803e-06,
  0.0001832372, 0.0004175425, 0.0007989063, 0.0008815113, 0.0002302487, 
    9.820127e-06, 6.292525e-06, 8.368396e-06, 5.441232e-06, 4.29181e-06, 
    1.808287e-06, 1.466937e-06, 1.196661e-06, 1.551448e-06, 1.483415e-06,
  1.072117e-05, 1.182884e-05, 9.537312e-06, 9.267013e-06, 1.080101e-05, 
    1.266408e-05, 1.098206e-05, 1.278258e-05, 1.656831e-05, 1.746488e-05, 
    1.713848e-05, 1.782634e-05, 1.607877e-05, 1.471399e-05, 1.030846e-05,
  1.825142e-05, 1.494518e-05, 8.980655e-06, 9.349052e-06, 1.050253e-05, 
    1.15778e-05, 9.279462e-06, 1.046129e-05, 1.33675e-05, 1.486324e-05, 
    1.794445e-05, 1.892634e-05, 1.994459e-05, 1.894679e-05, 1.399445e-05,
  2.492902e-05, 1.94888e-05, 1.534167e-05, 1.223365e-05, 9.854231e-06, 
    1.029888e-05, 7.948137e-06, 7.621092e-06, 1.020727e-05, 9.993582e-06, 
    1.132544e-05, 1.355887e-05, 1.50018e-05, 1.592432e-05, 1.302464e-05,
  3.647926e-05, 2.833849e-05, 2.064498e-05, 1.368517e-05, 1.112463e-05, 
    1.079547e-05, 1.002822e-05, 6.115174e-06, 6.17968e-06, 7.512522e-06, 
    8.752722e-06, 8.059151e-06, 1.020127e-05, 1.230546e-05, 1.032403e-05,
  4.883995e-05, 3.735815e-05, 2.551241e-05, 1.897361e-05, 1.406384e-05, 
    1.095518e-05, 8.603226e-06, 9.231649e-06, 7.644299e-06, 7.877415e-06, 
    6.82579e-06, 7.351402e-06, 7.61042e-06, 8.552e-06, 1.034721e-05,
  6.430708e-05, 5.023838e-05, 3.330268e-05, 2.55339e-05, 1.930961e-05, 
    1.240327e-05, 8.149943e-06, 1.107543e-05, 6.842897e-06, 5.629523e-06, 
    8.270539e-06, 5.586601e-06, 6.603202e-06, 8.725955e-06, 1.033217e-05,
  8.329598e-05, 6.20631e-05, 3.778173e-05, 3.069455e-05, 2.53121e-05, 
    1.510305e-05, 1.026745e-05, 9.539811e-06, 6.958644e-06, 5.518491e-06, 
    6.583698e-06, 6.326945e-06, 6.314808e-06, 7.663823e-06, 9.151691e-06,
  8.605101e-05, 7.746828e-05, 5.035429e-05, 3.432023e-05, 2.331262e-05, 
    1.886286e-05, 1.313949e-05, 1.0143e-05, 7.175979e-06, 5.993172e-06, 
    5.186088e-06, 4.819925e-06, 6.674341e-06, 7.145234e-06, 6.625435e-06,
  8.340042e-05, 9.186674e-05, 6.534038e-05, 4.098721e-05, 2.078137e-05, 
    1.747156e-05, 1.572234e-05, 1.196018e-05, 9.191271e-06, 6.071367e-06, 
    5.694357e-06, 5.380948e-06, 5.619492e-06, 7.502195e-06, 8.20783e-06,
  4.391629e-05, 7.338291e-05, 9.557512e-05, 4.486818e-05, 2.453132e-05, 
    1.023522e-05, 1.223802e-05, 1.262725e-05, 1.168945e-05, 6.858885e-06, 
    5.640609e-06, 4.682469e-06, 5.619081e-06, 9.097029e-06, 9.78256e-06,
  2.652944e-05, 2.540923e-05, 2.081321e-05, 2.03759e-05, 1.816417e-05, 
    1.681267e-05, 1.628699e-05, 1.307831e-05, 1.548726e-05, 1.570043e-05, 
    1.298513e-05, 1.376798e-05, 1.189586e-05, 1.108938e-05, 9.932219e-06,
  2.94278e-05, 2.953057e-05, 2.500021e-05, 2.33817e-05, 2.240671e-05, 
    2.113622e-05, 1.666259e-05, 1.582588e-05, 1.851646e-05, 1.696947e-05, 
    1.705348e-05, 1.675818e-05, 1.427524e-05, 1.491039e-05, 1.298797e-05,
  3.66552e-05, 3.30186e-05, 2.62702e-05, 1.930651e-05, 2.153488e-05, 
    2.52066e-05, 1.952194e-05, 1.7628e-05, 2.060237e-05, 1.822971e-05, 
    1.797401e-05, 1.832692e-05, 1.825173e-05, 1.796163e-05, 1.442257e-05,
  3.866573e-05, 3.680199e-05, 2.774556e-05, 2.249816e-05, 2.932447e-05, 
    2.64725e-05, 1.912897e-05, 2.241304e-05, 2.054184e-05, 1.976704e-05, 
    2.214522e-05, 1.80566e-05, 1.746092e-05, 1.781232e-05, 1.642926e-05,
  4.480297e-05, 3.819973e-05, 3.301341e-05, 3.771807e-05, 2.861409e-05, 
    2.575294e-05, 2.017814e-05, 1.991103e-05, 2.177474e-05, 2.2104e-05, 
    1.84385e-05, 1.910324e-05, 1.87854e-05, 1.513499e-05, 1.58245e-05,
  5.145586e-05, 4.838361e-05, 4.128701e-05, 4.44667e-05, 3.661949e-05, 
    3.521348e-05, 2.571918e-05, 2.010866e-05, 3.000361e-05, 2.501745e-05, 
    2.165855e-05, 1.752911e-05, 1.362912e-05, 1.577749e-05, 1.594213e-05,
  5.832479e-05, 5.883124e-05, 3.810999e-05, 4.105817e-05, 3.68923e-05, 
    4.060974e-05, 2.855953e-05, 3.119248e-05, 3.718763e-05, 3.1283e-05, 
    2.452491e-05, 1.859447e-05, 1.824416e-05, 1.5298e-05, 1.461791e-05,
  4.746613e-05, 4.863518e-05, 5.476022e-05, 4.363247e-05, 4.713355e-05, 
    3.569829e-05, 3.767203e-05, 3.672629e-05, 3.760338e-05, 3.656041e-05, 
    2.591476e-05, 2.365841e-05, 2.059889e-05, 1.97538e-05, 1.859805e-05,
  6.936338e-05, 5.837739e-05, 5.73105e-05, 4.582956e-05, 5.341393e-05, 
    3.383907e-05, 3.242677e-05, 3.182213e-05, 3.800542e-05, 2.640046e-05, 
    3.184903e-05, 2.696137e-05, 3.048047e-05, 2.648361e-05, 2.553696e-05,
  0.0001554669, 0.0001015712, 6.461525e-05, 5.556159e-05, 5.3471e-05, 
    5.169983e-05, 5.570152e-05, 4.794851e-05, 3.621505e-05, 4.349164e-05, 
    3.361281e-05, 3.509238e-05, 3.279791e-05, 3.597227e-05, 3.485872e-05,
  1.524692e-05, 1.795282e-05, 1.614593e-05, 1.559084e-05, 1.690799e-05, 
    1.900165e-05, 1.580435e-05, 1.488403e-05, 1.667132e-05, 1.44322e-05, 
    1.326767e-05, 1.512311e-05, 1.169138e-05, 1.286997e-05, 1.192098e-05,
  1.598298e-05, 1.642243e-05, 1.768784e-05, 1.856548e-05, 1.88031e-05, 
    2.104326e-05, 1.793986e-05, 2.084113e-05, 2.036124e-05, 2.057324e-05, 
    1.971533e-05, 1.76855e-05, 1.584422e-05, 1.342322e-05, 1.16014e-05,
  1.595282e-05, 2.067708e-05, 1.90477e-05, 1.20986e-05, 1.810052e-05, 
    2.057532e-05, 1.836384e-05, 1.877926e-05, 1.89798e-05, 2.4011e-05, 
    2.148283e-05, 2.123512e-05, 1.807742e-05, 1.459703e-05, 1.30517e-05,
  1.737609e-05, 2.14702e-05, 1.839437e-05, 1.766244e-05, 2.360567e-05, 
    1.931696e-05, 1.627661e-05, 1.902585e-05, 2.218932e-05, 1.979758e-05, 
    1.876167e-05, 2.063941e-05, 1.890649e-05, 1.869222e-05, 1.633066e-05,
  2.204301e-05, 2.394839e-05, 2.493219e-05, 2.665117e-05, 2.156855e-05, 
    2.013727e-05, 2.149545e-05, 1.992058e-05, 2.097565e-05, 2.157835e-05, 
    2.029767e-05, 1.782979e-05, 2.034346e-05, 1.990713e-05, 2.097199e-05,
  2.450051e-05, 2.797811e-05, 2.785652e-05, 2.650849e-05, 2.616793e-05, 
    2.517461e-05, 2.470634e-05, 2.459055e-05, 2.291432e-05, 2.158431e-05, 
    2.075929e-05, 1.926372e-05, 2.017698e-05, 2.226471e-05, 2.225566e-05,
  2.885796e-05, 3.008182e-05, 3.107476e-05, 3.135126e-05, 2.982149e-05, 
    2.712061e-05, 2.474822e-05, 2.437005e-05, 2.805174e-05, 2.533725e-05, 
    2.204356e-05, 2.114434e-05, 2.395713e-05, 2.500964e-05, 2.442202e-05,
  3.285678e-05, 3.259107e-05, 3.224845e-05, 3.047183e-05, 3.117543e-05, 
    3.020237e-05, 2.448148e-05, 2.173129e-05, 2.675114e-05, 2.389337e-05, 
    2.431582e-05, 2.457614e-05, 3.188573e-05, 3.043374e-05, 2.647616e-05,
  3.070431e-05, 3.379633e-05, 2.820139e-05, 2.911042e-05, 3.377144e-05, 
    3.436044e-05, 2.659992e-05, 2.621075e-05, 2.317001e-05, 2.222114e-05, 
    2.282946e-05, 2.945233e-05, 3.256219e-05, 3.264345e-05, 2.770887e-05,
  4.450671e-05, 3.774812e-05, 2.617328e-05, 2.904479e-05, 3.019391e-05, 
    2.820195e-05, 2.606738e-05, 2.398437e-05, 2.405174e-05, 2.560241e-05, 
    2.808454e-05, 3.258403e-05, 3.214548e-05, 3.594637e-05, 3.850917e-05,
  2.120664e-05, 2.050537e-05, 1.97445e-05, 1.719266e-05, 1.680251e-05, 
    1.408114e-05, 1.159257e-05, 1.198525e-05, 1.124926e-05, 8.387966e-06, 
    7.089914e-06, 6.198042e-06, 4.129095e-06, 4.921953e-06, 4.263447e-06,
  2.801326e-05, 2.601003e-05, 2.067052e-05, 1.799789e-05, 1.771822e-05, 
    1.64875e-05, 1.332023e-05, 1.088595e-05, 1.145989e-05, 9.580548e-06, 
    8.191671e-06, 7.328719e-06, 8.128015e-06, 6.562012e-06, 4.616023e-06,
  3.549872e-05, 2.989177e-05, 2.462631e-05, 2.125293e-05, 2.067442e-05, 
    1.554811e-05, 1.483407e-05, 1.431748e-05, 1.294965e-05, 1.350435e-05, 
    1.08475e-05, 1.096397e-05, 1.170763e-05, 8.541032e-06, 8.591916e-06,
  3.238747e-05, 3.011238e-05, 2.366121e-05, 2.091652e-05, 1.848901e-05, 
    1.763984e-05, 1.81198e-05, 1.437445e-05, 1.494736e-05, 1.406689e-05, 
    1.346957e-05, 1.698894e-05, 1.204916e-05, 1.149231e-05, 1.163647e-05,
  3.544206e-05, 2.828183e-05, 2.361394e-05, 2.139073e-05, 2.131905e-05, 
    2.120906e-05, 1.528612e-05, 1.743262e-05, 1.874225e-05, 1.775893e-05, 
    1.782978e-05, 1.756036e-05, 1.829469e-05, 1.268836e-05, 1.446826e-05,
  3.525681e-05, 2.994704e-05, 2.549229e-05, 2.544552e-05, 2.596738e-05, 
    2.323804e-05, 2.01782e-05, 2.142667e-05, 2.37091e-05, 2.236201e-05, 
    2.631205e-05, 2.3397e-05, 2.258521e-05, 1.847558e-05, 1.386654e-05,
  3.906349e-05, 3.056627e-05, 2.724744e-05, 2.961293e-05, 2.959017e-05, 
    2.948637e-05, 2.415084e-05, 2.366428e-05, 2.871465e-05, 2.953255e-05, 
    3.190829e-05, 3.202401e-05, 2.953383e-05, 1.842784e-05, 1.788143e-05,
  4.021635e-05, 3.21491e-05, 3.214699e-05, 3.613685e-05, 2.869326e-05, 
    3.444397e-05, 2.796526e-05, 2.938873e-05, 3.570653e-05, 3.276074e-05, 
    3.585239e-05, 3.715175e-05, 2.882286e-05, 2.306932e-05, 2.298607e-05,
  4.182626e-05, 3.671161e-05, 3.86444e-05, 3.726307e-05, 3.269033e-05, 
    3.911816e-05, 3.361258e-05, 3.694888e-05, 3.435212e-05, 4.063406e-05, 
    4.271267e-05, 3.58559e-05, 3.294798e-05, 2.998589e-05, 2.943214e-05,
  4.510748e-05, 4.069957e-05, 4.471449e-05, 4.338859e-05, 4.103703e-05, 
    4.602093e-05, 3.637809e-05, 3.86088e-05, 4.702593e-05, 4.764608e-05, 
    3.705298e-05, 4.131525e-05, 3.095489e-05, 3.551457e-05, 3.766371e-05,
  4.740726e-06, 3.615025e-06, 2.835193e-06, 4.196779e-06, 4.250864e-06, 
    4.137095e-06, 3.490201e-06, 4.843704e-06, 5.021172e-06, 4.532419e-06, 
    5.071776e-06, 3.594247e-06, 3.832301e-06, 4.758753e-06, 5.681814e-06,
  5.176787e-06, 6.008563e-06, 6.327712e-06, 5.777381e-06, 3.967294e-06, 
    3.633476e-06, 4.185232e-06, 5.367929e-06, 6.082792e-06, 6.382522e-06, 
    4.769607e-06, 5.304409e-06, 4.069464e-06, 4.865184e-06, 5.291305e-06,
  4.473478e-06, 6.859768e-06, 7.465684e-06, 6.454e-06, 4.722554e-06, 
    5.190868e-06, 5.00801e-06, 4.783662e-06, 6.650995e-06, 6.52512e-06, 
    6.186857e-06, 5.33395e-06, 4.859134e-06, 5.721139e-06, 7.5147e-06,
  6.588851e-06, 6.853807e-06, 6.764189e-06, 5.834858e-06, 6.618039e-06, 
    6.342902e-06, 5.292694e-06, 7.122605e-06, 7.212802e-06, 7.301318e-06, 
    5.712305e-06, 6.562758e-06, 7.098006e-06, 6.983899e-06, 8.429086e-06,
  7.479004e-06, 8.417393e-06, 7.86023e-06, 6.816856e-06, 7.069268e-06, 
    6.341662e-06, 7.253613e-06, 6.887473e-06, 9.203525e-06, 8.697189e-06, 
    7.736936e-06, 8.218269e-06, 7.546304e-06, 8.397104e-06, 4.480947e-06,
  8.471236e-06, 1.002346e-05, 9.056003e-06, 8.620807e-06, 8.860441e-06, 
    8.264063e-06, 7.389438e-06, 9.043852e-06, 1.200657e-05, 1.357947e-05, 
    1.017355e-05, 9.974136e-06, 9.203333e-06, 7.321857e-06, 6.18211e-06,
  1.006856e-05, 9.425135e-06, 1.147896e-05, 1.150308e-05, 1.096177e-05, 
    9.687684e-06, 1.014583e-05, 1.282543e-05, 1.615424e-05, 1.602389e-05, 
    1.369195e-05, 1.361925e-05, 1.223982e-05, 9.091927e-06, 7.964341e-06,
  1.247636e-05, 1.378424e-05, 1.091728e-05, 1.235398e-05, 1.490105e-05, 
    1.504833e-05, 1.411178e-05, 1.594436e-05, 2.074267e-05, 2.125011e-05, 
    1.979015e-05, 1.753052e-05, 1.502644e-05, 1.19538e-05, 9.978595e-06,
  1.416889e-05, 1.560247e-05, 1.676499e-05, 1.528701e-05, 1.860811e-05, 
    2.332119e-05, 2.219267e-05, 2.238747e-05, 2.408257e-05, 2.828729e-05, 
    2.66679e-05, 1.957439e-05, 1.75289e-05, 1.95003e-05, 1.482398e-05,
  1.612236e-05, 1.906337e-05, 1.977029e-05, 1.937778e-05, 1.97296e-05, 
    2.597101e-05, 3.222449e-05, 2.740179e-05, 2.73654e-05, 3.152897e-05, 
    2.760006e-05, 2.559867e-05, 2.176869e-05, 2.031771e-05, 1.742169e-05,
  7.772516e-06, 8.687576e-06, 5.939773e-06, 4.746375e-06, 6.956891e-06, 
    6.640647e-06, 4.861749e-06, 7.462516e-06, 1.650091e-05, 1.513701e-05, 
    9.305184e-06, 6.979818e-06, 1.038702e-05, 9.432266e-06, 8.252578e-06,
  7.509336e-06, 7.665768e-06, 5.088888e-06, 5.567448e-06, 5.84377e-06, 
    7.336986e-06, 9.282442e-06, 1.115761e-05, 1.360735e-05, 4.86513e-06, 
    7.458996e-06, 6.036709e-06, 5.760293e-06, 7.422626e-06, 7.869759e-06,
  5.832977e-06, 6.186542e-06, 4.159926e-06, 6.350042e-06, 8.51538e-06, 
    1.024981e-05, 1.229924e-05, 1.173723e-05, 7.447398e-06, 4.835714e-06, 
    5.213286e-06, 4.98069e-06, 3.376663e-06, 4.022031e-06, 7.639696e-06,
  5.539451e-06, 5.485317e-06, 6.054267e-06, 8.253459e-06, 1.161916e-05, 
    1.047496e-05, 6.52443e-06, 1.413428e-06, 3.848926e-07, 1.617134e-06, 
    2.384623e-07, 1.984966e-07, 2.173263e-07, 2.827935e-06, 3.68457e-06,
  5.443974e-06, 3.316846e-06, 2.491751e-06, 3.057671e-06, 3.998364e-06, 
    2.237522e-06, 3.190799e-06, 1.908486e-06, 1.126752e-06, 1.011109e-06, 
    9.411408e-07, 4.71312e-07, 4.096731e-07, 9.600702e-07, 3.009204e-06,
  4.627205e-06, 3.024996e-06, 3.301541e-06, 4.772182e-06, 2.885692e-06, 
    4.200583e-06, 1.730967e-06, 2.835707e-07, 1.29434e-06, 9.705058e-07, 
    1.022776e-06, 1.008855e-06, 7.911699e-07, 8.575713e-07, 1.272801e-06,
  2.878683e-06, 3.805748e-06, 3.147514e-06, 4.082562e-06, 2.86668e-06, 
    2.241592e-06, 2.962772e-06, 1.748966e-06, 1.067747e-06, 1.036964e-06, 
    9.607401e-07, 1.357988e-06, 6.878127e-07, 1.160723e-06, 7.200093e-07,
  3.729127e-06, 3.501377e-06, 2.801618e-06, 2.768797e-06, 3.05498e-06, 
    2.169398e-06, 1.558072e-06, 9.912421e-07, 1.212467e-06, 2.064994e-06, 
    2.863698e-06, 1.145858e-07, 7.990465e-07, 8.204589e-07, 8.066729e-07,
  3.648188e-06, 4.217561e-06, 3.571866e-06, 3.923708e-06, 2.696451e-06, 
    2.133053e-06, 1.319716e-06, 2.827811e-06, 1.34735e-06, 1.762263e-06, 
    1.626854e-06, 1.369371e-06, 2.111633e-06, 9.773449e-07, 1.78239e-06,
  2.98514e-06, 4.143197e-06, 3.440804e-06, 2.933498e-06, 2.306212e-06, 
    2.207972e-06, 1.873467e-06, 1.559048e-06, 1.543664e-06, 2.082962e-06, 
    3.043959e-06, 3.09767e-06, 1.909661e-06, 1.89202e-06, 9.090551e-07,
  1.208246e-05, 1.072573e-05, 7.194528e-06, 7.013947e-06, 7.929018e-06, 
    8.258065e-06, 8.008638e-06, 8.222113e-06, 9.139098e-06, 8.84144e-06, 
    6.742852e-06, 7.419618e-06, 6.317989e-06, 4.118966e-06, 3.203958e-06,
  1.172933e-05, 1.210087e-05, 1.05791e-05, 9.587392e-06, 9.350913e-06, 
    1.025587e-05, 6.980396e-06, 7.832112e-06, 9.390882e-06, 9.459135e-06, 
    7.312649e-06, 7.971364e-06, 6.086242e-06, 5.861016e-06, 5.665449e-06,
  1.266101e-05, 1.195225e-05, 1.071359e-05, 1.301549e-05, 1.058047e-05, 
    8.35146e-06, 8.337682e-06, 9.884752e-06, 1.235838e-05, 1.100199e-05, 
    9.289575e-06, 9.388589e-06, 8.974925e-06, 7.267581e-06, 8.037166e-06,
  5.290068e-06, 6.73785e-06, 5.739689e-06, 4.328256e-06, 5.07399e-06, 
    3.926263e-06, 5.723521e-06, 9.011093e-06, 1.000343e-05, 1.012741e-05, 
    1.255512e-05, 9.742203e-06, 1.02899e-05, 8.282083e-06, 1.045214e-05,
  3.864838e-06, 2.841246e-06, 3.246155e-06, 3.305544e-06, 3.509685e-06, 
    4.080626e-06, 5.050177e-06, 7.005103e-06, 9.678507e-06, 9.911203e-06, 
    1.032881e-05, 9.773726e-06, 9.577565e-06, 1.080155e-05, 1.155978e-05,
  2.864484e-06, 1.570738e-06, 2.899024e-06, 4.9772e-06, 3.67419e-06, 
    3.111706e-06, 4.738507e-06, 6.504872e-06, 8.781622e-06, 1.016597e-05, 
    1.050976e-05, 1.222703e-05, 1.103679e-05, 1.13227e-05, 9.586299e-06,
  1.731643e-06, 1.013216e-06, 3.540482e-06, 7.130825e-06, 3.798129e-06, 
    2.390695e-06, 3.386996e-06, 6.552955e-06, 1.11917e-05, 1.177707e-05, 
    1.175093e-05, 1.386338e-05, 1.181454e-05, 1.060109e-05, 1.145991e-05,
  1.792916e-06, 3.651291e-07, 2.222985e-06, 2.045207e-06, 2.440413e-06, 
    2.259684e-06, 3.031069e-06, 6.368944e-06, 9.535876e-06, 1.305789e-05, 
    1.1718e-05, 1.109754e-05, 1.438583e-05, 1.742724e-05, 1.316046e-05,
  1.702282e-06, 1.134976e-07, 2.911257e-07, 7.945919e-07, 2.267181e-06, 
    1.999947e-06, 2.680567e-06, 6.039005e-06, 8.891121e-06, 1.438138e-05, 
    1.170174e-05, 1.091675e-05, 1.677368e-05, 1.561897e-05, 1.665672e-05,
  2.452434e-07, 2.355795e-08, 8.263952e-08, 6.539933e-07, 1.338238e-06, 
    1.213056e-06, 3.300044e-06, 6.632991e-06, 9.865512e-06, 1.291275e-05, 
    1.302336e-05, 1.469301e-05, 1.471145e-05, 1.622623e-05, 1.673099e-05,
  1.05846e-05, 1.001245e-05, 1.051887e-05, 9.03238e-06, 8.921752e-06, 
    8.538897e-06, 7.210887e-06, 6.830708e-06, 9.163189e-06, 8.893891e-06, 
    7.478697e-06, 8.343787e-06, 7.180775e-06, 5.756132e-06, 6.712966e-06,
  1.130836e-05, 1.002362e-05, 8.812904e-06, 7.983978e-06, 8.591169e-06, 
    7.697824e-06, 7.30442e-06, 9.48255e-06, 9.642515e-06, 1.081943e-05, 
    9.254373e-06, 1.08989e-05, 1.037549e-05, 8.693518e-06, 7.161957e-06,
  1.37396e-05, 1.163056e-05, 1.169522e-05, 8.292347e-06, 1.009051e-05, 
    8.813107e-06, 8.733946e-06, 9.418898e-06, 1.080039e-05, 1.122247e-05, 
    1.082354e-05, 1.008189e-05, 1.071113e-05, 1.067607e-05, 9.223227e-06,
  1.51772e-05, 1.307071e-05, 1.287543e-05, 1.017122e-05, 9.668114e-06, 
    1.171944e-05, 1.071055e-05, 1.140523e-05, 1.311866e-05, 1.2962e-05, 
    1.292904e-05, 1.182911e-05, 1.061802e-05, 1.110545e-05, 1.270991e-05,
  1.196883e-05, 1.154424e-05, 1.499532e-05, 1.32897e-05, 1.510255e-05, 
    1.349308e-05, 1.381254e-05, 1.508708e-05, 1.625188e-05, 1.705153e-05, 
    1.49906e-05, 1.357912e-05, 1.211605e-05, 1.264146e-05, 1.202226e-05,
  1.358841e-05, 1.55213e-05, 1.627055e-05, 1.677854e-05, 1.731956e-05, 
    1.535795e-05, 1.403149e-05, 1.54112e-05, 1.808422e-05, 1.822132e-05, 
    1.73892e-05, 1.380585e-05, 1.454967e-05, 1.308026e-05, 1.228879e-05,
  1.41272e-05, 1.827228e-05, 1.854761e-05, 1.749264e-05, 1.906803e-05, 
    1.776568e-05, 1.657912e-05, 1.760154e-05, 1.655292e-05, 1.642332e-05, 
    1.451741e-05, 1.48231e-05, 1.487612e-05, 1.23073e-05, 1.014141e-05,
  1.782957e-05, 1.93246e-05, 2.131493e-05, 2.082091e-05, 2.155214e-05, 
    2.010404e-05, 1.78897e-05, 1.735004e-05, 1.490441e-05, 1.615122e-05, 
    1.614641e-05, 1.40456e-05, 1.178139e-05, 1.309477e-05, 1.378672e-05,
  2.178575e-05, 2.132614e-05, 2.298241e-05, 2.1908e-05, 1.954485e-05, 
    2.324063e-05, 1.826846e-05, 1.402513e-05, 2.154362e-05, 1.746807e-05, 
    1.966896e-05, 1.738591e-05, 1.581178e-05, 1.429236e-05, 1.363697e-05,
  2.273118e-05, 2.236423e-05, 2.200939e-05, 2.063167e-05, 2.288852e-05, 
    2.091385e-05, 1.768256e-05, 1.975953e-05, 1.830394e-05, 1.942068e-05, 
    1.81233e-05, 1.815227e-05, 1.644436e-05, 1.590272e-05, 1.747684e-05,
  2.481589e-06, 4.529695e-06, 5.542661e-06, 6.588683e-06, 6.295156e-06, 
    6.774302e-06, 5.379039e-06, 6.720868e-06, 7.129569e-06, 7.051123e-06, 
    4.412932e-06, 5.617161e-06, 2.523469e-06, 3.651623e-06, 3.303928e-06,
  1.056119e-05, 1.55333e-05, 1.673732e-05, 1.886511e-05, 1.737123e-05, 
    1.294789e-05, 1.286141e-05, 9.366408e-06, 7.717647e-06, 9.610775e-06, 
    7.933269e-06, 5.542158e-06, 3.738289e-06, 3.806032e-06, 3.621205e-06,
  1.547881e-05, 1.462503e-05, 1.597731e-05, 1.613819e-05, 1.439179e-05, 
    1.301728e-05, 1.082592e-05, 9.680026e-06, 7.932978e-06, 8.215852e-06, 
    6.827964e-06, 5.381698e-06, 5.052792e-06, 5.204333e-06, 4.929301e-06,
  8.206511e-06, 7.628689e-06, 4.784596e-06, 5.039074e-06, 5.344877e-06, 
    4.85434e-06, 3.916921e-06, 4.977306e-06, 5.203137e-06, 5.647761e-06, 
    6.615999e-06, 6.141803e-06, 6.756535e-06, 7.006031e-06, 7.453849e-06,
  5.513173e-06, 5.910409e-06, 4.89712e-06, 3.671061e-06, 3.167279e-06, 
    1.863163e-06, 1.613012e-06, 2.883263e-06, 4.720719e-06, 5.773496e-06, 
    6.798536e-06, 6.620596e-06, 5.969109e-06, 8.637631e-06, 6.798482e-06,
  6.780756e-06, 5.085855e-06, 3.396452e-06, 3.47238e-06, 3.012778e-06, 
    3.065737e-06, 3.593664e-06, 5.517453e-06, 6.874036e-06, 6.862736e-06, 
    6.377206e-06, 7.218204e-06, 8.379962e-06, 8.346433e-06, 8.28659e-06,
  6.346617e-06, 5.979955e-06, 2.445934e-06, 1.883282e-06, 4.11423e-06, 
    4.132125e-06, 5.938961e-06, 5.907982e-06, 6.930921e-06, 6.831144e-06, 
    8.392345e-06, 8.003562e-06, 9.898124e-06, 8.733588e-06, 7.642277e-06,
  6.853201e-06, 5.010603e-06, 2.513257e-06, 4.093199e-06, 4.865675e-06, 
    5.5173e-06, 6.496918e-06, 7.711805e-06, 9.523007e-06, 8.98798e-06, 
    8.94414e-06, 8.951341e-06, 9.178411e-06, 8.729149e-06, 7.783651e-06,
  5.850245e-06, 4.106508e-06, 4.541724e-06, 4.786869e-06, 6.099678e-06, 
    7.131757e-06, 7.699119e-06, 7.575613e-06, 8.823926e-06, 8.876294e-06, 
    1.035853e-05, 9.9525e-06, 8.915048e-06, 9.635537e-06, 7.454872e-06,
  4.375741e-06, 5.092498e-06, 4.89481e-06, 6.044556e-06, 6.462351e-06, 
    8.767182e-06, 1.023421e-05, 9.802886e-06, 8.431848e-06, 9.033694e-06, 
    9.498163e-06, 1.06412e-05, 9.598053e-06, 7.796371e-06, 8.816195e-06,
  9.773928e-08, 3.956657e-08, 3.046878e-08, 6.167498e-08, 9.687745e-08, 
    1.592901e-07, 2.224335e-07, 5.860946e-07, 6.661579e-07, 8.309307e-07, 
    9.814657e-07, 1.012687e-06, 1.171205e-06, 1.494387e-06, 2.113174e-06,
  3.117425e-06, 5.396183e-06, 3.358198e-06, 2.048489e-06, 1.693805e-06, 
    7.159333e-07, 8.13593e-07, 1.536389e-06, 2.116279e-06, 2.520005e-06, 
    1.351715e-06, 1.847111e-06, 3.840071e-06, 3.651109e-06, 2.606177e-06,
  1.251327e-05, 1.493999e-05, 1.324062e-05, 8.242176e-06, 5.226144e-06, 
    3.300172e-06, 2.251707e-06, 4.784121e-06, 6.015767e-06, 3.877677e-06, 
    3.83121e-06, 5.356213e-06, 6.895209e-06, 7.704765e-06, 6.70475e-06,
  1.516108e-05, 1.261087e-05, 1.160513e-05, 1.241228e-05, 9.175512e-06, 
    5.506725e-06, 4.579479e-06, 6.869651e-06, 8.677358e-06, 9.304495e-06, 
    9.065586e-06, 9.78728e-06, 9.038325e-06, 7.035326e-06, 5.471212e-06,
  1.158422e-05, 1.056659e-05, 1.26127e-05, 1.289579e-05, 8.140935e-06, 
    5.3848e-06, 4.746057e-06, 9.238957e-06, 1.05257e-05, 9.425454e-06, 
    1.00986e-05, 9.498691e-06, 6.561635e-06, 4.881177e-06, 4.182009e-06,
  9.270168e-06, 1.05068e-05, 9.954887e-06, 1.263898e-05, 1.000179e-05, 
    5.434501e-06, 7.246504e-06, 1.374886e-05, 1.540005e-05, 1.257443e-05, 
    1.097776e-05, 6.992176e-06, 4.995087e-06, 4.698802e-06, 4.870395e-06,
  3.590573e-06, 5.624874e-06, 7.296256e-06, 1.435174e-05, 1.429573e-05, 
    9.274461e-06, 1.28776e-05, 1.779431e-05, 1.73752e-05, 1.308925e-05, 
    8.866671e-06, 6.50635e-06, 4.772196e-06, 5.703544e-06, 7.369415e-06,
  3.751871e-06, 4.995965e-06, 7.337129e-06, 1.233653e-05, 1.448349e-05, 
    1.314859e-05, 1.846774e-05, 2.032662e-05, 1.598893e-05, 1.108544e-05, 
    8.120435e-06, 5.153075e-06, 6.16156e-06, 7.046934e-06, 8.047137e-06,
  3.836841e-06, 5.7911e-06, 7.909486e-06, 1.244793e-05, 1.582705e-05, 
    1.941834e-05, 2.132137e-05, 1.855482e-05, 1.324316e-05, 1.079447e-05, 
    8.803901e-06, 6.94654e-06, 7.696973e-06, 7.543157e-06, 6.217695e-06,
  8.125679e-06, 8.301984e-06, 7.391896e-06, 1.347105e-05, 1.657644e-05, 
    2.209417e-05, 2.016849e-05, 1.413155e-05, 1.027725e-05, 9.971671e-06, 
    8.294101e-06, 5.981255e-06, 6.18141e-06, 8.77421e-06, 8.192626e-06,
  8.882391e-06, 1.124004e-05, 2.415733e-05, 4.431911e-05, 7.094626e-05, 
    9.340319e-05, 8.798762e-05, 7.005101e-05, 5.580085e-05, 4.379443e-05, 
    2.966439e-05, 1.760951e-05, 1.01466e-05, 4.619978e-06, 3.69102e-06,
  5.654817e-07, 1.323653e-06, 3.944181e-06, 9.384509e-06, 1.527023e-05, 
    2.12771e-05, 3.056927e-05, 2.540163e-05, 3.020919e-05, 2.497549e-05, 
    1.415766e-05, 1.019628e-05, 7.573209e-06, 5.938896e-06, 6.48578e-06,
  6.003627e-07, 1.006103e-07, 1.717862e-07, 2.235052e-07, 2.803459e-07, 
    4.023098e-07, 1.416595e-06, 2.086192e-06, 3.257172e-06, 1.95541e-06, 
    4.543369e-06, 2.634205e-06, 3.48723e-06, 2.461943e-06, 2.560682e-06,
  6.124171e-07, 8.139201e-08, 4.894085e-08, 2.624097e-08, 5.870081e-08, 
    2.627303e-08, 7.515842e-08, 7.783706e-08, 3.116342e-07, 1.528428e-06, 
    2.078992e-06, 1.557859e-06, 1.379491e-06, 1.305448e-06, 1.110946e-06,
  6.000387e-07, 9.121347e-08, 1.386327e-07, 2.898708e-07, 4.182443e-07, 
    3.884006e-07, 1.770826e-06, 1.447529e-06, 1.639248e-06, 1.04872e-06, 
    1.291541e-06, 4.924476e-07, 1.212183e-06, 4.31042e-07, 5.146594e-07,
  3.523349e-06, 1.054111e-06, 1.051169e-06, 1.234243e-06, 1.067929e-06, 
    1.209548e-06, 2.602865e-06, 4.747724e-06, 3.817265e-06, 1.930123e-06, 
    5.91898e-07, 9.228882e-07, 4.821414e-07, 2.331473e-06, 3.928644e-06,
  1.134957e-05, 5.367724e-06, 3.420837e-06, 3.180385e-06, 2.202465e-06, 
    3.112467e-06, 5.829144e-06, 4.353015e-06, 2.36661e-06, 1.260125e-06, 
    7.518012e-07, 1.662538e-06, 3.248268e-06, 5.156218e-06, 2.986742e-06,
  2.051596e-05, 1.289857e-05, 1.21738e-05, 6.68111e-06, 2.778469e-06, 
    4.116315e-06, 8.016906e-06, 2.873301e-06, 1.137754e-06, 1.367945e-06, 
    1.073926e-06, 5.77105e-06, 3.998757e-06, 1.962632e-06, 1.575801e-06,
  2.697567e-05, 1.647882e-05, 1.618769e-05, 1.099127e-05, 3.780699e-06, 
    5.93154e-06, 4.028521e-06, 8.877172e-07, 6.637468e-07, 2.532722e-06, 
    6.243307e-06, 2.779597e-06, 2.057356e-06, 1.775044e-06, 1.780357e-06,
  3.063281e-05, 3.056235e-05, 2.483739e-05, 1.879096e-05, 7.491909e-06, 
    5.170513e-06, 1.522617e-06, 3.652461e-07, 2.651482e-06, 5.857589e-06, 
    4.235885e-06, 2.000759e-06, 1.508379e-06, 1.618713e-06, 1.320355e-06,
  0.0004790044, 0.0004242506, 0.0003569519, 0.0003115751, 0.000305537, 
    0.0002520712, 9.3653e-05, 2.116528e-05, 1.595635e-05, 1.785308e-05, 
    2.627891e-05, 3.798168e-05, 4.263541e-05, 2.538787e-05, 8.783915e-06,
  0.0004740677, 0.0004314163, 0.0003915418, 0.000357003, 0.0003462248, 
    0.0002498523, 0.0001032404, 2.085523e-05, 1.293623e-05, 1.858062e-05, 
    3.070986e-05, 5.029456e-05, 6.093377e-05, 4.353696e-05, 2.580794e-05,
  0.0004479897, 0.0004060523, 0.0003602432, 0.0003344339, 0.0003020553, 
    0.0002140021, 7.359392e-05, 1.58657e-05, 8.016289e-06, 9.349905e-06, 
    1.77722e-05, 3.458756e-05, 6.020672e-05, 5.581427e-05, 3.660125e-05,
  0.0004098036, 0.0003622146, 0.000346247, 0.000320187, 0.0002809222, 
    0.0001840762, 6.605614e-05, 1.492507e-05, 3.540908e-06, 3.58199e-06, 
    5.615083e-06, 1.316568e-05, 2.187142e-05, 2.732183e-05, 2.537827e-05,
  0.0003961785, 0.0003747825, 0.0003600873, 0.0003190035, 0.000233903, 
    0.0001136306, 4.29287e-05, 9.066986e-06, 2.792241e-06, 9.306372e-07, 
    3.80662e-07, 1.933793e-07, 1.379274e-06, 2.586101e-06, 5.488624e-06,
  0.0003023232, 0.0003111436, 0.0002966643, 0.0002481628, 0.0001440996, 
    4.938721e-05, 1.267776e-05, 1.014022e-05, 3.544903e-06, 1.131281e-06, 
    2.734547e-07, 9.648035e-07, 4.671674e-07, 1.045735e-06, 2.68122e-06,
  0.0001373369, 0.0001562175, 0.0001373989, 0.0001009608, 4.88313e-05, 
    1.433548e-05, 3.421892e-06, 4.181499e-06, 4.190807e-06, 2.135125e-06, 
    2.313652e-06, 1.581252e-06, 1.224329e-06, 4.69965e-07, 1.728005e-06,
  5.409778e-05, 5.449022e-05, 3.457128e-05, 2.685022e-05, 2.058306e-05, 
    1.002414e-05, 2.42221e-06, 2.087112e-06, 3.620036e-06, 3.729678e-06, 
    3.147257e-06, 1.600399e-06, 7.589662e-07, 8.901674e-07, 1.283546e-06,
  2.250787e-05, 1.847403e-05, 1.103235e-05, 1.026069e-05, 1.264353e-05, 
    1.637193e-05, 3.052149e-06, 3.116903e-06, 3.356811e-06, 7.178795e-06, 
    2.956975e-06, 1.319448e-06, 1.561479e-06, 1.735617e-06, 1.968348e-06,
  1.857534e-05, 1.832642e-05, 5.716507e-06, 7.256618e-06, 1.090575e-05, 
    1.948514e-05, 1.745653e-06, 3.575558e-06, 3.025312e-06, 3.613113e-06, 
    2.430057e-06, 2.155002e-06, 1.439261e-06, 2.002012e-06, 2.072762e-06,
  1.373025e-05, 1.525708e-05, 2.062559e-05, 2.361758e-05, 2.239067e-05, 
    2.330579e-05, 1.702308e-05, 1.579028e-05, 1.519925e-05, 1.355058e-05, 
    8.272137e-06, 2.874482e-06, 1.992112e-06, 3.303445e-06, 2.782775e-06,
  1.898282e-05, 2.636615e-05, 3.322094e-05, 3.481746e-05, 3.340789e-05, 
    3.194228e-05, 2.169639e-05, 2.016656e-05, 1.536272e-05, 1.306785e-05, 
    8.944844e-06, 4.299151e-06, 2.049371e-06, 2.189006e-06, 1.877293e-06,
  3.618743e-05, 5.547695e-05, 6.949151e-05, 7.593934e-05, 6.991485e-05, 
    4.688765e-05, 2.997932e-05, 2.558949e-05, 1.787182e-05, 1.284779e-05, 
    1.165258e-05, 7.335856e-06, 4.092103e-06, 2.720446e-06, 2.461166e-06,
  7.431359e-05, 0.0001008169, 0.0001121454, 0.0001192476, 0.000108944, 
    6.555138e-05, 3.599365e-05, 3.093765e-05, 2.228319e-05, 1.376366e-05, 
    1.304235e-05, 6.47285e-06, 4.530079e-06, 3.61087e-06, 2.176003e-06,
  0.000125095, 0.0001530171, 0.0001545395, 0.0001616798, 0.0001529645, 
    9.010761e-05, 5.028173e-05, 4.40589e-05, 3.204735e-05, 1.767322e-05, 
    1.365657e-05, 9.11801e-06, 5.955079e-06, 3.815706e-06, 3.266755e-06,
  0.0001871053, 0.0002107622, 0.0001989711, 0.0001906424, 0.0001790652, 
    0.0001166577, 7.506517e-05, 6.110415e-05, 4.657106e-05, 2.386017e-05, 
    1.32652e-05, 1.278336e-05, 8.438431e-06, 3.216567e-06, 1.633388e-06,
  0.0002587326, 0.0002593172, 0.0002180742, 0.0001986868, 0.0001729715, 
    0.000123616, 8.750282e-05, 7.753055e-05, 6.31698e-05, 3.567032e-05, 
    2.469127e-05, 2.134185e-05, 1.255498e-05, 3.111936e-06, 1.867714e-06,
  0.0002749847, 0.0002534846, 0.0002028699, 0.0001583371, 0.0001329189, 
    0.0001035611, 8.572922e-05, 8.350298e-05, 7.537209e-05, 6.034782e-05, 
    4.709635e-05, 3.319895e-05, 2.120913e-05, 6.795623e-06, 2.612304e-06,
  0.0002687611, 0.0002134756, 0.0001570394, 0.0001317517, 0.0001080628, 
    7.366482e-05, 6.681949e-05, 7.491952e-05, 8.066981e-05, 9.066921e-05, 
    8.498927e-05, 5.548788e-05, 3.080711e-05, 1.205387e-05, 3.563583e-06,
  0.0002503279, 0.0002006347, 0.0001651948, 0.0001241287, 8.9243e-05, 
    5.315548e-05, 3.5952e-05, 4.031818e-05, 6.105417e-05, 0.0001000546, 
    0.0001184953, 9.409305e-05, 4.397503e-05, 1.969983e-05, 7.053766e-06,
  4.944051e-06, 4.311934e-06, 7.5836e-06, 4.740765e-06, 1.727275e-05, 
    5.625823e-05, 0.0001212244, 0.0001666832, 0.0002012112, 0.0002542034, 
    0.0002440158, 0.0002045046, 0.0001652854, 0.0001301111, 0.0001488284,
  7.648985e-06, 6.885528e-06, 5.694664e-06, 5.993513e-06, 1.291403e-05, 
    2.575549e-05, 9.831336e-05, 0.0001578662, 0.0002017026, 0.0002231456, 
    0.0002174027, 0.0001680891, 0.0001418251, 0.0001349953, 0.000157315,
  6.250681e-06, 1.015732e-05, 6.223614e-06, 5.561853e-06, 8.065674e-06, 
    1.384819e-05, 4.642808e-05, 0.0001207395, 0.0001794383, 0.000202666, 
    0.0001877783, 0.0001602361, 0.0001286665, 0.0001106728, 0.0001181696,
  9.978506e-06, 1.185943e-05, 7.381604e-06, 5.759866e-06, 4.563132e-06, 
    7.050357e-06, 2.003918e-05, 6.354347e-05, 0.0001240071, 0.0001625921, 
    0.0001522562, 0.0001171851, 8.888721e-05, 7.129774e-05, 9.13308e-05,
  1.028889e-05, 1.282913e-05, 1.156806e-05, 8.795446e-06, 4.588621e-06, 
    3.432259e-06, 6.512515e-06, 3.487709e-05, 7.710644e-05, 0.0001023256, 
    0.0001205553, 9.385641e-05, 6.369854e-05, 5.456058e-05, 6.262761e-05,
  1.235934e-05, 1.367773e-05, 1.19309e-05, 8.86664e-06, 6.01671e-06, 
    3.579476e-06, 5.111398e-06, 1.294688e-05, 4.553086e-05, 6.194454e-05, 
    7.876192e-05, 7.679731e-05, 5.212986e-05, 5.725621e-05, 6.14653e-05,
  1.464721e-05, 1.127357e-05, 8.814137e-06, 3.587758e-06, 5.312717e-06, 
    3.981096e-06, 3.968573e-06, 4.817648e-06, 1.65546e-05, 3.501398e-05, 
    6.095009e-05, 6.274932e-05, 5.15309e-05, 7.78096e-05, 8.156512e-05,
  9.575268e-06, 1.008475e-05, 8.347804e-06, 5.652462e-06, 3.544956e-06, 
    3.268906e-06, 5.267444e-06, 6.03962e-06, 8.891567e-06, 2.54082e-05, 
    4.231371e-05, 4.047458e-05, 4.186262e-05, 7.673209e-05, 0.0001035004,
  1.177312e-05, 9.680345e-06, 8.01997e-06, 5.330224e-06, 3.4378e-06, 
    2.413479e-06, 6.577634e-06, 7.955864e-06, 1.18942e-05, 1.707195e-05, 
    3.688638e-05, 2.09853e-05, 2.148078e-05, 5.004789e-05, 9.80104e-05,
  1.224883e-05, 1.207009e-05, 7.783908e-06, 3.167674e-06, 1.244644e-06, 
    3.238673e-06, 5.602375e-06, 7.195279e-06, 1.213074e-05, 1.976208e-05, 
    3.500174e-05, 1.404926e-05, 8.267834e-06, 2.863568e-05, 6.979591e-05,
  0.0002044647, 0.0001955318, 0.0001338241, 4.175025e-05, 2.516365e-05, 
    3.436954e-05, 1.515691e-05, 1.410592e-05, 1.822108e-05, 8.791159e-06, 
    8.091302e-06, 8.778088e-06, 1.020776e-05, 1.0613e-05, 2.396058e-05,
  0.0002161528, 0.0002195045, 0.0001593587, 5.551151e-05, 2.875125e-05, 
    6.552472e-05, 5.358867e-05, 3.916704e-05, 3.427511e-05, 1.529001e-05, 
    5.443636e-06, 9.580137e-06, 7.680985e-06, 1.301081e-05, 2.323194e-05,
  0.0002055767, 0.0002221286, 0.0001776956, 6.415698e-05, 3.971671e-05, 
    9.087389e-05, 0.0001095912, 9.0067e-05, 5.921357e-05, 2.5355e-05, 
    9.69691e-06, 6.4251e-06, 4.100598e-06, 1.173035e-05, 2.085997e-05,
  0.0001594179, 0.00017919, 0.0001727465, 8.035579e-05, 4.155664e-05, 
    9.958809e-05, 0.0001372555, 0.0001322657, 9.763863e-05, 4.523884e-05, 
    1.018866e-05, 6.273274e-06, 4.389899e-06, 8.519175e-06, 1.947218e-05,
  0.0001083309, 0.0001334649, 0.0001428394, 8.04359e-05, 3.868182e-05, 
    0.0001023823, 0.0001266445, 0.0001435836, 0.0001192094, 7.421494e-05, 
    1.875483e-05, 6.888047e-06, 6.364108e-06, 8.044857e-06, 1.499346e-05,
  7.894708e-05, 0.0001092057, 0.0001254841, 7.877405e-05, 3.279753e-05, 
    7.546616e-05, 0.0001028938, 0.0001182431, 0.0001166263, 8.372439e-05, 
    2.996956e-05, 9.471607e-06, 1.011649e-05, 1.259207e-05, 1.593455e-05,
  6.558072e-05, 8.713079e-05, 0.0001033388, 6.98728e-05, 2.553532e-05, 
    5.380115e-05, 7.703959e-05, 8.237599e-05, 0.00010448, 8.001728e-05, 
    4.020216e-05, 1.417692e-05, 1.722889e-05, 2.542555e-05, 2.766985e-05,
  5.651197e-05, 6.904424e-05, 9.4684e-05, 6.285595e-05, 2.602751e-05, 
    5.575594e-05, 6.818416e-05, 6.554454e-05, 8.565461e-05, 8.287025e-05, 
    5.244242e-05, 2.420419e-05, 2.678852e-05, 4.331027e-05, 4.484604e-05,
  4.550747e-05, 5.5457e-05, 7.404948e-05, 6.322155e-05, 2.893436e-05, 
    6.612213e-05, 7.659542e-05, 6.024258e-05, 7.396017e-05, 8.393812e-05, 
    7.502751e-05, 5.740234e-05, 5.661918e-05, 6.931966e-05, 6.113794e-05,
  3.618322e-05, 4.890534e-05, 6.185214e-05, 6.390228e-05, 3.697076e-05, 
    7.981403e-05, 7.476028e-05, 5.516282e-05, 5.700475e-05, 7.477175e-05, 
    0.0001055129, 9.816813e-05, 9.204142e-05, 0.0001016994, 0.0001049693,
  9.25497e-05, 2.260013e-05, 6.722118e-06, 1.632968e-06, 5.215052e-06, 
    2.427459e-06, 7.754543e-06, 3.935475e-06, 1.798304e-05, 1.162373e-05, 
    2.121745e-05, 1.942391e-05, 2.907832e-05, 2.045517e-05, 1.836807e-05,
  0.0001803782, 5.447192e-05, 1.508728e-05, 1.105402e-05, 4.705077e-06, 
    5.807172e-06, 9.341212e-06, 1.960019e-05, 2.909332e-05, 1.756862e-05, 
    3.081824e-05, 2.35838e-05, 4.218066e-05, 3.715305e-05, 2.0708e-05,
  0.0002329874, 8.080695e-05, 2.03783e-05, 1.052748e-05, 8.541263e-06, 
    1.200519e-05, 1.830473e-05, 1.599316e-05, 3.299551e-05, 2.124836e-05, 
    3.315169e-05, 1.947452e-05, 2.789564e-05, 3.886161e-05, 1.692188e-05,
  0.0002526965, 9.82985e-05, 2.935294e-05, 1.000793e-05, 9.824116e-06, 
    8.816948e-06, 1.645564e-05, 8.652748e-06, 1.122203e-05, 1.389673e-05, 
    2.090277e-05, 2.820095e-05, 2.20895e-05, 2.692343e-05, 1.76848e-05,
  0.0002623712, 0.0001147814, 4.654893e-05, 8.00031e-06, 1.054558e-05, 
    9.709638e-06, 1.146396e-05, 1.089409e-05, 6.875446e-06, 1.111611e-05, 
    2.000755e-05, 2.015916e-05, 1.408205e-05, 1.865571e-05, 2.761856e-05,
  0.0002540643, 0.0001194717, 3.619729e-05, 8.950274e-06, 1.440858e-05, 
    8.036281e-06, 5.775707e-06, 8.687944e-06, 5.244491e-06, 1.607549e-05, 
    1.516342e-05, 1.127273e-05, 1.48785e-05, 1.452835e-05, 1.962144e-05,
  0.0002252281, 0.0001318636, 6.20109e-05, 1.047654e-05, 1.17961e-05, 
    1.015149e-05, 6.001414e-06, 5.76108e-06, 2.674917e-06, 6.882536e-06, 
    1.396896e-05, 1.771333e-05, 1.177896e-05, 1.526225e-05, 1.976259e-05,
  0.0001892522, 0.0001215045, 5.719241e-05, 6.700439e-06, 1.441456e-05, 
    1.118096e-05, 6.712681e-06, 7.590553e-06, 3.105885e-06, 1.118636e-05, 
    1.448269e-05, 7.886681e-06, 1.159033e-05, 1.384519e-05, 2.953692e-05,
  0.0001509941, 0.0001069792, 5.848899e-05, 4.236437e-06, 1.785331e-05, 
    9.699649e-06, 6.935302e-06, 8.667816e-06, 3.77784e-06, 5.977231e-06, 
    1.174149e-05, 1.094996e-05, 1.232212e-05, 2.745594e-05, 3.301121e-05,
  0.0001289836, 9.655391e-05, 5.030148e-05, 6.751402e-06, 2.527237e-05, 
    1.402447e-05, 8.839384e-06, 1.118337e-05, 5.854036e-06, 1.462487e-06, 
    1.539057e-05, 1.333766e-05, 1.650953e-05, 3.761182e-05, 2.229091e-05,
  2.592993e-05, 3.422895e-06, 1.263798e-06, 1.35639e-06, 2.16027e-06, 
    2.257755e-06, 2.464422e-06, 2.772746e-06, 3.755611e-06, 5.266361e-06, 
    8.144591e-06, 2.105049e-05, 0.00011383, 0.0001364255, 9.589405e-05,
  2.436155e-05, 1.405943e-06, 4.830391e-07, 1.071012e-06, 1.414873e-06, 
    1.525817e-06, 1.692165e-06, 2.328796e-06, 3.260578e-06, 4.436943e-06, 
    5.637421e-06, 1.127573e-05, 4.720649e-05, 8.56198e-05, 9.911275e-05,
  1.44032e-05, 1.123717e-06, 2.954041e-07, 9.695801e-07, 1.062228e-06, 
    1.454956e-06, 1.867196e-06, 1.864137e-06, 2.471523e-06, 4.764225e-06, 
    3.451053e-06, 5.570382e-06, 3.132221e-05, 7.389623e-05, 6.820872e-05,
  1.950247e-05, 1.601169e-06, 3.095428e-07, 1.522083e-06, 1.753735e-06, 
    8.752269e-07, 1.27683e-06, 2.3202e-06, 2.829792e-06, 3.344332e-06, 
    3.164004e-06, 3.05986e-06, 1.527905e-05, 5.577635e-05, 6.783023e-05,
  2.240422e-05, 2.339175e-06, 4.105399e-07, 1.641271e-06, 1.833858e-06, 
    7.517437e-07, 9.369945e-07, 1.826303e-06, 2.444737e-06, 2.949734e-06, 
    3.406108e-06, 2.781936e-06, 6.187294e-06, 3.609593e-05, 5.945072e-05,
  1.905725e-05, 1.72521e-06, 1.801845e-07, 1.010855e-06, 1.395141e-06, 
    1.535288e-06, 6.990567e-07, 9.5106e-07, 2.041056e-06, 3.119219e-06, 
    2.597317e-06, 1.904293e-06, 1.080827e-06, 1.644181e-05, 4.778397e-05,
  1.824729e-05, 1.596668e-06, 1.552277e-06, 9.414464e-07, 1.644865e-06, 
    1.340443e-06, 1.53137e-06, 1.668462e-06, 2.554946e-06, 3.588608e-06, 
    3.965246e-06, 1.946254e-06, 1.2549e-06, 3.785805e-06, 2.830293e-05,
  1.4397e-05, 8.438062e-07, 3.297667e-07, 7.437822e-07, 1.135207e-06, 
    1.01458e-06, 1.161527e-06, 1.442324e-06, 2.12676e-06, 2.410078e-06, 
    2.675595e-06, 1.557983e-06, 5.467976e-07, 3.396966e-07, 7.749348e-06,
  1.319448e-05, 1.089808e-06, 7.315373e-07, 1.060943e-06, 9.321681e-07, 
    1.359202e-06, 5.161532e-07, 8.74605e-07, 1.443741e-06, 2.906113e-06, 
    2.143816e-06, 2.191956e-06, 1.524444e-06, 2.902557e-07, 6.742951e-07,
  1.387666e-05, 1.182497e-06, 3.540665e-07, 8.578332e-07, 1.49325e-06, 
    2.359522e-06, 1.336471e-06, 1.105263e-06, 1.061997e-06, 1.581708e-06, 
    2.303632e-06, 3.309653e-06, 3.683005e-07, 7.303642e-08, 5.555342e-08,
  3.473019e-05, 3.143059e-05, 2.733448e-05, 5.046314e-05, 7.810252e-05, 
    6.989958e-05, 9.345816e-05, 0.0001160665, 0.0001285138, 0.0001610777, 
    0.0001393942, 0.0001638807, 7.575579e-05, 5.915999e-05, 5.580991e-05,
  4.542769e-05, 4.216053e-05, 4.732791e-05, 5.436933e-05, 8.33802e-05, 
    9.63769e-05, 0.0001102737, 0.0001301346, 0.0001306619, 0.0001486603, 
    0.0001830992, 0.0002104809, 9.850466e-05, 6.237679e-05, 6.525189e-05,
  6.815531e-05, 3.820716e-05, 7.664823e-05, 7.832211e-05, 7.229466e-05, 
    9.351707e-05, 0.0001086053, 0.0001435535, 0.0001482051, 0.0001297264, 
    0.0001795085, 0.0001838297, 0.0001585161, 7.096671e-05, 6.96187e-05,
  3.677085e-05, 2.386528e-05, 5.756974e-05, 7.604602e-05, 8.891578e-05, 
    0.0001079396, 0.0001414253, 0.0001348271, 0.0001552292, 0.0001407503, 
    0.0002073691, 0.0002037259, 0.0001822422, 0.0001297129, 7.939022e-05,
  3.138531e-05, 3.470487e-05, 9.297502e-05, 6.470691e-05, 8.549063e-05, 
    9.40205e-05, 0.0001076748, 0.0001183862, 0.0001295068, 0.0001631716, 
    0.0001914654, 0.0001960812, 0.0001587549, 0.0001002298, 7.837454e-05,
  3.195474e-05, 4.27812e-05, 4.234552e-05, 6.9934e-05, 7.414098e-05, 
    7.462061e-05, 0.0001043007, 0.0001192688, 9.281908e-05, 0.0001154756, 
    0.0001421514, 0.0001828874, 0.0001515874, 0.0001171236, 4.461326e-05,
  3.757018e-05, 4.241068e-05, 5.073006e-05, 7.049791e-05, 7.347136e-05, 
    8.42657e-05, 0.0001009223, 9.436246e-05, 9.835356e-05, 0.0001172817, 
    0.0001386899, 0.0002012179, 0.0001302028, 0.0001367652, 0.0001013549,
  3.788326e-05, 4.348532e-05, 5.211236e-05, 5.977413e-05, 5.939473e-05, 
    7.923054e-05, 9.40555e-05, 9.457746e-05, 8.651869e-05, 0.000123885, 
    0.0001397419, 0.0001873991, 0.0001447963, 0.0001091821, 7.009738e-05,
  2.660726e-05, 4.400946e-05, 5.747579e-05, 6.188308e-05, 5.458115e-05, 
    7.025745e-05, 8.135979e-05, 9.565438e-05, 9.04192e-05, 0.0001114487, 
    0.0001245657, 0.0001413153, 0.0001693958, 0.000119792, 8.728314e-05,
  1.71942e-05, 4.148688e-05, 5.416453e-05, 6.633954e-05, 6.535287e-05, 
    7.016878e-05, 7.630567e-05, 9.328619e-05, 8.687688e-05, 9.838689e-05, 
    0.000112465, 0.0001258462, 0.000157128, 0.0001154916, 9.509872e-05,
  1.431963e-05, 1.534567e-05, 1.416143e-05, 2.236249e-05, 2.943701e-05, 
    3.313318e-05, 3.579652e-05, 4.082571e-05, 4.881911e-05, 4.537959e-05, 
    3.340174e-05, 2.220531e-05, 2.220816e-05, 2.326846e-05, 2.147485e-05,
  1.488573e-05, 1.739162e-05, 1.966489e-05, 2.565659e-05, 3.59639e-05, 
    3.839418e-05, 4.748398e-05, 5.492808e-05, 6.270426e-05, 5.493598e-05, 
    3.739353e-05, 2.69182e-05, 2.83074e-05, 2.824878e-05, 2.359255e-05,
  1.799952e-05, 1.900445e-05, 2.265529e-05, 2.989314e-05, 4.849916e-05, 
    5.007149e-05, 8.248998e-05, 8.586707e-05, 9.638533e-05, 8.755211e-05, 
    5.084638e-05, 3.205449e-05, 3.88668e-05, 3.875499e-05, 3.191025e-05,
  1.945755e-05, 2.11011e-05, 2.811289e-05, 5.258351e-05, 6.897283e-05, 
    6.667792e-05, 8.858931e-05, 0.0001026389, 0.0001165574, 0.0001128513, 
    4.857633e-05, 3.516457e-05, 4.337912e-05, 5.025425e-05, 4.318414e-05,
  2.262826e-05, 2.485193e-05, 3.917957e-05, 7.32081e-05, 7.001522e-05, 
    8.060645e-05, 6.03201e-05, 0.0001012713, 7.7132e-05, 0.0001208544, 
    6.756544e-05, 4.896466e-05, 4.476722e-05, 5.361753e-05, 5.521296e-05,
  2.180917e-05, 2.869245e-05, 5.735394e-05, 7.553821e-05, 8.178966e-05, 
    7.696416e-05, 8.607764e-05, 0.0001098191, 0.0001167, 0.0001382363, 
    9.984577e-05, 6.688828e-05, 6.882045e-05, 6.599539e-05, 6.395709e-05,
  3.026129e-05, 3.231154e-05, 4.514949e-05, 7.649071e-05, 6.260331e-05, 
    9.515986e-05, 6.708243e-05, 7.792771e-05, 0.0001284895, 0.000105203, 
    0.0001360439, 7.709629e-05, 8.333785e-05, 8.491496e-05, 7.840931e-05,
  3.310338e-05, 6.076662e-05, 7.324643e-05, 5.793148e-05, 4.646613e-05, 
    6.514908e-05, 9.940502e-05, 9.583337e-05, 8.147835e-05, 0.0001177035, 
    0.000130925, 8.799059e-05, 9.059412e-05, 8.25448e-05, 8.364855e-05,
  4.757785e-05, 4.500069e-05, 4.906674e-05, 5.156979e-05, 7.591013e-05, 
    0.0001274155, 8.415832e-05, 8.205276e-05, 0.0001062231, 9.939518e-05, 
    0.0001030803, 9.082126e-05, 9.820777e-05, 7.731467e-05, 5.85262e-05,
  5.336965e-05, 3.915914e-05, 3.016368e-05, 4.944447e-05, 5.2633e-05, 
    8.3568e-05, 7.716507e-05, 6.748924e-05, 9.834622e-05, 0.0001019874, 
    7.996339e-05, 9.393814e-05, 0.0001172454, 7.269061e-05, 8.436652e-05,
  7.322763e-06, 7.791499e-06, 6.060613e-06, 5.649307e-06, 5.823201e-06, 
    6.369419e-06, 4.69078e-06, 4.963848e-06, 7.698233e-06, 5.16661e-06, 
    5.458467e-06, 4.131408e-06, 4.216692e-06, 2.180219e-06, 1.941044e-06,
  8.684389e-06, 7.5717e-06, 6.830423e-06, 8.383509e-06, 8.59862e-06, 
    7.935912e-06, 7.901047e-06, 7.406355e-06, 8.35533e-06, 8.736914e-06, 
    8.134643e-06, 6.882075e-06, 4.599666e-06, 3.903442e-06, 3.228475e-06,
  1.216754e-05, 1.145398e-05, 1.118068e-05, 1.069635e-05, 1.18188e-05, 
    1.350464e-05, 1.027703e-05, 1.061037e-05, 1.423866e-05, 1.179607e-05, 
    1.127942e-05, 1.063851e-05, 7.679313e-06, 6.244451e-06, 4.106038e-06,
  1.553657e-05, 1.595214e-05, 1.53311e-05, 1.679125e-05, 1.737447e-05, 
    1.653773e-05, 1.58686e-05, 1.771986e-05, 1.777032e-05, 1.741992e-05, 
    1.42762e-05, 1.038453e-05, 9.116603e-06, 6.778293e-06, 4.983302e-06,
  2.065868e-05, 2.027349e-05, 2.005375e-05, 2.335292e-05, 2.311776e-05, 
    2.160043e-05, 2.408199e-05, 2.427186e-05, 2.608943e-05, 2.57392e-05, 
    1.962297e-05, 1.563334e-05, 1.050807e-05, 7.035965e-06, 3.80994e-06,
  3.009697e-05, 2.691624e-05, 2.583337e-05, 2.867864e-05, 3.281609e-05, 
    3.030923e-05, 3.097671e-05, 3.451944e-05, 3.574356e-05, 3.37824e-05, 
    2.579088e-05, 1.559949e-05, 1.169036e-05, 7.180986e-06, 6.09364e-06,
  4.111726e-05, 3.466814e-05, 3.252614e-05, 3.749979e-05, 3.994766e-05, 
    3.927243e-05, 3.991834e-05, 4.31286e-05, 4.523927e-05, 3.440719e-05, 
    2.488082e-05, 1.449924e-05, 1.134976e-05, 8.068781e-06, 7.270361e-06,
  4.740939e-05, 3.830362e-05, 3.582612e-05, 3.969517e-05, 4.919555e-05, 
    4.560508e-05, 4.873429e-05, 4.785359e-05, 4.591772e-05, 3.645794e-05, 
    2.441242e-05, 1.552143e-05, 1.083733e-05, 9.214529e-06, 7.071005e-06,
  5.015381e-05, 3.907152e-05, 4.214697e-05, 4.232608e-05, 4.757012e-05, 
    5.200561e-05, 5.041571e-05, 6.23134e-05, 4.22043e-05, 4.123408e-05, 
    3.110793e-05, 1.910842e-05, 1.316805e-05, 1.079523e-05, 9.829682e-06,
  5.509864e-05, 4.513923e-05, 4.543347e-05, 4.398721e-05, 4.990538e-05, 
    6.026552e-05, 7.080691e-05, 6.092063e-05, 6.788491e-05, 5.045222e-05, 
    4.844147e-05, 3.078059e-05, 2.06246e-05, 2.117753e-05, 1.36934e-05,
  8.497707e-07, 5.211887e-07, 1.128265e-06, 1.378402e-06, 1.654908e-06, 
    2.387264e-06, 1.963188e-06, 2.86184e-06, 2.970476e-06, 5.266304e-06, 
    1.21307e-05, 2.008903e-05, 2.21959e-05, 3.289039e-05, 4.315161e-05,
  1.758594e-06, 2.217675e-06, 1.213528e-06, 1.6056e-06, 2.387158e-06, 
    1.060126e-06, 1.704637e-06, 2.646829e-06, 3.151508e-06, 2.851604e-06, 
    9.564539e-06, 2.159392e-05, 2.905138e-05, 3.911313e-05, 4.989729e-05,
  1.349607e-06, 1.823006e-06, 1.535626e-06, 1.447267e-06, 1.844158e-06, 
    1.218799e-06, 1.512008e-06, 1.63244e-06, 1.74704e-06, 2.246105e-06, 
    5.854944e-06, 1.846396e-05, 3.420559e-05, 4.212205e-05, 5.156043e-05,
  1.518086e-06, 1.715796e-06, 1.534808e-06, 1.637278e-06, 1.993422e-06, 
    1.155081e-06, 1.18172e-06, 1.451263e-06, 2.035754e-06, 2.05995e-06, 
    4.726518e-06, 1.752916e-05, 3.185227e-05, 4.332606e-05, 5.31545e-05,
  1.756467e-06, 1.814397e-06, 1.464407e-06, 1.305805e-06, 1.785636e-06, 
    1.424556e-06, 1.154719e-06, 1.946161e-06, 1.313659e-06, 3.310867e-06, 
    7.949619e-06, 2.010995e-05, 3.643155e-05, 4.681814e-05, 5.877755e-05,
  2.083981e-06, 1.89642e-06, 1.71763e-06, 2.262181e-06, 1.948745e-06, 
    1.106383e-06, 9.086778e-07, 1.501003e-06, 1.940477e-06, 3.807341e-06, 
    7.258558e-06, 1.799089e-05, 3.370913e-05, 4.804849e-05, 5.168017e-05,
  2.592858e-06, 2.411429e-06, 1.687237e-06, 2.444258e-06, 1.686501e-06, 
    2.013026e-06, 1.72979e-06, 2.279397e-06, 3.771135e-06, 3.138864e-06, 
    6.617534e-06, 1.475374e-05, 2.907594e-05, 4.734502e-05, 4.819017e-05,
  3.480695e-06, 2.870547e-06, 2.6442e-06, 2.962336e-06, 3.865439e-06, 
    3.39815e-06, 3.130733e-06, 2.688294e-06, 2.181445e-06, 2.88555e-06, 
    7.592144e-06, 1.484878e-05, 2.60044e-05, 3.908648e-05, 4.263678e-05,
  4.274352e-06, 3.92121e-06, 4.268863e-06, 3.591971e-06, 3.973656e-06, 
    3.604843e-06, 3.103937e-06, 2.615938e-06, 2.617519e-06, 2.279401e-06, 
    6.230825e-06, 1.305428e-05, 2.197191e-05, 3.233353e-05, 3.926914e-05,
  4.937212e-06, 5.577869e-06, 4.394456e-06, 4.604468e-06, 4.735646e-06, 
    6.130915e-06, 5.790348e-06, 3.625778e-06, 3.380486e-06, 3.578299e-06, 
    5.032384e-06, 1.118312e-05, 1.859612e-05, 2.827855e-05, 3.908063e-05,
  6.496969e-06, 5.255182e-06, 4.129182e-06, 6.105494e-06, 3.92027e-06, 
    1.710113e-06, 1.810727e-06, 1.393631e-05, 5.294811e-05, 8.526646e-05, 
    8.498626e-05, 5.563907e-05, 2.652839e-05, 1.729484e-05, 2.175799e-05,
  8.788228e-06, 6.425459e-06, 6.069462e-06, 3.268643e-06, 2.638505e-06, 
    1.251149e-06, 4.912796e-06, 2.261565e-05, 8.015987e-05, 0.0001136855, 
    8.33131e-05, 3.744485e-05, 3.517524e-05, 2.111864e-05, 2.073274e-05,
  7.620626e-06, 5.422962e-06, 3.91482e-06, 2.703973e-06, 3.022421e-06, 
    1.697441e-06, 3.648123e-06, 3.465099e-05, 0.0001127026, 0.0001267305, 
    7.276944e-05, 4.171539e-05, 3.917195e-05, 3.799935e-05, 2.755842e-05,
  6.007558e-06, 4.421425e-06, 4.326123e-06, 4.071997e-06, 1.243387e-06, 
    2.376415e-06, 3.101932e-06, 4.398773e-05, 0.0001353745, 0.0001302905, 
    5.003243e-05, 5.145556e-05, 3.921134e-05, 4.003941e-05, 3.276103e-05,
  5.239246e-06, 4.244469e-06, 4.696263e-06, 2.220474e-06, 1.248464e-06, 
    2.375633e-06, 2.724476e-06, 5.697062e-05, 0.0001326291, 9.737574e-05, 
    4.631095e-05, 4.24266e-05, 5.37504e-05, 6.290043e-05, 4.302077e-05,
  6.132479e-06, 4.886564e-06, 3.440231e-06, 2.310439e-06, 9.532604e-07, 
    1.528611e-06, 2.95058e-06, 5.654806e-05, 0.0001159097, 6.304542e-05, 
    4.567533e-05, 5.56669e-05, 7.72139e-05, 6.33753e-05, 5.697305e-05,
  4.067257e-06, 5.055763e-06, 2.713745e-06, 1.844891e-06, 1.059814e-06, 
    5.257669e-07, 6.449838e-06, 5.153185e-05, 8.811872e-05, 5.551237e-05, 
    5.159044e-05, 8.691953e-05, 5.733934e-05, 5.392748e-05, 4.353002e-05,
  4.181289e-06, 4.176316e-06, 2.814036e-06, 1.214587e-06, 1.36744e-06, 
    8.559292e-07, 1.439202e-05, 5.985115e-05, 7.392959e-05, 5.332326e-05, 
    5.727846e-05, 6.698118e-05, 8.523987e-05, 7.468391e-05, 5.900492e-05,
  3.961151e-06, 3.59182e-06, 1.295842e-06, 1.278181e-06, 1.502551e-06, 
    7.969048e-06, 2.913007e-05, 6.403174e-05, 6.725425e-05, 5.937635e-05, 
    6.171724e-05, 6.534322e-05, 7.445931e-05, 6.195065e-05, 6.421625e-05,
  4.627483e-06, 3.167633e-06, 1.845807e-06, 1.065958e-06, 1.912535e-06, 
    1.299117e-05, 4.770686e-05, 6.462842e-05, 6.14296e-05, 6.251377e-05, 
    6.746225e-05, 6.282047e-05, 6.330144e-05, 6.048854e-05, 6.85496e-05,
  3.896703e-05, 4.510076e-05, 5.550132e-05, 7.378834e-05, 0.0001085836, 
    6.786697e-05, 7.161564e-05, 6.296136e-05, 3.249944e-05, 6.062653e-06, 
    2.546833e-06, 3.117504e-07, 2.547003e-09, 3.258854e-09, 1.801721e-08,
  5.603384e-05, 4.2434e-05, 4.371077e-05, 8.417825e-05, 9.048535e-05, 
    7.619688e-05, 8.470082e-05, 7.117403e-05, 2.813355e-05, 2.436318e-06, 
    1.213834e-06, 2.449568e-09, 1.593394e-09, 3.471645e-09, 1.876973e-08,
  6.502681e-05, 4.611573e-05, 7.125951e-05, 8.22462e-05, 8.789767e-05, 
    8.603024e-05, 9.610618e-05, 7.828596e-05, 2.677399e-05, 3.349013e-06, 
    1.950695e-06, 5.898602e-07, 5.036593e-08, 1.285385e-07, 1.067887e-07,
  5.570944e-05, 5.234479e-05, 6.093537e-05, 8.432919e-05, 7.302691e-05, 
    9.094945e-05, 0.0001037432, 8.87701e-05, 3.154019e-05, 3.981347e-06, 
    2.838726e-06, 1.982543e-06, 6.490154e-07, 4.325142e-07, 2.324926e-07,
  5.471109e-05, 4.669086e-05, 6.934347e-05, 6.944084e-05, 7.851324e-05, 
    9.948204e-05, 0.0001150113, 0.0001095714, 4.549954e-05, 6.096448e-06, 
    9.923781e-06, 3.793347e-06, 4.210759e-06, 4.745901e-06, 1.23976e-06,
  6.552535e-05, 5.071489e-05, 7.133175e-05, 7.635252e-05, 8.838243e-05, 
    0.0001037275, 0.0001305567, 0.0001238824, 6.049444e-05, 1.410049e-05, 
    1.429997e-05, 9.297607e-06, 7.768662e-06, 5.796921e-06, 7.232321e-06,
  7.412345e-05, 6.246458e-05, 7.633675e-05, 7.837715e-05, 0.0001181249, 
    0.0001152511, 0.0001434792, 0.0001425827, 6.279409e-05, 2.200143e-05, 
    2.100044e-05, 1.57593e-05, 1.332554e-05, 1.085257e-05, 1.119453e-05,
  8.089469e-05, 7.62714e-05, 9.098365e-05, 8.858809e-05, 0.0001185191, 
    0.0001425117, 0.0001743288, 0.0001544128, 8.113479e-05, 3.962034e-05, 
    3.505323e-05, 3.037337e-05, 2.051428e-05, 1.990918e-05, 1.907607e-05,
  8.174028e-05, 9.21239e-05, 9.79768e-05, 0.0001096591, 0.0001361413, 
    0.0001529023, 0.0002029222, 0.0001809253, 9.483958e-05, 4.926034e-05, 
    4.661181e-05, 3.895308e-05, 3.078291e-05, 2.706495e-05, 2.797337e-05,
  9.362358e-05, 0.0001049087, 0.0001163603, 0.0001226669, 0.0001353817, 
    0.0001676246, 0.0002314877, 0.0001984609, 0.0001008108, 7.131751e-05, 
    6.561068e-05, 6.026686e-05, 5.097227e-05, 3.31219e-05, 3.320128e-05,
  5.067309e-06, 7.482342e-06, 7.019633e-06, 5.732216e-06, 9.910178e-06, 
    1.500674e-05, 1.883143e-05, 2.386667e-05, 3.562328e-05, 6.194326e-05, 
    9.005159e-05, 0.0001014201, 9.311732e-05, 8.07137e-05, 8.698428e-05,
  5.173511e-06, 1.141503e-05, 1.499962e-05, 1.017243e-05, 6.731594e-06, 
    8.6102e-06, 1.453809e-05, 2.979958e-05, 5.186021e-05, 8.162016e-05, 
    0.0001121317, 0.0001246733, 0.0001327531, 0.0001314864, 0.0001389122,
  3.843615e-06, 1.498109e-05, 2.78606e-05, 2.915654e-05, 2.324238e-05, 
    1.597993e-05, 1.320083e-05, 2.25727e-05, 4.1197e-05, 6.569916e-05, 
    8.836278e-05, 0.0001042006, 0.0001229964, 0.0001261271, 0.0001447935,
  1.274851e-06, 9.777732e-06, 2.863084e-05, 3.996171e-05, 4.852838e-05, 
    5.111332e-05, 4.541588e-05, 4.903978e-05, 6.014587e-05, 6.09161e-05, 
    6.346803e-05, 7.076555e-05, 7.797831e-05, 9.308611e-05, 0.0001242629,
  4.173512e-06, 4.817151e-06, 8.683273e-06, 1.849237e-05, 3.22894e-05, 
    4.480168e-05, 5.256806e-05, 7.17455e-05, 9.353639e-05, 0.0001089604, 
    0.0001045005, 0.0001014634, 0.0001023034, 0.0001102129, 0.0001436313,
  5.095809e-06, 6.758461e-06, 5.471309e-06, 6.523684e-06, 7.269257e-06, 
    1.332654e-05, 2.780849e-05, 5.188993e-05, 8.268655e-05, 0.0001208963, 
    0.0001354452, 0.0001502099, 0.0001642118, 0.0001810659, 0.0002053834,
  6.909503e-06, 7.96955e-06, 8.18676e-06, 6.760563e-06, 7.513522e-06, 
    7.061677e-06, 1.253444e-05, 3.309723e-05, 7.112842e-05, 0.0001020262, 
    0.0001220376, 0.000142271, 0.0001650969, 0.0001897019, 0.0002139926,
  9.304055e-06, 9.55133e-06, 8.951895e-06, 9.449345e-06, 8.526486e-06, 
    7.929802e-06, 1.007588e-05, 2.873316e-05, 6.344084e-05, 9.873801e-05, 
    0.0001191083, 0.0001297921, 0.0001446416, 0.000160845, 0.0001767798,
  9.946441e-06, 1.182813e-05, 1.059095e-05, 8.548993e-06, 8.556437e-06, 
    8.838049e-06, 8.437494e-06, 1.475841e-05, 4.100894e-05, 7.294606e-05, 
    0.0001046532, 0.0001303901, 0.000148152, 0.0001581739, 0.0001598285,
  1.266441e-05, 1.460137e-05, 1.208308e-05, 1.003937e-05, 8.169824e-06, 
    8.696739e-06, 8.389501e-06, 6.938116e-06, 1.744537e-05, 3.806833e-05, 
    7.294065e-05, 0.0001149985, 0.0001493555, 0.0001847198, 0.0001897824,
  8.706075e-06, 9.850874e-06, 2.772826e-05, 5.593886e-05, 8.170056e-05, 
    8.600276e-05, 5.131133e-05, 4.14549e-05, 1.834942e-05, 1.560529e-05, 
    2.157466e-05, 2.858604e-05, 3.860067e-05, 7.010253e-05, 0.0001068088,
  1.257017e-05, 2.453788e-05, 5.146511e-05, 7.792126e-05, 0.000101332, 
    8.135389e-05, 7.004209e-05, 6.143438e-05, 4.135536e-05, 3.684165e-05, 
    3.934032e-05, 4.566179e-05, 6.860676e-05, 0.000115632, 0.0001392218,
  1.586692e-05, 3.020713e-05, 4.902177e-05, 5.974459e-05, 5.941168e-05, 
    6.166012e-05, 7.25822e-05, 6.633332e-05, 5.989167e-05, 5.337285e-05, 
    5.128156e-05, 5.141473e-05, 9.129546e-05, 0.0001384039, 0.0001298487,
  2.075143e-05, 3.634408e-05, 4.700191e-05, 3.934478e-05, 5.178283e-05, 
    5.935124e-05, 6.932612e-05, 7.013155e-05, 5.997987e-05, 4.792278e-05, 
    4.75417e-05, 5.463165e-05, 0.0001025283, 0.0001243985, 8.945025e-05,
  1.983662e-05, 3.911306e-05, 4.56289e-05, 4.807023e-05, 5.678588e-05, 
    6.629853e-05, 7.348951e-05, 6.823978e-05, 4.970547e-05, 4.261917e-05, 
    4.661104e-05, 6.258264e-05, 0.0001022484, 9.081961e-05, 5.933421e-05,
  1.755254e-05, 3.921063e-05, 6.056955e-05, 7.482402e-05, 7.423686e-05, 
    7.097899e-05, 6.832524e-05, 5.734036e-05, 4.255015e-05, 4.623421e-05, 
    5.047532e-05, 7.747635e-05, 8.667503e-05, 6.502757e-05, 5.543162e-05,
  4.257705e-05, 6.941978e-05, 9.028692e-05, 9.586117e-05, 9.238307e-05, 
    7.501247e-05, 6.290757e-05, 5.869726e-05, 5.440413e-05, 4.682452e-05, 
    6.161128e-05, 8.006933e-05, 6.255244e-05, 5.297413e-05, 4.636145e-05,
  7.927471e-05, 9.513492e-05, 0.0001049385, 9.908811e-05, 8.655607e-05, 
    7.153269e-05, 6.924857e-05, 7.649223e-05, 7.525715e-05, 7.65708e-05, 
    9.563247e-05, 8.058664e-05, 5.682926e-05, 4.580065e-05, 2.615773e-05,
  8.891376e-05, 9.876792e-05, 9.901452e-05, 8.543789e-05, 7.349734e-05, 
    6.991982e-05, 7.572036e-05, 9.349501e-05, 0.0001075491, 0.0001347928, 
    0.0001367371, 0.0001053817, 5.773438e-05, 2.703056e-05, 1.633058e-05,
  7.472255e-05, 7.764259e-05, 8.130038e-05, 8.177355e-05, 9.105397e-05, 
    9.527858e-05, 0.0001021616, 0.0001252332, 0.0001518057, 0.0001788817, 
    0.0001717969, 0.0001244047, 6.547189e-05, 1.81434e-05, 8.867983e-06,
  3.462199e-05, 4.19496e-05, 4.507309e-05, 3.094988e-05, 1.614345e-05, 
    9.532209e-06, 7.821623e-06, 7.032105e-06, 1.211014e-05, 2.672428e-05, 
    2.102036e-05, 4.038252e-05, 2.185886e-05, 1.896917e-05, 1.127301e-05,
  5.748174e-05, 6.230719e-05, 5.643632e-05, 4.109781e-05, 1.723384e-05, 
    7.523716e-06, 7.734945e-06, 7.108247e-06, 2.694406e-05, 1.803948e-05, 
    1.986198e-05, 1.872669e-05, 2.492743e-05, 2.855746e-05, 1.907615e-05,
  6.067567e-05, 5.802459e-05, 5.203834e-05, 2.376342e-05, 1.168946e-05, 
    9.508652e-06, 1.056825e-05, 1.144543e-05, 1.244797e-05, 2.321764e-05, 
    3.049542e-05, 2.230876e-05, 3.136863e-05, 3.700073e-05, 1.98822e-05,
  6.753253e-05, 5.180012e-05, 2.120684e-05, 1.017007e-05, 9.642437e-06, 
    1.004141e-05, 1.034907e-05, 1.557556e-05, 2.260527e-05, 2.920349e-05, 
    2.876532e-05, 2.140864e-05, 2.003772e-05, 2.18335e-05, 1.485699e-05,
  5.231565e-05, 1.575012e-05, 4.758314e-06, 6.365452e-06, 1.087232e-05, 
    1.322754e-05, 1.104473e-05, 1.455718e-05, 1.74781e-05, 3.727436e-05, 
    2.926895e-05, 2.039213e-05, 1.914484e-05, 1.842658e-05, 1.63818e-05,
  1.79335e-05, 6.266895e-06, 1.14999e-05, 1.270084e-05, 1.277118e-05, 
    1.621946e-05, 1.456596e-05, 1.5596e-05, 1.895705e-05, 1.013542e-05, 
    2.935861e-05, 1.693703e-05, 1.425804e-05, 1.8082e-05, 1.817341e-05,
  7.64742e-06, 5.496173e-06, 7.686447e-06, 1.037004e-05, 1.095059e-05, 
    1.85103e-05, 1.456641e-05, 1.015443e-05, 8.244781e-06, 8.829425e-06, 
    1.463176e-05, 9.036441e-06, 1.153162e-05, 1.849517e-05, 1.916046e-05,
  7.376807e-06, 6.056051e-06, 5.949991e-06, 9.031639e-06, 1.102457e-05, 
    1.168997e-05, 1.759616e-05, 2.350291e-05, 2.658295e-05, 1.680758e-05, 
    1.070444e-05, 1.521137e-05, 1.380319e-05, 2.671727e-05, 3.264182e-05,
  7.95926e-06, 7.634527e-06, 8.106203e-06, 7.044124e-06, 6.972603e-06, 
    1.197631e-05, 1.20151e-05, 1.450563e-05, 2.220103e-05, 2.03512e-05, 
    1.750797e-05, 2.036147e-05, 2.386743e-05, 4.132877e-05, 5.41929e-05,
  8.723561e-06, 7.315561e-06, 7.468632e-06, 5.461674e-06, 6.226785e-06, 
    5.183254e-06, 6.965994e-06, 3.76545e-06, 3.919653e-06, 7.513244e-06, 
    1.703512e-05, 2.691183e-05, 4.008644e-05, 4.914914e-05, 6.170251e-05,
  8.388677e-06, 6.701761e-06, 1.032347e-05, 7.639379e-06, 1.5242e-05, 
    1.971945e-05, 1.286156e-05, 1.669645e-05, 2.939292e-05, 2.965359e-05, 
    3.104749e-05, 2.356553e-05, 2.299337e-05, 1.899021e-05, 1.603923e-05,
  1.39312e-05, 1.33154e-05, 1.848515e-05, 1.553864e-05, 3.911967e-05, 
    3.642197e-05, 3.17051e-05, 2.999112e-05, 3.158317e-05, 5.405866e-05, 
    3.772685e-05, 3.272372e-05, 2.54889e-05, 2.034345e-05, 2.32177e-05,
  1.959118e-05, 2.068274e-05, 2.580932e-05, 3.712028e-05, 4.783858e-05, 
    4.843221e-05, 2.902428e-05, 2.48284e-05, 3.093682e-05, 5.158964e-05, 
    3.091828e-05, 6.20211e-05, 7.199444e-05, 3.301565e-05, 1.488284e-05,
  2.388494e-05, 2.900303e-05, 3.88782e-05, 3.221706e-05, 4.634824e-05, 
    3.313312e-05, 1.219803e-05, 1.753328e-05, 4.173877e-05, 5.11503e-05, 
    3.312614e-05, 2.632866e-05, 2.222864e-05, 2.815432e-05, 2.134244e-05,
  2.959122e-05, 2.070299e-05, 2.662212e-05, 3.442758e-05, 3.858426e-05, 
    2.558322e-05, 1.892099e-05, 2.150871e-05, 5.806121e-05, 8.037102e-05, 
    5.936594e-05, 3.64218e-05, 2.833533e-05, 2.833403e-05, 5.188731e-05,
  3.337047e-05, 2.647682e-05, 5.003356e-05, 4.675286e-05, 5.390976e-05, 
    6.007979e-05, 3.208836e-05, 3.647382e-05, 8.199854e-05, 9.040383e-05, 
    8.635507e-05, 3.328476e-05, 2.55876e-05, 3.627078e-05, 1.690794e-05,
  4.145233e-05, 5.017481e-05, 5.68935e-05, 6.710162e-05, 5.594152e-05, 
    5.4604e-05, 4.630215e-05, 5.869127e-05, 4.732145e-05, 8.050475e-05, 
    3.961389e-05, 2.354272e-05, 2.328686e-05, 2.400266e-05, 2.356291e-05,
  7.508787e-05, 8.055743e-05, 7.965701e-05, 7.999848e-05, 6.408948e-05, 
    5.25105e-05, 3.334707e-05, 1.205944e-05, 3.760855e-05, 7.300927e-05, 
    6.145761e-05, 7.170581e-05, 3.027753e-05, 3.508149e-05, 1.537652e-05,
  0.000113068, 0.0001726928, 0.0001509685, 6.30943e-05, 6.605803e-05, 
    7.482383e-05, 3.201914e-05, 2.990558e-05, 2.200324e-05, 4.596359e-05, 
    9.031909e-05, 4.707756e-05, 1.763447e-05, 1.743946e-05, 1.402283e-05,
  8.381446e-05, 9.311659e-05, 8.042352e-05, 0.0001307663, 0.0001186129, 
    0.0001086975, 6.25695e-05, 5.033648e-05, 9.07138e-06, 7.018064e-06, 
    2.696363e-05, 2.39256e-05, 2.704797e-05, 2.55293e-05, 2.442555e-05,
  4.498138e-06, 4.260837e-06, 3.287658e-06, 2.330009e-06, 2.090504e-06, 
    2.062055e-06, 1.710144e-06, 2.178757e-06, 1.969515e-06, 2.633305e-06, 
    2.633417e-06, 2.844534e-06, 4.41067e-06, 4.046215e-06, 4.236111e-06,
  5.965974e-06, 5.172017e-06, 3.624124e-06, 4.235546e-06, 3.597358e-06, 
    3.139955e-06, 2.923893e-06, 2.863473e-06, 2.741721e-06, 3.159132e-06, 
    2.939625e-06, 3.522021e-06, 3.62628e-06, 3.607465e-06, 3.127455e-06,
  1.14659e-05, 6.547505e-06, 5.328289e-06, 5.537554e-06, 4.948822e-06, 
    3.283566e-06, 4.284547e-06, 3.702787e-06, 5.065544e-06, 3.874432e-06, 
    4.05737e-06, 4.155821e-06, 4.402063e-06, 3.525322e-06, 3.395782e-06,
  1.823007e-05, 1.180349e-05, 1.12881e-05, 7.514268e-06, 5.17702e-06, 
    4.183138e-06, 4.236328e-06, 3.92125e-06, 5.748775e-06, 6.623206e-06, 
    6.578654e-06, 4.657038e-06, 4.160663e-06, 2.649814e-06, 4.195048e-06,
  2.597929e-05, 2.333388e-05, 1.976154e-05, 1.518008e-05, 9.94692e-06, 
    6.196154e-06, 4.987273e-06, 6.247268e-06, 7.419434e-06, 8.034058e-06, 
    7.721166e-06, 7.644081e-06, 7.827335e-06, 6.138779e-06, 5.326102e-06,
  3.355018e-05, 2.764349e-05, 3.488725e-05, 2.955078e-05, 2.840504e-05, 
    1.087153e-05, 4.431541e-06, 7.161155e-06, 1.370434e-05, 1.180026e-05, 
    9.481316e-06, 9.827135e-06, 1.208065e-05, 1.077902e-05, 1.083816e-05,
  3.590962e-05, 4.636661e-05, 3.877017e-05, 2.412811e-05, 5.343761e-05, 
    4.443886e-05, 1.288706e-05, 1.162044e-05, 3.002965e-05, 2.581854e-05, 
    1.624508e-05, 1.783241e-05, 9.229148e-06, 6.302052e-06, 5.75327e-06,
  1.904075e-05, 2.003924e-05, 3.2433e-05, 1.574663e-05, 3.368979e-05, 
    4.198177e-05, 9.464606e-06, 1.179931e-05, 3.322029e-05, 2.00901e-05, 
    2.705537e-05, 2.3547e-05, 1.722105e-05, 1.539623e-05, 7.162395e-06,
  3.034195e-05, 3.683876e-05, 3.330476e-05, 1.388194e-05, 9.872069e-06, 
    1.699453e-05, 2.392834e-05, 2.546011e-05, 3.837021e-05, 2.585131e-05, 
    3.012771e-05, 4.419948e-05, 1.145093e-05, 1.52318e-05, 8.95329e-06,
  0.0001295382, 0.0001313731, 8.723985e-05, 4.763129e-05, 3.276127e-05, 
    2.601018e-05, 1.75464e-05, 1.308174e-05, 1.995988e-05, 2.651012e-05, 
    3.32289e-05, 2.070036e-05, 2.263476e-05, 2.15358e-05, 1.177818e-05,
  4.051827e-06, 3.550698e-06, 3.277849e-06, 3.000679e-06, 3.604495e-06, 
    3.876349e-06, 3.352631e-06, 4.846278e-06, 2.065254e-05, 7.055486e-05, 
    0.0001471032, 0.0002235307, 0.0002618989, 0.0002870112, 0.0003104184,
  4.521848e-06, 3.006299e-06, 2.294985e-06, 2.238119e-06, 2.223745e-06, 
    3.186032e-06, 3.980561e-06, 2.479799e-06, 2.082469e-06, 3.05001e-06, 
    1.141306e-05, 4.7147e-05, 0.0001129368, 0.0001776499, 0.0002349059,
  5.14529e-06, 3.804588e-06, 2.165471e-06, 2.161477e-06, 2.222865e-06, 
    2.019504e-06, 2.453861e-06, 2.542991e-06, 3.075198e-06, 4.962261e-06, 
    8.663453e-06, 7.672524e-06, 2.331076e-05, 7.202686e-05, 0.0001439146,
  7.34794e-06, 4.075877e-06, 3.167757e-06, 3.15887e-06, 1.804391e-06, 
    1.12317e-06, 1.050703e-06, 1.029599e-06, 1.66773e-06, 1.143571e-06, 
    3.54442e-06, 5.774677e-06, 1.444918e-05, 3.11699e-05, 7.343018e-05,
  7.924068e-06, 5.397164e-06, 4.38865e-06, 3.608647e-06, 2.052542e-06, 
    2.262914e-06, 1.330419e-06, 6.407146e-07, 2.524839e-07, 3.736887e-07, 
    8.631679e-07, 2.931822e-06, 5.61158e-06, 1.01989e-05, 2.570308e-05,
  1.100784e-05, 6.848105e-06, 4.830088e-06, 3.971009e-06, 3.168141e-06, 
    2.202218e-06, 1.570409e-06, 5.849773e-07, 2.668401e-07, 1.497331e-07, 
    3.495142e-07, 3.98711e-07, 1.312558e-06, 2.721961e-06, 4.750542e-06,
  1.058213e-05, 9.492049e-06, 8.049645e-06, 5.045637e-06, 5.166927e-06, 
    3.50894e-06, 1.57722e-06, 9.944305e-07, 5.069941e-07, 3.916102e-07, 
    4.207976e-07, 6.088693e-07, 2.817897e-07, 4.992489e-07, 8.428123e-07,
  1.806953e-05, 1.262273e-05, 9.573752e-06, 6.945302e-06, 7.178865e-06, 
    8.320745e-06, 4.245185e-06, 2.50423e-06, 1.997588e-06, 1.949395e-06, 
    1.263532e-06, 1.031105e-06, 9.494393e-07, 6.730916e-07, 4.84064e-07,
  2.048296e-05, 1.379714e-05, 9.587761e-06, 8.064415e-06, 8.291132e-06, 
    8.211769e-06, 6.589609e-06, 5.200118e-06, 2.241901e-06, 2.461792e-06, 
    2.26157e-06, 1.303982e-06, 1.035096e-06, 8.443139e-07, 6.814609e-07,
  2.823249e-05, 2.330774e-05, 1.592189e-05, 1.18185e-05, 9.458419e-06, 
    1.022829e-05, 9.863366e-06, 5.76201e-06, 8.150824e-06, 2.960641e-06, 
    2.586034e-06, 2.385476e-06, 1.64199e-06, 1.193395e-06, 6.435149e-07,
  7.408797e-05, 0.0001205701, 0.0001799992, 0.0002826532, 0.0004042927, 
    0.0005149455, 0.0007273526, 0.001074923, 0.001120381, 0.0007243397, 
    0.0005211917, 0.000407679, 0.0002998024, 0.0001637479, 5.053101e-05,
  6.170427e-05, 8.098369e-05, 0.0001199108, 0.0001841572, 0.0002689092, 
    0.0003643779, 0.0005593468, 0.000960919, 0.001096659, 0.0008240907, 
    0.0006057415, 0.0005048788, 0.0004269553, 0.0002970254, 0.0001316551,
  3.682518e-05, 5.81335e-05, 9.264913e-05, 0.0001472662, 0.000205317, 
    0.000275858, 0.0003971041, 0.0007026911, 0.0008958643, 0.0008106089, 
    0.0006182775, 0.0004876259, 0.0004440458, 0.0003738084, 0.0002398915,
  1.165135e-05, 2.499945e-05, 4.906115e-05, 8.731907e-05, 0.0001497683, 
    0.0002392886, 0.0003180349, 0.000511448, 0.0006701908, 0.0006872079, 
    0.0005790928, 0.0004870621, 0.0004290005, 0.0004061165, 0.0003136051,
  1.047545e-06, 2.112234e-06, 6.500654e-06, 1.895409e-05, 4.794654e-05, 
    0.0001059946, 0.000203307, 0.0003277498, 0.0004621816, 0.0005275304, 
    0.0005463673, 0.000516193, 0.000487407, 0.0004280458, 0.0003812392,
  2.600263e-07, 1.768345e-07, 2.982453e-07, 1.433695e-06, 5.360586e-06, 
    1.673254e-05, 7.659182e-05, 0.0001797804, 0.0002842976, 0.0003626444, 
    0.0004111052, 0.0004683447, 0.0005064743, 0.00048904, 0.0004488072,
  3.440717e-07, 8.970748e-08, 8.282744e-08, 2.284401e-07, 3.394392e-07, 
    8.728741e-07, 7.753099e-06, 5.010231e-05, 0.0001403355, 0.0002259927, 
    0.0002762526, 0.0003379313, 0.0004236895, 0.0004794823, 0.0004467491,
  2.299143e-06, 1.815968e-07, 1.065221e-07, 1.062301e-07, 1.005033e-07, 
    1.661801e-07, 8.159332e-07, 6.608182e-06, 3.104185e-05, 9.788464e-05, 
    0.0001446372, 0.0002091379, 0.0002845221, 0.0003382012, 0.0003902582,
  5.386197e-06, 1.368898e-06, 2.308087e-07, 7.428063e-08, 1.410792e-07, 
    7.088413e-08, 1.228456e-07, 4.902662e-07, 2.372909e-06, 1.660378e-05, 
    4.357813e-05, 9.674155e-05, 0.000154076, 0.0002030815, 0.0002744571,
  8.640734e-06, 5.729228e-06, 1.00757e-06, 2.198953e-07, 8.893493e-08, 
    1.083319e-07, 2.545838e-08, 6.8544e-08, 2.656014e-07, 7.065597e-07, 
    4.355401e-06, 2.086314e-05, 4.427082e-05, 9.225238e-05, 0.00014677,
  7.245574e-05, 7.953868e-05, 8.140947e-05, 6.700328e-05, 3.574699e-05, 
    1.425644e-05, 9.476536e-06, 1.157169e-05, 1.596475e-05, 2.257633e-05, 
    2.525744e-05, 3.273925e-05, 3.494156e-05, 4.549262e-05, 4.564875e-05,
  7.241339e-05, 8.121647e-05, 9.744289e-05, 9.496193e-05, 7.696899e-05, 
    5.688026e-05, 4.576489e-05, 4.962969e-05, 2.667965e-05, 2.951799e-05, 
    2.829594e-05, 3.564418e-05, 4.527296e-05, 5.152704e-05, 5.619155e-05,
  7.219423e-05, 8.266047e-05, 9.347897e-05, 8.7926e-05, 9.166435e-05, 
    8.760206e-05, 8.299606e-05, 9.782887e-05, 9.902754e-05, 3.864301e-05, 
    3.265464e-05, 4.063647e-05, 4.18653e-05, 5.839549e-05, 6.477802e-05,
  7.826004e-05, 8.775706e-05, 8.44925e-05, 8.779082e-05, 9.322975e-05, 
    9.993673e-05, 0.000102441, 0.0001304601, 0.000172067, 0.0001128566, 
    4.758684e-05, 4.525617e-05, 5.532049e-05, 5.857956e-05, 5.918928e-05,
  6.787876e-05, 8.523511e-05, 9.968896e-05, 0.0001087526, 0.0001182306, 
    0.0001402177, 0.0001401598, 0.0001637172, 0.0002077952, 0.000192721, 
    0.0001267508, 5.061858e-05, 4.629899e-05, 5.733382e-05, 5.124407e-05,
  6.643998e-05, 9.396441e-05, 0.0001051436, 0.0001149974, 0.0001388664, 
    0.0001692603, 0.0002190521, 0.0002272775, 0.0002422143, 0.0002473078, 
    0.0002026442, 0.0001011909, 3.983112e-05, 3.621836e-05, 3.844719e-05,
  6.325975e-05, 8.787148e-05, 9.170363e-05, 9.799487e-05, 0.0001209316, 
    0.0001647304, 0.0002243483, 0.0002831334, 0.0002819644, 0.0003064614, 
    0.0002684898, 0.0001793086, 9.272004e-05, 4.99487e-05, 3.952493e-05,
  6.23205e-05, 7.77071e-05, 7.939725e-05, 7.728849e-05, 9.812002e-05, 
    0.0001466792, 0.0001983306, 0.0002450751, 0.0003132898, 0.0003454717, 
    0.0003268729, 0.0002696207, 0.0001833953, 0.0001328058, 7.601439e-05,
  6.692547e-05, 7.940183e-05, 7.899738e-05, 7.024817e-05, 7.231708e-05, 
    0.0001079815, 0.0001611318, 0.0002020557, 0.0002300512, 0.0003055236, 
    0.0003471303, 0.0003424241, 0.0002851511, 0.0002080338, 0.0001352167,
  8.137905e-05, 8.919875e-05, 7.904854e-05, 6.503928e-05, 6.053818e-05, 
    6.868424e-05, 0.0001031349, 0.0001440693, 0.0001844766, 0.0002160185, 
    0.0002816804, 0.0003427147, 0.0003325516, 0.0002936732, 0.0002083448,
  2.319909e-06, 2.130847e-06, 3.152306e-06, 2.769369e-06, 3.334058e-06, 
    4.912478e-06, 5.772536e-06, 7.616583e-06, 9.1239e-06, 1.091136e-05, 
    1.050216e-05, 1.409246e-05, 1.735196e-05, 2.771128e-05, 3.784928e-05,
  2.662782e-06, 2.425588e-06, 2.587192e-06, 4.112325e-06, 4.771617e-06, 
    5.535267e-06, 6.655243e-06, 8.047566e-06, 1.01518e-05, 1.304847e-05, 
    8.995403e-06, 9.287523e-06, 1.710626e-05, 3.160628e-05, 4.627246e-05,
  4.024216e-06, 3.948217e-06, 3.036843e-06, 4.660363e-06, 5.830905e-06, 
    7.510191e-06, 7.477688e-06, 7.07796e-06, 9.643755e-06, 9.907319e-06, 
    8.357461e-06, 8.628325e-06, 1.741979e-05, 3.541205e-05, 4.830968e-05,
  2.663316e-06, 3.139366e-06, 3.882906e-06, 5.317201e-06, 6.356343e-06, 
    5.735624e-06, 7.746919e-06, 7.910102e-06, 8.823319e-06, 9.550104e-06, 
    8.11747e-06, 6.933906e-06, 1.498678e-05, 2.94849e-05, 3.660638e-05,
  2.264384e-06, 3.700799e-06, 3.673807e-06, 5.137065e-06, 5.865376e-06, 
    6.232523e-06, 5.560776e-06, 7.024327e-06, 9.426023e-06, 1.118191e-05, 
    1.080779e-05, 9.131318e-06, 8.232328e-06, 1.067388e-05, 1.477805e-05,
  2.883255e-06, 3.630558e-06, 4.021085e-06, 7.372165e-06, 9.014026e-06, 
    5.41576e-06, 5.218024e-06, 9.455464e-06, 1.919868e-05, 2.244379e-05, 
    2.569713e-05, 2.230626e-05, 1.607542e-05, 1.958099e-05, 1.829423e-05,
  3.038331e-06, 4.142947e-06, 8.817996e-06, 9.401653e-06, 1.322647e-05, 
    6.123925e-06, 3.159945e-06, 1.290956e-05, 2.546346e-05, 3.911127e-05, 
    3.747987e-05, 3.433181e-05, 3.704146e-05, 2.804743e-05, 3.379726e-05,
  5.25454e-06, 4.521324e-06, 9.617211e-06, 9.156427e-06, 1.481142e-05, 
    8.258209e-06, 6.303072e-06, 1.962227e-05, 3.600784e-05, 4.558815e-05, 
    4.028725e-05, 4.743882e-05, 3.529837e-05, 3.59828e-05, 2.983863e-05,
  3.305507e-06, 2.666563e-06, 4.195177e-06, 7.176671e-06, 2.495523e-05, 
    3.023226e-05, 1.94106e-05, 1.194523e-05, 2.485053e-05, 4.460669e-05, 
    5.296259e-05, 4.928594e-05, 3.156379e-05, 3.034992e-05, 1.993441e-05,
  4.220257e-06, 5.006131e-06, 4.244921e-06, 4.806977e-06, 2.153262e-05, 
    3.208708e-05, 2.458664e-05, 1.740825e-05, 2.386747e-05, 4.261123e-05, 
    5.356633e-05, 5.270818e-05, 3.46318e-05, 2.061645e-05, 1.792392e-05,
  2.920066e-06, 3.895681e-06, 2.367899e-06, 3.832549e-06, 6.653804e-06, 
    2.65009e-05, 7.561437e-05, 0.00014336, 0.000215506, 0.0003174705, 
    0.0004136766, 0.000376125, 0.0001944927, 4.716737e-05, 1.014658e-05,
  3.233909e-06, 3.374549e-06, 2.938755e-06, 4.405517e-06, 7.222674e-06, 
    3.288983e-05, 8.259616e-05, 0.0001483283, 0.0002456135, 0.0003382555, 
    0.0004161042, 0.0003565779, 0.0001835797, 2.913636e-05, 8.429814e-06,
  2.426496e-06, 2.812177e-06, 4.56515e-06, 3.58764e-06, 1.135116e-05, 
    3.356113e-05, 7.699458e-05, 0.0001483762, 0.0002371006, 0.0003202541, 
    0.0003790706, 0.0003202268, 0.0001656475, 2.202584e-05, 1.140781e-05,
  4.098465e-06, 5.085341e-06, 3.255785e-06, 2.709211e-06, 9.003913e-06, 
    2.408122e-05, 5.405558e-05, 0.0001258309, 0.000193371, 0.0002660828, 
    0.000311686, 0.0002825945, 0.0001628072, 3.584354e-05, 2.395897e-05,
  3.527083e-06, 2.409595e-06, 2.940797e-06, 2.252088e-06, 7.925088e-06, 
    1.890399e-05, 5.054162e-05, 0.0001070629, 0.0001672711, 0.0002392392, 
    0.0002767213, 0.0002591065, 0.0001552719, 4.992314e-05, 3.066098e-05,
  3.663034e-06, 2.559239e-06, 2.907298e-06, 5.07244e-06, 9.406711e-06, 
    1.961817e-05, 5.734121e-05, 0.0001091547, 0.0001809203, 0.0002555891, 
    0.000272335, 0.0002349004, 0.0001262409, 3.170875e-05, 1.80189e-05,
  2.530991e-06, 1.995993e-06, 4.039134e-06, 7.795319e-06, 1.144334e-05, 
    1.749656e-05, 5.49482e-05, 0.0001122636, 0.0002061275, 0.0002832961, 
    0.0002546913, 0.000182247, 7.700153e-05, 1.474406e-05, 1.204136e-05,
  3.617411e-06, 3.374837e-06, 3.113286e-06, 7.240787e-06, 9.216097e-06, 
    1.572795e-05, 5.447725e-05, 0.0001237228, 0.0002400343, 0.0002781054, 
    0.0002113777, 0.0001214761, 3.045091e-05, 7.062929e-06, 8.30287e-06,
  4.376316e-06, 3.176231e-06, 3.322729e-06, 5.357484e-06, 5.82228e-06, 
    6.618601e-06, 4.807024e-05, 0.0001394182, 0.0002276871, 0.0002235233, 
    0.0001515875, 6.956296e-05, 1.196723e-05, 5.792603e-06, 6.712695e-06,
  3.38923e-06, 5.562378e-06, 2.240172e-06, 3.033512e-06, 2.559248e-06, 
    6.714379e-06, 5.55529e-05, 0.0001344189, 0.000173721, 0.0001407862, 
    8.675524e-05, 3.188994e-05, 4.927394e-06, 4.724269e-06, 6.175345e-06,
  3.351893e-05, 3.406493e-05, 4.701544e-05, 5.388599e-05, 3.558495e-05, 
    2.046291e-05, 2.161174e-05, 1.948406e-05, 2.109291e-05, 1.919814e-05, 
    3.001787e-05, 2.055657e-05, 3.724737e-05, 2.077414e-05, 1.185585e-05,
  4.358873e-05, 4.02419e-05, 5.988421e-05, 6.463403e-05, 4.749549e-05, 
    2.577806e-05, 2.080018e-05, 2.569756e-05, 1.854883e-05, 1.891278e-05, 
    1.869784e-05, 1.665811e-05, 1.892983e-05, 1.014317e-05, 1.390378e-05,
  5.151414e-05, 4.390895e-05, 6.935123e-05, 7.701672e-05, 4.622099e-05, 
    2.737632e-05, 3.343042e-05, 3.165934e-05, 2.553427e-05, 2.281498e-05, 
    1.568172e-05, 1.073173e-05, 1.06434e-05, 5.720657e-06, 5.504201e-06,
  5.326516e-05, 4.800273e-05, 7.773089e-05, 8.291425e-05, 4.288691e-05, 
    4.51901e-05, 5.204001e-05, 5.53268e-05, 4.279599e-05, 3.961688e-05, 
    3.348031e-05, 1.485714e-05, 7.458513e-06, 6.203139e-06, 6.769405e-06,
  5.498147e-05, 4.413302e-05, 8.619169e-05, 9.171331e-05, 5.104679e-05, 
    5.165337e-05, 7.046729e-05, 7.590438e-05, 6.634245e-05, 5.897985e-05, 
    3.908326e-05, 8.156685e-06, 1.508674e-05, 7.94167e-06, 8.989708e-06,
  5.954828e-05, 5.285477e-05, 9.476718e-05, 0.0001009091, 5.671892e-05, 
    6.330875e-05, 8.067187e-05, 8.833697e-05, 6.647634e-05, 5.460213e-05, 
    4.638865e-05, 2.109437e-05, 8.561629e-06, 6.042514e-06, 7.297013e-06,
  6.515575e-05, 5.884478e-05, 0.0001010475, 0.0001074852, 5.932688e-05, 
    6.348042e-05, 9.248772e-05, 9.792435e-05, 6.570694e-05, 5.431042e-05, 
    6.078945e-05, 3.74376e-05, 1.838946e-05, 8.866445e-06, 1.069998e-05,
  6.971111e-05, 6.821498e-05, 0.0001030765, 0.0001107491, 5.882094e-05, 
    6.722028e-05, 9.218061e-05, 0.000103024, 5.747933e-05, 6.763345e-05, 
    7.777251e-05, 6.279426e-05, 3.216881e-05, 1.265486e-05, 1.556015e-05,
  7.355034e-05, 6.335408e-05, 0.0001017361, 0.0001074672, 5.459802e-05, 
    6.822797e-05, 0.0001087736, 0.0001088006, 6.993554e-05, 0.0001071891, 
    0.0001089932, 7.49816e-05, 3.08546e-05, 9.298114e-06, 1.468361e-05,
  8.98725e-05, 6.244249e-05, 8.824206e-05, 0.0001021451, 4.994685e-05, 
    6.610435e-05, 0.0001240791, 0.0001235244, 9.960585e-05, 0.0001540608, 
    0.0001471727, 8.499439e-05, 2.456833e-05, 1.006597e-05, 8.879108e-06,
  1.200945e-06, 1.215306e-06, 3.68717e-06, 2.405818e-06, 4.945616e-06, 
    7.029601e-06, 7.043496e-06, 7.587415e-06, 6.033556e-06, 9.066599e-06, 
    1.156515e-05, 7.21005e-06, 3.65806e-06, 4.416358e-07, 2.444777e-06,
  4.684552e-06, 2.210076e-06, 1.298979e-06, 4.685235e-06, 7.284249e-06, 
    1.214023e-05, 8.277565e-06, 5.78354e-06, 4.849807e-06, 9.28902e-06, 
    8.754363e-06, 5.107649e-06, 1.234778e-06, 2.731972e-09, 4.359923e-09,
  8.337705e-06, 3.925602e-06, 4.176587e-06, 4.757527e-06, 5.753233e-06, 
    9.585289e-06, 6.419451e-06, 5.477037e-06, 9.059534e-06, 1.178617e-05, 
    1.215694e-05, 5.258382e-06, 5.068407e-06, 7.386632e-07, 3.151006e-06,
  1.497139e-05, 1.027026e-05, 8.375157e-06, 6.758119e-06, 8.156058e-06, 
    4.315084e-06, 2.822499e-06, 5.67054e-06, 1.151512e-05, 1.186825e-05, 
    1.055656e-05, 5.266444e-06, 1.814759e-06, 3.891751e-06, 3.425894e-06,
  1.537525e-05, 1.077578e-05, 8.509186e-06, 8.04388e-06, 1.008575e-05, 
    2.609626e-06, 2.951213e-06, 7.180729e-06, 1.200851e-05, 1.589356e-05, 
    7.836348e-06, 4.0418e-06, 3.094431e-06, 8.477133e-06, 3.074617e-06,
  8.134943e-06, 5.819258e-06, 6.093143e-06, 3.495436e-06, 6.450739e-06, 
    1.857138e-06, 1.227984e-05, 1.907762e-05, 7.157427e-06, 1.156147e-05, 
    1.547681e-05, 1.375204e-05, 3.198639e-06, 7.220999e-06, 1.251392e-05,
  3.268798e-06, 5.061012e-06, 5.44593e-06, 4.113686e-06, 8.929772e-06, 
    2.168218e-06, 1.888123e-06, 6.123318e-06, 1.840302e-05, 1.771013e-05, 
    4.587724e-05, 1.979678e-05, 1.625629e-05, 1.011381e-05, 1.150578e-05,
  2.202066e-06, 6.183855e-06, 6.274252e-06, 2.845307e-06, 3.59394e-06, 
    1.820974e-05, 4.606657e-07, 9.161062e-07, 1.146139e-05, 8.534223e-06, 
    4.588516e-06, 5.760889e-06, 1.752715e-05, 2.022689e-05, 2.899738e-05,
  1.037163e-06, 2.401703e-06, 2.592089e-06, 5.158733e-06, 8.78952e-06, 
    9.077094e-06, 4.369004e-06, 3.639758e-06, 7.579219e-06, 1.605145e-05, 
    1.377057e-05, 7.401787e-06, 1.542962e-05, 1.879127e-05, 5.317689e-06,
  1.087483e-06, 1.488482e-06, 1.251618e-06, 1.435306e-06, 2.813451e-06, 
    5.049398e-06, 3.22332e-06, 4.851991e-06, 8.85282e-06, 1.287649e-05, 
    1.898075e-05, 2.958275e-05, 1.768456e-05, 7.572908e-06, 5.69653e-06,
  2.162379e-06, 2.766683e-06, 3.483074e-06, 5.476368e-06, 4.424968e-06, 
    6.382046e-06, 1.048623e-05, 1.001171e-05, 9.165457e-06, 7.240012e-06, 
    4.415755e-06, 2.887899e-06, 2.098521e-06, 3.689069e-06, 7.371657e-06,
  9.97122e-07, 1.091862e-06, 7.537296e-07, 3.761023e-07, 1.15597e-06, 
    3.834873e-06, 3.508894e-06, 5.489708e-06, 9.205295e-06, 1.390957e-06, 
    1.035193e-06, 5.440002e-07, 2.958743e-06, 7.651712e-06, 1.014349e-05,
  1.383076e-06, 1.067047e-06, 7.607537e-07, 6.105166e-07, 3.117614e-07, 
    1.56671e-06, 1.837892e-06, 2.585183e-06, 4.207153e-06, 4.668584e-06, 
    1.621564e-06, 4.202944e-06, 7.084449e-06, 8.583123e-06, 9.922427e-06,
  1.553444e-06, 1.215e-06, 7.403594e-07, 5.281689e-07, 8.541426e-08, 
    1.282111e-06, 6.974901e-07, 1.618342e-06, 8.441308e-07, 6.265403e-06, 
    5.825136e-06, 8.860269e-06, 8.08821e-06, 6.745046e-06, 9.29932e-06,
  1.650821e-06, 9.226461e-07, 8.610817e-07, 1.064196e-06, 3.916261e-07, 
    3.096648e-07, 4.476768e-07, 8.125937e-08, 3.423278e-06, 7.782913e-06, 
    7.368942e-06, 8.804128e-06, 7.62043e-06, 9.85885e-06, 1.513447e-05,
  1.527201e-06, 8.766755e-07, 1.100294e-06, 1.480022e-06, 1.394432e-06, 
    8.106728e-08, 1.287154e-07, 1.029365e-06, 4.198874e-06, 6.307649e-06, 
    1.012076e-05, 1.109472e-05, 1.457912e-05, 1.401464e-05, 1.602011e-05,
  1.345084e-06, 1.434311e-06, 2.23198e-06, 3.23337e-06, 3.386262e-06, 
    5.340866e-07, 7.968185e-07, 2.882821e-06, 4.857421e-06, 7.040629e-06, 
    8.599403e-06, 1.182446e-05, 1.186174e-05, 1.235207e-05, 1.072513e-05,
  1.40758e-06, 3.204124e-06, 4.478727e-06, 3.805522e-06, 2.617347e-06, 
    2.451824e-06, 2.424863e-06, 3.60749e-06, 5.311451e-06, 6.309634e-06, 
    6.890426e-06, 8.083345e-06, 1.202507e-05, 1.291823e-05, 1.368198e-05,
  9.454282e-07, 1.3766e-06, 5.415539e-06, 4.015987e-06, 5.298036e-06, 
    4.709328e-06, 3.691923e-06, 4.668273e-06, 6.745083e-06, 5.037991e-06, 
    8.5004e-06, 7.281314e-06, 1.332692e-05, 1.379643e-05, 1.648526e-05,
  5.546341e-07, 2.009052e-06, 5.96537e-06, 2.220964e-06, 2.391073e-06, 
    7.000086e-06, 9.44531e-06, 6.516878e-06, 7.143411e-06, 5.734349e-06, 
    6.71595e-06, 1.096224e-05, 1.449909e-05, 1.687454e-05, 1.815484e-05,
  1.367788e-07, 3.655367e-07, 1.194272e-06, 1.026502e-06, 1.405114e-06, 
    8.302079e-07, 1.550495e-06, 5.402848e-07, 1.518716e-06, 9.941654e-07, 
    3.898425e-07, 7.127631e-09, 1.302296e-08, 3.437969e-07, 3.697469e-05,
  6.068898e-09, 1.469883e-07, 7.048102e-07, 1.172246e-06, 5.703085e-07, 
    1.276186e-06, 1.117136e-06, 7.361646e-07, 1.345575e-06, 9.737793e-07, 
    4.234328e-07, 3.126464e-07, 6.24147e-08, 1.964303e-06, 8.934393e-06,
  1.709138e-07, 2.571142e-07, 7.629714e-07, 5.57218e-07, 1.266944e-06, 
    1.086792e-06, 8.496611e-07, 8.788118e-07, 4.528067e-07, 7.279548e-07, 
    2.70504e-06, 5.584227e-06, 1.679094e-06, 3.581644e-06, 4.044646e-06,
  2.559586e-07, 1.409143e-07, 3.324573e-07, 5.448288e-07, 1.044572e-06, 
    1.037861e-06, 1.05009e-06, 1.838953e-06, 3.583875e-06, 4.692447e-06, 
    6.24711e-06, 7.410994e-06, 7.66501e-06, 6.900756e-06, 3.897321e-06,
  3.635172e-07, 8.900529e-07, 7.90269e-07, 6.183716e-07, 9.380202e-07, 
    1.608555e-06, 7.688218e-06, 4.912642e-06, 7.11552e-06, 1.08852e-05, 
    1.066817e-05, 9.323035e-06, 9.408064e-06, 7.420276e-06, 2.623561e-06,
  2.401734e-07, 7.485713e-07, 1.483954e-06, 2.114881e-06, 3.886708e-06, 
    3.753742e-06, 9.595722e-06, 1.112187e-05, 9.000713e-06, 5.711446e-06, 
    3.550297e-06, 8.455764e-06, 6.30249e-06, 6.047284e-06, 3.516178e-06,
  7.547384e-07, 1.250882e-06, 2.750572e-06, 7.661764e-06, 9.466593e-06, 
    1.166788e-05, 1.159766e-05, 1.260971e-05, 1.117264e-05, 3.241812e-06, 
    3.451429e-06, 4.933312e-06, 5.043629e-06, 5.848942e-06, 5.29064e-06,
  3.498488e-06, 3.91316e-06, 6.69093e-06, 6.595816e-06, 8.880326e-06, 
    1.212641e-05, 7.216118e-06, 5.841116e-06, 6.996907e-06, 4.992212e-06, 
    3.042074e-06, 5.158509e-06, 6.508155e-06, 6.692756e-06, 6.934496e-06,
  5.882597e-06, 5.863115e-06, 7.486555e-06, 6.017611e-06, 7.601553e-06, 
    8.07987e-06, 5.000398e-06, 7.417454e-06, 4.947252e-06, 3.913604e-06, 
    4.614669e-06, 8.598805e-06, 7.248959e-06, 6.041458e-06, 7.383615e-06,
  5.382798e-06, 8.402234e-06, 1.045121e-05, 1.045288e-05, 1.215055e-05, 
    1.055025e-05, 9.759707e-06, 6.586238e-06, 3.456656e-06, 8.114373e-06, 
    6.359431e-06, 3.011276e-06, 4.639133e-06, 4.583301e-06, 5.768899e-06 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
