netcdf atmos_daily.00010101-00010701.pv350K.tile2 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pv350K(time, grid_yt, grid_xt) ;
		pv350K:_FillValue = -1.e+10f ;
		pv350K:missing_value = -1.e+10f ;
		pv350K:units = "(K m**2) / (kg s)" ;
		pv350K:long_name = "350-K potential vorticity; needs x350 scaling" ;
		pv350K:cell_methods = "time: mean" ;
		pv350K:time_avg_info = "average_T1,average_T2,average_DT" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:53:56 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile2.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile2.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pv350K =
  -1.152597e-08, -1.242575e-08, -1.311111e-08, -1.362801e-08, -1.427807e-08, 
    -1.531632e-08, -1.571502e-08, -1.679802e-08, -1.768108e-08, 
    -1.770433e-08, -1.755651e-08, -1.736157e-08, -1.694493e-08, 
    -1.652093e-08, -1.607771e-08,
  -9.942039e-09, -1.097235e-08, -1.18535e-08, -1.247177e-08, -1.315546e-08, 
    -1.380663e-08, -1.468359e-08, -1.509875e-08, -1.575749e-08, 
    -1.639434e-08, -1.617013e-08, -1.586742e-08, -1.552977e-08, 
    -1.507326e-08, -1.46677e-08,
  -8.327726e-09, -9.278547e-09, -1.032448e-08, -1.11856e-08, -1.190493e-08, 
    -1.259758e-08, -1.333462e-08, -1.402435e-08, -1.426862e-08, 
    -1.469151e-08, -1.503246e-08, -1.473402e-08, -1.438969e-08, -1.38926e-08, 
    -1.346963e-08,
  -7.020802e-09, -7.700704e-09, -8.629867e-09, -9.67623e-09, -1.056414e-08, 
    -1.132559e-08, -1.198218e-08, -1.283065e-08, -1.322992e-08, -1.33578e-08, 
    -1.360355e-08, -1.366414e-08, -1.342542e-08, -1.306781e-08, -1.260943e-08,
  -5.244819e-09, -6.039624e-09, -6.844372e-09, -7.813499e-09, -9.003505e-09, 
    -1.004621e-08, -1.073797e-08, -1.143491e-08, -1.215647e-08, 
    -1.247187e-08, -1.24606e-08, -1.249531e-08, -1.245805e-08, -1.228813e-08, 
    -1.199928e-08,
  -3.487547e-09, -4.54028e-09, -5.242782e-09, -5.956367e-09, -6.825223e-09, 
    -8.067653e-09, -9.256897e-09, -1.010068e-08, -1.079468e-08, 
    -1.151488e-08, -1.171929e-08, -1.162417e-08, -1.154902e-08, 
    -1.145671e-08, -1.132708e-08,
  -2.199789e-09, -2.932914e-09, -3.79252e-09, -4.419265e-09, -5.113743e-09, 
    -5.846315e-09, -7.024714e-09, -8.393589e-09, -9.355908e-09, 
    -1.006322e-08, -1.066025e-08, -1.089131e-08, -1.083678e-08, 
    -1.068295e-08, -1.056823e-08,
  -1.410875e-09, -1.746793e-09, -2.385333e-09, -3.039489e-09, -3.55787e-09, 
    -4.116112e-09, -4.903992e-09, -6.149473e-09, -7.600808e-09, 
    -8.604677e-09, -9.180953e-09, -9.695343e-09, -9.945365e-09, 
    -9.881857e-09, -9.710114e-09,
  -1.238036e-09, -1.27962e-09, -1.422865e-09, -1.922654e-09, -2.454418e-09, 
    -2.895453e-09, -3.320068e-09, -3.97669e-09, -5.178145e-09, -6.73264e-09, 
    -7.781828e-09, -8.332671e-09, -8.848391e-09, -9.036319e-09, -9.037117e-09,
  -1.176383e-09, -1.143625e-09, -1.221623e-09, -1.434992e-09, -1.780073e-09, 
    -2.172308e-09, -2.533448e-09, -2.850154e-09, -3.363319e-09, 
    -4.515408e-09, -5.947426e-09, -6.977368e-09, -7.664052e-09, 
    -8.251912e-09, -8.419059e-09,
  -1.199831e-08, -1.185244e-08, -1.142727e-08, -1.000614e-08, -9.989741e-09, 
    -1.073041e-08, -1.114057e-08, -1.131262e-08, -1.244264e-08, 
    -1.351136e-08, -1.452225e-08, -1.586259e-08, -1.750312e-08, 
    -1.840523e-08, -1.95125e-08,
  -1.133006e-08, -1.19165e-08, -1.19862e-08, -1.14418e-08, -1.040147e-08, 
    -1.049594e-08, -1.095951e-08, -1.137615e-08, -1.183432e-08, 
    -1.282031e-08, -1.398038e-08, -1.499029e-08, -1.629827e-08, 
    -1.750711e-08, -1.843236e-08,
  -1.14812e-08, -1.156661e-08, -1.219543e-08, -1.211942e-08, -1.141729e-08, 
    -1.082523e-08, -1.088914e-08, -1.117322e-08, -1.159282e-08, 
    -1.212621e-08, -1.320079e-08, -1.455602e-08, -1.563994e-08, 
    -1.675077e-08, -1.77159e-08,
  -1.203952e-08, -1.147295e-08, -1.16236e-08, -1.233741e-08, -1.227362e-08, 
    -1.161963e-08, -1.120719e-08, -1.121933e-08, -1.146985e-08, 
    -1.187808e-08, -1.251375e-08, -1.377346e-08, -1.519307e-08, 
    -1.617248e-08, -1.702602e-08,
  -1.297624e-08, -1.219208e-08, -1.15721e-08, -1.183505e-08, -1.247507e-08, 
    -1.245935e-08, -1.182516e-08, -1.143832e-08, -1.149658e-08, 
    -1.181624e-08, -1.226383e-08, -1.308788e-08, -1.438584e-08, 
    -1.564342e-08, -1.644199e-08,
  -1.338577e-08, -1.292611e-08, -1.226756e-08, -1.189865e-08, -1.216997e-08, 
    -1.260481e-08, -1.259101e-08, -1.208663e-08, -1.172969e-08, 
    -1.189698e-08, -1.232204e-08, -1.272746e-08, -1.35974e-08, -1.486572e-08, 
    -1.59568e-08,
  -1.316979e-08, -1.333091e-08, -1.275759e-08, -1.229465e-08, -1.215643e-08, 
    -1.239691e-08, -1.269501e-08, -1.265991e-08, -1.236627e-08, 
    -1.226458e-08, -1.269454e-08, -1.29629e-08, -1.333283e-08, -1.40859e-08, 
    -1.513642e-08,
  -1.258753e-08, -1.332479e-08, -1.327039e-08, -1.260577e-08, -1.237481e-08, 
    -1.245189e-08, -1.265785e-08, -1.284052e-08, -1.284476e-08, 
    -1.266883e-08, -1.29179e-08, -1.333686e-08, -1.368051e-08, -1.408751e-08, 
    -1.468966e-08,
  -1.247014e-08, -1.269985e-08, -1.314227e-08, -1.30202e-08, -1.251253e-08, 
    -1.240235e-08, -1.248847e-08, -1.280063e-08, -1.303387e-08, -1.31238e-08, 
    -1.331193e-08, -1.360069e-08, -1.388127e-08, -1.423476e-08, -1.459136e-08,
  -1.067157e-08, -1.248197e-08, -1.252964e-08, -1.274493e-08, -1.271569e-08, 
    -1.247858e-08, -1.242808e-08, -1.251329e-08, -1.28752e-08, -1.303716e-08, 
    -1.345072e-08, -1.381502e-08, -1.393871e-08, -1.439624e-08, -1.476775e-08,
  -8.787681e-09, -8.609041e-09, -8.560748e-09, -8.830355e-09, -8.867562e-09, 
    -8.781359e-09, -8.503936e-09, -8.423308e-09, -8.521984e-09, 
    -8.653641e-09, -9.010302e-09, -9.398334e-09, -1.007244e-08, 
    -1.161625e-08, -1.33177e-08,
  -9.349169e-09, -9.234014e-09, -8.977599e-09, -8.874501e-09, -8.942087e-09, 
    -8.976568e-09, -8.993533e-09, -8.704252e-09, -8.616742e-09, 
    -8.563076e-09, -8.54557e-09, -8.809315e-09, -9.335573e-09, -9.981127e-09, 
    -1.080632e-08,
  -9.534208e-09, -9.616483e-09, -9.559459e-09, -9.330424e-09, -9.193886e-09, 
    -9.094124e-09, -9.134433e-09, -9.109462e-09, -8.86111e-09, -8.77905e-09, 
    -8.667813e-09, -8.529931e-09, -8.604506e-09, -9.01885e-09, -9.633643e-09,
  -9.540092e-09, -9.603809e-09, -9.765214e-09, -9.806528e-09, -9.686981e-09, 
    -9.451766e-09, -9.270991e-09, -9.284593e-09, -9.277715e-09, 
    -9.078235e-09, -8.987215e-09, -8.760221e-09, -8.626336e-09, 
    -8.677031e-09, -9.018006e-09,
  -9.653973e-09, -9.618468e-09, -9.603509e-09, -9.815578e-09, -9.951246e-09, 
    -9.936022e-09, -9.67295e-09, -9.423874e-09, -9.3574e-09, -9.326379e-09, 
    -9.284578e-09, -9.206532e-09, -8.95211e-09, -8.708297e-09, -8.692546e-09,
  -9.757166e-09, -9.628394e-09, -9.554619e-09, -9.489972e-09, -9.784076e-09, 
    -1.004362e-08, -1.01901e-08, -9.94394e-09, -9.706664e-09, -9.511047e-09, 
    -9.362327e-09, -9.410533e-09, -9.390257e-09, -9.224173e-09, -9.035768e-09,
  -1.023601e-08, -9.859751e-09, -9.630353e-09, -9.521608e-09, -9.526206e-09, 
    -9.824523e-09, -1.022397e-08, -1.040714e-08, -1.022865e-08, 
    -1.003824e-08, -9.74743e-09, -9.555376e-09, -9.471461e-09, -9.452759e-09, 
    -9.465211e-09,
  -1.050531e-08, -1.028568e-08, -9.935135e-09, -9.645822e-09, -9.581605e-09, 
    -9.683941e-09, -9.940703e-09, -1.029666e-08, -1.041736e-08, 
    -1.028099e-08, -1.007965e-08, -9.873875e-09, -9.733547e-09, 
    -9.595395e-09, -9.646345e-09,
  -1.046658e-08, -1.057374e-08, -1.041863e-08, -1.006229e-08, -9.740121e-09, 
    -9.610332e-09, -9.748526e-09, -9.995195e-09, -1.026172e-08, 
    -1.027961e-08, -1.004414e-08, -9.798803e-09, -9.686111e-09, -9.57995e-09, 
    -9.564985e-09,
  -1.037532e-08, -1.045954e-08, -1.067293e-08, -1.040117e-08, -9.949598e-09, 
    -9.747797e-09, -9.569068e-09, -9.73775e-09, -1.000194e-08, -1.016011e-08, 
    -1.002524e-08, -9.702616e-09, -9.485472e-09, -9.349232e-09, -9.237188e-09,
  -7.067799e-09, -7.282364e-09, -7.883546e-09, -8.762414e-09, -9.223413e-09, 
    -9.353284e-09, -9.546133e-09, -9.974923e-09, -1.068641e-08, -1.18209e-08, 
    -1.268247e-08, -1.321613e-08, -1.372132e-08, -1.409271e-08, -1.437362e-08,
  -6.801098e-09, -6.978726e-09, -7.220506e-09, -7.795133e-09, -8.502039e-09, 
    -8.867897e-09, -9.057193e-09, -9.285558e-09, -9.623181e-09, 
    -1.007346e-08, -1.089426e-08, -1.159557e-08, -1.202433e-08, 
    -1.235562e-08, -1.262473e-08,
  -6.689524e-09, -6.786105e-09, -6.914639e-09, -7.128885e-09, -7.668036e-09, 
    -8.219358e-09, -8.508726e-09, -8.712001e-09, -8.945816e-09, 
    -9.197791e-09, -9.514406e-09, -1.000257e-08, -1.048256e-08, 
    -1.077303e-08, -1.097659e-08,
  -6.693046e-09, -6.718734e-09, -6.752005e-09, -6.875246e-09, -7.076923e-09, 
    -7.522157e-09, -7.984587e-09, -8.244029e-09, -8.416515e-09, 
    -8.621909e-09, -8.757889e-09, -8.959684e-09, -9.249375e-09, 
    -9.510568e-09, -9.664096e-09,
  -6.890217e-09, -6.798001e-09, -6.764048e-09, -6.787828e-09, -6.909826e-09, 
    -7.092793e-09, -7.435267e-09, -7.79724e-09, -8.038372e-09, -8.233016e-09, 
    -8.40276e-09, -8.496324e-09, -8.608882e-09, -8.740415e-09, -8.834267e-09,
  -7.124387e-09, -7.120428e-09, -7.021514e-09, -6.921022e-09, -6.898618e-09, 
    -6.997094e-09, -7.161124e-09, -7.431677e-09, -7.683023e-09, 
    -7.905464e-09, -8.070852e-09, -8.223998e-09, -8.277006e-09, -8.34862e-09, 
    -8.392961e-09,
  -7.104886e-09, -7.183862e-09, -7.263195e-09, -7.18982e-09, -7.062803e-09, 
    -7.009359e-09, -7.073392e-09, -7.257901e-09, -7.482524e-09, -7.68848e-09, 
    -7.857997e-09, -7.987233e-09, -8.097555e-09, -8.147522e-09, -8.204125e-09,
  -7.375715e-09, -7.293034e-09, -7.278201e-09, -7.292014e-09, -7.194657e-09, 
    -7.141387e-09, -7.156554e-09, -7.291106e-09, -7.466342e-09, 
    -7.678306e-09, -7.87303e-09, -8.046238e-09, -8.187341e-09, -8.299494e-09, 
    -8.355458e-09,
  -7.570118e-09, -7.522908e-09, -7.379213e-09, -7.299896e-09, -7.342903e-09, 
    -7.367407e-09, -7.433591e-09, -7.548382e-09, -7.664299e-09, 
    -7.784625e-09, -7.959764e-09, -8.140979e-09, -8.336711e-09, -8.47726e-09, 
    -8.62101e-09,
  -7.590714e-09, -7.823424e-09, -7.703535e-09, -7.489964e-09, -7.408523e-09, 
    -7.545891e-09, -7.660879e-09, -7.822449e-09, -7.949573e-09, 
    -8.018812e-09, -8.153164e-09, -8.337426e-09, -8.518496e-09, 
    -8.736594e-09, -8.97516e-09,
  -6.658278e-09, -6.727318e-09, -6.808565e-09, -6.919183e-09, -7.023923e-09, 
    -7.197501e-09, -7.340927e-09, -7.503007e-09, -7.753693e-09, 
    -8.032488e-09, -8.427343e-09, -9.08217e-09, -9.808637e-09, -1.050055e-08, 
    -1.11592e-08,
  -6.631881e-09, -6.727104e-09, -6.841296e-09, -6.971556e-09, -7.116358e-09, 
    -7.323552e-09, -7.523975e-09, -7.619185e-09, -7.730666e-09, 
    -7.926696e-09, -8.185426e-09, -8.584375e-09, -9.14955e-09, -9.815929e-09, 
    -1.056744e-08,
  -6.651302e-09, -6.769238e-09, -6.890887e-09, -7.011046e-09, -7.121757e-09, 
    -7.291492e-09, -7.520274e-09, -7.681264e-09, -7.74171e-09, -7.845028e-09, 
    -8.004393e-09, -8.285232e-09, -8.752592e-09, -9.328962e-09, -9.88786e-09,
  -6.498176e-09, -6.662937e-09, -6.832742e-09, -6.95602e-09, -7.077316e-09, 
    -7.200471e-09, -7.3872e-09, -7.616414e-09, -7.749726e-09, -7.883329e-09, 
    -8.009324e-09, -8.181044e-09, -8.438325e-09, -8.889038e-09, -9.477328e-09,
  -6.422538e-09, -6.590978e-09, -6.726421e-09, -6.827022e-09, -6.943937e-09, 
    -7.066954e-09, -7.221605e-09, -7.447551e-09, -7.648458e-09, 
    -7.822461e-09, -8.009111e-09, -8.2206e-09, -8.442598e-09, -8.739575e-09, 
    -9.100535e-09,
  -6.203711e-09, -6.415557e-09, -6.602331e-09, -6.711423e-09, -6.803432e-09, 
    -6.916058e-09, -7.06285e-09, -7.248836e-09, -7.506062e-09, -7.739683e-09, 
    -7.977489e-09, -8.236169e-09, -8.45362e-09, -8.695386e-09, -8.956894e-09,
  -6.051836e-09, -6.303941e-09, -6.590869e-09, -6.751646e-09, -6.798102e-09, 
    -6.809715e-09, -6.903411e-09, -7.075824e-09, -7.3523e-09, -7.680861e-09, 
    -7.93977e-09, -8.201612e-09, -8.374873e-09, -8.522446e-09, -8.662965e-09,
  -5.917894e-09, -6.264887e-09, -6.492863e-09, -6.679944e-09, -6.791256e-09, 
    -6.833456e-09, -6.818188e-09, -6.866292e-09, -7.076586e-09, 
    -7.407278e-09, -7.743165e-09, -8.007174e-09, -8.201073e-09, 
    -8.322366e-09, -8.424713e-09,
  -5.609876e-09, -6.159591e-09, -6.459023e-09, -6.551806e-09, -6.444295e-09, 
    -6.567883e-09, -6.754117e-09, -6.882999e-09, -6.946293e-09, 
    -7.120084e-09, -7.389958e-09, -7.677193e-09, -7.863551e-09, 
    -8.031874e-09, -8.140887e-09,
  -5.036761e-09, -5.59881e-09, -5.834099e-09, -5.967299e-09, -6.370152e-09, 
    -6.546756e-09, -6.743993e-09, -6.785553e-09, -6.861052e-09, 
    -7.000696e-09, -7.176441e-09, -7.389742e-09, -7.582457e-09, 
    -7.736651e-09, -7.85703e-09,
  -1.136881e-08, -1.117924e-08, -1.092254e-08, -1.068959e-08, -1.046506e-08, 
    -1.018699e-08, -9.883305e-09, -9.67521e-09, -9.466456e-09, -9.335816e-09, 
    -9.19601e-09, -9.085477e-09, -8.937958e-09, -8.773757e-09, -8.534015e-09,
  -9.555237e-09, -9.31682e-09, -9.044836e-09, -8.763177e-09, -8.507718e-09, 
    -8.24542e-09, -8.003664e-09, -7.853626e-09, -7.778971e-09, -7.760183e-09, 
    -7.71051e-09, -7.650485e-09, -7.578032e-09, -7.466048e-09, -7.298015e-09,
  -7.482467e-09, -7.50947e-09, -7.382168e-09, -7.202885e-09, -6.972181e-09, 
    -6.707349e-09, -6.500679e-09, -6.385732e-09, -6.396329e-09, 
    -6.437827e-09, -6.415417e-09, -6.410769e-09, -6.406494e-09, -6.36411e-09, 
    -6.257187e-09,
  -4.749565e-09, -4.922775e-09, -4.96863e-09, -4.972191e-09, -4.933761e-09, 
    -4.837314e-09, -4.701622e-09, -4.678162e-09, -4.746146e-09, 
    -4.871877e-09, -4.941615e-09, -4.986587e-09, -5.054665e-09, 
    -5.129498e-09, -5.137143e-09,
  -2.500983e-09, -2.692298e-09, -2.85295e-09, -3.019203e-09, -3.179322e-09, 
    -3.285473e-09, -3.354826e-09, -3.409348e-09, -3.47937e-09, -3.533357e-09, 
    -3.596767e-09, -3.692988e-09, -3.775335e-09, -3.900347e-09, -4.039997e-09,
  -1.485057e-09, -1.577416e-09, -1.733781e-09, -1.952974e-09, -2.184332e-09, 
    -2.414921e-09, -2.643676e-09, -2.849635e-09, -2.988038e-09, 
    -3.071791e-09, -3.122195e-09, -3.18042e-09, -3.283719e-09, -3.4466e-09, 
    -3.657794e-09,
  -1.373301e-09, -1.430665e-09, -1.556371e-09, -1.739221e-09, -1.97533e-09, 
    -2.17409e-09, -2.378628e-09, -2.584237e-09, -2.766548e-09, -2.911198e-09, 
    -3.015538e-09, -3.093701e-09, -3.239699e-09, -3.423586e-09, -3.636793e-09,
  -1.32091e-09, -1.383799e-09, -1.462928e-09, -1.615944e-09, -1.780663e-09, 
    -1.952215e-09, -2.11728e-09, -2.315024e-09, -2.510503e-09, -2.703029e-09, 
    -2.876312e-09, -3.022347e-09, -3.220761e-09, -3.447764e-09, -3.698688e-09,
  -1.407479e-09, -1.410555e-09, -1.454615e-09, -1.54086e-09, -1.663086e-09, 
    -1.839062e-09, -1.992336e-09, -2.147782e-09, -2.313625e-09, 
    -2.470587e-09, -2.637241e-09, -2.82925e-09, -3.063124e-09, -3.323085e-09, 
    -3.585852e-09,
  -1.425126e-09, -1.386862e-09, -1.386848e-09, -1.391937e-09, -1.4787e-09, 
    -1.708327e-09, -1.941959e-09, -2.119216e-09, -2.243395e-09, 
    -2.371075e-09, -2.550868e-09, -2.789685e-09, -3.049447e-09, 
    -3.326047e-09, -3.590867e-09,
  -1.004914e-08, -9.867713e-09, -9.315571e-09, -8.869373e-09, -8.503548e-09, 
    -8.143624e-09, -8.03472e-09, -8.065917e-09, -8.206513e-09, -8.426725e-09, 
    -8.816872e-09, -9.470986e-09, -1.034065e-08, -1.133108e-08, -1.219279e-08,
  -1.032082e-08, -1.06225e-08, -1.051436e-08, -9.986173e-09, -9.518398e-09, 
    -9.112651e-09, -8.600618e-09, -8.155106e-09, -7.784069e-09, 
    -7.734188e-09, -7.866058e-09, -8.404975e-09, -9.107914e-09, 
    -1.001415e-08, -1.100896e-08,
  -8.315766e-09, -9.719575e-09, -1.07985e-08, -1.134696e-08, -1.111245e-08, 
    -1.055503e-08, -9.962183e-09, -9.447507e-09, -8.897416e-09, 
    -8.396349e-09, -7.89029e-09, -7.746911e-09, -8.183179e-09, -8.830415e-09, 
    -9.7827e-09,
  -5.403448e-09, -6.722074e-09, -8.138907e-09, -9.654629e-09, -1.100968e-08, 
    -1.172681e-08, -1.176226e-08, -1.115312e-08, -1.045885e-08, 
    -9.826795e-09, -9.278386e-09, -8.50705e-09, -8.076725e-09, -8.293104e-09, 
    -8.963149e-09,
  -2.774472e-09, -3.696845e-09, -4.899713e-09, -6.332655e-09, -7.796748e-09, 
    -9.376399e-09, -1.077452e-08, -1.175818e-08, -1.204845e-08, 
    -1.150265e-08, -1.080315e-08, -9.776043e-09, -9.062994e-09, 
    -8.556994e-09, -8.575137e-09,
  -1.874946e-09, -2.034068e-09, -2.359834e-09, -3.029754e-09, -4.087703e-09, 
    -5.561279e-09, -7.09357e-09, -8.64955e-09, -9.932893e-09, -1.117742e-08, 
    -1.177194e-08, -1.164476e-08, -1.111855e-08, -1.004225e-08, -8.870459e-09,
  -1.907134e-09, -1.867963e-09, -1.848211e-09, -1.907337e-09, -2.116089e-09, 
    -2.608522e-09, -3.49567e-09, -4.807783e-09, -6.253035e-09, -7.626019e-09, 
    -8.898306e-09, -9.979559e-09, -1.069409e-08, -1.100668e-08, -1.070143e-08,
  -2.10801e-09, -2.029351e-09, -1.929553e-09, -1.849685e-09, -1.84243e-09, 
    -1.885015e-09, -2.040813e-09, -2.404624e-09, -3.169694e-09, 
    -4.259472e-09, -5.629222e-09, -6.874037e-09, -8.079903e-09, 
    -8.920815e-09, -9.518475e-09,
  -2.463916e-09, -2.330278e-09, -2.195467e-09, -2.048404e-09, -1.901935e-09, 
    -1.800515e-09, -1.766117e-09, -1.757701e-09, -1.889032e-09, 
    -2.233305e-09, -2.978794e-09, -4.043542e-09, -5.290616e-09, -6.50145e-09, 
    -7.494039e-09,
  -2.637542e-09, -2.561056e-09, -2.501388e-09, -2.410382e-09, -2.278158e-09, 
    -2.118119e-09, -1.90373e-09, -1.740923e-09, -1.674385e-09, -1.776104e-09, 
    -1.915165e-09, -2.272145e-09, -2.881609e-09, -3.7745e-09, -4.847521e-09,
  -1.212733e-08, -1.271781e-08, -1.327192e-08, -1.374817e-08, -1.406273e-08, 
    -1.435023e-08, -1.44804e-08, -1.457186e-08, -1.457731e-08, -1.455046e-08, 
    -1.426229e-08, -1.365119e-08, -1.285829e-08, -1.20285e-08, -1.133329e-08,
  -1.003511e-08, -1.063812e-08, -1.127925e-08, -1.187715e-08, -1.236349e-08, 
    -1.27277e-08, -1.295398e-08, -1.30647e-08, -1.308319e-08, -1.309819e-08, 
    -1.30282e-08, -1.27574e-08, -1.216026e-08, -1.148407e-08, -1.086573e-08,
  -7.940812e-09, -8.517752e-09, -9.097576e-09, -9.658368e-09, -1.021057e-08, 
    -1.06287e-08, -1.097264e-08, -1.115855e-08, -1.125977e-08, -1.136163e-08, 
    -1.150913e-08, -1.158148e-08, -1.12986e-08, -1.079467e-08, -1.030384e-08,
  -5.448257e-09, -6.142951e-09, -6.713551e-09, -7.262953e-09, -7.766727e-09, 
    -8.217462e-09, -8.557437e-09, -8.866192e-09, -9.104464e-09, 
    -9.308756e-09, -9.587168e-09, -9.981092e-09, -1.014938e-08, 
    -9.990063e-09, -9.660126e-09,
  -3.549373e-09, -4.024608e-09, -4.52265e-09, -4.963425e-09, -5.393988e-09, 
    -5.771603e-09, -6.140872e-09, -6.474989e-09, -6.851956e-09, 
    -7.152635e-09, -7.492075e-09, -7.943687e-09, -8.49129e-09, -8.909905e-09, 
    -8.892711e-09,
  -2.462066e-09, -2.745242e-09, -3.062066e-09, -3.328955e-09, -3.603732e-09, 
    -3.861737e-09, -4.138758e-09, -4.426197e-09, -4.786838e-09, 
    -5.200144e-09, -5.58196e-09, -6.107264e-09, -6.724798e-09, -7.464358e-09, 
    -8.038088e-09,
  -2.10164e-09, -2.241661e-09, -2.443063e-09, -2.633437e-09, -2.776362e-09, 
    -2.926827e-09, -3.081658e-09, -3.261052e-09, -3.518139e-09, 
    -3.871262e-09, -4.284336e-09, -4.746086e-09, -5.351593e-09, 
    -6.038622e-09, -6.981766e-09,
  -1.926543e-09, -2.017584e-09, -2.143152e-09, -2.298581e-09, -2.421583e-09, 
    -2.535246e-09, -2.625039e-09, -2.743852e-09, -2.857216e-09, 
    -3.095677e-09, -3.401066e-09, -3.784157e-09, -4.300228e-09, 
    -4.917817e-09, -5.730665e-09,
  -1.80554e-09, -1.862199e-09, -1.947254e-09, -2.030285e-09, -2.120515e-09, 
    -2.211155e-09, -2.317624e-09, -2.402981e-09, -2.516625e-09, 
    -2.591678e-09, -2.786744e-09, -3.015902e-09, -3.424122e-09, 
    -3.949471e-09, -4.698359e-09,
  -1.657006e-09, -1.671073e-09, -1.73314e-09, -1.797152e-09, -1.863599e-09, 
    -1.91276e-09, -1.978527e-09, -2.061166e-09, -2.201769e-09, -2.332938e-09, 
    -2.489961e-09, -2.616179e-09, -2.815984e-09, -3.155455e-09, -3.669775e-09,
  -6.607806e-09, -6.510198e-09, -6.220078e-09, -5.734333e-09, -5.525351e-09, 
    -5.553365e-09, -5.670302e-09, -6.098957e-09, -6.561351e-09, 
    -7.263576e-09, -7.904289e-09, -8.638332e-09, -9.420707e-09, -1.03149e-08, 
    -1.10803e-08,
  -8.085598e-09, -8.265468e-09, -8.163193e-09, -7.621114e-09, -7.012003e-09, 
    -6.75386e-09, -7.041333e-09, -7.321447e-09, -7.752897e-09, -8.298419e-09, 
    -8.895856e-09, -9.658553e-09, -1.054979e-08, -1.143454e-08, -1.204636e-08,
  -8.775217e-09, -8.863895e-09, -8.887637e-09, -8.960646e-09, -8.708663e-09, 
    -8.311502e-09, -8.347576e-09, -8.713167e-09, -9.013803e-09, 
    -9.435754e-09, -9.917823e-09, -1.06954e-08, -1.148652e-08, -1.225679e-08, 
    -1.288854e-08,
  -9.736197e-09, -9.880507e-09, -9.859003e-09, -9.651452e-09, -9.375689e-09, 
    -9.170101e-09, -9.270268e-09, -9.315359e-09, -9.696881e-09, 
    -1.015678e-08, -1.07129e-08, -1.148909e-08, -1.217103e-08, -1.287263e-08, 
    -1.378551e-08,
  -1.121543e-08, -1.081088e-08, -1.058834e-08, -1.079659e-08, -1.072736e-08, 
    -1.052498e-08, -1.028237e-08, -1.044841e-08, -1.068194e-08, 
    -1.091646e-08, -1.133733e-08, -1.212647e-08, -1.307585e-08, 
    -1.392865e-08, -1.490065e-08,
  -8.351755e-09, -1.133344e-08, -1.259515e-08, -1.166883e-08, -1.12702e-08, 
    -1.136212e-08, -1.126525e-08, -1.126826e-08, -1.141226e-08, 
    -1.168302e-08, -1.211661e-08, -1.284009e-08, -1.371783e-08, 
    -1.469302e-08, -1.592039e-08,
  -4.293849e-09, -6.63495e-09, -9.80562e-09, -1.26197e-08, -1.308152e-08, 
    -1.206488e-08, -1.14642e-08, -1.164056e-08, -1.190287e-08, -1.200284e-08, 
    -1.223295e-08, -1.285869e-08, -1.387217e-08, -1.49769e-08, -1.635242e-08,
  -2.106e-09, -3.419975e-09, -5.470246e-09, -7.853663e-09, -1.101466e-08, 
    -1.31029e-08, -1.269659e-08, -1.181971e-08, -1.15914e-08, -1.204227e-08, 
    -1.212428e-08, -1.250754e-08, -1.331731e-08, -1.469127e-08, -1.634567e-08,
  -1.751096e-09, -1.922489e-09, -2.900921e-09, -4.513287e-09, -6.427184e-09, 
    -8.718332e-09, -1.113836e-08, -1.243648e-08, -1.181504e-08, 
    -1.144545e-08, -1.147214e-08, -1.191998e-08, -1.245573e-08, 
    -1.365663e-08, -1.56268e-08,
  -1.541654e-09, -1.599498e-09, -1.759373e-09, -2.442555e-09, -3.779533e-09, 
    -5.320961e-09, -6.993382e-09, -8.874674e-09, -1.052939e-08, 
    -1.143119e-08, -1.117599e-08, -1.086927e-08, -1.120149e-08, 
    -1.206689e-08, -1.364169e-08,
  -5.720582e-09, -6.458531e-09, -7.179332e-09, -7.814602e-09, -8.17977e-09, 
    -8.314339e-09, -8.262523e-09, -8.025069e-09, -7.606105e-09, 
    -7.130569e-09, -6.524853e-09, -5.888116e-09, -5.162272e-09, 
    -4.457368e-09, -3.898909e-09,
  -4.389379e-09, -5.14974e-09, -5.987765e-09, -6.789533e-09, -7.35038e-09, 
    -7.627326e-09, -7.74406e-09, -7.730346e-09, -7.474781e-09, -6.977014e-09, 
    -6.293126e-09, -5.639152e-09, -4.954351e-09, -4.395576e-09, -4.169012e-09,
  -3.481574e-09, -4.081042e-09, -4.824994e-09, -5.69925e-09, -6.492598e-09, 
    -6.948059e-09, -7.13653e-09, -7.279027e-09, -7.198377e-09, -6.856737e-09, 
    -6.248608e-09, -5.607536e-09, -5.048755e-09, -4.570795e-09, -4.30696e-09,
  -2.881838e-09, -3.310417e-09, -3.893211e-09, -4.684876e-09, -5.522998e-09, 
    -6.130133e-09, -6.508538e-09, -6.697457e-09, -6.630403e-09, 
    -6.434333e-09, -6.030396e-09, -5.536448e-09, -5.017707e-09, 
    -4.537821e-09, -4.285238e-09,
  -2.694482e-09, -2.869452e-09, -3.274486e-09, -3.926937e-09, -4.736749e-09, 
    -5.416052e-09, -5.807882e-09, -6.147917e-09, -6.123937e-09, 
    -5.852729e-09, -5.503527e-09, -5.257947e-09, -4.836592e-09, 
    -4.367427e-09, -4.299295e-09,
  -2.653644e-09, -2.657023e-09, -2.870074e-09, -3.370452e-09, -4.089171e-09, 
    -4.79104e-09, -5.414901e-09, -5.618185e-09, -5.612343e-09, -5.520855e-09, 
    -5.183206e-09, -4.833222e-09, -4.572667e-09, -4.343469e-09, -4.34382e-09,
  -2.622464e-09, -2.629264e-09, -2.679573e-09, -2.987674e-09, -3.602839e-09, 
    -4.32506e-09, -4.882273e-09, -5.382692e-09, -5.543262e-09, -5.213166e-09, 
    -4.99805e-09, -4.768866e-09, -4.462729e-09, -4.337645e-09, -4.523899e-09,
  -2.205017e-09, -2.480285e-09, -2.615743e-09, -2.746593e-09, -3.202345e-09, 
    -4.014022e-09, -4.633776e-09, -5.051538e-09, -5.315666e-09, 
    -5.430024e-09, -4.982886e-09, -4.672901e-09, -4.478022e-09, 
    -4.387924e-09, -4.738898e-09,
  -1.729804e-09, -2.106735e-09, -2.448975e-09, -2.595705e-09, -2.894324e-09, 
    -3.588952e-09, -4.693869e-09, -5.431697e-09, -5.411625e-09, 
    -5.405224e-09, -5.331327e-09, -4.979365e-09, -4.625137e-09, 
    -4.486383e-09, -4.958464e-09,
  -1.281027e-09, -1.644597e-09, -2.086646e-09, -2.4169e-09, -2.606353e-09, 
    -3.116861e-09, -3.999308e-09, -5.413889e-09, -6.232411e-09, 
    -6.220555e-09, -5.603039e-09, -5.134301e-09, -4.915988e-09, 
    -4.843776e-09, -5.155079e-09,
  -4.248926e-09, -4.745461e-09, -5.230566e-09, -5.985862e-09, -6.976887e-09, 
    -7.845195e-09, -8.658272e-09, -9.412545e-09, -1.004587e-08, 
    -1.066145e-08, -1.11739e-08, -1.154768e-08, -1.188179e-08, -1.207804e-08, 
    -1.200824e-08,
  -3.471106e-09, -4.239668e-09, -4.84722e-09, -5.34766e-09, -6.035012e-09, 
    -6.906065e-09, -7.714666e-09, -8.617001e-09, -9.444737e-09, 
    -1.011313e-08, -1.066072e-08, -1.101718e-08, -1.134737e-08, 
    -1.153577e-08, -1.146037e-08,
  -2.733703e-09, -3.565114e-09, -4.296568e-09, -4.946498e-09, -5.412088e-09, 
    -6.06451e-09, -6.854286e-09, -7.684797e-09, -8.60592e-09, -9.439961e-09, 
    -1.013316e-08, -1.065476e-08, -1.100185e-08, -1.115261e-08, -1.098715e-08,
  -2.423145e-09, -3.036017e-09, -3.695107e-09, -4.399819e-09, -5.073306e-09, 
    -5.532585e-09, -6.184703e-09, -6.897007e-09, -7.752762e-09, 
    -8.619527e-09, -9.416362e-09, -1.010063e-08, -1.058378e-08, -1.08241e-08, 
    -1.066649e-08,
  -2.279586e-09, -2.536659e-09, -3.232225e-09, -3.860026e-09, -4.583808e-09, 
    -5.232716e-09, -5.709671e-09, -6.369635e-09, -7.073973e-09, 
    -7.900526e-09, -8.698924e-09, -9.459138e-09, -1.004859e-08, 
    -1.037361e-08, -1.026961e-08,
  -2.215805e-09, -2.27066e-09, -2.767869e-09, -3.454931e-09, -4.075344e-09, 
    -4.796154e-09, -5.410624e-09, -5.860427e-09, -6.513682e-09, 
    -7.258214e-09, -8.041094e-09, -8.777499e-09, -9.484228e-09, 
    -9.855102e-09, -9.878285e-09,
  -2.080568e-09, -2.107036e-09, -2.413831e-09, -3.047468e-09, -3.664994e-09, 
    -4.367656e-09, -5.020271e-09, -5.630092e-09, -6.091183e-09, 
    -6.701748e-09, -7.391912e-09, -8.084016e-09, -8.733438e-09, -9.24444e-09, 
    -9.353279e-09,
  -1.799395e-09, -1.986816e-09, -2.142426e-09, -2.691103e-09, -3.261332e-09, 
    -3.966223e-09, -4.633639e-09, -5.262697e-09, -5.772741e-09, 
    -6.291018e-09, -6.904281e-09, -7.551447e-09, -8.116238e-09, 
    -8.596837e-09, -8.81599e-09,
  -1.393665e-09, -1.753597e-09, -1.991348e-09, -2.364274e-09, -2.897335e-09, 
    -3.602233e-09, -4.216052e-09, -4.875182e-09, -5.438623e-09, -5.84314e-09, 
    -6.36732e-09, -6.993834e-09, -7.614005e-09, -8.061677e-09, -8.275101e-09,
  -1.060026e-09, -1.463808e-09, -1.819545e-09, -2.070139e-09, -2.531106e-09, 
    -3.191243e-09, -3.870359e-09, -4.415186e-09, -5.150648e-09, 
    -5.536313e-09, -5.924467e-09, -6.461636e-09, -7.023663e-09, 
    -7.567972e-09, -7.735526e-09,
  -5.2688e-09, -7.10532e-09, -9.573887e-09, -1.148338e-08, -1.348595e-08, 
    -1.51536e-08, -1.581088e-08, -1.650251e-08, -1.752122e-08, -1.865731e-08, 
    -1.959096e-08, -1.982396e-08, -2.016458e-08, -2.049528e-08, -2.071599e-08,
  -3.352627e-09, -4.596733e-09, -6.294762e-09, -8.465459e-09, -1.03418e-08, 
    -1.246502e-08, -1.447313e-08, -1.528179e-08, -1.568946e-08, 
    -1.669314e-08, -1.820124e-08, -1.954281e-08, -2.029316e-08, 
    -2.088202e-08, -2.132678e-08,
  -2.252257e-09, -2.809078e-09, -3.845841e-09, -5.501189e-09, -7.37283e-09, 
    -9.298632e-09, -1.135455e-08, -1.322952e-08, -1.468069e-08, 
    -1.533416e-08, -1.653263e-08, -1.815983e-08, -1.987083e-08, 
    -2.107035e-08, -2.151515e-08,
  -2.072758e-09, -2.087228e-09, -2.506223e-09, -3.428257e-09, -4.852652e-09, 
    -6.476228e-09, -8.261511e-09, -1.009762e-08, -1.196314e-08, 
    -1.365521e-08, -1.491768e-08, -1.643938e-08, -1.802568e-08, 
    -1.890818e-08, -1.882744e-08,
  -1.673577e-09, -1.792705e-09, -1.861055e-09, -2.281703e-09, -3.119818e-09, 
    -4.334431e-09, -5.731491e-09, -7.309773e-09, -8.967079e-09, 
    -1.083027e-08, -1.266065e-08, -1.396143e-08, -1.544607e-08, 
    -1.635283e-08, -1.675805e-08,
  -1.300067e-09, -1.522079e-09, -1.637982e-09, -1.775015e-09, -2.161938e-09, 
    -2.917352e-09, -3.926444e-09, -5.176413e-09, -6.543299e-09, 
    -8.095344e-09, -9.909978e-09, -1.154057e-08, -1.292368e-08, 
    -1.395505e-08, -1.472346e-08,
  -1.032213e-09, -1.203172e-09, -1.413227e-09, -1.561116e-09, -1.721925e-09, 
    -2.098909e-09, -2.743115e-09, -3.613802e-09, -4.691051e-09, 
    -5.932939e-09, -7.434324e-09, -9.015694e-09, -1.061715e-08, 
    -1.204145e-08, -1.317371e-08,
  -9.158707e-10, -9.809914e-10, -1.211588e-09, -1.420382e-09, -1.561601e-09, 
    -1.751083e-09, -2.108438e-09, -2.713874e-09, -3.447256e-09, 
    -4.320934e-09, -5.42608e-09, -6.833196e-09, -8.435176e-09, -1.005499e-08, 
    -1.160613e-08,
  -8.384644e-10, -8.617947e-10, -1.035632e-09, -1.273877e-09, -1.433312e-09, 
    -1.571728e-09, -1.791543e-09, -2.150351e-09, -2.65864e-09, -3.258706e-09, 
    -3.990635e-09, -5.036696e-09, -6.520259e-09, -8.195332e-09, -9.824766e-09,
  -7.297507e-10, -7.598291e-10, -8.839785e-10, -1.1192e-09, -1.30426e-09, 
    -1.445681e-09, -1.61349e-09, -1.867857e-09, -2.154641e-09, -2.614013e-09, 
    -3.218365e-09, -3.995071e-09, -5.163646e-09, -6.722709e-09, -8.25443e-09,
  -1.359299e-08, -1.502319e-08, -1.656676e-08, -1.785092e-08, -1.894959e-08, 
    -1.977134e-08, -2.051552e-08, -2.112621e-08, -2.168578e-08, 
    -2.214238e-08, -2.238104e-08, -2.246593e-08, -2.247497e-08, 
    -2.242484e-08, -2.261662e-08,
  -1.025082e-08, -1.197796e-08, -1.350662e-08, -1.494216e-08, -1.629089e-08, 
    -1.741133e-08, -1.846285e-08, -1.941263e-08, -2.022809e-08, 
    -2.089574e-08, -2.147307e-08, -2.193107e-08, -2.231117e-08, 
    -2.247308e-08, -2.262721e-08,
  -6.742402e-09, -8.472799e-09, -1.020399e-08, -1.17792e-08, -1.328893e-08, 
    -1.464793e-08, -1.590695e-08, -1.692397e-08, -1.787834e-08, 
    -1.875841e-08, -1.946714e-08, -2.015635e-08, -2.067705e-08, 
    -2.110546e-08, -2.146122e-08,
  -3.936867e-09, -5.279666e-09, -6.807471e-09, -8.385703e-09, -1.002334e-08, 
    -1.155033e-08, -1.298571e-08, -1.432036e-08, -1.537478e-08, 
    -1.635132e-08, -1.720481e-08, -1.79102e-08, -1.858002e-08, -1.905119e-08, 
    -1.957446e-08,
  -2.000262e-09, -2.827149e-09, -3.90307e-09, -5.173945e-09, -6.663274e-09, 
    -8.240698e-09, -9.797657e-09, -1.125211e-08, -1.265694e-08, 
    -1.382325e-08, -1.481368e-08, -1.558409e-08, -1.636353e-08, -1.70869e-08, 
    -1.769022e-08,
  -1.15388e-09, -1.451244e-09, -1.921626e-09, -2.651391e-09, -3.703139e-09, 
    -5.022852e-09, -6.521692e-09, -7.992969e-09, -9.520787e-09, 
    -1.088946e-08, -1.226478e-08, -1.326575e-08, -1.415017e-08, 
    -1.495847e-08, -1.577504e-08,
  -1.054404e-09, -1.047598e-09, -1.094626e-09, -1.276261e-09, -1.721328e-09, 
    -2.480572e-09, -3.591202e-09, -4.924197e-09, -6.402992e-09, 
    -7.837748e-09, -9.156983e-09, -1.04862e-08, -1.160524e-08, -1.267445e-08, 
    -1.357729e-08,
  -1.107921e-09, -1.019263e-09, -9.465667e-10, -9.012047e-10, -9.931307e-10, 
    -1.305036e-09, -1.879133e-09, -2.68026e-09, -3.750459e-09, -5.033435e-09, 
    -6.37161e-09, -7.752109e-09, -9.090567e-09, -1.027561e-08, -1.135493e-08,
  -1.234862e-09, -1.153419e-09, -1.073892e-09, -9.793738e-10, -9.549082e-10, 
    -1.01503e-09, -1.221784e-09, -1.594987e-09, -2.11498e-09, -2.839099e-09, 
    -3.855483e-09, -5.110115e-09, -6.353904e-09, -7.672759e-09, -8.943218e-09,
  -1.276233e-09, -1.22205e-09, -1.206925e-09, -1.197263e-09, -1.165335e-09, 
    -1.11007e-09, -1.091487e-09, -1.177457e-09, -1.380091e-09, -1.738556e-09, 
    -2.309847e-09, -3.247202e-09, -4.329999e-09, -5.489067e-09, -6.746725e-09,
  -1.573826e-08, -1.625974e-08, -1.664143e-08, -1.714891e-08, -1.774777e-08, 
    -1.826777e-08, -1.869258e-08, -1.908855e-08, -1.960768e-08, 
    -2.006387e-08, -2.026991e-08, -2.053459e-08, -2.119422e-08, 
    -2.204441e-08, -2.26577e-08,
  -1.493035e-08, -1.564763e-08, -1.628062e-08, -1.668522e-08, -1.717846e-08, 
    -1.773439e-08, -1.838585e-08, -1.909258e-08, -1.974993e-08, 
    -2.019868e-08, -2.076442e-08, -2.121021e-08, -2.147185e-08, 
    -2.185371e-08, -2.210059e-08,
  -1.302439e-08, -1.411801e-08, -1.508929e-08, -1.582888e-08, -1.643026e-08, 
    -1.691306e-08, -1.748906e-08, -1.821421e-08, -1.912738e-08, 
    -1.988177e-08, -2.057315e-08, -2.110132e-08, -2.146741e-08, 
    -2.187735e-08, -2.225873e-08,
  -1.027466e-08, -1.167575e-08, -1.292754e-08, -1.402297e-08, -1.497367e-08, 
    -1.57592e-08, -1.641682e-08, -1.704271e-08, -1.775362e-08, -1.859584e-08, 
    -1.936962e-08, -2.006965e-08, -2.052227e-08, -2.084248e-08, -2.112752e-08,
  -7.025562e-09, -8.579041e-09, -1.004873e-08, -1.134605e-08, -1.253321e-08, 
    -1.363213e-08, -1.455039e-08, -1.541119e-08, -1.614465e-08, 
    -1.686595e-08, -1.75758e-08, -1.817443e-08, -1.869718e-08, -1.902067e-08, 
    -1.931676e-08,
  -4.087396e-09, -5.319745e-09, -6.734834e-09, -8.142004e-09, -9.499686e-09, 
    -1.071894e-08, -1.183226e-08, -1.282128e-08, -1.373774e-08, 
    -1.455625e-08, -1.530412e-08, -1.591777e-08, -1.650073e-08, 
    -1.690357e-08, -1.721341e-08,
  -2.516916e-09, -3.091242e-09, -3.91723e-09, -4.974156e-09, -6.205488e-09, 
    -7.461481e-09, -8.641145e-09, -9.721956e-09, -1.070257e-08, -1.15894e-08, 
    -1.236967e-08, -1.303193e-08, -1.358847e-08, -1.406377e-08, -1.444958e-08,
  -2.082588e-09, -2.26135e-09, -2.535562e-09, -2.983363e-09, -3.604145e-09, 
    -4.416823e-09, -5.360057e-09, -6.353593e-09, -7.306476e-09, 
    -8.191241e-09, -9.012133e-09, -9.720661e-09, -1.034176e-08, 
    -1.089422e-08, -1.138306e-08,
  -1.918403e-09, -1.996148e-09, -2.105152e-09, -2.264418e-09, -2.484088e-09, 
    -2.782675e-09, -3.191189e-09, -3.706735e-09, -4.311836e-09, 
    -4.961314e-09, -5.594146e-09, -6.225236e-09, -6.806994e-09, 
    -7.366299e-09, -7.861606e-09,
  -1.825028e-09, -1.854054e-09, -1.888635e-09, -1.940611e-09, -2.013133e-09, 
    -2.117642e-09, -2.261077e-09, -2.442779e-09, -2.679285e-09, 
    -2.966638e-09, -3.296796e-09, -3.653282e-09, -4.042398e-09, -4.45506e-09, 
    -4.871246e-09,
  -6.231607e-09, -6.810973e-09, -7.53063e-09, -8.253457e-09, -8.901947e-09, 
    -9.491263e-09, -1.00378e-08, -1.063928e-08, -1.119015e-08, -1.171413e-08, 
    -1.212113e-08, -1.258046e-08, -1.303532e-08, -1.341865e-08, -1.37168e-08,
  -5.749278e-09, -6.300422e-09, -6.956041e-09, -7.754403e-09, -8.553399e-09, 
    -9.301154e-09, -9.848661e-09, -1.029007e-08, -1.07022e-08, -1.116531e-08, 
    -1.156363e-08, -1.193172e-08, -1.230002e-08, -1.269175e-08, -1.316146e-08,
  -5.300223e-09, -5.874031e-09, -6.453885e-09, -7.13599e-09, -7.927328e-09, 
    -8.79114e-09, -9.568662e-09, -1.004511e-08, -1.038899e-08, -1.076719e-08, 
    -1.120889e-08, -1.174546e-08, -1.227708e-08, -1.260028e-08, -1.288749e-08,
  -4.683907e-09, -5.345822e-09, -5.964676e-09, -6.65365e-09, -7.385887e-09, 
    -8.167644e-09, -9.011408e-09, -9.790582e-09, -1.029392e-08, 
    -1.056547e-08, -1.077268e-08, -1.11338e-08, -1.174663e-08, -1.24921e-08, 
    -1.31389e-08,
  -3.811102e-09, -4.57908e-09, -5.264547e-09, -5.95778e-09, -6.688886e-09, 
    -7.519235e-09, -8.369736e-09, -9.233534e-09, -1.008406e-08, 
    -1.070475e-08, -1.100619e-08, -1.118754e-08, -1.135882e-08, 
    -1.176048e-08, -1.235102e-08,
  -2.66908e-09, -3.465902e-09, -4.302701e-09, -5.128118e-09, -5.920454e-09, 
    -6.679227e-09, -7.49917e-09, -8.403487e-09, -9.280263e-09, -1.016222e-08, 
    -1.08505e-08, -1.135625e-08, -1.182513e-08, -1.204376e-08, -1.220925e-08,
  -1.921241e-09, -2.294876e-09, -2.965122e-09, -3.783737e-09, -4.742882e-09, 
    -5.664986e-09, -6.524993e-09, -7.381252e-09, -8.261456e-09, 
    -9.092451e-09, -9.865825e-09, -1.056183e-08, -1.114068e-08, -1.17255e-08, 
    -1.21734e-08,
  -1.809677e-09, -1.863921e-09, -2.068084e-09, -2.499901e-09, -3.187128e-09, 
    -4.09934e-09, -5.101198e-09, -6.131175e-09, -7.104794e-09, -8.003556e-09, 
    -8.744843e-09, -9.449821e-09, -1.002655e-08, -1.060043e-08, -1.106843e-08,
  -1.659845e-09, -1.750969e-09, -1.838131e-09, -1.937774e-09, -2.162823e-09, 
    -2.621085e-09, -3.343189e-09, -4.267184e-09, -5.350572e-09, 
    -6.406349e-09, -7.303018e-09, -8.049338e-09, -8.649826e-09, 
    -9.167079e-09, -9.672957e-09,
  -1.456848e-09, -1.567793e-09, -1.693527e-09, -1.792031e-09, -1.841369e-09, 
    -1.933119e-09, -2.206374e-09, -2.780687e-09, -3.558053e-09, 
    -4.539349e-09, -5.46889e-09, -6.304654e-09, -6.981511e-09, -7.49268e-09, 
    -7.94456e-09,
  -4.833491e-09, -5.14933e-09, -5.594266e-09, -6.052946e-09, -6.531638e-09, 
    -7.008353e-09, -7.409788e-09, -7.704958e-09, -7.902619e-09, 
    -8.131045e-09, -8.393128e-09, -8.615928e-09, -8.773191e-09, 
    -8.879639e-09, -8.943306e-09,
  -3.769557e-09, -4.100656e-09, -4.430953e-09, -4.792657e-09, -5.157304e-09, 
    -5.520431e-09, -5.87342e-09, -6.271039e-09, -6.581364e-09, -6.932809e-09, 
    -7.375353e-09, -7.744353e-09, -8.0628e-09, -8.286752e-09, -8.490772e-09,
  -2.974524e-09, -3.197478e-09, -3.45317e-09, -3.755191e-09, -4.048097e-09, 
    -4.338694e-09, -4.625409e-09, -4.981675e-09, -5.385328e-09, -5.79407e-09, 
    -6.27532e-09, -6.735614e-09, -7.168246e-09, -7.60938e-09, -7.981805e-09,
  -2.264047e-09, -2.452908e-09, -2.667398e-09, -2.91644e-09, -3.158838e-09, 
    -3.395308e-09, -3.605869e-09, -3.876409e-09, -4.229402e-09, 
    -4.680593e-09, -5.199107e-09, -5.69029e-09, -6.195352e-09, -6.745136e-09, 
    -7.281986e-09,
  -1.693537e-09, -1.852862e-09, -2.034732e-09, -2.236065e-09, -2.453397e-09, 
    -2.662971e-09, -2.830435e-09, -3.004933e-09, -3.265931e-09, 
    -3.641756e-09, -4.171368e-09, -4.728542e-09, -5.246754e-09, 
    -5.792038e-09, -6.464437e-09,
  -1.355121e-09, -1.425018e-09, -1.548924e-09, -1.69607e-09, -1.838447e-09, 
    -2.002212e-09, -2.140549e-09, -2.263113e-09, -2.435984e-09, 
    -2.733043e-09, -3.198816e-09, -3.775696e-09, -4.365751e-09, 
    -4.978379e-09, -5.630569e-09,
  -1.284189e-09, -1.277492e-09, -1.330982e-09, -1.391295e-09, -1.451954e-09, 
    -1.525093e-09, -1.641453e-09, -1.702678e-09, -1.798088e-09, 
    -2.017002e-09, -2.441883e-09, -2.936648e-09, -3.495408e-09, 
    -4.182046e-09, -4.979597e-09,
  -1.175873e-09, -1.184682e-09, -1.232475e-09, -1.27391e-09, -1.288075e-09, 
    -1.291095e-09, -1.320496e-09, -1.365898e-09, -1.415571e-09, 
    -1.582886e-09, -1.931336e-09, -2.494062e-09, -3.05853e-09, -3.70168e-09, 
    -4.465892e-09,
  -1.022324e-09, -1.042181e-09, -1.098763e-09, -1.146732e-09, -1.208769e-09, 
    -1.24491e-09, -1.254513e-09, -1.244515e-09, -1.251412e-09, -1.367669e-09, 
    -1.626156e-09, -2.130576e-09, -2.764626e-09, -3.44794e-09, -4.146555e-09,
  -1.014359e-09, -1.019967e-09, -1.056339e-09, -1.077868e-09, -1.101778e-09, 
    -1.14771e-09, -1.185233e-09, -1.210338e-09, -1.220149e-09, -1.321394e-09, 
    -1.51092e-09, -1.926484e-09, -2.518268e-09, -3.196221e-09, -3.958891e-09,
  -4.007469e-09, -4.245527e-09, -4.493376e-09, -4.761441e-09, -5.142752e-09, 
    -5.703269e-09, -6.606435e-09, -7.467358e-09, -8.159941e-09, 
    -8.853003e-09, -9.443614e-09, -1.005016e-08, -1.062805e-08, 
    -1.137236e-08, -1.207985e-08,
  -3.828236e-09, -4.047401e-09, -4.312403e-09, -4.554056e-09, -4.815367e-09, 
    -5.214726e-09, -5.731259e-09, -6.70508e-09, -7.570732e-09, -8.304608e-09, 
    -8.991955e-09, -9.677574e-09, -1.032353e-08, -1.100794e-08, -1.179538e-08,
  -3.639385e-09, -3.927502e-09, -4.187041e-09, -4.438312e-09, -4.642511e-09, 
    -4.873326e-09, -5.247856e-09, -5.784384e-09, -6.817747e-09, -7.70108e-09, 
    -8.448293e-09, -9.210092e-09, -9.955225e-09, -1.067135e-08, -1.140662e-08,
  -3.168404e-09, -3.658226e-09, -4.035543e-09, -4.335095e-09, -4.574644e-09, 
    -4.753053e-09, -5.03692e-09, -5.367943e-09, -5.932126e-09, -6.871564e-09, 
    -7.789208e-09, -8.630849e-09, -9.45095e-09, -1.020125e-08, -1.098757e-08,
  -2.744826e-09, -3.190099e-09, -3.72342e-09, -4.166365e-09, -4.516134e-09, 
    -4.745447e-09, -4.976421e-09, -5.245719e-09, -5.592409e-09, 
    -6.170899e-09, -7.068977e-09, -7.945331e-09, -8.822123e-09, 
    -9.599667e-09, -1.039983e-08,
  -2.311962e-09, -2.812269e-09, -3.280982e-09, -3.794256e-09, -4.286656e-09, 
    -4.68987e-09, -5.001088e-09, -5.277841e-09, -5.566478e-09, -5.96401e-09, 
    -6.569455e-09, -7.331384e-09, -8.176574e-09, -8.989631e-09, -9.779487e-09,
  -2.027554e-09, -2.341844e-09, -2.812266e-09, -3.306043e-09, -3.860145e-09, 
    -4.428891e-09, -4.863056e-09, -5.238417e-09, -5.508896e-09, 
    -5.822155e-09, -6.298628e-09, -6.833112e-09, -7.478832e-09, 
    -8.273488e-09, -8.994569e-09,
  -1.848811e-09, -2.018924e-09, -2.297094e-09, -2.736483e-09, -3.272789e-09, 
    -3.895042e-09, -4.490321e-09, -4.942292e-09, -5.369972e-09, 
    -5.612916e-09, -5.973592e-09, -6.405989e-09, -6.843988e-09, 
    -7.439245e-09, -8.020824e-09,
  -1.899968e-09, -1.860368e-09, -1.9755e-09, -2.281997e-09, -2.736427e-09, 
    -3.261992e-09, -3.844437e-09, -4.381425e-09, -4.893651e-09, 
    -5.333856e-09, -5.669571e-09, -5.968286e-09, -6.27562e-09, -6.700075e-09, 
    -7.062048e-09,
  -2.002806e-09, -1.862847e-09, -1.826949e-09, -1.953618e-09, -2.27021e-09, 
    -2.727098e-09, -3.220267e-09, -3.748897e-09, -4.23506e-09, -4.740128e-09, 
    -5.204878e-09, -5.579868e-09, -5.873328e-09, -6.092564e-09, -6.222726e-09,
  -1.020917e-08, -1.078223e-08, -1.138053e-08, -1.187579e-08, -1.218052e-08, 
    -1.241285e-08, -1.260187e-08, -1.266488e-08, -1.267754e-08, 
    -1.249694e-08, -1.226171e-08, -1.197414e-08, -1.168303e-08, 
    -1.135754e-08, -1.093504e-08,
  -9.369174e-09, -9.984271e-09, -1.063691e-08, -1.119342e-08, -1.155614e-08, 
    -1.180104e-08, -1.200378e-08, -1.208736e-08, -1.214166e-08, 
    -1.200018e-08, -1.177319e-08, -1.154783e-08, -1.125879e-08, 
    -1.086877e-08, -1.046518e-08,
  -8.733226e-09, -9.257043e-09, -9.808602e-09, -1.035398e-08, -1.079553e-08, 
    -1.107648e-08, -1.129117e-08, -1.144245e-08, -1.149955e-08, 
    -1.144155e-08, -1.131196e-08, -1.110806e-08, -1.080278e-08, -1.04262e-08, 
    -1.000898e-08,
  -8.023529e-09, -8.534401e-09, -9.053839e-09, -9.619962e-09, -1.009151e-08, 
    -1.045523e-08, -1.071932e-08, -1.083449e-08, -1.096335e-08, 
    -1.101043e-08, -1.097647e-08, -1.088109e-08, -1.066757e-08, -1.02578e-08, 
    -9.783094e-09,
  -7.409736e-09, -7.780719e-09, -8.345163e-09, -8.908396e-09, -9.393803e-09, 
    -9.768568e-09, -1.004471e-08, -1.025618e-08, -1.046261e-08, -1.06359e-08, 
    -1.068389e-08, -1.066605e-08, -1.047699e-08, -1.006629e-08, -9.326802e-09,
  -7.036141e-09, -7.307901e-09, -7.784527e-09, -8.24087e-09, -8.658311e-09, 
    -9.008721e-09, -9.35955e-09, -9.714126e-09, -1.001207e-08, -1.032737e-08, 
    -1.049398e-08, -1.050321e-08, -1.020205e-08, -9.44224e-09, -8.22777e-09,
  -6.610779e-09, -6.904062e-09, -7.292284e-09, -7.658344e-09, -7.961647e-09, 
    -8.296965e-09, -8.717886e-09, -9.191664e-09, -9.623522e-09, 
    -1.003712e-08, -1.020507e-08, -9.992678e-09, -9.451138e-09, 
    -8.212598e-09, -6.586683e-09,
  -6.290346e-09, -6.535825e-09, -6.823154e-09, -7.136728e-09, -7.37842e-09, 
    -7.715721e-09, -8.174342e-09, -8.684627e-09, -9.221548e-09, 
    -9.496243e-09, -9.375664e-09, -8.966841e-09, -7.938866e-09, 
    -6.396078e-09, -4.899804e-09,
  -6.066656e-09, -6.206568e-09, -6.382602e-09, -6.617212e-09, -6.860176e-09, 
    -7.213338e-09, -7.655896e-09, -8.093179e-09, -8.457527e-09, 
    -8.382642e-09, -8.088607e-09, -7.434644e-09, -6.158918e-09, 
    -4.854055e-09, -3.544299e-09,
  -5.918073e-09, -5.965337e-09, -6.039537e-09, -6.173992e-09, -6.394912e-09, 
    -6.612833e-09, -6.946848e-09, -7.184853e-09, -7.206354e-09, 
    -7.024921e-09, -6.57785e-09, -5.703361e-09, -4.600749e-09, -3.442141e-09, 
    -2.600161e-09,
  -1.431653e-09, -1.599525e-09, -1.717507e-09, -1.881648e-09, -2.091031e-09, 
    -2.281828e-09, -2.488766e-09, -2.709323e-09, -2.815602e-09, 
    -2.852904e-09, -2.845294e-09, -2.928567e-09, -3.038474e-09, 
    -3.158855e-09, -3.319924e-09,
  -1.303822e-09, -1.489898e-09, -1.665276e-09, -1.844342e-09, -2.067121e-09, 
    -2.235371e-09, -2.399412e-09, -2.508821e-09, -2.661683e-09, 
    -2.774786e-09, -2.852022e-09, -2.910082e-09, -3.078469e-09, 
    -3.332786e-09, -3.655312e-09,
  -1.259404e-09, -1.421714e-09, -1.656264e-09, -1.870072e-09, -2.034792e-09, 
    -2.219622e-09, -2.336544e-09, -2.399577e-09, -2.505161e-09, 
    -2.645034e-09, -2.771906e-09, -2.995132e-09, -3.387735e-09, 
    -3.950376e-09, -4.589077e-09,
  -1.200978e-09, -1.327985e-09, -1.500379e-09, -1.745266e-09, -1.984475e-09, 
    -2.180363e-09, -2.237845e-09, -2.326829e-09, -2.466169e-09, 
    -2.740872e-09, -3.138284e-09, -3.729986e-09, -4.412591e-09, 
    -5.264648e-09, -5.932462e-09,
  -1.279276e-09, -1.309813e-09, -1.420955e-09, -1.717495e-09, -2.054803e-09, 
    -2.223099e-09, -2.358566e-09, -2.464206e-09, -2.769862e-09, 
    -3.206024e-09, -3.947941e-09, -4.904011e-09, -5.745335e-09, -6.39886e-09, 
    -6.893575e-09,
  -1.376576e-09, -1.377634e-09, -1.515247e-09, -1.838946e-09, -2.162218e-09, 
    -2.408142e-09, -2.617178e-09, -2.797621e-09, -3.3833e-09, -4.242661e-09, 
    -5.170243e-09, -6.122032e-09, -7.066432e-09, -7.848197e-09, -8.848183e-09,
  -1.592836e-09, -1.529467e-09, -1.6861e-09, -2.012197e-09, -2.332395e-09, 
    -2.624788e-09, -2.888356e-09, -3.305063e-09, -4.159924e-09, 
    -5.160022e-09, -6.403519e-09, -7.875857e-09, -9.687147e-09, 
    -1.139133e-08, -1.271573e-08,
  -1.918029e-09, -1.883574e-09, -2.03218e-09, -2.299974e-09, -2.615802e-09, 
    -2.834702e-09, -3.331085e-09, -4.140045e-09, -4.975908e-09, 
    -6.526465e-09, -8.397754e-09, -1.096381e-08, -1.32726e-08, -1.493698e-08, 
    -1.577491e-08,
  -2.309904e-09, -2.30328e-09, -2.454736e-09, -2.610628e-09, -2.848767e-09, 
    -3.369601e-09, -4.077623e-09, -4.734086e-09, -6.211036e-09, 
    -8.239322e-09, -1.140695e-08, -1.441391e-08, -1.688114e-08, 
    -1.820361e-08, -1.584602e-08,
  -2.710281e-09, -2.687477e-09, -2.834019e-09, -3.075622e-09, -3.576022e-09, 
    -3.983806e-09, -4.628737e-09, -5.801458e-09, -7.697844e-09, 
    -1.092276e-08, -1.436016e-08, -1.823363e-08, -2.040018e-08, 
    -1.789013e-08, -1.23888e-08,
  -2.377713e-09, -2.072736e-09, -1.907827e-09, -1.924937e-09, -1.912109e-09, 
    -1.883567e-09, -1.873884e-09, -1.898134e-09, -1.891005e-09, 
    -1.905455e-09, -1.893947e-09, -1.890195e-09, -1.857245e-09, 
    -1.863809e-09, -1.895631e-09,
  -1.738139e-09, -1.775703e-09, -1.97405e-09, -1.929653e-09, -1.769463e-09, 
    -1.651305e-09, -1.493229e-09, -1.356753e-09, -1.230177e-09, 
    -1.225649e-09, -1.19009e-09, -1.286964e-09, -1.429046e-09, -1.653199e-09, 
    -1.868373e-09,
  -1.901715e-09, -2.342865e-09, -2.201461e-09, -1.596172e-09, -1.236103e-09, 
    -1.043046e-09, -8.440472e-10, -7.991759e-10, -7.788841e-10, 
    -8.208624e-10, -9.755873e-10, -1.268578e-09, -1.555952e-09, 
    -1.714033e-09, -1.800218e-09,
  -2.282211e-09, -2.835412e-09, -1.725047e-09, -1.162931e-09, -1.00493e-09, 
    -9.830552e-10, -1.013255e-09, -1.060524e-09, -1.205148e-09, 
    -1.431445e-09, -1.881469e-09, -2.027075e-09, -1.96716e-09, -1.75688e-09, 
    -1.533417e-09,
  -3.297918e-09, -2.788671e-09, -1.469007e-09, -1.280383e-09, -1.395529e-09, 
    -1.398399e-09, -1.540236e-09, -1.613389e-09, -2.120981e-09, 
    -2.644422e-09, -3.153726e-09, -3.030587e-09, -2.588747e-09, -2.14214e-09, 
    -1.907764e-09,
  -3.878843e-09, -2.513073e-09, -1.741193e-09, -1.684432e-09, -1.780204e-09, 
    -1.943067e-09, -2.526354e-09, -3.36672e-09, -4.100663e-09, -3.944375e-09, 
    -4.046236e-09, -3.509242e-09, -2.767893e-09, -2.073528e-09, -1.589597e-09,
  -3.962607e-09, -3.032761e-09, -2.409185e-09, -2.165784e-09, -2.484998e-09, 
    -2.815326e-09, -3.543535e-09, -4.353529e-09, -4.795918e-09, 
    -5.023664e-09, -4.532438e-09, -2.878265e-09, -1.574363e-09, 
    -1.251997e-09, -1.248764e-09,
  -4.372893e-09, -3.801865e-09, -3.21055e-09, -2.931761e-09, -3.044011e-09, 
    -3.643662e-09, -4.177302e-09, -4.532126e-09, -4.213225e-09, 
    -3.747983e-09, -2.644732e-09, -1.789361e-09, -1.424389e-09, 
    -1.948431e-09, -1.617468e-09,
  -4.847245e-09, -4.654255e-09, -4.116087e-09, -3.838586e-09, -4.144655e-09, 
    -4.568083e-09, -4.830397e-09, -5.24259e-09, -4.892478e-09, -3.97141e-09, 
    -2.741971e-09, -2.224353e-09, -2.851658e-09, -2.528438e-09, -2.061796e-09,
  -5.215266e-09, -5.583609e-09, -5.587793e-09, -5.255158e-09, -5.410659e-09, 
    -5.86659e-09, -6.083236e-09, -6.098833e-09, -5.679439e-09, -5.044301e-09, 
    -3.725205e-09, -3.367203e-09, -4.427437e-09, -3.666447e-09, -3.234805e-09,
  -6.711612e-09, -6.618182e-09, -6.412832e-09, -6.191039e-09, -5.982701e-09, 
    -5.761345e-09, -5.500094e-09, -5.231758e-09, -4.946553e-09, 
    -4.661673e-09, -4.332132e-09, -3.978606e-09, -3.595179e-09, 
    -3.219332e-09, -2.897392e-09,
  -6.33572e-09, -6.116945e-09, -6.083322e-09, -6.065343e-09, -5.908951e-09, 
    -5.50962e-09, -5.064107e-09, -4.591028e-09, -4.133671e-09, -3.582918e-09, 
    -3.025054e-09, -2.45365e-09, -1.906035e-09, -1.452233e-09, -1.129647e-09,
  -5.854805e-09, -5.907971e-09, -6.07284e-09, -5.734004e-09, -5.151653e-09, 
    -4.403985e-09, -3.673549e-09, -3.003944e-09, -2.318403e-09, 
    -1.544857e-09, -8.808644e-10, -4.392331e-10, -2.328555e-10, -1.64917e-10, 
    -1.352629e-10,
  -6.289206e-09, -6.567248e-09, -5.934357e-09, -4.894274e-09, -4.210762e-09, 
    -3.577997e-09, -2.794533e-09, -1.729404e-09, -7.710079e-10, 
    -3.027457e-10, -1.73598e-10, -2.133323e-10, -2.727661e-10, -4.319365e-10, 
    -6.518446e-10,
  -6.898638e-09, -6.308154e-09, -5.018375e-09, -4.17297e-09, -3.610093e-09, 
    -2.685494e-09, -1.53692e-09, -7.083394e-10, -1.480305e-10, 8.481596e-11, 
    -8.435181e-11, -4.779064e-10, -9.670772e-10, -1.496676e-09, -2.059519e-09,
  -6.846445e-09, -5.205648e-09, -4.24088e-09, -3.817105e-09, -2.673865e-09, 
    -1.541538e-09, -9.551784e-10, -8.467547e-10, -7.666676e-10, 
    -1.323559e-09, -1.934044e-09, -2.387111e-09, -2.582958e-09, 
    -2.593819e-09, -2.768944e-09,
  -5.654426e-09, -4.510091e-09, -4.396965e-09, -3.172166e-09, -1.798165e-09, 
    -1.158095e-09, -9.888083e-10, -1.264191e-09, -2.416056e-09, 
    -2.857336e-09, -2.283064e-09, -2.04085e-09, -1.710959e-09, -2.610684e-09, 
    -3.705569e-09,
  -5.442876e-09, -4.577904e-09, -3.920617e-09, -2.915115e-09, -1.624947e-09, 
    -1.020141e-09, -7.95138e-10, -1.096188e-09, -1.574462e-09, -1.677638e-09, 
    -1.142662e-09, -1.475235e-09, -3.473022e-09, -5.617904e-09, -5.348586e-09,
  -5.168895e-09, -4.311047e-09, -3.843385e-09, -2.996313e-09, -2.10565e-09, 
    -1.084677e-09, -1.222496e-09, -1.578495e-09, -1.612335e-09, 
    -1.894243e-09, -2.140908e-09, -1.99254e-09, -4.716556e-09, -5.343787e-09, 
    -5.155618e-09,
  -5.528411e-09, -4.625182e-09, -4.145134e-09, -3.985115e-09, -3.881029e-09, 
    -3.283393e-09, -3.618378e-09, -3.187916e-09, -3.316245e-09, 
    -3.520719e-09, -3.289151e-09, -3.027244e-09, -4.726409e-09, 
    -5.726439e-09, -5.296252e-09,
  -2.205517e-09, -2.558084e-09, -2.951225e-09, -3.214981e-09, -3.526754e-09, 
    -3.762283e-09, -4.070399e-09, -4.387362e-09, -4.640718e-09, -4.87937e-09, 
    -5.123423e-09, -5.194277e-09, -5.113688e-09, -4.887637e-09, -4.632914e-09,
  -2.760548e-09, -2.935259e-09, -3.280382e-09, -3.585449e-09, -3.843817e-09, 
    -4.069415e-09, -4.258429e-09, -4.474745e-09, -4.707888e-09, 
    -4.904796e-09, -5.017107e-09, -5.005601e-09, -4.788578e-09, -4.57464e-09, 
    -4.391082e-09,
  -3.641899e-09, -3.894062e-09, -4.089427e-09, -4.322005e-09, -4.483584e-09, 
    -4.588777e-09, -4.706716e-09, -4.882337e-09, -5.073489e-09, 
    -5.215765e-09, -5.158894e-09, -4.926658e-09, -4.644758e-09, -4.39031e-09, 
    -4.186425e-09,
  -4.84503e-09, -4.9422e-09, -5.105453e-09, -5.279704e-09, -5.433773e-09, 
    -5.507365e-09, -5.655653e-09, -5.874013e-09, -5.985979e-09, 
    -5.843767e-09, -5.438284e-09, -5.021573e-09, -4.67091e-09, -4.466333e-09, 
    -4.208641e-09,
  -6.485096e-09, -6.573178e-09, -6.637429e-09, -6.696856e-09, -6.670008e-09, 
    -6.644077e-09, -6.69267e-09, -6.652e-09, -6.38318e-09, -5.914158e-09, 
    -5.486828e-09, -5.119256e-09, -4.94722e-09, -4.731541e-09, -4.588743e-09,
  -7.400097e-09, -7.524327e-09, -7.613511e-09, -7.446333e-09, -7.275319e-09, 
    -7.227833e-09, -7.029904e-09, -6.754088e-09, -6.396971e-09, 
    -5.907046e-09, -5.596887e-09, -5.403198e-09, -5.217572e-09, 
    -5.147955e-09, -5.590237e-09,
  -7.726045e-09, -7.84666e-09, -7.784214e-09, -7.662695e-09, -7.535393e-09, 
    -7.274309e-09, -6.922486e-09, -6.55232e-09, -6.120823e-09, -5.856784e-09, 
    -5.766455e-09, -5.544673e-09, -5.267639e-09, -5.632268e-09, -5.943672e-09,
  -8.060903e-09, -7.956013e-09, -7.888897e-09, -7.681638e-09, -7.442582e-09, 
    -7.028942e-09, -6.699519e-09, -6.23753e-09, -5.97763e-09, -5.853841e-09, 
    -5.854036e-09, -5.544925e-09, -5.566436e-09, -5.95431e-09, -5.864857e-09,
  -8.217727e-09, -7.958188e-09, -7.633066e-09, -7.367612e-09, -6.964082e-09, 
    -6.520264e-09, -6.319687e-09, -6.070154e-09, -5.980522e-09, 
    -6.006977e-09, -5.950859e-09, -5.878654e-09, -6.206022e-09, 
    -5.996114e-09, -6.038432e-09,
  -7.974218e-09, -7.502465e-09, -7.030456e-09, -6.632227e-09, -6.140211e-09, 
    -6.040382e-09, -6.137643e-09, -6.095386e-09, -6.105869e-09, 
    -6.112591e-09, -6.234576e-09, -6.490507e-09, -6.396909e-09, -6.45705e-09, 
    -6.483344e-09,
  -3.369809e-09, -3.605467e-09, -4.007107e-09, -4.483213e-09, -5.065077e-09, 
    -5.742279e-09, -6.688075e-09, -7.949827e-09, -9.617888e-09, 
    -1.124152e-08, -1.265776e-08, -1.418856e-08, -1.528066e-08, 
    -1.584217e-08, -1.575623e-08,
  -2.75733e-09, -2.763561e-09, -2.858097e-09, -3.067745e-09, -3.313071e-09, 
    -3.645489e-09, -4.12446e-09, -4.780585e-09, -5.509879e-09, -6.251821e-09, 
    -7.00014e-09, -7.584098e-09, -8.063305e-09, -8.404237e-09, -8.420417e-09,
  -2.385683e-09, -2.304348e-09, -2.22527e-09, -2.19449e-09, -2.19103e-09, 
    -2.24999e-09, -2.403892e-09, -2.690627e-09, -2.983839e-09, -3.288014e-09, 
    -3.632595e-09, -3.961913e-09, -4.265746e-09, -4.323824e-09, -4.373005e-09,
  -2.35445e-09, -2.205763e-09, -2.076304e-09, -1.97013e-09, -1.892758e-09, 
    -1.886261e-09, -1.934233e-09, -1.951545e-09, -1.98003e-09, -2.01882e-09, 
    -2.171031e-09, -2.464392e-09, -2.627478e-09, -2.794744e-09, -2.988692e-09,
  -2.844815e-09, -2.677119e-09, -2.466192e-09, -2.290282e-09, -2.196044e-09, 
    -2.175166e-09, -2.178723e-09, -2.076368e-09, -2.052025e-09, 
    -1.964783e-09, -2.044071e-09, -2.268731e-09, -2.52217e-09, -2.943361e-09, 
    -3.644783e-09,
  -4.097167e-09, -3.893398e-09, -3.599331e-09, -3.315793e-09, -3.180133e-09, 
    -3.115392e-09, -3.055162e-09, -2.947437e-09, -2.848396e-09, -2.75615e-09, 
    -2.760625e-09, -2.803095e-09, -2.948539e-09, -3.422263e-09, -4.381679e-09,
  -6.00047e-09, -6.034614e-09, -5.968058e-09, -5.786377e-09, -5.523687e-09, 
    -5.31086e-09, -5.058268e-09, -4.783537e-09, -4.534316e-09, -4.306897e-09, 
    -4.11769e-09, -4.018918e-09, -4.084912e-09, -4.278176e-09, -4.780291e-09,
  -7.664125e-09, -7.665949e-09, -7.598965e-09, -7.554834e-09, -7.348796e-09, 
    -7.060662e-09, -6.763407e-09, -6.468898e-09, -6.143951e-09, 
    -5.804056e-09, -5.51399e-09, -5.391444e-09, -5.400998e-09, -5.497098e-09, 
    -5.545046e-09,
  -8.500466e-09, -8.517888e-09, -8.305705e-09, -8.443668e-09, -8.668673e-09, 
    -8.79134e-09, -8.562049e-09, -8.30328e-09, -8.006049e-09, -7.678225e-09, 
    -7.165959e-09, -6.899145e-09, -6.689994e-09, -6.557902e-09, -6.403597e-09,
  -8.569395e-09, -8.696032e-09, -8.878608e-09, -9.289606e-09, -9.569607e-09, 
    -9.392642e-09, -9.093608e-09, -8.671951e-09, -8.481346e-09, 
    -8.413349e-09, -7.874447e-09, -7.773647e-09, -7.652573e-09, 
    -7.560408e-09, -7.266725e-09,
  -3.979462e-09, -4.055889e-09, -4.21388e-09, -4.374989e-09, -4.534664e-09, 
    -4.828166e-09, -5.497318e-09, -6.490153e-09, -7.750375e-09, 
    -8.648817e-09, -1.021732e-08, -1.220319e-08, -1.490342e-08, 
    -1.686704e-08, -1.803029e-08,
  -3.053275e-09, -3.17805e-09, -3.330699e-09, -3.530512e-09, -3.686122e-09, 
    -3.800644e-09, -4.039412e-09, -4.505956e-09, -5.279945e-09, 
    -6.500724e-09, -7.794053e-09, -9.707275e-09, -1.148535e-08, 
    -1.419872e-08, -1.637014e-08,
  -2.897994e-09, -2.915127e-09, -3.013195e-09, -3.198814e-09, -3.423392e-09, 
    -3.566466e-09, -3.557231e-09, -3.624952e-09, -3.914864e-09, 
    -4.551067e-09, -5.34813e-09, -6.797062e-09, -8.657206e-09, -1.069674e-08, 
    -1.321544e-08,
  -2.891971e-09, -2.964157e-09, -3.01608e-09, -3.154022e-09, -3.400962e-09, 
    -3.642594e-09, -3.702526e-09, -3.63119e-09, -3.55607e-09, -3.758655e-09, 
    -4.25267e-09, -4.958141e-09, -5.993109e-09, -7.803348e-09, -9.731021e-09,
  -2.90342e-09, -3.113505e-09, -3.184577e-09, -3.256514e-09, -3.318606e-09, 
    -3.497391e-09, -3.699306e-09, -3.850221e-09, -3.84983e-09, -3.782947e-09, 
    -3.753942e-09, -4.098483e-09, -4.683331e-09, -5.549516e-09, -7.195689e-09,
  -2.75895e-09, -2.955751e-09, -2.9927e-09, -3.170185e-09, -3.243372e-09, 
    -3.295653e-09, -3.438204e-09, -3.70464e-09, -3.92466e-09, -4.188998e-09, 
    -4.144882e-09, -3.962662e-09, -4.068801e-09, -4.494659e-09, -5.327951e-09,
  -2.792928e-09, -2.831196e-09, -2.938097e-09, -3.108691e-09, -3.2166e-09, 
    -3.238884e-09, -3.313747e-09, -3.460663e-09, -3.688807e-09, 
    -3.957647e-09, -4.270999e-09, -4.392492e-09, -4.500108e-09, 
    -4.500428e-09, -4.894452e-09,
  -2.889045e-09, -2.944833e-09, -3.089033e-09, -3.148012e-09, -3.263173e-09, 
    -3.348643e-09, -3.368158e-09, -3.3507e-09, -3.400371e-09, -3.563412e-09, 
    -3.894316e-09, -4.208088e-09, -4.509093e-09, -4.604294e-09, -4.885089e-09,
  -3.241405e-09, -3.371272e-09, -3.530531e-09, -3.642179e-09, -3.636883e-09, 
    -3.5207e-09, -3.536493e-09, -3.465098e-09, -3.439052e-09, -3.366922e-09, 
    -3.474411e-09, -3.683196e-09, -4.016334e-09, -4.324358e-09, -4.475982e-09,
  -3.850461e-09, -4.052606e-09, -4.144867e-09, -4.225752e-09, -5.217067e-09, 
    -5.786704e-09, -5.297325e-09, -4.425682e-09, -3.724174e-09, 
    -3.336623e-09, -3.211432e-09, -3.240966e-09, -3.346554e-09, 
    -3.568893e-09, -3.788747e-09,
  -1.017129e-08, -1.005594e-08, -9.895163e-09, -9.765099e-09, -9.639597e-09, 
    -9.654652e-09, -9.631482e-09, -9.667133e-09, -9.63057e-09, -9.715665e-09, 
    -9.747985e-09, -9.932406e-09, -1.022072e-08, -1.058299e-08, -1.104401e-08,
  -1.01757e-08, -9.998234e-09, -9.901387e-09, -9.799958e-09, -9.74464e-09, 
    -9.675899e-09, -9.584338e-09, -9.483384e-09, -9.458279e-09, 
    -9.439455e-09, -9.51762e-09, -9.665433e-09, -9.965371e-09, -1.026033e-08, 
    -1.049232e-08,
  -9.395319e-09, -9.278041e-09, -9.161754e-09, -9.056293e-09, -8.949602e-09, 
    -8.862552e-09, -8.794638e-09, -8.769323e-09, -8.713106e-09, -8.67421e-09, 
    -8.653212e-09, -8.690305e-09, -8.848514e-09, -9.180075e-09, -9.280389e-09,
  -8.241405e-09, -8.227586e-09, -8.170913e-09, -8.077632e-09, -7.982672e-09, 
    -7.911243e-09, -7.848344e-09, -7.805411e-09, -7.727807e-09, 
    -7.667856e-09, -7.626227e-09, -7.620178e-09, -7.675188e-09, 
    -7.771474e-09, -7.886268e-09,
  -6.539336e-09, -6.590371e-09, -6.596245e-09, -6.563396e-09, -6.550657e-09, 
    -6.534289e-09, -6.528298e-09, -6.528327e-09, -6.538644e-09, 
    -6.499826e-09, -6.444254e-09, -6.356792e-09, -6.277387e-09, 
    -6.186497e-09, -6.175913e-09,
  -5.026561e-09, -5.126342e-09, -5.136999e-09, -5.113616e-09, -5.100707e-09, 
    -5.085917e-09, -5.049212e-09, -5.013058e-09, -4.982619e-09, 
    -4.915414e-09, -4.865488e-09, -4.730845e-09, -4.539301e-09, 
    -4.399614e-09, -4.325698e-09,
  -3.633672e-09, -3.776163e-09, -3.820269e-09, -3.809199e-09, -3.834475e-09, 
    -3.795967e-09, -3.729539e-09, -3.721333e-09, -3.753528e-09, 
    -3.747277e-09, -3.702389e-09, -3.636092e-09, -3.533149e-09, 
    -3.490152e-09, -3.429475e-09,
  -2.967623e-09, -3.053364e-09, -3.043008e-09, -3.007293e-09, -3.016916e-09, 
    -3.047349e-09, -3.07006e-09, -3.123578e-09, -3.158751e-09, -3.166895e-09, 
    -3.117915e-09, -3.117697e-09, -3.084936e-09, -3.058521e-09, -3.035447e-09,
  -2.991021e-09, -2.8986e-09, -2.852469e-09, -2.799768e-09, -2.833309e-09, 
    -2.864687e-09, -2.935242e-09, -3.040766e-09, -3.070666e-09, 
    -3.086909e-09, -3.049973e-09, -3.022523e-09, -2.992765e-09, 
    -3.002803e-09, -3.094524e-09,
  -3.062369e-09, -2.951382e-09, -2.942524e-09, -2.947742e-09, -2.872859e-09, 
    -2.858004e-09, -2.912018e-09, -3.056275e-09, -3.190091e-09, 
    -3.297299e-09, -3.35235e-09, -3.384657e-09, -3.337609e-09, -3.281539e-09, 
    -3.243784e-09,
  -5.109781e-09, -4.958519e-09, -4.842713e-09, -4.744154e-09, -4.674352e-09, 
    -4.712605e-09, -4.941199e-09, -5.22919e-09, -5.588034e-09, -6.081263e-09, 
    -6.533984e-09, -6.889121e-09, -7.18213e-09, -7.390216e-09, -7.55461e-09,
  -5.39614e-09, -5.045277e-09, -4.779597e-09, -4.625258e-09, -4.574193e-09, 
    -4.535732e-09, -4.560761e-09, -4.686632e-09, -4.9072e-09, -5.194358e-09, 
    -5.569969e-09, -5.969135e-09, -6.341138e-09, -6.687836e-09, -7.024669e-09,
  -5.809815e-09, -5.271209e-09, -4.855229e-09, -4.588828e-09, -4.545287e-09, 
    -4.565658e-09, -4.591234e-09, -4.632818e-09, -4.717926e-09, 
    -4.859643e-09, -5.067368e-09, -5.361551e-09, -5.730481e-09, 
    -6.167015e-09, -6.621605e-09,
  -6.516081e-09, -5.873864e-09, -5.336281e-09, -4.980838e-09, -4.804766e-09, 
    -4.788669e-09, -4.812044e-09, -4.887022e-09, -4.973593e-09, 
    -5.084702e-09, -5.238341e-09, -5.454676e-09, -5.785929e-09, 
    -6.193114e-09, -6.67509e-09,
  -7.889513e-09, -7.064458e-09, -6.378797e-09, -5.927736e-09, -5.696733e-09, 
    -5.620001e-09, -5.614047e-09, -5.635803e-09, -5.710367e-09, 
    -5.822238e-09, -5.986413e-09, -6.18969e-09, -6.434816e-09, -6.732897e-09, 
    -7.072544e-09,
  -9.363716e-09, -8.621557e-09, -7.736558e-09, -7.202912e-09, -6.902768e-09, 
    -6.776813e-09, -6.731629e-09, -6.701806e-09, -6.769872e-09, 
    -6.851928e-09, -7.029751e-09, -7.196544e-09, -7.440303e-09, -7.63117e-09, 
    -7.831588e-09,
  -1.050367e-08, -1.009893e-08, -9.366915e-09, -8.804367e-09, -8.548108e-09, 
    -8.506004e-09, -8.429963e-09, -8.298866e-09, -8.179396e-09, 
    -8.110883e-09, -8.112364e-09, -8.147866e-09, -8.139307e-09, 
    -8.178034e-09, -8.177664e-09,
  -9.640899e-09, -1.049968e-08, -1.073418e-08, -1.046327e-08, -1.050902e-08, 
    -1.060123e-08, -1.065384e-08, -1.054446e-08, -1.033695e-08, 
    -1.004732e-08, -9.695323e-09, -9.34687e-09, -9.065559e-09, -8.793462e-09, 
    -8.56415e-09,
  -7.790035e-09, -9.341496e-09, -1.013366e-08, -1.056065e-08, -1.070839e-08, 
    -1.082013e-08, -1.087929e-08, -1.078396e-08, -1.071668e-08, 
    -1.054268e-08, -1.029363e-08, -1.000248e-08, -9.700368e-09, 
    -9.424239e-09, -9.150075e-09,
  -5.572809e-09, -7.67801e-09, -8.816221e-09, -9.442614e-09, -9.713561e-09, 
    -9.839268e-09, -9.553769e-09, -9.336886e-09, -9.217164e-09, 
    -8.986722e-09, -8.696697e-09, -8.443245e-09, -8.195668e-09, 
    -7.993772e-09, -7.857842e-09,
  -6.135902e-09, -6.193425e-09, -6.262692e-09, -6.386092e-09, -6.520854e-09, 
    -6.668913e-09, -6.816643e-09, -6.94922e-09, -7.08949e-09, -7.260119e-09, 
    -7.398264e-09, -7.380803e-09, -7.280585e-09, -7.120116e-09, -6.948337e-09,
  -6.468119e-09, -6.55365e-09, -6.742896e-09, -6.979922e-09, -7.146447e-09, 
    -7.304302e-09, -7.450479e-09, -7.580955e-09, -7.731697e-09, 
    -7.792302e-09, -7.622591e-09, -7.346432e-09, -7.016308e-09, 
    -6.676587e-09, -6.339389e-09,
  -6.797945e-09, -6.987538e-09, -7.188083e-09, -7.388036e-09, -7.463156e-09, 
    -7.576174e-09, -7.640188e-09, -7.744127e-09, -7.734922e-09, 
    -7.497283e-09, -7.118566e-09, -6.712176e-09, -6.264873e-09, 
    -5.831355e-09, -5.41235e-09,
  -7.018929e-09, -7.253706e-09, -7.491844e-09, -7.683947e-09, -7.762798e-09, 
    -7.779791e-09, -7.820769e-09, -7.790585e-09, -7.509085e-09, 
    -7.062412e-09, -6.586075e-09, -6.145807e-09, -5.733585e-09, 
    -5.383432e-09, -5.072661e-09,
  -7.138409e-09, -7.404675e-09, -7.666969e-09, -7.888109e-09, -7.939438e-09, 
    -7.940771e-09, -7.897795e-09, -7.637282e-09, -7.191345e-09, 
    -6.691295e-09, -6.280761e-09, -5.864548e-09, -5.57746e-09, -5.396218e-09, 
    -5.468892e-09,
  -7.073787e-09, -7.463058e-09, -7.795861e-09, -8.056279e-09, -8.086568e-09, 
    -8.047126e-09, -7.931603e-09, -7.491076e-09, -6.987342e-09, 
    -6.520807e-09, -6.229329e-09, -6.084764e-09, -6.124101e-09, 
    -6.357407e-09, -6.753222e-09,
  -6.797237e-09, -7.291601e-09, -7.698385e-09, -7.954142e-09, -8.048353e-09, 
    -7.964183e-09, -7.715722e-09, -7.226973e-09, -6.943802e-09, 
    -6.869322e-09, -7.07309e-09, -7.378699e-09, -7.82032e-09, -8.157961e-09, 
    -8.501584e-09,
  -6.318965e-09, -6.779145e-09, -7.340172e-09, -7.737663e-09, -7.840387e-09, 
    -7.903014e-09, -7.838e-09, -7.982386e-09, -8.402231e-09, -8.940551e-09, 
    -9.378039e-09, -9.80336e-09, -1.011122e-08, -1.035553e-08, -1.040078e-08,
  -5.602611e-09, -5.97526e-09, -6.553808e-09, -7.181174e-09, -7.591766e-09, 
    -7.89788e-09, -8.199785e-09, -8.683821e-09, -9.128249e-09, -9.492104e-09, 
    -9.94497e-09, -1.038087e-08, -1.083911e-08, -1.125665e-08, -1.1156e-08,
  -4.852337e-09, -5.084587e-09, -5.634591e-09, -6.234179e-09, -6.853212e-09, 
    -7.349492e-09, -7.951605e-09, -8.390069e-09, -8.812047e-09, -9.16118e-09, 
    -9.672716e-09, -1.001538e-08, -1.052533e-08, -1.059556e-08, -9.706196e-09,
  -1.790696e-08, -1.878302e-08, -1.9586e-08, -2.092138e-08, -2.189917e-08, 
    -2.231414e-08, -2.182106e-08, -2.105797e-08, -1.974841e-08, 
    -1.788407e-08, -1.601201e-08, -1.42358e-08, -1.234692e-08, -1.082698e-08, 
    -9.594994e-09,
  -1.68639e-08, -1.691149e-08, -1.721214e-08, -1.741547e-08, -1.781258e-08, 
    -1.899531e-08, -1.943639e-08, -1.900643e-08, -1.758702e-08, -1.6015e-08, 
    -1.437544e-08, -1.26586e-08, -1.107124e-08, -9.961491e-09, -8.90991e-09,
  -1.604143e-08, -1.597073e-08, -1.596339e-08, -1.568162e-08, -1.539802e-08, 
    -1.530278e-08, -1.53569e-08, -1.561042e-08, -1.470997e-08, -1.380216e-08, 
    -1.26967e-08, -1.137916e-08, -1.022554e-08, -9.176397e-09, -8.109198e-09,
  -1.516805e-08, -1.518758e-08, -1.499503e-08, -1.486598e-08, -1.43954e-08, 
    -1.370964e-08, -1.316694e-08, -1.273437e-08, -1.225752e-08, 
    -1.195398e-08, -1.118132e-08, -1.036366e-08, -9.435262e-09, 
    -8.546197e-09, -7.707039e-09,
  -1.470904e-08, -1.449389e-08, -1.409844e-08, -1.37749e-08, -1.32316e-08, 
    -1.292768e-08, -1.237613e-08, -1.151749e-08, -1.100353e-08, 
    -1.043693e-08, -9.94693e-09, -9.240751e-09, -8.547677e-09, -7.795141e-09, 
    -7.277531e-09,
  -1.381633e-08, -1.353437e-08, -1.298948e-08, -1.247954e-08, -1.182159e-08, 
    -1.121746e-08, -1.055968e-08, -1.027221e-08, -9.837012e-09, 
    -9.466685e-09, -8.875378e-09, -8.287475e-09, -7.773919e-09, 
    -7.419039e-09, -7.535462e-09,
  -1.161567e-08, -1.12875e-08, -1.085994e-08, -1.041689e-08, -9.951618e-09, 
    -9.441088e-09, -8.970942e-09, -8.714566e-09, -8.614234e-09, 
    -8.262554e-09, -7.917866e-09, -7.665282e-09, -7.502539e-09, 
    -7.417031e-09, -7.798707e-09,
  -8.458956e-09, -8.369667e-09, -8.227276e-09, -8.001878e-09, -7.679592e-09, 
    -7.386738e-09, -7.046372e-09, -6.910834e-09, -6.881135e-09, 
    -6.806429e-09, -7.023875e-09, -7.267052e-09, -7.267734e-09, 
    -7.422615e-09, -7.389747e-09,
  -5.949638e-09, -5.965094e-09, -6.029385e-09, -6.036807e-09, -6.00271e-09, 
    -5.98342e-09, -5.989497e-09, -6.209038e-09, -6.375839e-09, -6.857277e-09, 
    -7.109125e-09, -7.102347e-09, -7.128647e-09, -7.139958e-09, -6.50777e-09,
  -4.976865e-09, -5.131519e-09, -5.222196e-09, -5.357499e-09, -5.398548e-09, 
    -5.605322e-09, -5.821263e-09, -6.226667e-09, -6.540792e-09, 
    -6.956222e-09, -6.980583e-09, -6.908978e-09, -6.826237e-09, 
    -6.369174e-09, -6.037632e-09,
  -5.553356e-09, -5.744724e-09, -5.947235e-09, -6.27544e-09, -6.766705e-09, 
    -7.577636e-09, -8.649361e-09, -9.936537e-09, -1.143066e-08, 
    -1.270903e-08, -1.397986e-08, -1.540193e-08, -1.727222e-08, 
    -1.872451e-08, -2.002096e-08,
  -5.486054e-09, -5.606217e-09, -5.772314e-09, -6.076562e-09, -6.576299e-09, 
    -7.283615e-09, -8.192976e-09, -9.405766e-09, -1.081943e-08, 
    -1.202923e-08, -1.335482e-08, -1.456773e-08, -1.604155e-08, 
    -1.723714e-08, -1.832836e-08,
  -5.489164e-09, -5.624444e-09, -5.72467e-09, -5.9492e-09, -6.363567e-09, 
    -7.076848e-09, -7.760768e-09, -8.614371e-09, -1.005198e-08, 
    -1.112693e-08, -1.235538e-08, -1.352536e-08, -1.462546e-08, 
    -1.574696e-08, -1.678513e-08,
  -5.405075e-09, -5.617379e-09, -5.763737e-09, -5.926482e-09, -6.185544e-09, 
    -6.751873e-09, -7.603632e-09, -8.255722e-09, -9.13892e-09, -1.018701e-08, 
    -1.135812e-08, -1.226376e-08, -1.330406e-08, -1.40521e-08, -1.467962e-08,
  -5.479314e-09, -5.549101e-09, -5.699489e-09, -5.888461e-09, -6.077161e-09, 
    -6.42963e-09, -7.086511e-09, -7.971766e-09, -8.651742e-09, -9.496651e-09, 
    -1.028258e-08, -1.112221e-08, -1.194238e-08, -1.278914e-08, -1.314574e-08,
  -5.713839e-09, -5.798996e-09, -5.840458e-09, -5.861406e-09, -6.106876e-09, 
    -6.378317e-09, -6.681398e-09, -7.490824e-09, -8.201011e-09, 
    -8.979564e-09, -9.840226e-09, -1.049757e-08, -1.109188e-08, 
    -1.158361e-08, -1.138392e-08,
  -6.450406e-09, -6.436596e-09, -6.513332e-09, -6.44194e-09, -6.456932e-09, 
    -6.700128e-09, -6.997992e-09, -7.415866e-09, -8.371196e-09, 
    -9.196789e-09, -9.999889e-09, -1.066201e-08, -1.094063e-08, 
    -1.080683e-08, -1.012885e-08,
  -8.131199e-09, -8.024513e-09, -8.004542e-09, -7.953012e-09, -7.85119e-09, 
    -7.861676e-09, -8.075364e-09, -8.262588e-09, -8.694404e-09, 
    -9.308348e-09, -9.641428e-09, -1.003252e-08, -9.863629e-09, 
    -9.491722e-09, -9.097766e-09,
  -1.011201e-08, -9.833478e-09, -9.83291e-09, -9.873689e-09, -9.642447e-09, 
    -9.549542e-09, -9.378149e-09, -9.48075e-09, -9.176035e-09, -9.253346e-09, 
    -9.058038e-09, -9.047321e-09, -8.801528e-09, -8.615281e-09, -8.336897e-09,
  -1.240769e-08, -1.216062e-08, -1.156724e-08, -1.134211e-08, -1.095958e-08, 
    -1.069573e-08, -1.004105e-08, -9.847366e-09, -9.423079e-09, 
    -9.316926e-09, -9.039973e-09, -8.775933e-09, -8.590738e-09, 
    -8.506872e-09, -8.311157e-09,
  -3.428516e-09, -3.68044e-09, -3.905629e-09, -4.084136e-09, -4.309257e-09, 
    -4.455666e-09, -4.574683e-09, -4.676861e-09, -4.782742e-09, 
    -4.902288e-09, -5.034031e-09, -5.181257e-09, -5.33998e-09, -5.492755e-09, 
    -5.735471e-09,
  -3.222591e-09, -3.49346e-09, -3.726477e-09, -3.927125e-09, -4.116814e-09, 
    -4.246755e-09, -4.345863e-09, -4.460864e-09, -4.574883e-09, 
    -4.699908e-09, -4.862121e-09, -5.029146e-09, -5.21352e-09, -5.339666e-09, 
    -5.569028e-09,
  -2.927778e-09, -3.299236e-09, -3.618776e-09, -3.870884e-09, -4.015418e-09, 
    -4.098886e-09, -4.210864e-09, -4.337684e-09, -4.500059e-09, -4.65441e-09, 
    -4.812432e-09, -4.91244e-09, -5.074903e-09, -5.189476e-09, -5.384657e-09,
  -2.711279e-09, -3.061227e-09, -3.45088e-09, -3.743863e-09, -3.964205e-09, 
    -4.118415e-09, -4.244562e-09, -4.390026e-09, -4.51801e-09, -4.642146e-09, 
    -4.818106e-09, -4.965024e-09, -5.192335e-09, -5.338187e-09, -5.50047e-09,
  -2.709486e-09, -3.063519e-09, -3.458591e-09, -3.757287e-09, -4.039845e-09, 
    -4.306639e-09, -4.539484e-09, -4.682289e-09, -4.820933e-09, 
    -5.003202e-09, -5.155795e-09, -5.280363e-09, -5.384917e-09, -5.49637e-09, 
    -5.617853e-09,
  -2.761311e-09, -3.140678e-09, -3.535084e-09, -3.878678e-09, -4.210118e-09, 
    -4.521643e-09, -4.855535e-09, -5.181323e-09, -5.414893e-09, 
    -5.451732e-09, -5.467116e-09, -5.48805e-09, -5.650333e-09, -5.787872e-09, 
    -5.93569e-09,
  -3.00643e-09, -3.32782e-09, -3.849753e-09, -4.298151e-09, -4.740139e-09, 
    -5.105086e-09, -5.286297e-09, -5.410053e-09, -5.526561e-09, 
    -5.739714e-09, -5.887729e-09, -5.828908e-09, -5.853064e-09, -5.83859e-09, 
    -5.921897e-09,
  -3.378115e-09, -3.761663e-09, -4.207358e-09, -4.7031e-09, -5.04249e-09, 
    -5.311942e-09, -5.59696e-09, -5.817673e-09, -5.927624e-09, -5.991156e-09, 
    -6.068706e-09, -6.032433e-09, -6.031651e-09, -5.984724e-09, -6.03109e-09,
  -3.73847e-09, -4.304954e-09, -4.944837e-09, -5.259119e-09, -5.481443e-09, 
    -5.637628e-09, -5.816611e-09, -5.896482e-09, -5.967597e-09, 
    -6.057674e-09, -6.058188e-09, -6.0463e-09, -6.115031e-09, -6.197959e-09, 
    -6.148605e-09,
  -4.331519e-09, -4.836405e-09, -5.222157e-09, -5.47452e-09, -5.600872e-09, 
    -5.680283e-09, -5.762525e-09, -5.852065e-09, -5.9238e-09, -6.084487e-09, 
    -6.327324e-09, -6.37429e-09, -6.49532e-09, -6.748911e-09, -6.986146e-09,
  -1.816693e-09, -1.877334e-09, -1.915986e-09, -2.003924e-09, -2.120249e-09, 
    -2.282062e-09, -2.424686e-09, -2.65634e-09, -2.91724e-09, -3.160247e-09, 
    -3.360171e-09, -3.585098e-09, -3.802743e-09, -4.028027e-09, -4.242585e-09,
  -1.615539e-09, -1.646091e-09, -1.726979e-09, -1.865989e-09, -2.045955e-09, 
    -2.255619e-09, -2.454259e-09, -2.606051e-09, -2.764844e-09, 
    -2.981236e-09, -3.233767e-09, -3.515098e-09, -3.790002e-09, 
    -3.999049e-09, -4.189252e-09,
  -1.673752e-09, -1.714704e-09, -1.790647e-09, -1.929234e-09, -2.062182e-09, 
    -2.283954e-09, -2.495094e-09, -2.682589e-09, -2.869204e-09, 
    -3.093773e-09, -3.328459e-09, -3.621268e-09, -3.911062e-09, 
    -4.151201e-09, -4.303419e-09,
  -1.571935e-09, -1.668756e-09, -1.796425e-09, -1.950344e-09, -2.19274e-09, 
    -2.380261e-09, -2.583024e-09, -2.78367e-09, -3.00839e-09, -3.290508e-09, 
    -3.554717e-09, -3.775134e-09, -3.958954e-09, -4.167647e-09, -4.341107e-09,
  -1.651698e-09, -1.737625e-09, -1.843184e-09, -2.042651e-09, -2.260891e-09, 
    -2.472515e-09, -2.692192e-09, -2.99387e-09, -3.281573e-09, -3.550518e-09, 
    -3.718796e-09, -3.822248e-09, -3.927433e-09, -4.059792e-09, -4.319602e-09,
  -1.694441e-09, -1.815075e-09, -1.971417e-09, -2.184144e-09, -2.371909e-09, 
    -2.620592e-09, -2.851151e-09, -3.157565e-09, -3.426483e-09, 
    -3.521174e-09, -3.611797e-09, -3.733585e-09, -3.902715e-09, 
    -4.098262e-09, -4.345783e-09,
  -1.835671e-09, -1.97081e-09, -2.143796e-09, -2.306967e-09, -2.478214e-09, 
    -2.693763e-09, -2.967491e-09, -3.189716e-09, -3.419209e-09, 
    -3.593517e-09, -3.718013e-09, -3.840642e-09, -4.010233e-09, 
    -4.305687e-09, -4.685516e-09,
  -2.013383e-09, -2.220225e-09, -2.249381e-09, -2.363751e-09, -2.513855e-09, 
    -2.776611e-09, -3.006787e-09, -3.271013e-09, -3.506506e-09, 
    -3.721324e-09, -3.945048e-09, -4.144946e-09, -4.484638e-09, 
    -4.814053e-09, -5.089579e-09,
  -2.365382e-09, -2.327418e-09, -2.251258e-09, -2.352191e-09, -2.58184e-09, 
    -2.900625e-09, -3.206588e-09, -3.601958e-09, -3.968623e-09, 
    -4.294856e-09, -4.55216e-09, -4.71263e-09, -4.926109e-09, -5.126184e-09, 
    -5.215472e-09,
  -2.517567e-09, -2.349693e-09, -2.303407e-09, -2.45008e-09, -2.80951e-09, 
    -3.342015e-09, -3.749145e-09, -4.211991e-09, -4.548707e-09, 
    -4.720847e-09, -4.889603e-09, -4.963366e-09, -5.068546e-09, 
    -5.072436e-09, -5.07884e-09,
  -3.618884e-09, -3.808668e-09, -3.880859e-09, -3.846748e-09, -3.63013e-09, 
    -3.277702e-09, -2.821162e-09, -2.392894e-09, -2.051667e-09, 
    -1.783597e-09, -1.589561e-09, -1.466042e-09, -1.413928e-09, 
    -1.406684e-09, -1.464304e-09,
  -2.266627e-09, -2.455415e-09, -2.568302e-09, -2.64055e-09, -2.562134e-09, 
    -2.389371e-09, -2.136794e-09, -1.887795e-09, -1.665832e-09, 
    -1.484609e-09, -1.380626e-09, -1.32338e-09, -1.348537e-09, -1.38948e-09, 
    -1.482327e-09,
  -1.734277e-09, -1.830504e-09, -1.893214e-09, -1.950283e-09, -1.932923e-09, 
    -1.85279e-09, -1.737163e-09, -1.617549e-09, -1.480632e-09, -1.397327e-09, 
    -1.355832e-09, -1.370257e-09, -1.394896e-09, -1.475734e-09, -1.614244e-09,
  -1.621368e-09, -1.653438e-09, -1.647124e-09, -1.618511e-09, -1.597346e-09, 
    -1.551213e-09, -1.505047e-09, -1.438254e-09, -1.359089e-09, -1.33469e-09, 
    -1.344335e-09, -1.408546e-09, -1.524579e-09, -1.688308e-09, -1.892667e-09,
  -1.578523e-09, -1.603389e-09, -1.588491e-09, -1.559132e-09, -1.513851e-09, 
    -1.480036e-09, -1.435975e-09, -1.410283e-09, -1.376079e-09, 
    -1.411712e-09, -1.513747e-09, -1.648108e-09, -1.883128e-09, 
    -2.137451e-09, -2.361172e-09,
  -1.531274e-09, -1.547532e-09, -1.53897e-09, -1.522003e-09, -1.501817e-09, 
    -1.448903e-09, -1.421315e-09, -1.389718e-09, -1.469968e-09, 
    -1.594285e-09, -1.784423e-09, -2.004056e-09, -2.300656e-09, -2.67081e-09, 
    -3.070334e-09,
  -1.451783e-09, -1.494639e-09, -1.504221e-09, -1.506192e-09, -1.520098e-09, 
    -1.506287e-09, -1.463328e-09, -1.534779e-09, -1.640212e-09, 
    -1.844599e-09, -2.074735e-09, -2.372963e-09, -2.845686e-09, 
    -3.594011e-09, -4.343487e-09,
  -1.42441e-09, -1.468942e-09, -1.527199e-09, -1.541576e-09, -1.577792e-09, 
    -1.597873e-09, -1.620081e-09, -1.708734e-09, -1.928894e-09, 
    -2.159033e-09, -2.510238e-09, -2.942839e-09, -3.647395e-09, 
    -4.323558e-09, -4.886771e-09,
  -1.566431e-09, -1.575096e-09, -1.578381e-09, -1.631721e-09, -1.651471e-09, 
    -1.740056e-09, -1.807862e-09, -1.979541e-09, -2.249194e-09, 
    -2.578482e-09, -3.022644e-09, -3.617747e-09, -4.356988e-09, -4.94167e-09, 
    -5.113553e-09,
  -1.836283e-09, -1.746937e-09, -1.730127e-09, -1.733966e-09, -1.763189e-09, 
    -1.878981e-09, -2.050027e-09, -2.272541e-09, -2.592377e-09, 
    -2.985481e-09, -3.493595e-09, -4.171941e-09, -4.944519e-09, 
    -5.292391e-09, -5.161665e-09,
  -1.443125e-08, -1.498449e-08, -1.61255e-08, -1.7449e-08, -1.938255e-08, 
    -2.145492e-08, -2.327648e-08, -2.528474e-08, -2.688157e-08, 
    -2.745893e-08, -2.684974e-08, -2.500256e-08, -2.162409e-08, 
    -1.795916e-08, -1.432439e-08,
  -1.418666e-08, -1.50442e-08, -1.591551e-08, -1.724776e-08, -1.866971e-08, 
    -2.036019e-08, -2.265494e-08, -2.412942e-08, -2.561514e-08, 
    -2.576545e-08, -2.505445e-08, -2.339939e-08, -2.028654e-08, 
    -1.706918e-08, -1.342543e-08,
  -1.366983e-08, -1.445669e-08, -1.558542e-08, -1.681019e-08, -1.796469e-08, 
    -1.930897e-08, -2.12587e-08, -2.306915e-08, -2.38351e-08, -2.385303e-08, 
    -2.275351e-08, -2.104937e-08, -1.867027e-08, -1.566497e-08, -1.221089e-08,
  -1.261936e-08, -1.349181e-08, -1.454543e-08, -1.598676e-08, -1.725271e-08, 
    -1.857005e-08, -1.984581e-08, -2.148686e-08, -2.227891e-08, 
    -2.196411e-08, -2.062681e-08, -1.890098e-08, -1.653427e-08, 
    -1.387396e-08, -1.108424e-08,
  -1.220548e-08, -1.259172e-08, -1.350717e-08, -1.480601e-08, -1.606189e-08, 
    -1.752165e-08, -1.846871e-08, -1.952367e-08, -2.029431e-08, 
    -1.978724e-08, -1.850729e-08, -1.72472e-08, -1.495759e-08, -1.261886e-08, 
    -1.000809e-08,
  -1.113779e-08, -1.208271e-08, -1.253101e-08, -1.377414e-08, -1.482407e-08, 
    -1.620781e-08, -1.701278e-08, -1.76139e-08, -1.81298e-08, -1.780338e-08, 
    -1.664879e-08, -1.515131e-08, -1.352769e-08, -1.105245e-08, -8.788029e-09,
  -8.995538e-09, -1.057599e-08, -1.166167e-08, -1.271617e-08, -1.362607e-08, 
    -1.477462e-08, -1.53119e-08, -1.585689e-08, -1.589665e-08, -1.565484e-08, 
    -1.457351e-08, -1.308556e-08, -1.165048e-08, -9.581663e-09, -7.816129e-09,
  -7.286584e-09, -8.645527e-09, -1.017124e-08, -1.140633e-08, -1.220365e-08, 
    -1.328563e-08, -1.386742e-08, -1.445353e-08, -1.428914e-08, 
    -1.377255e-08, -1.274715e-08, -1.143378e-08, -1.012716e-08, 
    -8.233005e-09, -6.894767e-09,
  -5.568533e-09, -6.916958e-09, -8.434625e-09, -9.905619e-09, -1.077551e-08, 
    -1.175884e-08, -1.231124e-08, -1.287248e-08, -1.272661e-08, 
    -1.208595e-08, -1.10824e-08, -1.010941e-08, -8.764029e-09, -7.279022e-09, 
    -6.0229e-09,
  -3.762472e-09, -5.329625e-09, -6.718027e-09, -8.154227e-09, -9.306528e-09, 
    -1.029766e-08, -1.091811e-08, -1.119539e-08, -1.120843e-08, 
    -1.060684e-08, -9.906169e-09, -8.829733e-09, -7.541103e-09, 
    -6.502311e-09, -5.249861e-09,
  -9.991764e-09, -9.660253e-09, -9.058009e-09, -8.484392e-09, -8.136521e-09, 
    -8.107521e-09, -8.342223e-09, -8.700677e-09, -9.570348e-09, 
    -1.187083e-08, -1.627284e-08, -2.369758e-08, -3.086322e-08, 
    -3.558302e-08, -3.21306e-08,
  -9.492567e-09, -9.375243e-09, -8.942211e-09, -8.474767e-09, -8.115374e-09, 
    -8.108799e-09, -8.385737e-09, -8.865911e-09, -9.825966e-09, 
    -1.189654e-08, -1.603505e-08, -2.299035e-08, -3.005583e-08, 
    -3.447996e-08, -3.367799e-08,
  -9.049748e-09, -9.121567e-09, -8.76884e-09, -8.476761e-09, -8.132483e-09, 
    -8.080765e-09, -8.438495e-09, -8.974443e-09, -9.934204e-09, 
    -1.164282e-08, -1.563686e-08, -2.230706e-08, -2.810765e-08, 
    -3.277954e-08, -3.436475e-08,
  -8.772511e-09, -8.848931e-09, -8.595478e-09, -8.438345e-09, -8.151339e-09, 
    -8.039342e-09, -8.334288e-09, -8.922631e-09, -9.93801e-09, -1.124858e-08, 
    -1.498664e-08, -2.133535e-08, -2.546402e-08, -2.973489e-08, -3.34019e-08,
  -8.626814e-09, -8.733181e-09, -8.438578e-09, -8.395928e-09, -8.169962e-09, 
    -7.999075e-09, -8.235267e-09, -8.825869e-09, -9.728735e-09, 
    -1.074743e-08, -1.399094e-08, -1.961266e-08, -2.328575e-08, 
    -2.534553e-08, -2.990088e-08,
  -8.714907e-09, -8.654136e-09, -8.425149e-09, -8.374831e-09, -8.236781e-09, 
    -8.107833e-09, -8.217052e-09, -8.710825e-09, -9.836543e-09, 
    -1.050682e-08, -1.298068e-08, -1.800837e-08, -2.107028e-08, 
    -2.253561e-08, -2.647615e-08,
  -8.986079e-09, -8.769018e-09, -8.469322e-09, -8.378021e-09, -8.245341e-09, 
    -8.127559e-09, -8.213577e-09, -8.735833e-09, -9.767101e-09, 
    -1.046444e-08, -1.238704e-08, -1.622766e-08, -1.892379e-08, 
    -2.058845e-08, -2.261358e-08,
  -9.135291e-09, -9.005205e-09, -8.729269e-09, -8.613643e-09, -8.407651e-09, 
    -8.26154e-09, -8.376105e-09, -8.854339e-09, -9.916471e-09, -1.058189e-08, 
    -1.214177e-08, -1.527889e-08, -1.691637e-08, -1.81737e-08, -2.018116e-08,
  -9.470223e-09, -9.200186e-09, -9.058682e-09, -8.956826e-09, -8.737882e-09, 
    -8.574487e-09, -8.636663e-09, -9.298649e-09, -1.029251e-08, 
    -1.082981e-08, -1.175629e-08, -1.37659e-08, -1.557885e-08, -1.676644e-08, 
    -1.840863e-08,
  -1.014055e-08, -9.627822e-09, -9.394167e-09, -9.447711e-09, -9.205027e-09, 
    -9.128482e-09, -9.576013e-09, -1.012342e-08, -1.061786e-08, 
    -1.099316e-08, -1.185444e-08, -1.376879e-08, -1.54803e-08, -1.667767e-08, 
    -1.752807e-08,
  -8.448399e-09, -1.059505e-08, -1.282331e-08, -1.451479e-08, -1.566419e-08, 
    -1.64249e-08, -1.685781e-08, -1.73408e-08, -1.7387e-08, -1.761857e-08, 
    -1.761355e-08, -1.761121e-08, -1.806343e-08, -2.086216e-08, -2.437399e-08,
  -7.168696e-09, -9.139812e-09, -1.132537e-08, -1.335962e-08, -1.482935e-08, 
    -1.584833e-08, -1.626828e-08, -1.671812e-08, -1.702264e-08, -1.72246e-08, 
    -1.75467e-08, -1.772654e-08, -1.735499e-08, -1.853468e-08, -2.075772e-08,
  -5.846049e-09, -7.836216e-09, -9.834639e-09, -1.196909e-08, -1.376579e-08, 
    -1.503725e-08, -1.58731e-08, -1.610207e-08, -1.652444e-08, -1.678568e-08, 
    -1.699237e-08, -1.710401e-08, -1.697653e-08, -1.70266e-08, -1.802711e-08,
  -5.032381e-09, -6.580783e-09, -8.422784e-09, -1.056541e-08, -1.25456e-08, 
    -1.402368e-08, -1.518503e-08, -1.576751e-08, -1.597359e-08, 
    -1.636704e-08, -1.649577e-08, -1.653436e-08, -1.630031e-08, 
    -1.621278e-08, -1.620154e-08,
  -4.124537e-09, -5.479693e-09, -7.274521e-09, -9.14813e-09, -1.12074e-08, 
    -1.285916e-08, -1.415022e-08, -1.508529e-08, -1.5638e-08, -1.585621e-08, 
    -1.614212e-08, -1.595977e-08, -1.565028e-08, -1.536269e-08, -1.519412e-08,
  -3.257245e-09, -4.497688e-09, -6.172687e-09, -8.043809e-09, -9.904371e-09, 
    -1.165881e-08, -1.30524e-08, -1.41096e-08, -1.490575e-08, -1.543074e-08, 
    -1.566316e-08, -1.561108e-08, -1.51725e-08, -1.47646e-08, -1.435881e-08,
  -2.590273e-09, -3.550705e-09, -5.165421e-09, -7.026313e-09, -8.71061e-09, 
    -1.044908e-08, -1.18542e-08, -1.301728e-08, -1.387756e-08, -1.470887e-08, 
    -1.501367e-08, -1.515833e-08, -1.470668e-08, -1.423754e-08, -1.370044e-08,
  -2.16388e-09, -2.76193e-09, -4.243634e-09, -6.118368e-09, -7.836913e-09, 
    -9.362288e-09, -1.083056e-08, -1.187188e-08, -1.277398e-08, 
    -1.364493e-08, -1.420564e-08, -1.43538e-08, -1.403999e-08, -1.350502e-08, 
    -1.28663e-08,
  -1.864258e-09, -2.233654e-09, -3.448113e-09, -5.201394e-09, -6.936137e-09, 
    -8.397512e-09, -9.861133e-09, -1.089601e-08, -1.173691e-08, 
    -1.258799e-08, -1.315573e-08, -1.341669e-08, -1.309473e-08, 
    -1.253341e-08, -1.182929e-08,
  -1.625191e-09, -1.888766e-09, -2.79709e-09, -4.420719e-09, -6.119123e-09, 
    -7.658842e-09, -9.029385e-09, -1.012198e-08, -1.085521e-08, 
    -1.157913e-08, -1.20167e-08, -1.209531e-08, -1.167904e-08, -1.101866e-08, 
    -1.019642e-08,
  -6.153908e-09, -8.00228e-09, -9.856503e-09, -1.179466e-08, -1.49607e-08, 
    -1.756798e-08, -1.997235e-08, -2.248868e-08, -2.383156e-08, 
    -2.424026e-08, -2.384048e-08, -2.400375e-08, -2.401615e-08, 
    -2.392067e-08, -2.357215e-08,
  -3.94182e-09, -5.7066e-09, -7.748307e-09, -9.661519e-09, -1.168209e-08, 
    -1.448895e-08, -1.724059e-08, -1.969161e-08, -2.186966e-08, 
    -2.341175e-08, -2.381988e-08, -2.393889e-08, -2.401369e-08, -2.41097e-08, 
    -2.413288e-08,
  -3.007191e-09, -3.94139e-09, -5.620212e-09, -7.700284e-09, -9.522781e-09, 
    -1.15776e-08, -1.42868e-08, -1.697139e-08, -1.933766e-08, -2.114602e-08, 
    -2.280255e-08, -2.325314e-08, -2.367519e-08, -2.389157e-08, -2.404119e-08,
  -2.207621e-09, -2.945936e-09, -3.927669e-09, -5.723308e-09, -7.687866e-09, 
    -9.552918e-09, -1.159934e-08, -1.417615e-08, -1.675435e-08, 
    -1.871087e-08, -2.054751e-08, -2.207759e-08, -2.292583e-08, 
    -2.354149e-08, -2.377085e-08,
  -1.819673e-09, -2.284324e-09, -3.010656e-09, -4.162401e-09, -5.839312e-09, 
    -7.7536e-09, -9.746736e-09, -1.178635e-08, -1.425258e-08, -1.634019e-08, 
    -1.817422e-08, -1.99077e-08, -2.143712e-08, -2.255204e-08, -2.311686e-08,
  -1.717279e-09, -1.958092e-09, -2.371425e-09, -3.258341e-09, -4.476858e-09, 
    -6.001238e-09, -7.902652e-09, -9.95075e-09, -1.208703e-08, -1.410789e-08, 
    -1.592102e-08, -1.770195e-08, -1.944737e-08, -2.088351e-08, -2.193695e-08,
  -1.86979e-09, -1.930488e-09, -2.163567e-09, -2.634555e-09, -3.600171e-09, 
    -4.817962e-09, -6.280113e-09, -8.150695e-09, -1.025135e-08, 
    -1.212504e-08, -1.383392e-08, -1.555625e-08, -1.722598e-08, 
    -1.890683e-08, -2.033115e-08,
  -2.084864e-09, -1.992948e-09, -2.165009e-09, -2.476939e-09, -2.997533e-09, 
    -3.951435e-09, -5.162342e-09, -6.670044e-09, -8.51609e-09, -1.041218e-08, 
    -1.214612e-08, -1.37408e-08, -1.522635e-08, -1.673464e-08, -1.814718e-08,
  -2.049393e-09, -2.08933e-09, -2.215381e-09, -2.42892e-09, -2.805315e-09, 
    -3.382174e-09, -4.366711e-09, -5.643171e-09, -7.121511e-09, 
    -8.695951e-09, -1.046711e-08, -1.218307e-08, -1.366328e-08, 
    -1.495608e-08, -1.617197e-08,
  -1.811757e-09, -1.967075e-09, -2.218796e-09, -2.461764e-09, -2.730728e-09, 
    -3.121397e-09, -3.761985e-09, -4.841787e-09, -6.116972e-09, 
    -7.434788e-09, -8.847066e-09, -1.048373e-08, -1.202347e-08, 
    -1.335464e-08, -1.446617e-08,
  -1.19381e-08, -9.84584e-09, -1.14171e-08, -1.265229e-08, -1.436002e-08, 
    -1.576848e-08, -1.663684e-08, -1.759641e-08, -1.856529e-08, 
    -1.887624e-08, -1.910972e-08, -1.949841e-08, -2.024297e-08, 
    -2.118098e-08, -2.170927e-08,
  -1.181945e-08, -1.121449e-08, -1.105572e-08, -1.19309e-08, -1.301822e-08, 
    -1.415223e-08, -1.529981e-08, -1.604684e-08, -1.723678e-08, -1.85839e-08, 
    -1.939194e-08, -1.985912e-08, -2.009614e-08, -2.040001e-08, -2.120844e-08,
  -9.361142e-09, -1.014438e-08, -1.006015e-08, -1.017778e-08, -1.119133e-08, 
    -1.21781e-08, -1.33211e-08, -1.461304e-08, -1.563845e-08, -1.660334e-08, 
    -1.826567e-08, -1.972423e-08, -2.039379e-08, -2.076252e-08, -2.083064e-08,
  -7.23523e-09, -8.337369e-09, -9.352625e-09, -9.269126e-09, -9.563636e-09, 
    -1.047558e-08, -1.139029e-08, -1.272089e-08, -1.440348e-08, 
    -1.547927e-08, -1.691166e-08, -1.811996e-08, -1.984697e-08, 
    -2.086006e-08, -2.141448e-08,
  -4.456212e-09, -5.77691e-09, -7.188841e-09, -8.255105e-09, -8.472468e-09, 
    -9.034675e-09, -9.740293e-09, -1.059365e-08, -1.194674e-08, 
    -1.368601e-08, -1.527529e-08, -1.657191e-08, -1.844536e-08, 
    -2.000976e-08, -2.127159e-08,
  -2.155007e-09, -2.989913e-09, -4.258119e-09, -5.874861e-09, -7.025512e-09, 
    -7.508804e-09, -8.114462e-09, -8.736202e-09, -9.62832e-09, -1.112133e-08, 
    -1.282903e-08, -1.488054e-08, -1.659112e-08, -1.842471e-08, -1.99692e-08,
  -1.132609e-09, -1.44577e-09, -2.070173e-09, -3.150296e-09, -4.706935e-09, 
    -5.927137e-09, -6.654141e-09, -7.12788e-09, -7.621022e-09, -8.759763e-09, 
    -1.016875e-08, -1.188111e-08, -1.378853e-08, -1.604235e-08, -1.806405e-08,
  -9.577272e-10, -9.974376e-10, -1.182221e-09, -1.638083e-09, -2.524257e-09, 
    -3.843812e-09, -5.107776e-09, -6.220421e-09, -6.728726e-09, 
    -7.196795e-09, -8.10005e-09, -9.467819e-09, -1.128842e-08, -1.336442e-08, 
    -1.553737e-08,
  -8.893047e-10, -9.012657e-10, -9.643112e-10, -1.145724e-09, -1.570607e-09, 
    -2.341208e-09, -3.399591e-09, -4.602079e-09, -5.823166e-09, 
    -6.687348e-09, -7.270584e-09, -7.968667e-09, -9.074871e-09, 
    -1.075759e-08, -1.249177e-08,
  -7.862692e-10, -8.135964e-10, -8.552312e-10, -9.53651e-10, -1.158367e-09, 
    -1.537727e-09, -2.129278e-09, -2.988641e-09, -4.212149e-09, 
    -5.530306e-09, -6.543354e-09, -6.984854e-09, -7.523398e-09, 
    -8.958141e-09, -1.076047e-08,
  -4.787968e-09, -5.22556e-09, -5.742345e-09, -6.268619e-09, -6.850534e-09, 
    -7.492499e-09, -8.127329e-09, -8.815598e-09, -9.559706e-09, 
    -1.016853e-08, -1.05353e-08, -1.085882e-08, -1.097351e-08, -1.112263e-08, 
    -1.127575e-08,
  -4.226445e-09, -4.753579e-09, -5.229284e-09, -5.771744e-09, -6.278563e-09, 
    -6.862621e-09, -7.519075e-09, -8.255234e-09, -9.01774e-09, -9.725106e-09, 
    -1.019611e-08, -1.064679e-08, -1.079698e-08, -1.096513e-08, -1.118312e-08,
  -4.155556e-09, -4.541534e-09, -4.924461e-09, -5.362962e-09, -5.852256e-09, 
    -6.383791e-09, -7.01918e-09, -7.708562e-09, -8.456647e-09, -9.182981e-09, 
    -9.745221e-09, -1.026883e-08, -1.051691e-08, -1.07773e-08, -1.092141e-08,
  -4.176167e-09, -4.518919e-09, -4.874568e-09, -5.238903e-09, -5.665659e-09, 
    -6.174059e-09, -6.772743e-09, -7.420113e-09, -8.147044e-09, 
    -8.815136e-09, -9.382465e-09, -9.805913e-09, -1.013557e-08, 
    -1.029262e-08, -1.050946e-08,
  -4.150987e-09, -4.578284e-09, -4.948238e-09, -5.300852e-09, -5.660638e-09, 
    -6.092033e-09, -6.611665e-09, -7.233705e-09, -7.922812e-09, -8.61105e-09, 
    -9.233349e-09, -9.763922e-09, -1.027104e-08, -1.066693e-08, -1.075212e-08,
  -3.85508e-09, -4.308436e-09, -4.780351e-09, -5.247603e-09, -5.695122e-09, 
    -6.152799e-09, -6.693511e-09, -7.182837e-09, -7.735211e-09, 
    -8.280867e-09, -8.844874e-09, -9.432695e-09, -1.002543e-08, 
    -1.061216e-08, -1.110519e-08,
  -3.660486e-09, -4.038823e-09, -4.45054e-09, -4.914908e-09, -5.416611e-09, 
    -5.900602e-09, -6.407348e-09, -6.970466e-09, -7.420259e-09, 
    -7.853567e-09, -8.2174e-09, -8.645118e-09, -9.15428e-09, -9.702402e-09, 
    -1.029191e-08,
  -3.334333e-09, -3.693325e-09, -4.03986e-09, -4.495263e-09, -4.992124e-09, 
    -5.612832e-09, -6.187817e-09, -6.694123e-09, -7.240944e-09, 
    -7.685784e-09, -8.138122e-09, -8.48084e-09, -8.771596e-09, -8.989514e-09, 
    -9.301584e-09,
  -2.943131e-09, -3.27728e-09, -3.557359e-09, -3.959284e-09, -4.382191e-09, 
    -4.88075e-09, -5.494763e-09, -5.975926e-09, -6.574764e-09, -7.158139e-09, 
    -7.745354e-09, -8.14947e-09, -8.445987e-09, -8.558477e-09, -8.804165e-09,
  -2.534142e-09, -2.776515e-09, -3.005288e-09, -3.324656e-09, -3.69188e-09, 
    -4.102325e-09, -4.639636e-09, -5.176876e-09, -5.656399e-09, 
    -6.146988e-09, -6.690593e-09, -7.201971e-09, -7.543919e-09, 
    -7.756995e-09, -8.019126e-09,
  -2.370917e-09, -2.291283e-09, -2.240421e-09, -2.189982e-09, -2.18381e-09, 
    -2.223493e-09, -2.310605e-09, -2.360242e-09, -2.457677e-09, 
    -2.738628e-09, -3.192822e-09, -3.798942e-09, -4.519415e-09, 
    -5.127121e-09, -5.821393e-09,
  -2.220292e-09, -2.127962e-09, -2.049872e-09, -1.995408e-09, -1.956625e-09, 
    -1.937077e-09, -1.947505e-09, -2.002948e-09, -2.05573e-09, -2.216257e-09, 
    -2.612713e-09, -3.049648e-09, -3.655364e-09, -4.217611e-09, -4.805979e-09,
  -2.131711e-09, -2.019749e-09, -1.925745e-09, -1.845721e-09, -1.772257e-09, 
    -1.718765e-09, -1.670955e-09, -1.650376e-09, -1.683733e-09, 
    -1.768625e-09, -2.0402e-09, -2.453469e-09, -2.957912e-09, -3.473435e-09, 
    -3.980055e-09,
  -1.987119e-09, -1.893165e-09, -1.795145e-09, -1.686977e-09, -1.593761e-09, 
    -1.513276e-09, -1.445496e-09, -1.392193e-09, -1.355239e-09, 
    -1.373856e-09, -1.548845e-09, -1.843964e-09, -2.269548e-09, -2.78141e-09, 
    -3.348425e-09,
  -1.846133e-09, -1.756756e-09, -1.675393e-09, -1.575737e-09, -1.474293e-09, 
    -1.381956e-09, -1.300228e-09, -1.246916e-09, -1.207247e-09, 
    -1.181569e-09, -1.275644e-09, -1.490007e-09, -1.820806e-09, 
    -2.255715e-09, -2.78702e-09,
  -1.806804e-09, -1.726204e-09, -1.612418e-09, -1.524956e-09, -1.438005e-09, 
    -1.338526e-09, -1.241903e-09, -1.159223e-09, -1.093199e-09, 
    -1.063124e-09, -1.124756e-09, -1.307771e-09, -1.577842e-09, 
    -1.920395e-09, -2.370488e-09,
  -1.74855e-09, -1.722538e-09, -1.644427e-09, -1.524762e-09, -1.420968e-09, 
    -1.300359e-09, -1.182846e-09, -1.081727e-09, -9.851232e-10, 
    -9.651777e-10, -1.036516e-09, -1.186977e-09, -1.399402e-09, 
    -1.690866e-09, -2.066185e-09,
  -1.623345e-09, -1.69443e-09, -1.693885e-09, -1.608274e-09, -1.458634e-09, 
    -1.291586e-09, -1.122253e-09, -9.825279e-10, -8.875226e-10, 
    -8.616758e-10, -9.171061e-10, -1.050202e-09, -1.242359e-09, 
    -1.526518e-09, -1.891434e-09,
  -1.735295e-09, -1.77228e-09, -1.829637e-09, -1.818744e-09, -1.678257e-09, 
    -1.45776e-09, -1.21072e-09, -9.909582e-10, -8.446126e-10, -7.723227e-10, 
    -8.06203e-10, -9.533486e-10, -1.184737e-09, -1.493491e-09, -1.821796e-09,
  -2.002421e-09, -1.796152e-09, -1.840526e-09, -1.91967e-09, -1.921499e-09, 
    -1.723801e-09, -1.44473e-09, -1.182442e-09, -1.003121e-09, -8.956283e-10, 
    -8.983572e-10, -1.01971e-09, -1.219618e-09, -1.493516e-09, -1.769387e-09,
  -6.172982e-09, -6.995388e-09, -8.073605e-09, -9.547177e-09, -1.137833e-08, 
    -1.258677e-08, -1.267856e-08, -1.250558e-08, -1.283464e-08, 
    -1.290915e-08, -1.327963e-08, -1.334379e-08, -1.323077e-08, 
    -1.316933e-08, -1.309011e-08,
  -4.597492e-09, -5.329693e-09, -6.120112e-09, -7.051109e-09, -8.125924e-09, 
    -9.372334e-09, -1.085463e-08, -1.179932e-08, -1.175016e-08, 
    -1.196026e-08, -1.217636e-08, -1.244927e-08, -1.237941e-08, 
    -1.219575e-08, -1.199119e-08,
  -3.481528e-09, -4.073868e-09, -4.725712e-09, -5.393517e-09, -6.185315e-09, 
    -7.071369e-09, -7.953442e-09, -9.068039e-09, -1.019457e-08, 
    -1.106987e-08, -1.130511e-08, -1.160339e-08, -1.199088e-08, 
    -1.194336e-08, -1.164639e-08,
  -2.018159e-09, -2.756506e-09, -3.416077e-09, -4.082372e-09, -4.724474e-09, 
    -5.39348e-09, -6.097233e-09, -6.948393e-09, -7.840973e-09, -8.775449e-09, 
    -9.729108e-09, -1.038096e-08, -1.086797e-08, -1.120587e-08, -1.127932e-08,
  -7.945382e-10, -1.264093e-09, -1.899327e-09, -2.568121e-09, -3.179729e-09, 
    -3.771104e-09, -4.373635e-09, -4.982597e-09, -5.671371e-09, 
    -6.452304e-09, -7.209582e-09, -8.00134e-09, -8.710009e-09, -9.27792e-09, 
    -9.757632e-09,
  -5.842326e-10, -5.668103e-10, -8.3361e-10, -1.330026e-09, -1.959504e-09, 
    -2.566553e-09, -3.166083e-09, -3.716956e-09, -4.215604e-09, 
    -4.773475e-09, -5.316084e-09, -5.8862e-09, -6.454182e-09, -7.065259e-09, 
    -7.561957e-09,
  -6.600445e-10, -5.397915e-10, -4.585832e-10, -5.716675e-10, -9.362628e-10, 
    -1.494582e-09, -2.073667e-09, -2.63317e-09, -3.12585e-09, -3.544573e-09, 
    -3.860601e-09, -4.17393e-09, -4.496256e-09, -4.792825e-09, -5.076453e-09,
  -7.593239e-10, -7.730465e-10, -7.720343e-10, -6.705765e-10, -6.756945e-10, 
    -8.959119e-10, -1.325547e-09, -1.826297e-09, -2.287776e-09, 
    -2.669764e-09, -2.957501e-09, -3.188352e-09, -3.417276e-09, 
    -3.657487e-09, -3.928267e-09,
  -7.269808e-10, -7.247349e-10, -7.975449e-10, -8.672975e-10, -8.597713e-10, 
    -9.109363e-10, -1.098797e-09, -1.438654e-09, -1.795622e-09, 
    -2.141784e-09, -2.509885e-09, -2.78388e-09, -3.000233e-09, -3.124064e-09, 
    -3.214289e-09,
  -7.574929e-10, -7.56667e-10, -7.727609e-10, -8.244133e-10, -9.012977e-10, 
    -1.041017e-09, -1.183548e-09, -1.346472e-09, -1.592721e-09, 
    -1.895627e-09, -2.216948e-09, -2.470058e-09, -2.643195e-09, 
    -2.752566e-09, -2.800594e-09,
  -5.746826e-09, -7.005165e-09, -9.017711e-09, -1.133595e-08, -1.373115e-08, 
    -1.582017e-08, -1.609633e-08, -1.551713e-08, -1.480618e-08, 
    -1.400169e-08, -1.304277e-08, -1.231251e-08, -1.213437e-08, 
    -1.260013e-08, -1.317096e-08,
  -4.546693e-09, -5.573125e-09, -6.693343e-09, -8.555082e-09, -1.064703e-08, 
    -1.298811e-08, -1.538429e-08, -1.5853e-08, -1.549942e-08, -1.50818e-08, 
    -1.460461e-08, -1.372802e-08, -1.299739e-08, -1.260484e-08, -1.260007e-08,
  -3.473068e-09, -4.517247e-09, -5.435291e-09, -6.479612e-09, -8.169962e-09, 
    -1.02111e-08, -1.249351e-08, -1.485869e-08, -1.570127e-08, -1.517098e-08, 
    -1.495035e-08, -1.458629e-08, -1.395629e-08, -1.340933e-08, -1.303497e-08,
  -2.41937e-09, -3.352417e-09, -4.444619e-09, -5.335445e-09, -6.300019e-09, 
    -7.796994e-09, -9.846035e-09, -1.192639e-08, -1.430837e-08, 
    -1.548295e-08, -1.516458e-08, -1.48588e-08, -1.457632e-08, -1.4042e-08, 
    -1.352267e-08,
  -1.711599e-09, -2.301713e-09, -3.203411e-09, -4.34932e-09, -5.259686e-09, 
    -6.131543e-09, -7.471419e-09, -9.373283e-09, -1.127978e-08, 
    -1.350311e-08, -1.499093e-08, -1.51383e-08, -1.493178e-08, -1.454227e-08, 
    -1.39751e-08,
  -1.462758e-09, -1.727685e-09, -2.210003e-09, -3.083636e-09, -4.25262e-09, 
    -5.184095e-09, -6.011167e-09, -7.22442e-09, -8.836104e-09, -1.064785e-08, 
    -1.252957e-08, -1.419182e-08, -1.496783e-08, -1.503963e-08, -1.461851e-08,
  -1.256654e-09, -1.486063e-09, -1.751166e-09, -2.16825e-09, -2.958692e-09, 
    -4.127569e-09, -5.069569e-09, -5.926233e-09, -7.004009e-09, 
    -8.344773e-09, -9.987134e-09, -1.158758e-08, -1.311923e-08, -1.42799e-08, 
    -1.488338e-08,
  -1.022157e-09, -1.220086e-09, -1.457882e-09, -1.729657e-09, -2.105463e-09, 
    -2.79886e-09, -3.877013e-09, -4.840288e-09, -5.760832e-09, -6.695286e-09, 
    -7.856384e-09, -9.163711e-09, -1.065318e-08, -1.195006e-08, -1.323583e-08,
  -6.782517e-10, -9.617785e-10, -1.175225e-09, -1.407348e-09, -1.675085e-09, 
    -2.015961e-09, -2.66415e-09, -3.566673e-09, -4.584705e-09, -5.477024e-09, 
    -6.391816e-09, -7.250407e-09, -8.281069e-09, -9.39028e-09, -1.057206e-08,
  -3.934773e-10, -6.589024e-10, -9.265538e-10, -1.121642e-09, -1.353035e-09, 
    -1.586461e-09, -1.881703e-09, -2.416159e-09, -3.225554e-09, 
    -4.212056e-09, -5.157948e-09, -6.014225e-09, -6.772964e-09, 
    -7.547637e-09, -8.380785e-09,
  -3.786373e-09, -4.351888e-09, -5.580675e-09, -7.582657e-09, -9.985334e-09, 
    -1.218612e-08, -1.374561e-08, -1.457183e-08, -1.430038e-08, 
    -1.359389e-08, -1.32749e-08, -1.298168e-08, -1.302804e-08, -1.310428e-08, 
    -1.321916e-08,
  -3.091894e-09, -3.504026e-09, -4.105737e-09, -5.293049e-09, -7.106819e-09, 
    -9.478965e-09, -1.178974e-08, -1.353031e-08, -1.46075e-08, -1.467237e-08, 
    -1.414873e-08, -1.382684e-08, -1.348671e-08, -1.338336e-08, -1.339493e-08,
  -2.750067e-09, -2.973527e-09, -3.31258e-09, -3.912076e-09, -4.968217e-09, 
    -6.747928e-09, -9.151841e-09, -1.162166e-08, -1.343129e-08, 
    -1.466884e-08, -1.498385e-08, -1.463754e-08, -1.437261e-08, 
    -1.410671e-08, -1.406245e-08,
  -2.45433e-09, -2.66471e-09, -2.880355e-09, -3.227735e-09, -3.767369e-09, 
    -4.729821e-09, -6.400287e-09, -8.848231e-09, -1.144242e-08, -1.33905e-08, 
    -1.473782e-08, -1.527044e-08, -1.515466e-08, -1.495624e-08, -1.484396e-08,
  -2.009372e-09, -2.309331e-09, -2.52507e-09, -2.775296e-09, -3.167385e-09, 
    -3.685997e-09, -4.597422e-09, -6.193318e-09, -8.619242e-09, 
    -1.127728e-08, -1.334358e-08, -1.476605e-08, -1.542147e-08, 
    -1.551064e-08, -1.560388e-08,
  -1.630807e-09, -1.951828e-09, -2.214005e-09, -2.41717e-09, -2.683397e-09, 
    -3.130566e-09, -3.661453e-09, -4.575678e-09, -6.141886e-09, -8.55793e-09, 
    -1.122035e-08, -1.334801e-08, -1.479184e-08, -1.553241e-08, -1.582094e-08,
  -1.207643e-09, -1.544488e-09, -1.866507e-09, -2.135251e-09, -2.341723e-09, 
    -2.64252e-09, -3.107791e-09, -3.65655e-09, -4.564581e-09, -6.162143e-09, 
    -8.594938e-09, -1.121424e-08, -1.338523e-08, -1.485178e-08, -1.566172e-08,
  -8.362171e-10, -1.164599e-09, -1.489032e-09, -1.84263e-09, -2.130043e-09, 
    -2.348586e-09, -2.68249e-09, -3.175345e-09, -3.732194e-09, -4.641622e-09, 
    -6.280427e-09, -8.656936e-09, -1.125561e-08, -1.342207e-08, -1.486931e-08,
  -5.707898e-10, -7.801881e-10, -1.106475e-09, -1.43246e-09, -1.801091e-09, 
    -2.09555e-09, -2.361336e-09, -2.735186e-09, -3.258647e-09, -3.836166e-09, 
    -4.812205e-09, -6.483523e-09, -8.805598e-09, -1.135504e-08, -1.336133e-08,
  -5.419661e-10, -5.723053e-10, -7.699918e-10, -1.090637e-09, -1.4242e-09, 
    -1.768878e-09, -2.067623e-09, -2.380639e-09, -2.817764e-09, 
    -3.330918e-09, -3.95789e-09, -4.973558e-09, -6.659858e-09, -8.948749e-09, 
    -1.137947e-08,
  -1.102181e-08, -1.225807e-08, -1.19881e-08, -1.180115e-08, -1.167592e-08, 
    -1.251362e-08, -1.331146e-08, -1.394804e-08, -1.443988e-08, 
    -1.509446e-08, -1.603128e-08, -1.705805e-08, -1.800434e-08, 
    -1.828606e-08, -1.838e-08,
  -9.121917e-09, -1.080781e-08, -1.168199e-08, -1.214027e-08, -1.174823e-08, 
    -1.199971e-08, -1.262902e-08, -1.318434e-08, -1.392988e-08, 
    -1.465237e-08, -1.532485e-08, -1.591557e-08, -1.694356e-08, 
    -1.761777e-08, -1.804812e-08,
  -6.834709e-09, -8.930326e-09, -1.073887e-08, -1.149848e-08, -1.174288e-08, 
    -1.189001e-08, -1.232767e-08, -1.29243e-08, -1.328847e-08, -1.408499e-08, 
    -1.495848e-08, -1.553679e-08, -1.611571e-08, -1.689316e-08, -1.743472e-08,
  -4.737856e-09, -6.383508e-09, -8.381727e-09, -1.045963e-08, -1.164629e-08, 
    -1.161752e-08, -1.195929e-08, -1.272313e-08, -1.335493e-08, 
    -1.361264e-08, -1.424708e-08, -1.491108e-08, -1.546135e-08, 
    -1.616026e-08, -1.661787e-08,
  -3.402402e-09, -4.487787e-09, -6.078087e-09, -7.816488e-09, -9.943673e-09, 
    -1.138467e-08, -1.170179e-08, -1.186756e-08, -1.276961e-08, 
    -1.370024e-08, -1.432981e-08, -1.48342e-08, -1.521873e-08, -1.574066e-08, 
    -1.612482e-08,
  -2.922462e-09, -3.365012e-09, -4.364767e-09, -5.668606e-09, -7.419076e-09, 
    -9.317687e-09, -1.09489e-08, -1.180531e-08, -1.222467e-08, -1.272478e-08, 
    -1.362238e-08, -1.473383e-08, -1.539244e-08, -1.574689e-08, -1.589755e-08,
  -2.637533e-09, -2.819514e-09, -3.283671e-09, -4.126426e-09, -5.320385e-09, 
    -7.033513e-09, -8.625725e-09, -1.017031e-08, -1.140557e-08, 
    -1.229603e-08, -1.284608e-08, -1.361409e-08, -1.463699e-08, 
    -1.548087e-08, -1.591703e-08,
  -2.405852e-09, -2.502765e-09, -2.735977e-09, -3.200074e-09, -3.877946e-09, 
    -5.073645e-09, -6.532356e-09, -8.061958e-09, -9.451609e-09, 
    -1.068339e-08, -1.176153e-08, -1.269652e-08, -1.350035e-08, 
    -1.424646e-08, -1.488106e-08,
  -2.056698e-09, -2.266771e-09, -2.373391e-09, -2.649589e-09, -3.063749e-09, 
    -3.727842e-09, -4.724666e-09, -5.885082e-09, -7.1912e-09, -8.523987e-09, 
    -9.747975e-09, -1.089208e-08, -1.187623e-08, -1.285835e-08, -1.355772e-08,
  -1.516997e-09, -1.909757e-09, -2.119773e-09, -2.253596e-09, -2.487384e-09, 
    -2.909464e-09, -3.606647e-09, -4.527152e-09, -5.505099e-09, 
    -6.546749e-09, -7.583996e-09, -8.670906e-09, -9.735914e-09, 
    -1.071091e-08, -1.168998e-08,
  -4.312056e-09, -5.017497e-09, -5.794854e-09, -6.544855e-09, -7.399429e-09, 
    -7.986556e-09, -8.152591e-09, -7.630938e-09, -7.318405e-09, 
    -7.425474e-09, -7.812205e-09, -8.227199e-09, -8.704875e-09, 
    -8.845407e-09, -8.826819e-09,
  -3.855178e-09, -4.457998e-09, -5.235371e-09, -6.100166e-09, -6.903793e-09, 
    -7.677023e-09, -8.392568e-09, -8.17771e-09, -7.644643e-09, -7.408913e-09, 
    -7.651943e-09, -8.061351e-09, -8.421857e-09, -8.833507e-09, -9.057861e-09,
  -3.232867e-09, -4.059444e-09, -4.686906e-09, -5.580361e-09, -6.524506e-09, 
    -7.309986e-09, -8.136013e-09, -8.797262e-09, -8.093047e-09, 
    -7.591876e-09, -7.604317e-09, -8.123305e-09, -8.421346e-09, 
    -8.719702e-09, -9.016832e-09,
  -2.885103e-09, -3.532879e-09, -4.334044e-09, -5.025609e-09, -6.081402e-09, 
    -6.976687e-09, -7.756856e-09, -8.739532e-09, -9.220824e-09, 
    -8.185825e-09, -7.780588e-09, -7.914481e-09, -8.450075e-09, 
    -8.737016e-09, -9.062974e-09,
  -2.720167e-09, -3.177645e-09, -3.917215e-09, -4.656478e-09, -5.524067e-09, 
    -6.665823e-09, -7.493806e-09, -8.353448e-09, -9.38681e-09, -9.465221e-09, 
    -8.411428e-09, -8.438858e-09, -8.554436e-09, -8.909888e-09, -9.255573e-09,
  -2.734752e-09, -3.015525e-09, -3.527255e-09, -4.309889e-09, -5.070677e-09, 
    -6.184401e-09, -7.301653e-09, -8.149975e-09, -9.195992e-09, 
    -1.006125e-08, -9.418883e-09, -8.983015e-09, -9.211988e-09, 
    -9.406901e-09, -9.502958e-09,
  -2.724945e-09, -3.005202e-09, -3.409503e-09, -3.876632e-09, -4.705308e-09, 
    -5.71325e-09, -7.026927e-09, -8.147626e-09, -9.097151e-09, -1.026549e-08, 
    -1.050459e-08, -9.845855e-09, -9.9277e-09, -1.058096e-08, -1.08244e-08,
  -2.520017e-09, -3.047799e-09, -3.382788e-09, -3.732437e-09, -4.227773e-09, 
    -5.182444e-09, -6.607299e-09, -8.008182e-09, -9.13376e-09, -1.01534e-08, 
    -1.107646e-08, -1.104899e-08, -1.091062e-08, -1.128414e-08, -1.196956e-08,
  -2.263002e-09, -2.869864e-09, -3.378486e-09, -3.717561e-09, -4.077567e-09, 
    -4.654223e-09, -5.943456e-09, -7.658053e-09, -9.032227e-09, 
    -1.029207e-08, -1.128029e-08, -1.140788e-08, -1.137426e-08, 
    -1.177573e-08, -1.242782e-08,
  -1.965869e-09, -2.677233e-09, -3.244067e-09, -3.687492e-09, -4.009861e-09, 
    -4.411428e-09, -5.192712e-09, -6.968499e-09, -8.677061e-09, 
    -1.018843e-08, -1.173299e-08, -1.261136e-08, -1.250277e-08, 
    -1.244449e-08, -1.300349e-08,
  -3.115271e-09, -3.596855e-09, -4.047793e-09, -4.428726e-09, -4.848439e-09, 
    -5.351959e-09, -5.920389e-09, -6.522091e-09, -7.022613e-09, -7.44887e-09, 
    -7.807611e-09, -8.068839e-09, -8.280847e-09, -8.37594e-09, -8.394406e-09,
  -2.409025e-09, -2.871896e-09, -3.355446e-09, -3.750439e-09, -4.094199e-09, 
    -4.484424e-09, -4.990625e-09, -5.485322e-09, -6.023602e-09, 
    -6.457848e-09, -6.828158e-09, -7.13582e-09, -7.326588e-09, -7.486989e-09, 
    -7.56898e-09,
  -1.738967e-09, -2.149076e-09, -2.589333e-09, -3.041069e-09, -3.431919e-09, 
    -3.759057e-09, -4.12231e-09, -4.592276e-09, -5.054695e-09, -5.554286e-09, 
    -5.946493e-09, -6.27084e-09, -6.507777e-09, -6.673377e-09, -6.815415e-09,
  -1.080307e-09, -1.468592e-09, -1.892626e-09, -2.323467e-09, -2.708193e-09, 
    -3.087238e-09, -3.437538e-09, -3.797064e-09, -4.220969e-09, 
    -4.692853e-09, -5.121246e-09, -5.482252e-09, -5.769909e-09, 
    -5.984725e-09, -6.159345e-09,
  -7.503516e-10, -1.015662e-09, -1.346626e-09, -1.747672e-09, -2.159082e-09, 
    -2.547555e-09, -2.894677e-09, -3.221873e-09, -3.572228e-09, 
    -3.997062e-09, -4.436879e-09, -4.775486e-09, -5.082415e-09, 
    -5.344734e-09, -5.586723e-09,
  -5.87383e-10, -7.159731e-10, -9.593439e-10, -1.230328e-09, -1.598806e-09, 
    -2.032368e-09, -2.449817e-09, -2.802067e-09, -3.105878e-09, 
    -3.452537e-09, -3.859229e-09, -4.219646e-09, -4.512126e-09, 
    -4.782427e-09, -5.087565e-09,
  -5.819059e-10, -6.21549e-10, -7.45337e-10, -9.46959e-10, -1.160775e-09, 
    -1.539426e-09, -1.987746e-09, -2.421176e-09, -2.769222e-09, 
    -3.061758e-09, -3.405878e-09, -3.723658e-09, -4.092721e-09, 
    -4.388654e-09, -4.767682e-09,
  -5.959402e-10, -6.137562e-10, -6.799262e-10, -7.718396e-10, -9.056556e-10, 
    -1.165368e-09, -1.551636e-09, -2.01048e-09, -2.454781e-09, -2.800718e-09, 
    -3.079448e-09, -3.38446e-09, -3.671887e-09, -4.086301e-09, -4.557994e-09,
  -5.724369e-10, -5.794707e-10, -6.491105e-10, -7.195575e-10, -7.713661e-10, 
    -9.274012e-10, -1.244932e-09, -1.679813e-09, -2.145831e-09, 
    -2.569565e-09, -2.867033e-09, -3.133998e-09, -3.434194e-09, 
    -3.889181e-09, -4.474372e-09,
  -6.694641e-10, -5.692208e-10, -5.829188e-10, -6.354933e-10, -7.019261e-10, 
    -8.125434e-10, -1.073131e-09, -1.47213e-09, -1.931209e-09, -2.357321e-09, 
    -2.666857e-09, -2.926903e-09, -3.25701e-09, -3.830171e-09, -4.429587e-09,
  -1.927982e-09, -2.344432e-09, -2.828146e-09, -3.395572e-09, -3.948337e-09, 
    -4.498726e-09, -5.191476e-09, -6.154864e-09, -7.121905e-09, 
    -8.019209e-09, -8.795271e-09, -9.430472e-09, -9.940117e-09, 
    -1.039355e-08, -1.070328e-08,
  -1.469835e-09, -1.872164e-09, -2.278337e-09, -2.747882e-09, -3.269709e-09, 
    -3.80907e-09, -4.380678e-09, -5.048149e-09, -5.940537e-09, -6.884743e-09, 
    -7.780995e-09, -8.618108e-09, -9.303299e-09, -9.868481e-09, -1.035334e-08,
  -1.086002e-09, -1.461828e-09, -1.873679e-09, -2.276813e-09, -2.723204e-09, 
    -3.198727e-09, -3.711613e-09, -4.276086e-09, -4.897448e-09, 
    -5.743945e-09, -6.625966e-09, -7.512219e-09, -8.362103e-09, 
    -9.102246e-09, -9.700321e-09,
  -7.376482e-10, -1.049186e-09, -1.437731e-09, -1.855623e-09, -2.284724e-09, 
    -2.719487e-09, -3.142257e-09, -3.625374e-09, -4.175598e-09, 
    -4.768004e-09, -5.549641e-09, -6.392664e-09, -7.226214e-09, -8.06202e-09, 
    -8.817387e-09,
  -4.651106e-10, -7.450621e-10, -1.069537e-09, -1.462281e-09, -1.868802e-09, 
    -2.32794e-09, -2.758146e-09, -3.146815e-09, -3.601349e-09, -4.100955e-09, 
    -4.660022e-09, -5.371043e-09, -6.143963e-09, -6.934503e-09, -7.726946e-09,
  -2.702356e-10, -4.784702e-10, -7.725681e-10, -1.112236e-09, -1.497515e-09, 
    -1.911518e-09, -2.387641e-09, -2.815571e-09, -3.184572e-09, 
    -3.592911e-09, -4.049739e-09, -4.580747e-09, -5.210392e-09, 
    -5.911996e-09, -6.667464e-09,
  -2.318115e-10, -3.435443e-10, -5.258944e-10, -8.276803e-10, -1.181416e-09, 
    -1.574716e-09, -2.002194e-09, -2.467964e-09, -2.880662e-09, -3.23274e-09, 
    -3.588442e-09, -3.996936e-09, -4.48949e-09, -5.05951e-09, -5.684794e-09,
  -2.529388e-10, -3.044664e-10, -3.9813e-10, -5.826833e-10, -9.04144e-10, 
    -1.283955e-09, -1.699767e-09, -2.13818e-09, -2.582248e-09, -2.972938e-09, 
    -3.300152e-09, -3.635001e-09, -3.998395e-09, -4.429737e-09, -4.910675e-09,
  -1.453168e-10, -2.305804e-10, -2.996523e-10, -4.284388e-10, -6.58741e-10, 
    -1.011229e-09, -1.402565e-09, -1.848351e-09, -2.29706e-09, -2.728382e-09, 
    -3.043459e-09, -3.356549e-09, -3.657606e-09, -3.977727e-09, -4.333796e-09,
  -9.723495e-12, -7.944662e-11, -1.804554e-10, -2.914368e-10, -4.751257e-10, 
    -7.560789e-10, -1.129067e-09, -1.546456e-09, -1.998322e-09, 
    -2.473265e-09, -2.849238e-09, -3.148249e-09, -3.418835e-09, 
    -3.679314e-09, -3.94046e-09,
  -4.486842e-10, -6.035071e-10, -8.843049e-10, -1.284942e-09, -1.765593e-09, 
    -2.459636e-09, -3.495356e-09, -4.730496e-09, -6.592475e-09, 
    -9.216627e-09, -1.209972e-08, -1.473125e-08, -1.756029e-08, 
    -2.011793e-08, -2.058751e-08,
  -3.466498e-10, -4.542468e-10, -6.123946e-10, -9.017904e-10, -1.325192e-09, 
    -1.832041e-09, -2.548015e-09, -3.486341e-09, -4.761838e-09, 
    -6.542003e-09, -9.013802e-09, -1.17892e-08, -1.430041e-08, -1.680544e-08, 
    -1.920219e-08,
  -3.029583e-10, -3.78931e-10, -4.841767e-10, -6.490138e-10, -9.491065e-10, 
    -1.371605e-09, -1.893549e-09, -2.576624e-09, -3.509206e-09, 
    -4.834564e-09, -6.527966e-09, -8.879625e-09, -1.144277e-08, 
    -1.395925e-08, -1.630761e-08,
  -3.069454e-10, -3.273982e-10, -4.091533e-10, -5.141639e-10, -6.800439e-10, 
    -9.762616e-10, -1.414821e-09, -1.939995e-09, -2.593685e-09, 
    -3.541978e-09, -4.883938e-09, -6.536534e-09, -8.718609e-09, 
    -1.110821e-08, -1.348213e-08,
  -2.723108e-10, -3.180655e-10, -3.586756e-10, -4.397526e-10, -5.442924e-10, 
    -7.241442e-10, -1.038453e-09, -1.476066e-09, -1.991796e-09, 
    -2.649811e-09, -3.61601e-09, -4.989924e-09, -6.586164e-09, -8.654409e-09, 
    -1.082895e-08,
  -2.41512e-10, -2.733905e-10, -3.326187e-10, -3.92194e-10, -4.665519e-10, 
    -5.683198e-10, -7.718771e-10, -1.119355e-09, -1.548491e-09, 
    -2.063006e-09, -2.744897e-09, -3.755302e-09, -5.088265e-09, 
    -6.633222e-09, -8.593742e-09,
  -1.736032e-10, -2.305768e-10, -2.862593e-10, -3.592698e-10, -4.266052e-10, 
    -5.005931e-10, -6.027889e-10, -8.263042e-10, -1.17821e-09, -1.61477e-09, 
    -2.1491e-09, -2.895882e-09, -3.944184e-09, -5.213515e-09, -6.696991e-09,
  -1.526005e-10, -2.072053e-10, -2.487952e-10, -3.137237e-10, -3.946199e-10, 
    -4.69302e-10, -5.386523e-10, -6.668979e-10, -9.000756e-10, -1.237899e-09, 
    -1.692614e-09, -2.228497e-09, -3.040258e-09, -4.120042e-09, -5.319115e-09,
  -1.404514e-10, -1.678808e-10, -2.321069e-10, -2.794035e-10, -3.480677e-10, 
    -4.375096e-10, -5.102541e-10, -5.971679e-10, -7.65262e-10, -1.013357e-09, 
    -1.358468e-09, -1.804244e-09, -2.365569e-09, -3.251075e-09, -4.251433e-09,
  -1.719646e-10, -1.652988e-10, -1.951174e-10, -2.669113e-10, -3.32613e-10, 
    -4.005599e-10, -4.814036e-10, -5.698695e-10, -6.922813e-10, 
    -9.050166e-10, -1.180489e-09, -1.547167e-09, -1.961335e-09, -2.60388e-09, 
    -3.450984e-09,
  -4.141796e-10, -5.013159e-10, -4.189914e-10, -2.778517e-10, -2.52707e-10, 
    -1.819827e-10, -7.637645e-11, -2.40895e-10, -4.836436e-10, -6.89385e-10, 
    -1.097287e-09, -1.856615e-09, -3.030476e-09, -4.444274e-09, -6.150513e-09,
  -4.00953e-10, -4.490718e-10, -4.78069e-10, -3.334159e-10, -2.841752e-10, 
    -2.305393e-10, -1.282221e-10, -8.027899e-11, -2.775138e-10, 
    -5.278952e-10, -8.364477e-10, -1.351204e-09, -2.263072e-09, 
    -3.622785e-09, -5.249565e-09,
  -3.637751e-10, -4.376111e-10, -4.722329e-10, -4.343813e-10, -3.005298e-10, 
    -2.74341e-10, -2.144418e-10, -1.041698e-10, -1.214574e-10, -3.460609e-10, 
    -6.209127e-10, -1.035377e-09, -1.709025e-09, -2.8454e-09, -4.41238e-09,
  -2.665933e-10, -3.845889e-10, -4.897937e-10, -5.233637e-10, -4.28527e-10, 
    -2.916819e-10, -3.026402e-10, -1.291042e-10, -5.298183e-11, 
    -1.427269e-10, -4.03616e-10, -7.429515e-10, -1.317202e-09, -2.199193e-09, 
    -3.637714e-09,
  -1.650109e-10, -2.729489e-10, -4.246613e-10, -5.325477e-10, -5.253648e-10, 
    -4.184601e-10, -3.75268e-10, -2.708143e-10, 2.257179e-11, 1.784961e-11, 
    -1.929704e-10, -5.039101e-10, -9.901464e-10, -1.712423e-09, -2.916101e-09,
  -1.542583e-10, -1.760726e-10, -2.802125e-10, -4.393173e-10, -5.544095e-10, 
    -4.721465e-10, -4.113442e-10, -3.569393e-10, -1.551002e-10, 8.166487e-11, 
    -1.324588e-11, -2.940332e-10, -7.05767e-10, -1.341854e-09, -2.30698e-09,
  -2.256181e-10, -1.764335e-10, -1.939952e-10, -2.972991e-10, -4.48681e-10, 
    -5.187427e-10, -4.301353e-10, -3.870875e-10, -2.483751e-10, 
    -6.774012e-11, -1.273029e-11, -1.472948e-10, -4.681779e-10, 
    -1.030427e-09, -1.88645e-09,
  -2.463676e-10, -1.93143e-10, -1.73598e-10, -2.015689e-10, -3.331141e-10, 
    -4.691658e-10, -4.528961e-10, -4.015665e-10, -3.038005e-10, 
    -1.663344e-10, -1.032544e-10, -1.410435e-10, -3.591388e-10, 
    -7.788445e-10, -1.525151e-09,
  -2.449134e-10, -2.393279e-10, -1.842019e-10, -1.755752e-10, -2.463502e-10, 
    -3.845411e-10, -4.590865e-10, -4.196323e-10, -3.371875e-10, 
    -2.360506e-10, -1.750277e-10, -1.859914e-10, -3.226238e-10, 
    -6.151384e-10, -1.205693e-09,
  -1.873115e-10, -2.74211e-10, -2.025735e-10, -2.028424e-10, -2.39689e-10, 
    -3.33798e-10, -4.271215e-10, -4.498691e-10, -3.603524e-10, -2.814726e-10, 
    -2.367189e-10, -2.186928e-10, -3.278754e-10, -5.226583e-10, -9.562606e-10,
  -2.865421e-10, -3.044857e-10, -3.318418e-10, -3.654432e-10, -4.063702e-10, 
    -4.458189e-10, -4.718967e-10, -4.555001e-10, -4.827888e-10, 
    -5.010799e-10, -4.85402e-10, -4.354141e-10, -3.882128e-10, -3.721737e-10, 
    -3.967147e-10,
  -2.048193e-10, -2.143989e-10, -2.2837e-10, -2.348776e-10, -2.45232e-10, 
    -2.6348e-10, -2.845061e-10, -2.946089e-10, -2.731004e-10, -2.943348e-10, 
    -3.13951e-10, -2.952586e-10, -2.678308e-10, -2.422717e-10, -2.518796e-10,
  -1.622724e-10, -1.604522e-10, -1.662529e-10, -1.673154e-10, -1.704582e-10, 
    -1.705535e-10, -1.848043e-10, -2.171822e-10, -1.900251e-10, -1.76908e-10, 
    -1.701152e-10, -1.665939e-10, -1.761347e-10, -1.481288e-10, -1.76135e-10,
  -1.665063e-10, -1.447202e-10, -1.34312e-10, -1.169768e-10, -1.001753e-10, 
    -1.232889e-10, -1.817538e-10, -2.011506e-10, -2.402349e-10, 
    -2.109184e-10, -1.960261e-10, -1.780611e-10, -1.633728e-10, 
    -1.465965e-10, -1.70519e-10,
  -2.517059e-10, -2.270307e-10, -2.172612e-10, -1.826504e-10, -1.455134e-10, 
    -1.71942e-10, -2.215515e-10, -4.283242e-10, -4.494058e-10, -2.915278e-10, 
    -2.180125e-10, -2.054212e-10, -2.336724e-10, -1.985077e-10, -1.970218e-10,
  -3.953868e-10, -3.421345e-10, -2.836979e-10, -2.819789e-10, -2.774157e-10, 
    -4.487462e-10, -4.855041e-10, -6.387437e-10, -8.545493e-10, 
    -5.943958e-10, -2.755055e-10, -2.501718e-10, -2.905415e-10, -2.76695e-10, 
    -2.465842e-10,
  -5.436588e-10, -4.969087e-10, -3.796765e-10, -3.453689e-10, -5.92686e-10, 
    -6.501652e-10, -4.33924e-10, -4.854273e-10, -7.528321e-10, -7.685798e-10, 
    -3.531663e-10, -2.985011e-10, -2.934595e-10, -2.865321e-10, -2.7492e-10,
  -5.182001e-10, -5.636039e-10, -4.253705e-10, -4.215335e-10, -6.71236e-10, 
    -6.847278e-10, -4.838591e-10, -4.263064e-10, -5.04567e-10, -8.160711e-10, 
    -5.091387e-10, -3.023446e-10, -2.904108e-10, -2.555111e-10, -2.389463e-10,
  -5.975486e-10, -5.90882e-10, -4.719589e-10, -4.014523e-10, -5.824499e-10, 
    -4.561579e-10, -3.640047e-10, -2.42318e-10, -3.196539e-10, -6.780103e-10, 
    -6.134477e-10, -3.524607e-10, -2.606025e-10, -2.109333e-10, -2.101611e-10,
  -6.988601e-10, -4.511178e-10, -3.354043e-10, -4.214237e-10, -4.923451e-10, 
    -4.904604e-10, -4.52056e-10, -3.28816e-10, -2.697352e-10, -5.758998e-10, 
    -6.863963e-10, -3.590064e-10, -2.431906e-10, -1.760524e-10, -1.980068e-10,
  -2.234349e-09, -2.549474e-09, -2.833591e-09, -3.192156e-09, -3.544324e-09, 
    -3.912178e-09, -4.215796e-09, -4.521192e-09, -4.879376e-09, 
    -5.351637e-09, -5.844656e-09, -6.336342e-09, -6.751868e-09, 
    -7.110411e-09, -7.395217e-09,
  -1.480564e-09, -1.868624e-09, -2.171643e-09, -2.416866e-09, -2.671286e-09, 
    -2.98081e-09, -3.312816e-09, -3.664849e-09, -3.95481e-09, -4.240287e-09, 
    -4.55029e-09, -4.859917e-09, -5.171261e-09, -5.469928e-09, -5.696193e-09,
  -7.790436e-10, -1.01164e-09, -1.356891e-09, -1.694448e-09, -1.9741e-09, 
    -2.225139e-09, -2.490257e-09, -2.789856e-09, -3.098738e-09, -3.39439e-09, 
    -3.623278e-09, -3.83077e-09, -4.013986e-09, -4.171986e-09, -4.305445e-09,
  -4.715484e-10, -5.291447e-10, -6.475213e-10, -8.497815e-10, -1.147899e-09, 
    -1.436297e-09, -1.712118e-09, -1.967969e-09, -2.239346e-09, 
    -2.543802e-09, -2.821707e-09, -3.052651e-09, -3.223682e-09, 
    -3.346139e-09, -3.41546e-09,
  -3.036561e-10, -3.061324e-10, -3.477884e-10, -4.143354e-10, -5.273735e-10, 
    -7.342418e-10, -9.684937e-10, -1.217211e-09, -1.439597e-09, 
    -1.652189e-09, -1.905107e-09, -2.183301e-09, -2.440905e-09, 
    -2.638693e-09, -2.761417e-09,
  -2.399992e-10, -2.034934e-10, -1.931295e-10, -2.207101e-10, -2.617921e-10, 
    -3.383145e-10, -4.710052e-10, -6.471614e-10, -8.794143e-10, 
    -1.081006e-09, -1.252377e-09, -1.390631e-09, -1.535828e-09, -1.7246e-09, 
    -1.91583e-09,
  -6.430164e-10, -5.148652e-10, -4.161601e-10, -3.139631e-10, -2.464647e-10, 
    -2.125413e-10, -2.257108e-10, -2.818068e-10, -3.780878e-10, 
    -5.400203e-10, -6.827715e-10, -9.178665e-10, -1.075257e-09, 
    -1.153448e-09, -1.263555e-09,
  -9.095764e-10, -8.383964e-10, -7.869793e-10, -6.739138e-10, -5.434302e-10, 
    -4.37063e-10, -3.894309e-10, -3.414427e-10, -3.279819e-10, -3.307959e-10, 
    -3.679438e-10, -4.757177e-10, -6.806749e-10, -8.414981e-10, -9.46857e-10,
  -1.056708e-09, -1.032865e-09, -1.001005e-09, -9.468462e-10, -9.053209e-10, 
    -8.352813e-10, -7.563253e-10, -6.846099e-10, -5.512537e-10, 
    -3.905447e-10, -2.899802e-10, -2.603694e-10, -3.222114e-10, 
    -4.401036e-10, -5.765174e-10,
  -1.07364e-09, -9.478145e-10, -8.531522e-10, -6.661707e-10, -5.476607e-10, 
    -4.707449e-10, -3.856133e-10, -4.075288e-10, -4.967405e-10, 
    -4.566688e-10, -4.114345e-10, -2.874009e-10, -2.167133e-10, 
    -2.183924e-10, -2.609885e-10,
  -4.443464e-09, -5.033637e-09, -5.887538e-09, -6.693072e-09, -7.290193e-09, 
    -8.04355e-09, -8.605899e-09, -8.959591e-09, -9.25708e-09, -9.538088e-09, 
    -9.860508e-09, -1.01761e-08, -1.044357e-08, -1.059363e-08, -1.069252e-08,
  -3.827811e-09, -4.083266e-09, -4.500073e-09, -5.232672e-09, -6.03903e-09, 
    -6.721852e-09, -7.252927e-09, -7.792343e-09, -8.25737e-09, -8.70376e-09, 
    -9.085406e-09, -9.474181e-09, -9.801544e-09, -1.009067e-08, -1.034349e-08,
  -3.284714e-09, -3.525537e-09, -3.754268e-09, -4.050665e-09, -4.527863e-09, 
    -5.237666e-09, -5.985743e-09, -6.59532e-09, -7.080032e-09, -7.524395e-09, 
    -7.938052e-09, -8.305599e-09, -8.7051e-09, -9.077685e-09, -9.437497e-09,
  -2.330133e-09, -2.908366e-09, -3.227338e-09, -3.462763e-09, -3.711176e-09, 
    -4.028021e-09, -4.468892e-09, -5.072128e-09, -5.681616e-09, 
    -6.234258e-09, -6.646272e-09, -7.046995e-09, -7.396558e-09, 
    -7.750658e-09, -8.107419e-09,
  -1.224343e-09, -1.810966e-09, -2.417686e-09, -2.859257e-09, -3.137581e-09, 
    -3.385368e-09, -3.6549e-09, -3.958702e-09, -4.33957e-09, -4.814227e-09, 
    -5.27926e-09, -5.690129e-09, -6.041338e-09, -6.335187e-09, -6.62124e-09,
  -6.72235e-10, -9.077264e-10, -1.342353e-09, -1.84198e-09, -2.337238e-09, 
    -2.657286e-09, -2.927322e-09, -3.18813e-09, -3.432284e-09, -3.705176e-09, 
    -4.024668e-09, -4.379932e-09, -4.72546e-09, -5.028171e-09, -5.28437e-09,
  -4.090444e-10, -5.215502e-10, -7.203049e-10, -1.00395e-09, -1.389837e-09, 
    -1.767562e-09, -2.091008e-09, -2.378565e-09, -2.658814e-09, 
    -2.906515e-09, -3.11903e-09, -3.3492e-09, -3.599786e-09, -3.858867e-09, 
    -4.114124e-09,
  -4.069605e-10, -4.47292e-10, -5.313516e-10, -6.838085e-10, -9.028736e-10, 
    -1.134615e-09, -1.34175e-09, -1.558989e-09, -1.796081e-09, -2.03069e-09, 
    -2.236678e-09, -2.408773e-09, -2.580639e-09, -2.731363e-09, -2.901204e-09,
  -6.508137e-10, -6.050205e-10, -6.196239e-10, -6.360724e-10, -7.162008e-10, 
    -8.197085e-10, -9.368988e-10, -1.053842e-09, -1.210675e-09, 
    -1.397216e-09, -1.595879e-09, -1.769186e-09, -1.888056e-09, 
    -1.983805e-09, -2.084569e-09,
  -1.050153e-09, -9.097341e-10, -8.147221e-10, -7.501231e-10, -7.111476e-10, 
    -7.082535e-10, -7.414193e-10, -7.900411e-10, -8.692412e-10, 
    -9.528599e-10, -1.052001e-09, -1.138457e-09, -1.207906e-09, 
    -1.254702e-09, -1.300971e-09,
  -4.473617e-09, -5.464252e-09, -6.543513e-09, -7.474837e-09, -8.395848e-09, 
    -9.255031e-09, -9.854376e-09, -1.003568e-08, -9.879788e-09, 
    -9.519894e-09, -9.279339e-09, -9.07292e-09, -8.989673e-09, -9.068923e-09, 
    -9.251975e-09,
  -4.058655e-09, -4.404977e-09, -5.340806e-09, -6.433269e-09, -7.384425e-09, 
    -8.253807e-09, -9.094112e-09, -9.740629e-09, -1.003121e-08, 
    -9.803607e-09, -9.442636e-09, -9.035166e-09, -8.815647e-09, 
    -8.671091e-09, -8.655828e-09,
  -3.900916e-09, -4.023072e-09, -4.335305e-09, -5.131776e-09, -6.215734e-09, 
    -7.302978e-09, -8.163799e-09, -9.004487e-09, -9.635395e-09, 
    -9.951465e-09, -9.839298e-09, -9.41426e-09, -8.865221e-09, -8.540504e-09, 
    -8.3666e-09,
  -3.509028e-09, -3.772501e-09, -3.992676e-09, -4.332021e-09, -4.95713e-09, 
    -6.011015e-09, -7.080244e-09, -8.008429e-09, -8.98331e-09, -9.625543e-09, 
    -1.001695e-08, -1.006968e-08, -9.709447e-09, -9.09233e-09, -8.54391e-09,
  -3.087874e-09, -3.322332e-09, -3.628635e-09, -3.923565e-09, -4.268059e-09, 
    -4.793445e-09, -5.752718e-09, -6.720499e-09, -7.691201e-09, 
    -8.637315e-09, -9.416814e-09, -9.955365e-09, -1.012947e-08, 
    -9.931224e-09, -9.400812e-09,
  -2.410566e-09, -2.79862e-09, -3.127827e-09, -3.438614e-09, -3.7635e-09, 
    -4.156948e-09, -4.662007e-09, -5.504344e-09, -6.309326e-09, 
    -7.323544e-09, -8.121712e-09, -8.993491e-09, -9.689992e-09, 
    -1.005205e-08, -1.009389e-08,
  -1.679464e-09, -2.110648e-09, -2.494378e-09, -2.851391e-09, -3.152724e-09, 
    -3.483473e-09, -3.831746e-09, -4.333637e-09, -4.98885e-09, -5.749469e-09, 
    -6.663128e-09, -7.420752e-09, -8.219801e-09, -8.866644e-09, -9.394609e-09,
  -1.216449e-09, -1.384734e-09, -1.677164e-09, -2.083236e-09, -2.424201e-09, 
    -2.804807e-09, -3.15224e-09, -3.528895e-09, -3.957168e-09, -4.463411e-09, 
    -5.096849e-09, -5.846272e-09, -6.586697e-09, -7.326476e-09, -7.853948e-09,
  -1.075757e-09, -1.142917e-09, -1.255741e-09, -1.458865e-09, -1.661225e-09, 
    -1.940197e-09, -2.249287e-09, -2.589364e-09, -2.969292e-09, 
    -3.385241e-09, -3.844371e-09, -4.393195e-09, -4.963056e-09, 
    -5.550693e-09, -6.149857e-09,
  -1.136265e-09, -1.101084e-09, -1.157553e-09, -1.253923e-09, -1.411945e-09, 
    -1.541459e-09, -1.729815e-09, -1.932644e-09, -2.154482e-09, 
    -2.407344e-09, -2.727872e-09, -3.105616e-09, -3.590987e-09, 
    -4.120193e-09, -4.671359e-09,
  -6.405181e-09, -7.615673e-09, -8.631951e-09, -9.501609e-09, -1.005634e-08, 
    -1.058596e-08, -1.109885e-08, -1.1529e-08, -1.16846e-08, -1.122538e-08, 
    -1.059561e-08, -1.018968e-08, -9.976015e-09, -9.795254e-09, -9.667024e-09,
  -4.942902e-09, -6.249764e-09, -7.446304e-09, -8.396988e-09, -9.218973e-09, 
    -9.878682e-09, -1.044009e-08, -1.102185e-08, -1.156318e-08, 
    -1.195155e-08, -1.197962e-08, -1.156306e-08, -1.109303e-08, 
    -1.067721e-08, -1.042662e-08,
  -3.776698e-09, -4.831819e-09, -6.087675e-09, -7.251098e-09, -8.141827e-09, 
    -8.964748e-09, -9.657797e-09, -1.021577e-08, -1.0817e-08, -1.13408e-08, 
    -1.186867e-08, -1.215295e-08, -1.218941e-08, -1.20236e-08, -1.172551e-08,
  -3.124914e-09, -3.791749e-09, -4.769542e-09, -5.961023e-09, -7.086226e-09, 
    -7.922808e-09, -8.758633e-09, -9.44287e-09, -9.981261e-09, -1.054844e-08, 
    -1.097921e-08, -1.138839e-08, -1.170054e-08, -1.190643e-08, -1.207472e-08,
  -2.510839e-09, -3.013322e-09, -3.733859e-09, -4.684587e-09, -5.86055e-09, 
    -6.916983e-09, -7.755087e-09, -8.565388e-09, -9.211782e-09, 
    -9.762534e-09, -1.033281e-08, -1.068801e-08, -1.099606e-08, 
    -1.121092e-08, -1.140444e-08,
  -2.0166e-09, -2.421638e-09, -2.94708e-09, -3.658566e-09, -4.611873e-09, 
    -5.719246e-09, -6.75692e-09, -7.618922e-09, -8.352882e-09, -8.800572e-09, 
    -9.275917e-09, -9.749528e-09, -1.010549e-08, -1.044733e-08, -1.072712e-08,
  -1.642298e-09, -1.96865e-09, -2.373528e-09, -2.87837e-09, -3.606268e-09, 
    -4.558608e-09, -5.56921e-09, -6.551044e-09, -7.472198e-09, -8.092365e-09, 
    -8.502475e-09, -8.885295e-09, -9.141925e-09, -9.428705e-09, -9.736689e-09,
  -1.483735e-09, -1.67067e-09, -1.975207e-09, -2.33967e-09, -2.813769e-09, 
    -3.534212e-09, -4.464902e-09, -5.365961e-09, -6.332469e-09, 
    -7.055263e-09, -7.634795e-09, -8.029537e-09, -8.416376e-09, 
    -8.682968e-09, -8.918105e-09,
  -1.327297e-09, -1.454281e-09, -1.663847e-09, -1.936748e-09, -2.301856e-09, 
    -2.752581e-09, -3.396231e-09, -4.198459e-09, -5.072152e-09, 
    -5.930123e-09, -6.597796e-09, -7.063788e-09, -7.432118e-09, 
    -7.717782e-09, -7.996986e-09,
  -1.180877e-09, -1.311789e-09, -1.471434e-09, -1.689224e-09, -1.955063e-09, 
    -2.247107e-09, -2.655595e-09, -3.219664e-09, -3.887094e-09, 
    -4.604582e-09, -5.283988e-09, -5.806273e-09, -6.195324e-09, 
    -6.461234e-09, -6.748456e-09,
  -3.572941e-09, -4.013303e-09, -4.141683e-09, -4.413353e-09, -4.589514e-09, 
    -4.78096e-09, -5.051132e-09, -5.417479e-09, -6.009417e-09, -6.467915e-09, 
    -6.768112e-09, -7.245093e-09, -8.048982e-09, -8.643159e-09, -1.023202e-08,
  -3.616947e-09, -4.264268e-09, -4.543224e-09, -4.753467e-09, -4.968528e-09, 
    -5.175274e-09, -5.371362e-09, -5.606338e-09, -6.034307e-09, -6.49366e-09, 
    -6.799378e-09, -7.07126e-09, -7.678446e-09, -8.249452e-09, -8.813715e-09,
  -3.623505e-09, -4.265122e-09, -4.789143e-09, -5.13127e-09, -5.343253e-09, 
    -5.547679e-09, -5.795918e-09, -6.03002e-09, -6.376118e-09, -6.760831e-09, 
    -7.102485e-09, -7.338997e-09, -7.722248e-09, -8.22067e-09, -8.567737e-09,
  -3.821445e-09, -4.235559e-09, -4.920834e-09, -5.372225e-09, -5.720892e-09, 
    -5.981282e-09, -6.232769e-09, -6.448549e-09, -6.784373e-09, 
    -7.128391e-09, -7.427637e-09, -7.618623e-09, -7.979726e-09, 
    -8.491943e-09, -8.91394e-09,
  -3.966109e-09, -4.326583e-09, -5.000165e-09, -5.61332e-09, -6.06354e-09, 
    -6.438349e-09, -6.822882e-09, -7.071738e-09, -7.348058e-09, 
    -7.657307e-09, -7.920026e-09, -8.067842e-09, -8.225932e-09, 
    -8.643091e-09, -9.123807e-09,
  -4.096236e-09, -4.445111e-09, -5.051655e-09, -5.760406e-09, -6.306062e-09, 
    -6.785707e-09, -7.197722e-09, -7.45711e-09, -7.708014e-09, -7.994905e-09, 
    -8.24329e-09, -8.440706e-09, -8.621384e-09, -8.854972e-09, -9.194558e-09,
  -4.134302e-09, -4.463812e-09, -5.09612e-09, -5.798982e-09, -6.428732e-09, 
    -7.046984e-09, -7.624462e-09, -7.90731e-09, -8.197124e-09, -8.512208e-09, 
    -8.793155e-09, -9.062425e-09, -9.261112e-09, -9.412951e-09, -9.586073e-09,
  -4.082241e-09, -4.476721e-09, -4.984474e-09, -5.800095e-09, -6.635815e-09, 
    -7.255184e-09, -7.790611e-09, -8.34646e-09, -8.884408e-09, -9.294285e-09, 
    -9.615192e-09, -9.875398e-09, -1.010356e-08, -1.029307e-08, -1.049951e-08,
  -3.894896e-09, -4.326767e-09, -5.000271e-09, -5.989064e-09, -6.855062e-09, 
    -7.607373e-09, -8.567871e-09, -9.325903e-09, -1.004136e-08, 
    -1.042191e-08, -1.039518e-08, -1.029556e-08, -1.0216e-08, -1.021639e-08, 
    -1.023011e-08,
  -3.700855e-09, -4.077406e-09, -4.945715e-09, -6.000133e-09, -6.802487e-09, 
    -7.689025e-09, -8.513264e-09, -8.884513e-09, -8.983241e-09, 
    -8.833924e-09, -8.546373e-09, -8.44614e-09, -8.32703e-09, -8.322808e-09, 
    -8.27958e-09,
  -1.288139e-09, -1.347391e-09, -1.437903e-09, -1.533635e-09, -1.615225e-09, 
    -1.671876e-09, -1.713678e-09, -1.741652e-09, -1.775026e-09, 
    -1.838029e-09, -1.903387e-09, -2.016259e-09, -2.083028e-09, 
    -2.181878e-09, -2.242038e-09,
  -1.046669e-09, -1.124748e-09, -1.230929e-09, -1.337906e-09, -1.466234e-09, 
    -1.564658e-09, -1.638592e-09, -1.706127e-09, -1.76798e-09, -1.839911e-09, 
    -1.909659e-09, -1.945908e-09, -2.031672e-09, -2.093493e-09, -2.219353e-09,
  -7.941047e-10, -8.562752e-10, -9.361831e-10, -1.02853e-09, -1.138286e-09, 
    -1.257211e-09, -1.351595e-09, -1.454601e-09, -1.562129e-09, 
    -1.698692e-09, -1.848507e-09, -1.97108e-09, -2.040178e-09, -2.133506e-09, 
    -2.220477e-09,
  -6.364214e-10, -6.828164e-10, -7.328425e-10, -7.971697e-10, -8.777204e-10, 
    -9.642405e-10, -1.026815e-09, -1.077781e-09, -1.153139e-09, 
    -1.279471e-09, -1.453992e-09, -1.680712e-09, -1.867009e-09, 
    -2.034447e-09, -2.220173e-09,
  -6.524692e-10, -7.067609e-10, -7.565398e-10, -8.174657e-10, -8.802932e-10, 
    -9.645587e-10, -1.043986e-09, -1.093996e-09, -1.151195e-09, 
    -1.225845e-09, -1.301554e-09, -1.391677e-09, -1.5387e-09, -1.732962e-09, 
    -1.988729e-09,
  -7.623456e-10, -8.485975e-10, -9.777574e-10, -1.122906e-09, -1.222884e-09, 
    -1.304128e-09, -1.349161e-09, -1.33627e-09, -1.33424e-09, -1.359435e-09, 
    -1.411036e-09, -1.46171e-09, -1.503255e-09, -1.593282e-09, -1.723962e-09,
  -1.353055e-09, -1.617007e-09, -1.872563e-09, -2.01005e-09, -2.118415e-09, 
    -2.161888e-09, -2.210456e-09, -2.173446e-09, -2.115202e-09, 
    -2.017901e-09, -1.912387e-09, -1.843935e-09, -1.745058e-09, 
    -1.751077e-09, -1.796095e-09,
  -2.384587e-09, -2.609261e-09, -2.86198e-09, -3.121597e-09, -3.272295e-09, 
    -3.316578e-09, -3.291888e-09, -3.245697e-09, -3.16336e-09, -3.019406e-09, 
    -2.780834e-09, -2.53125e-09, -2.372864e-09, -2.289427e-09, -2.248674e-09,
  -3.516677e-09, -3.65438e-09, -3.799874e-09, -3.868151e-09, -3.817419e-09, 
    -3.799932e-09, -3.844755e-09, -3.987609e-09, -4.27823e-09, -4.537021e-09, 
    -4.688477e-09, -4.572003e-09, -4.196011e-09, -3.691019e-09, -3.230336e-09,
  -4.469153e-09, -4.392176e-09, -4.32504e-09, -4.157283e-09, -4.122365e-09, 
    -4.279145e-09, -4.645363e-09, -4.80639e-09, -5.07082e-09, -5.264376e-09, 
    -5.450716e-09, -5.724903e-09, -6.228899e-09, -6.597833e-09, -6.671451e-09,
  -2.038818e-09, -2.065905e-09, -2.079027e-09, -2.085417e-09, -2.089217e-09, 
    -2.081888e-09, -2.073988e-09, -2.067954e-09, -2.064973e-09, 
    -2.065158e-09, -2.070255e-09, -2.076343e-09, -2.104134e-09, 
    -2.153378e-09, -2.224309e-09,
  -2.100378e-09, -2.118102e-09, -2.140576e-09, -2.164068e-09, -2.179386e-09, 
    -2.195971e-09, -2.209676e-09, -2.225406e-09, -2.236487e-09, 
    -2.237365e-09, -2.229791e-09, -2.206676e-09, -2.178006e-09, 
    -2.164616e-09, -2.164079e-09,
  -2.090155e-09, -2.098306e-09, -2.063602e-09, -2.043271e-09, -2.025691e-09, 
    -2.030279e-09, -2.037827e-09, -2.05823e-09, -2.08995e-09, -2.130577e-09, 
    -2.172301e-09, -2.209638e-09, -2.233913e-09, -2.251538e-09, -2.26506e-09,
  -1.680543e-09, -1.618346e-09, -1.613484e-09, -1.768241e-09, -1.951879e-09, 
    -2.071117e-09, -2.104797e-09, -2.088379e-09, -2.026401e-09, 
    -1.954758e-09, -1.90453e-09, -1.889769e-09, -1.905805e-09, -1.953401e-09, 
    -2.013843e-09,
  -1.804384e-09, -2.355789e-09, -3.042549e-09, -3.22243e-09, -3.120844e-09, 
    -2.955132e-09, -2.796934e-09, -2.702731e-09, -2.651205e-09, -2.61408e-09, 
    -2.593385e-09, -2.561521e-09, -2.492228e-09, -2.37846e-09, -2.225897e-09,
  -3.822842e-09, -4.48287e-09, -4.179853e-09, -3.608929e-09, -3.086633e-09, 
    -2.655141e-09, -2.368715e-09, -2.154055e-09, -2.046448e-09, 
    -1.992254e-09, -1.988845e-09, -2.026108e-09, -2.091641e-09, 
    -2.164781e-09, -2.28565e-09,
  -5.713249e-09, -4.614698e-09, -3.360825e-09, -2.406403e-09, -1.930343e-09, 
    -1.593513e-09, -1.440858e-09, -1.401417e-09, -1.420367e-09, 
    -1.442825e-09, -1.434037e-09, -1.440115e-09, -1.491073e-09, 
    -1.594717e-09, -1.750148e-09,
  -5.009009e-09, -3.383483e-09, -2.188071e-09, -1.545011e-09, -1.097668e-09, 
    -7.814902e-10, -6.674644e-10, -6.741842e-10, -7.755125e-10, 
    -9.289483e-10, -1.109933e-09, -1.239739e-09, -1.244392e-09, 
    -1.263358e-09, -1.308271e-09,
  -4.606004e-09, -2.802861e-09, -1.840927e-09, -1.14058e-09, -6.108398e-10, 
    -3.444271e-10, -2.280206e-10, -1.992508e-10, -2.140601e-10, -3.0841e-10, 
    -4.730527e-10, -7.42171e-10, -1.024285e-09, -1.262808e-09, -1.369909e-09,
  -4.050908e-09, -2.504413e-09, -1.594454e-09, -8.262388e-10, -2.689264e-10, 
    -7.242654e-11, -4.373185e-11, -8.40231e-11, -1.413603e-10, -2.235095e-10, 
    -3.699196e-10, -5.005144e-10, -6.392887e-10, -8.508438e-10, -1.125035e-09,
  -9.557709e-10, -1.040406e-09, -1.133712e-09, -1.241164e-09, -1.356374e-09, 
    -1.464402e-09, -1.560708e-09, -1.650727e-09, -1.755936e-09, 
    -1.906836e-09, -2.094142e-09, -2.32488e-09, -2.626816e-09, -3.02249e-09, 
    -3.509105e-09,
  -8.317972e-10, -8.942519e-10, -9.759807e-10, -1.064787e-09, -1.152213e-09, 
    -1.246798e-09, -1.346633e-09, -1.443539e-09, -1.531117e-09, 
    -1.612742e-09, -1.714579e-09, -1.841921e-09, -2.012673e-09, 
    -2.244341e-09, -2.550759e-09,
  -7.683623e-10, -8.026752e-10, -8.557059e-10, -9.235762e-10, -9.999641e-10, 
    -1.080536e-09, -1.165489e-09, -1.257254e-09, -1.351881e-09, 
    -1.441795e-09, -1.524359e-09, -1.602729e-09, -1.682363e-09, -1.78448e-09, 
    -1.930537e-09,
  -8.33374e-10, -8.52989e-10, -8.761585e-10, -9.138746e-10, -9.597468e-10, 
    -1.014002e-09, -1.074399e-09, -1.141806e-09, -1.220265e-09, 
    -1.302059e-09, -1.380917e-09, -1.456469e-09, -1.526152e-09, 
    -1.593426e-09, -1.657496e-09,
  -1.134414e-09, -1.144467e-09, -1.19147e-09, -1.281671e-09, -1.380434e-09, 
    -1.464598e-09, -1.524918e-09, -1.567974e-09, -1.607715e-09, 
    -1.654102e-09, -1.723827e-09, -1.802314e-09, -1.870296e-09, 
    -1.918427e-09, -1.90325e-09,
  -1.771431e-09, -1.985771e-09, -2.164133e-09, -2.281338e-09, -2.338453e-09, 
    -2.358133e-09, -2.3158e-09, -2.271147e-09, -2.220248e-09, -2.158061e-09, 
    -2.101515e-09, -2.048396e-09, -2.014712e-09, -1.989705e-09, -2.019024e-09,
  -3.036644e-09, -3.569982e-09, -3.726778e-09, -3.739892e-09, -3.654665e-09, 
    -3.434301e-09, -3.19672e-09, -2.993517e-09, -2.805665e-09, -2.636804e-09, 
    -2.477205e-09, -2.330615e-09, -2.217377e-09, -2.145434e-09, -2.117829e-09,
  -4.431763e-09, -4.621571e-09, -4.518729e-09, -4.272595e-09, -3.928278e-09, 
    -3.574561e-09, -3.298928e-09, -3.073753e-09, -2.88764e-09, -2.74993e-09, 
    -2.610514e-09, -2.453618e-09, -2.255206e-09, -2.077909e-09, -1.963415e-09,
  -4.095738e-09, -3.549827e-09, -3.005489e-09, -2.499876e-09, -2.116873e-09, 
    -1.849919e-09, -1.662561e-09, -1.496944e-09, -1.383921e-09, 
    -1.302511e-09, -1.285073e-09, -1.302422e-09, -1.343259e-09, -1.37988e-09, 
    -1.408088e-09,
  -2.317932e-09, -1.525296e-09, -9.403762e-10, -6.777371e-10, -5.477028e-10, 
    -4.506008e-10, -3.58293e-10, -2.925284e-10, -2.455532e-10, -2.370232e-10, 
    -2.468719e-10, -3.038103e-10, -3.697224e-10, -4.065848e-10, -4.702168e-10,
  -1.598777e-09, -1.558491e-09, -1.524114e-09, -1.489709e-09, -1.457079e-09, 
    -1.430838e-09, -1.41363e-09, -1.401841e-09, -1.388974e-09, -1.362166e-09, 
    -1.326963e-09, -1.274991e-09, -1.212198e-09, -1.141581e-09, -1.069938e-09,
  -1.82286e-09, -1.781521e-09, -1.733659e-09, -1.690427e-09, -1.643635e-09, 
    -1.609753e-09, -1.583082e-09, -1.564169e-09, -1.549957e-09, 
    -1.534549e-09, -1.511765e-09, -1.480191e-09, -1.428297e-09, 
    -1.367456e-09, -1.294038e-09,
  -2.007743e-09, -1.957626e-09, -1.908483e-09, -1.85019e-09, -1.790126e-09, 
    -1.732949e-09, -1.681759e-09, -1.639022e-09, -1.603773e-09, 
    -1.577355e-09, -1.55759e-09, -1.547321e-09, -1.542829e-09, -1.528295e-09, 
    -1.493873e-09,
  -2.034612e-09, -1.976231e-09, -1.913182e-09, -1.847497e-09, -1.786958e-09, 
    -1.726335e-09, -1.671323e-09, -1.622102e-09, -1.581721e-09, -1.54998e-09, 
    -1.527273e-09, -1.508694e-09, -1.502741e-09, -1.505155e-09, -1.515481e-09,
  -1.961205e-09, -1.912861e-09, -1.852456e-09, -1.7899e-09, -1.728834e-09, 
    -1.670145e-09, -1.617482e-09, -1.571641e-09, -1.528488e-09, 
    -1.483461e-09, -1.455633e-09, -1.444301e-09, -1.441966e-09, 
    -1.447205e-09, -1.456022e-09,
  -1.733881e-09, -1.70016e-09, -1.69248e-09, -1.693273e-09, -1.666631e-09, 
    -1.631168e-09, -1.57781e-09, -1.519394e-09, -1.465899e-09, -1.413138e-09, 
    -1.374342e-09, -1.336472e-09, -1.319622e-09, -1.321792e-09, -1.33762e-09,
  -1.545017e-09, -1.52889e-09, -1.569593e-09, -1.641807e-09, -1.717233e-09, 
    -1.769093e-09, -1.779325e-09, -1.739079e-09, -1.665368e-09, 
    -1.571273e-09, -1.476609e-09, -1.396204e-09, -1.32695e-09, -1.274039e-09, 
    -1.235081e-09,
  -1.30514e-09, -1.259426e-09, -1.251413e-09, -1.273939e-09, -1.370351e-09, 
    -1.516888e-09, -1.684714e-09, -1.860714e-09, -1.992749e-09, 
    -2.082561e-09, -2.07673e-09, -1.966366e-09, -1.757449e-09, -1.50437e-09, 
    -1.339607e-09,
  -9.844288e-10, -8.487768e-10, -7.246235e-10, -6.698461e-10, -6.681091e-10, 
    -7.376169e-10, -8.842819e-10, -1.078729e-09, -1.328968e-09, 
    -1.588314e-09, -1.86688e-09, -2.112296e-09, -2.231044e-09, -2.232162e-09, 
    -2.109239e-09,
  -6.108801e-10, -4.275452e-10, -3.516305e-10, -3.381573e-10, -3.462018e-10, 
    -3.738612e-10, -4.171247e-10, -4.894362e-10, -6.021538e-10, 
    -7.756613e-10, -1.023845e-09, -1.292119e-09, -1.595652e-09, 
    -1.871476e-09, -2.14963e-09,
  -3.946303e-09, -4.557902e-09, -5.820182e-09, -7.323145e-09, -8.601382e-09, 
    -9.531597e-09, -1.015505e-08, -1.052841e-08, -1.073431e-08, 
    -1.081772e-08, -1.068751e-08, -1.040029e-08, -1.003547e-08, 
    -9.613053e-09, -9.16237e-09,
  -3.279855e-09, -3.375814e-09, -3.639457e-09, -4.172335e-09, -5.011531e-09, 
    -5.909906e-09, -6.593289e-09, -7.09631e-09, -7.423242e-09, -7.658594e-09, 
    -7.722232e-09, -7.67617e-09, -7.481843e-09, -7.200958e-09, -6.823155e-09,
  -3.147115e-09, -3.096471e-09, -3.070686e-09, -3.099964e-09, -3.264188e-09, 
    -3.576105e-09, -4.038959e-09, -4.478881e-09, -4.805795e-09, 
    -5.018269e-09, -5.092514e-09, -5.087539e-09, -4.962216e-09, 
    -4.746497e-09, -4.469634e-09,
  -2.921586e-09, -3.003403e-09, -3.025607e-09, -3.005667e-09, -2.958304e-09, 
    -2.931941e-09, -2.970695e-09, -3.092593e-09, -3.221025e-09, 
    -3.341254e-09, -3.400802e-09, -3.420191e-09, -3.363528e-09, 
    -3.266666e-09, -3.139344e-09,
  -2.420191e-09, -2.595253e-09, -2.762042e-09, -2.839455e-09, -2.853652e-09, 
    -2.826747e-09, -2.787707e-09, -2.762533e-09, -2.756189e-09, 
    -2.774756e-09, -2.782665e-09, -2.791453e-09, -2.767298e-09, 
    -2.734757e-09, -2.68045e-09,
  -2.129176e-09, -2.223494e-09, -2.347639e-09, -2.469874e-09, -2.524778e-09, 
    -2.559299e-09, -2.580175e-09, -2.603872e-09, -2.606269e-09, 
    -2.606301e-09, -2.585573e-09, -2.575706e-09, -2.547656e-09, -2.50666e-09, 
    -2.460677e-09,
  -2.078656e-09, -2.073385e-09, -2.109966e-09, -2.167603e-09, -2.229942e-09, 
    -2.286944e-09, -2.32359e-09, -2.35134e-09, -2.369429e-09, -2.375579e-09, 
    -2.37083e-09, -2.352003e-09, -2.325238e-09, -2.286928e-09, -2.25048e-09,
  -2.129534e-09, -2.063033e-09, -2.024918e-09, -2.003767e-09, -1.99953e-09, 
    -1.994521e-09, -1.998889e-09, -2.005204e-09, -2.017391e-09, 
    -2.013356e-09, -2.009561e-09, -1.9865e-09, -1.974945e-09, -1.964543e-09, 
    -1.978617e-09,
  -2.057992e-09, -1.975333e-09, -1.893722e-09, -1.820721e-09, -1.764098e-09, 
    -1.726343e-09, -1.691866e-09, -1.661935e-09, -1.628172e-09, 
    -1.598872e-09, -1.567809e-09, -1.545155e-09, -1.521873e-09, 
    -1.531316e-09, -1.587809e-09,
  -1.820879e-09, -1.727748e-09, -1.623889e-09, -1.530238e-09, -1.462065e-09, 
    -1.4051e-09, -1.353946e-09, -1.309092e-09, -1.264348e-09, -1.219505e-09, 
    -1.167945e-09, -1.120068e-09, -1.06564e-09, -1.031179e-09, -1.012491e-09,
  -5.800993e-09, -8.152772e-09, -1.122764e-08, -1.334211e-08, -1.493061e-08, 
    -1.633812e-08, -1.749108e-08, -1.853105e-08, -1.932365e-08, 
    -1.978013e-08, -2.002324e-08, -1.994833e-08, -1.989657e-08, 
    -1.975367e-08, -1.967177e-08,
  -3.919735e-09, -5.285602e-09, -7.473752e-09, -1.002203e-08, -1.210511e-08, 
    -1.391635e-08, -1.523137e-08, -1.63173e-08, -1.745746e-08, -1.854184e-08, 
    -1.925956e-08, -1.976148e-08, -1.991664e-08, -2.003633e-08, -1.996912e-08,
  -3.330668e-09, -3.705188e-09, -4.894382e-09, -6.837822e-09, -8.997396e-09, 
    -1.10149e-08, -1.280965e-08, -1.421081e-08, -1.534108e-08, -1.640191e-08, 
    -1.731261e-08, -1.800874e-08, -1.839738e-08, -1.864861e-08, -1.878179e-08,
  -3.047943e-09, -3.170559e-09, -3.458972e-09, -4.438249e-09, -6.014395e-09, 
    -7.848974e-09, -9.626938e-09, -1.122985e-08, -1.257755e-08, 
    -1.374894e-08, -1.480329e-08, -1.564813e-08, -1.625011e-08, 
    -1.650964e-08, -1.671215e-08,
  -2.915908e-09, -2.969952e-09, -3.129499e-09, -3.354825e-09, -4.046494e-09, 
    -5.284458e-09, -6.796677e-09, -8.295301e-09, -9.609593e-09, 
    -1.073146e-08, -1.174599e-08, -1.261451e-08, -1.334916e-08, 
    -1.385343e-08, -1.409222e-08,
  -2.695405e-09, -2.70737e-09, -2.783083e-09, -2.952728e-09, -3.15924e-09, 
    -3.612253e-09, -4.48363e-09, -5.688636e-09, -6.865594e-09, -7.958242e-09, 
    -8.930802e-09, -9.738291e-09, -1.030962e-08, -1.07776e-08, -1.104223e-08,
  -2.578052e-09, -2.554126e-09, -2.567092e-09, -2.602339e-09, -2.714387e-09, 
    -2.913337e-09, -3.175832e-09, -3.730131e-09, -4.509454e-09, 
    -5.345937e-09, -6.179877e-09, -7.008216e-09, -7.612821e-09, 
    -8.066182e-09, -8.261826e-09,
  -2.590555e-09, -2.531446e-09, -2.475256e-09, -2.456831e-09, -2.419665e-09, 
    -2.486753e-09, -2.627924e-09, -2.810105e-09, -3.137614e-09, 
    -3.585569e-09, -4.125753e-09, -4.601045e-09, -5.088356e-09, 
    -5.524963e-09, -5.815096e-09,
  -2.488979e-09, -2.489582e-09, -2.487344e-09, -2.484549e-09, -2.457438e-09, 
    -2.416274e-09, -2.39247e-09, -2.426396e-09, -2.511978e-09, -2.628943e-09, 
    -2.768325e-09, -2.981882e-09, -3.228434e-09, -3.512798e-09, -3.793115e-09,
  -2.44983e-09, -2.404453e-09, -2.369912e-09, -2.365921e-09, -2.367192e-09, 
    -2.368475e-09, -2.353888e-09, -2.354182e-09, -2.340027e-09, -2.35315e-09, 
    -2.369645e-09, -2.403667e-09, -2.444071e-09, -2.510272e-09, -2.569433e-09,
  -4.209845e-09, -5.146091e-09, -6.443266e-09, -8.273788e-09, -1.087322e-08, 
    -1.266541e-08, -1.401729e-08, -1.520242e-08, -1.615104e-08, 
    -1.713395e-08, -1.824248e-08, -1.940514e-08, -2.033889e-08, 
    -2.116763e-08, -2.175174e-08,
  -3.34329e-09, -4.144109e-09, -5.090073e-09, -6.354951e-09, -8.149652e-09, 
    -1.057451e-08, -1.234477e-08, -1.371768e-08, -1.48933e-08, -1.594366e-08, 
    -1.699799e-08, -1.802449e-08, -1.909609e-08, -1.996067e-08, -2.077191e-08,
  -2.829189e-09, -3.305114e-09, -4.064899e-09, -5.023977e-09, -6.253247e-09, 
    -8.021171e-09, -1.033629e-08, -1.213783e-08, -1.349444e-08, 
    -1.468435e-08, -1.577183e-08, -1.686767e-08, -1.785397e-08, 
    -1.883367e-08, -1.973273e-08,
  -2.606564e-09, -2.785053e-09, -3.251655e-09, -3.993057e-09, -4.928008e-09, 
    -6.151008e-09, -7.893793e-09, -1.006368e-08, -1.190217e-08, -1.32965e-08, 
    -1.450129e-08, -1.558322e-08, -1.680924e-08, -1.772787e-08, -1.86496e-08,
  -2.425425e-09, -2.61283e-09, -2.804033e-09, -3.251651e-09, -3.941232e-09, 
    -4.822377e-09, -6.032441e-09, -7.715692e-09, -9.81085e-09, -1.173022e-08, 
    -1.315135e-08, -1.442349e-08, -1.545643e-08, -1.67549e-08, -1.764954e-08,
  -2.294251e-09, -2.434224e-09, -2.637373e-09, -2.831983e-09, -3.270085e-09, 
    -3.903086e-09, -4.70919e-09, -5.859921e-09, -7.458023e-09, -9.529118e-09, 
    -1.144914e-08, -1.300137e-08, -1.420408e-08, -1.536635e-08, -1.647767e-08,
  -2.179296e-09, -2.312382e-09, -2.454665e-09, -2.673833e-09, -2.873776e-09, 
    -3.300385e-09, -3.864813e-09, -4.590931e-09, -5.606539e-09, 
    -7.122443e-09, -9.106027e-09, -1.108802e-08, -1.275178e-08, 
    -1.399199e-08, -1.514644e-08,
  -2.167493e-09, -2.297321e-09, -2.395145e-09, -2.522585e-09, -2.678426e-09, 
    -2.900354e-09, -3.252812e-09, -3.75059e-09, -4.361036e-09, -5.273393e-09, 
    -6.63121e-09, -8.412338e-09, -1.04132e-08, -1.213332e-08, -1.346196e-08,
  -2.254384e-09, -2.279125e-09, -2.403813e-09, -2.533742e-09, -2.634338e-09, 
    -2.713775e-09, -2.911631e-09, -3.197688e-09, -3.604714e-09, 
    -4.106612e-09, -4.882468e-09, -5.958938e-09, -7.486768e-09, 
    -9.290622e-09, -1.093235e-08,
  -2.493776e-09, -2.442421e-09, -2.420093e-09, -2.506461e-09, -2.630357e-09, 
    -2.737676e-09, -2.80271e-09, -2.914319e-09, -3.10957e-09, -3.399331e-09, 
    -3.838121e-09, -4.455053e-09, -5.253712e-09, -6.340372e-09, -7.615268e-09,
  -3.099771e-09, -3.784408e-09, -4.837702e-09, -6.258075e-09, -7.84638e-09, 
    -1.009621e-08, -1.249547e-08, -1.448781e-08, -1.580508e-08, 
    -1.711127e-08, -1.856436e-08, -2.009035e-08, -2.12517e-08, -2.203702e-08, 
    -2.251505e-08,
  -2.448576e-09, -3.05219e-09, -3.829698e-09, -4.94631e-09, -6.289728e-09, 
    -7.9733e-09, -1.007578e-08, -1.250929e-08, -1.442234e-08, -1.586308e-08, 
    -1.719876e-08, -1.860145e-08, -1.997738e-08, -2.111119e-08, -2.186323e-08,
  -2.171223e-09, -2.570528e-09, -3.127598e-09, -3.93911e-09, -5.000687e-09, 
    -6.395649e-09, -8.052145e-09, -1.015855e-08, -1.258952e-08, 
    -1.446269e-08, -1.595017e-08, -1.722212e-08, -1.853158e-08, 
    -1.981553e-08, -2.09687e-08,
  -1.867901e-09, -2.227105e-09, -2.663713e-09, -3.252328e-09, -4.039733e-09, 
    -5.066679e-09, -6.496899e-09, -8.146523e-09, -1.025764e-08, -1.26612e-08, 
    -1.449737e-08, -1.597661e-08, -1.720856e-08, -1.838061e-08, -1.954822e-08,
  -1.573218e-09, -1.932449e-09, -2.328772e-09, -2.776706e-09, -3.395e-09, 
    -4.157122e-09, -5.172261e-09, -6.624874e-09, -8.281168e-09, 
    -1.046334e-08, -1.274205e-08, -1.449294e-08, -1.589853e-08, 
    -1.712803e-08, -1.822091e-08,
  -1.308641e-09, -1.614799e-09, -2.032143e-09, -2.457398e-09, -2.927101e-09, 
    -3.558887e-09, -4.298902e-09, -5.295606e-09, -6.681428e-09, 
    -8.434072e-09, -1.073049e-08, -1.282624e-08, -1.440094e-08, 
    -1.569547e-08, -1.68399e-08,
  -1.128566e-09, -1.31628e-09, -1.685394e-09, -2.145244e-09, -2.596412e-09, 
    -3.119339e-09, -3.730585e-09, -4.487581e-09, -5.449686e-09, -6.70563e-09, 
    -8.607398e-09, -1.097898e-08, -1.29415e-08, -1.43542e-08, -1.551935e-08,
  -1.025556e-09, -1.170121e-09, -1.452982e-09, -1.858419e-09, -2.294948e-09, 
    -2.76319e-09, -3.296055e-09, -3.907894e-09, -4.690382e-09, -5.627896e-09, 
    -6.786259e-09, -8.765127e-09, -1.103797e-08, -1.285636e-08, -1.416693e-08,
  -9.213167e-10, -1.067932e-09, -1.314174e-09, -1.68593e-09, -2.060569e-09, 
    -2.46469e-09, -2.897116e-09, -3.423828e-09, -4.059418e-09, -4.858405e-09, 
    -5.76086e-09, -7.039649e-09, -8.979216e-09, -1.09905e-08, -1.259002e-08,
  -7.962095e-10, -8.93681e-10, -1.148668e-09, -1.492744e-09, -1.877366e-09, 
    -2.244477e-09, -2.628759e-09, -3.022138e-09, -3.518212e-09, 
    -4.163184e-09, -4.920413e-09, -5.774447e-09, -7.164636e-09, 
    -8.994355e-09, -1.075822e-08,
  -1.027382e-09, -1.181714e-09, -1.470616e-09, -1.835914e-09, -2.267719e-09, 
    -2.78993e-09, -3.493878e-09, -4.368344e-09, -5.305918e-09, -5.971387e-09, 
    -6.806334e-09, -8.207419e-09, -1.002548e-08, -1.139443e-08, -1.226966e-08,
  -6.738685e-10, -7.653203e-10, -9.145986e-10, -1.131837e-09, -1.421578e-09, 
    -1.771818e-09, -2.24e-09, -2.859591e-09, -3.582897e-09, -4.480169e-09, 
    -5.320049e-09, -6.379375e-09, -7.894903e-09, -9.669184e-09, -1.117374e-08,
  -5.40277e-10, -5.57825e-10, -6.286712e-10, -7.503302e-10, -9.263413e-10, 
    -1.173354e-09, -1.493701e-09, -1.943208e-09, -2.531816e-09, 
    -3.195315e-09, -4.036279e-09, -5.035226e-09, -6.280589e-09, 
    -7.894081e-09, -9.625649e-09,
  -4.802468e-10, -4.807866e-10, -5.036224e-10, -5.581838e-10, -6.587404e-10, 
    -8.048788e-10, -1.025038e-09, -1.312985e-09, -1.764282e-09, 
    -2.324599e-09, -3.031905e-09, -3.867624e-09, -5.0403e-09, -6.483753e-09, 
    -8.174795e-09,
  -4.581036e-10, -4.685352e-10, -4.740664e-10, -4.953701e-10, -5.462651e-10, 
    -6.418088e-10, -7.78333e-10, -9.783556e-10, -1.269314e-09, -1.66249e-09, 
    -2.222276e-09, -2.997362e-09, -3.939642e-09, -5.253276e-09, -6.794483e-09,
  -4.611448e-10, -4.42587e-10, -4.446178e-10, -4.542379e-10, -4.922542e-10, 
    -5.476706e-10, -6.549185e-10, -7.783539e-10, -9.969301e-10, -1.29671e-09, 
    -1.658552e-09, -2.251054e-09, -3.108241e-09, -4.20754e-09, -5.550876e-09,
  -4.743669e-10, -4.662398e-10, -4.496893e-10, -4.440245e-10, -4.496106e-10, 
    -4.922647e-10, -5.836579e-10, -6.915506e-10, -8.279776e-10, -1.03789e-09, 
    -1.338252e-09, -1.750012e-09, -2.415605e-09, -3.417448e-09, -4.633069e-09,
  -4.179697e-10, -4.594433e-10, -4.653203e-10, -4.6317e-10, -4.516943e-10, 
    -4.541492e-10, -5.107076e-10, -6.162327e-10, -7.331509e-10, -8.92741e-10, 
    -1.106789e-09, -1.427299e-09, -1.928228e-09, -2.718413e-09, -3.874489e-09,
  -3.411742e-10, -4.174285e-10, -4.621936e-10, -4.90963e-10, -4.99265e-10, 
    -4.827859e-10, -4.905971e-10, -5.60877e-10, -6.674597e-10, -8.047773e-10, 
    -9.877952e-10, -1.231281e-09, -1.629503e-09, -2.246887e-09, -3.210703e-09,
  -2.774967e-10, -3.322481e-10, -4.060341e-10, -4.655432e-10, -5.178612e-10, 
    -5.399168e-10, -5.386975e-10, -5.616079e-10, -6.511379e-10, 
    -7.650755e-10, -9.318929e-10, -1.139653e-09, -1.430307e-09, 
    -1.939258e-09, -2.750489e-09,
  -4.851239e-09, -6.425754e-09, -8.178422e-09, -9.995954e-09, -1.168326e-08, 
    -1.297089e-08, -1.36871e-08, -1.392825e-08, -1.363659e-08, -1.31891e-08, 
    -1.296543e-08, -1.319068e-08, -1.362093e-08, -1.420765e-08, -1.492701e-08,
  -2.705995e-09, -4.06254e-09, -5.563231e-09, -7.175044e-09, -8.897148e-09, 
    -1.070681e-08, -1.218387e-08, -1.32609e-08, -1.370421e-08, -1.350972e-08, 
    -1.310014e-08, -1.276803e-08, -1.291725e-08, -1.330577e-08, -1.386136e-08,
  -1.087788e-09, -1.8351e-09, -3.013246e-09, -4.526829e-09, -6.165505e-09, 
    -7.87703e-09, -9.67299e-09, -1.117552e-08, -1.243786e-08, -1.306075e-08, 
    -1.311379e-08, -1.269232e-08, -1.232123e-08, -1.241234e-08, -1.273541e-08,
  -8.493891e-10, -9.524664e-10, -1.333144e-09, -2.190415e-09, -3.456624e-09, 
    -5.058021e-09, -6.823033e-09, -8.54007e-09, -1.009076e-08, -1.132659e-08, 
    -1.207089e-08, -1.237906e-08, -1.208524e-08, -1.170536e-08, -1.175233e-08,
  -8.469834e-10, -8.308857e-10, -8.90822e-10, -1.076709e-09, -1.621008e-09, 
    -2.581393e-09, -3.989295e-09, -5.777241e-09, -7.51324e-09, -9.033565e-09, 
    -1.024543e-08, -1.109954e-08, -1.152459e-08, -1.135707e-08, -1.102468e-08,
  -9.08473e-10, -8.757358e-10, -8.596961e-10, -8.669449e-10, -9.724167e-10, 
    -1.28346e-09, -1.910694e-09, -2.993862e-09, -4.690349e-09, -6.522938e-09, 
    -7.936716e-09, -9.154968e-09, -1.010071e-08, -1.057882e-08, -1.050289e-08,
  -8.484033e-10, -8.651957e-10, -8.701674e-10, -8.711237e-10, -8.638188e-10, 
    -9.160752e-10, -1.114362e-09, -1.457235e-09, -2.172524e-09, 
    -3.626778e-09, -5.442105e-09, -6.904763e-09, -7.981744e-09, 
    -9.006449e-09, -9.574712e-09,
  -7.22957e-10, -7.678146e-10, -8.006807e-10, -8.153552e-10, -8.272267e-10, 
    -8.242134e-10, -8.53024e-10, -9.602048e-10, -1.160424e-09, -1.627509e-09, 
    -2.663174e-09, -4.305367e-09, -5.750243e-09, -6.79818e-09, -7.738101e-09,
  -6.707743e-10, -6.716718e-10, -7.0111e-10, -7.371111e-10, -7.53988e-10, 
    -7.606777e-10, -7.482439e-10, -7.69202e-10, -8.154615e-10, -9.609465e-10, 
    -1.272771e-09, -1.983697e-09, -3.283524e-09, -4.584823e-09, -5.596201e-09,
  -7.155931e-10, -6.78223e-10, -6.533007e-10, -6.596983e-10, -6.804571e-10, 
    -6.961376e-10, -6.959691e-10, -6.737027e-10, -6.748315e-10, 
    -7.026795e-10, -7.97192e-10, -9.991539e-10, -1.470945e-09, -2.427357e-09, 
    -3.48534e-09,
  -2.267159e-09, -2.310921e-09, -2.346609e-09, -2.382352e-09, -2.445381e-09, 
    -2.63961e-09, -3.024152e-09, -3.524183e-09, -4.132302e-09, -4.846701e-09, 
    -5.540334e-09, -6.071201e-09, -6.597938e-09, -7.033195e-09, -7.434823e-09,
  -1.932907e-09, -2.036837e-09, -2.129048e-09, -2.200525e-09, -2.254397e-09, 
    -2.321242e-09, -2.518092e-09, -2.896239e-09, -3.417918e-09, 
    -4.052099e-09, -4.78704e-09, -5.441194e-09, -5.881564e-09, -6.299854e-09, 
    -6.740537e-09,
  -1.689729e-09, -1.732335e-09, -1.824632e-09, -1.931895e-09, -2.029119e-09, 
    -2.108276e-09, -2.201759e-09, -2.432784e-09, -2.865712e-09, 
    -3.446699e-09, -4.15242e-09, -4.953455e-09, -5.626996e-09, -5.919543e-09, 
    -6.282516e-09,
  -1.573559e-09, -1.588655e-09, -1.616085e-09, -1.68342e-09, -1.772998e-09, 
    -1.865184e-09, -1.959936e-09, -2.08214e-09, -2.378709e-09, -2.8705e-09, 
    -3.498827e-09, -4.287508e-09, -5.166457e-09, -5.87974e-09, -6.132038e-09,
  -1.635721e-09, -1.585101e-09, -1.568611e-09, -1.570721e-09, -1.620837e-09, 
    -1.692883e-09, -1.775333e-09, -1.867779e-09, -2.015412e-09, -2.3831e-09, 
    -2.946232e-09, -3.625923e-09, -4.481867e-09, -5.436625e-09, -6.20605e-09,
  -1.619859e-09, -1.606164e-09, -1.582594e-09, -1.575577e-09, -1.576585e-09, 
    -1.606331e-09, -1.653824e-09, -1.720518e-09, -1.809948e-09, 
    -1.979914e-09, -2.45339e-09, -3.109616e-09, -3.845501e-09, -4.745184e-09, 
    -5.782586e-09,
  -1.451382e-09, -1.46925e-09, -1.498239e-09, -1.511717e-09, -1.503641e-09, 
    -1.514682e-09, -1.56666e-09, -1.638206e-09, -1.712702e-09, -1.800139e-09, 
    -2.01457e-09, -2.5384e-09, -3.299943e-09, -4.069098e-09, -5.071811e-09,
  -1.117827e-09, -1.177603e-09, -1.25485e-09, -1.346429e-09, -1.409535e-09, 
    -1.43022e-09, -1.435747e-09, -1.484185e-09, -1.585742e-09, -1.71399e-09, 
    -1.835294e-09, -2.094578e-09, -2.684548e-09, -3.477994e-09, -4.346308e-09,
  -7.408377e-10, -8.233903e-10, -9.174062e-10, -1.034606e-09, -1.154515e-09, 
    -1.266511e-09, -1.349818e-09, -1.390183e-09, -1.441432e-09, 
    -1.544272e-09, -1.693145e-09, -1.833156e-09, -2.145989e-09, 
    -2.826116e-09, -3.664122e-09,
  -6.296347e-10, -6.893157e-10, -7.763503e-10, -8.560138e-10, -9.437999e-10, 
    -1.063453e-09, -1.186458e-09, -1.284948e-09, -1.354431e-09, 
    -1.426515e-09, -1.509692e-09, -1.676123e-09, -1.823397e-09, 
    -2.195163e-09, -2.923437e-09,
  -7.977536e-09, -8.475426e-09, -8.990986e-09, -9.535432e-09, -1.001108e-08, 
    -1.0529e-08, -1.099983e-08, -1.140153e-08, -1.169963e-08, -1.218959e-08, 
    -1.3068e-08, -1.407307e-08, -1.501732e-08, -1.588296e-08, -1.667159e-08,
  -6.090881e-09, -6.67019e-09, -7.171785e-09, -7.674961e-09, -8.173962e-09, 
    -8.715611e-09, -9.208826e-09, -9.687204e-09, -1.012079e-08, 
    -1.050669e-08, -1.083627e-08, -1.121669e-08, -1.183671e-08, 
    -1.254926e-08, -1.325266e-08,
  -4.264679e-09, -4.718464e-09, -5.24314e-09, -5.768413e-09, -6.249488e-09, 
    -6.712123e-09, -7.203923e-09, -7.718641e-09, -8.22598e-09, -8.688112e-09, 
    -9.131956e-09, -9.526122e-09, -9.859055e-09, -1.014691e-08, -1.057417e-08,
  -3.060177e-09, -3.32001e-09, -3.641291e-09, -4.020769e-09, -4.451662e-09, 
    -4.913264e-09, -5.346345e-09, -5.795501e-09, -6.257749e-09, 
    -6.746386e-09, -7.243426e-09, -7.734601e-09, -8.181623e-09, 
    -8.583116e-09, -8.89922e-09,
  -2.221719e-09, -2.388067e-09, -2.572623e-09, -2.78298e-09, -3.022925e-09, 
    -3.301016e-09, -3.618098e-09, -3.976656e-09, -4.366249e-09, 
    -4.777189e-09, -5.209044e-09, -5.658055e-09, -6.121734e-09, 
    -6.570603e-09, -6.982661e-09,
  -1.794759e-09, -1.858145e-09, -1.942514e-09, -2.061515e-09, -2.20181e-09, 
    -2.364621e-09, -2.548882e-09, -2.747574e-09, -2.986794e-09, 
    -3.249301e-09, -3.563963e-09, -3.909494e-09, -4.292115e-09, -4.69887e-09, 
    -5.112239e-09,
  -1.688452e-09, -1.692885e-09, -1.700302e-09, -1.725367e-09, -1.764481e-09, 
    -1.808159e-09, -1.872283e-09, -1.961698e-09, -2.087695e-09, 
    -2.247106e-09, -2.436501e-09, -2.655663e-09, -2.910321e-09, 
    -3.211104e-09, -3.54489e-09,
  -1.985584e-09, -1.948936e-09, -1.912088e-09, -1.877495e-09, -1.848641e-09, 
    -1.838016e-09, -1.827679e-09, -1.829269e-09, -1.843193e-09, -1.88058e-09, 
    -1.944619e-09, -2.025208e-09, -2.136069e-09, -2.269198e-09, -2.439535e-09,
  -2.037959e-09, -2.02295e-09, -2.01481e-09, -2.015153e-09, -2.008002e-09, 
    -2.01059e-09, -2.009075e-09, -2.003696e-09, -2.005912e-09, -2.012518e-09, 
    -2.029548e-09, -2.048042e-09, -2.065844e-09, -2.086229e-09, -2.114546e-09,
  -1.946273e-09, -1.833196e-09, -1.741145e-09, -1.678307e-09, -1.650225e-09, 
    -1.668693e-09, -1.71559e-09, -1.797944e-09, -1.891327e-09, -1.993373e-09, 
    -2.072494e-09, -2.132786e-09, -2.176458e-09, -2.207981e-09, -2.220954e-09,
  -1.665762e-08, -1.684678e-08, -1.692361e-08, -1.688791e-08, -1.676798e-08, 
    -1.663222e-08, -1.685328e-08, -1.689672e-08, -1.707907e-08, 
    -1.713903e-08, -1.743006e-08, -1.775006e-08, -1.8215e-08, -1.885331e-08, 
    -1.961358e-08,
  -1.540708e-08, -1.586572e-08, -1.62613e-08, -1.647728e-08, -1.661511e-08, 
    -1.652139e-08, -1.637312e-08, -1.62161e-08, -1.624207e-08, -1.623012e-08, 
    -1.631317e-08, -1.641261e-08, -1.660658e-08, -1.695548e-08, -1.729044e-08,
  -1.336527e-08, -1.419515e-08, -1.482307e-08, -1.536059e-08, -1.576857e-08, 
    -1.603826e-08, -1.617736e-08, -1.617193e-08, -1.603311e-08, 
    -1.584659e-08, -1.567803e-08, -1.560221e-08, -1.558494e-08, 
    -1.562736e-08, -1.573319e-08,
  -1.074211e-08, -1.165861e-08, -1.256984e-08, -1.330322e-08, -1.404487e-08, 
    -1.462109e-08, -1.507178e-08, -1.538363e-08, -1.560309e-08, 
    -1.573893e-08, -1.576413e-08, -1.565807e-08, -1.549893e-08, 
    -1.531261e-08, -1.51658e-08,
  -8.222072e-09, -8.995734e-09, -9.823955e-09, -1.062675e-08, -1.141475e-08, 
    -1.214097e-08, -1.288905e-08, -1.351046e-08, -1.406058e-08, 
    -1.448642e-08, -1.479415e-08, -1.502052e-08, -1.516247e-08, 
    -1.524122e-08, -1.524016e-08,
  -6.098454e-09, -6.63667e-09, -7.211306e-09, -7.824721e-09, -8.481718e-09, 
    -9.127819e-09, -9.81882e-09, -1.051399e-08, -1.122867e-08, -1.19315e-08, 
    -1.259548e-08, -1.319942e-08, -1.369871e-08, -1.411173e-08, -1.44428e-08,
  -4.48606e-09, -4.809198e-09, -5.159119e-09, -5.529555e-09, -5.92846e-09, 
    -6.351315e-09, -6.821092e-09, -7.347266e-09, -7.9151e-09, -8.522003e-09, 
    -9.142872e-09, -9.783142e-09, -1.042967e-08, -1.107114e-08, -1.168813e-08,
  -3.341563e-09, -3.505605e-09, -3.675464e-09, -3.872757e-09, -4.097269e-09, 
    -4.340052e-09, -4.61218e-09, -4.929813e-09, -5.301572e-09, -5.715893e-09, 
    -6.200692e-09, -6.71624e-09, -7.275557e-09, -7.855185e-09, -8.474624e-09,
  -2.742696e-09, -2.78042e-09, -2.822805e-09, -2.892129e-09, -2.990736e-09, 
    -3.120876e-09, -3.279406e-09, -3.481726e-09, -3.719726e-09, 
    -3.977958e-09, -4.264023e-09, -4.57716e-09, -4.940545e-09, -5.343433e-09, 
    -5.796746e-09,
  -2.531745e-09, -2.525876e-09, -2.510723e-09, -2.508868e-09, -2.532086e-09, 
    -2.562183e-09, -2.605992e-09, -2.671155e-09, -2.769864e-09, 
    -2.903371e-09, -3.068331e-09, -3.257854e-09, -3.479311e-09, 
    -3.746187e-09, -4.03277e-09,
  -2.337626e-08, -2.244218e-08, -2.063827e-08, -2.119788e-08, -1.831943e-08, 
    -1.574512e-08, -1.483636e-08, -1.489769e-08, -1.470209e-08, 
    -1.414685e-08, -1.364719e-08, -1.339568e-08, -1.349051e-08, 
    -1.379789e-08, -1.387274e-08,
  -2.256646e-08, -2.411736e-08, -2.394118e-08, -2.210036e-08, -2.114469e-08, 
    -1.969676e-08, -1.704481e-08, -1.576718e-08, -1.527792e-08, 
    -1.510415e-08, -1.447134e-08, -1.43466e-08, -1.423524e-08, -1.418786e-08, 
    -1.42813e-08,
  -1.79773e-08, -1.919885e-08, -2.197171e-08, -2.336686e-08, -2.290561e-08, 
    -2.287555e-08, -2.118744e-08, -1.813615e-08, -1.647798e-08, 
    -1.585994e-08, -1.530987e-08, -1.492391e-08, -1.467558e-08, -1.46161e-08, 
    -1.467386e-08,
  -1.577705e-08, -1.648245e-08, -1.775827e-08, -1.910666e-08, -2.106457e-08, 
    -2.257354e-08, -2.258064e-08, -2.289853e-08, -2.087278e-08, 
    -1.777925e-08, -1.625467e-08, -1.555993e-08, -1.535426e-08, 
    -1.535646e-08, -1.545906e-08,
  -1.370136e-08, -1.391377e-08, -1.479459e-08, -1.566207e-08, -1.719615e-08, 
    -1.856932e-08, -2.031055e-08, -2.173783e-08, -2.184964e-08, 
    -2.192669e-08, -2.063034e-08, -1.731367e-08, -1.612748e-08, 
    -1.554807e-08, -1.555931e-08,
  -1.118142e-08, -1.139265e-08, -1.190581e-08, -1.239813e-08, -1.350833e-08, 
    -1.465337e-08, -1.630049e-08, -1.810528e-08, -1.998851e-08, 
    -2.146649e-08, -2.14107e-08, -2.117996e-08, -1.966033e-08, -1.750105e-08, 
    -1.657339e-08,
  -8.552108e-09, -8.583695e-09, -8.717315e-09, -8.943489e-09, -9.468432e-09, 
    -1.018443e-08, -1.127543e-08, -1.269974e-08, -1.450187e-08, 
    -1.662287e-08, -1.87473e-08, -2.01868e-08, -2.048644e-08, -2.028022e-08, 
    -1.888696e-08,
  -6.538161e-09, -6.318418e-09, -6.206346e-09, -6.184071e-09, -6.383762e-09, 
    -6.805746e-09, -7.378662e-09, -8.282955e-09, -9.396794e-09, 
    -1.102222e-08, -1.302334e-08, -1.554398e-08, -1.774826e-08, 
    -1.910382e-08, -1.941081e-08,
  -4.591059e-09, -4.140145e-09, -3.791723e-09, -3.572024e-09, -3.515612e-09, 
    -3.579392e-09, -3.83052e-09, -4.275613e-09, -4.924692e-09, -5.941457e-09, 
    -7.186439e-09, -9.006897e-09, -1.127574e-08, -1.384922e-08, -1.648016e-08,
  -2.873887e-09, -2.432808e-09, -2.130255e-09, -1.966603e-09, -1.893612e-09, 
    -1.872646e-09, -1.948881e-09, -2.077141e-09, -2.322664e-09, 
    -2.712464e-09, -3.314609e-09, -4.19124e-09, -5.527505e-09, -7.414547e-09, 
    -9.704588e-09,
  -1.847881e-08, -1.927249e-08, -1.977843e-08, -2.047797e-08, -2.070439e-08, 
    -2.082531e-08, -2.023163e-08, -1.943422e-08, -1.880501e-08, 
    -1.799029e-08, -1.724341e-08, -1.632057e-08, -1.534731e-08, 
    -1.432699e-08, -1.319351e-08,
  -1.835535e-08, -1.885368e-08, -1.909724e-08, -1.956336e-08, -1.974077e-08, 
    -1.975772e-08, -1.943467e-08, -1.881852e-08, -1.792365e-08, 
    -1.762856e-08, -1.721264e-08, -1.653638e-08, -1.578613e-08, 
    -1.493139e-08, -1.409399e-08,
  -1.744536e-08, -1.782816e-08, -1.809814e-08, -1.858142e-08, -1.806053e-08, 
    -1.782304e-08, -1.803466e-08, -1.800756e-08, -1.73101e-08, -1.661548e-08, 
    -1.627364e-08, -1.585834e-08, -1.543017e-08, -1.491187e-08, -1.438697e-08,
  -1.677325e-08, -1.730461e-08, -1.784213e-08, -1.693527e-08, -1.584077e-08, 
    -1.518441e-08, -1.476345e-08, -1.46855e-08, -1.49729e-08, -1.513493e-08, 
    -1.472887e-08, -1.460092e-08, -1.440083e-08, -1.422056e-08, -1.42218e-08,
  -1.591857e-08, -1.609765e-08, -1.56455e-08, -1.360996e-08, -1.230615e-08, 
    -1.136957e-08, -1.103963e-08, -1.111969e-08, -1.186478e-08, 
    -1.277462e-08, -1.362773e-08, -1.352017e-08, -1.367111e-08, 
    -1.374708e-08, -1.348052e-08,
  -1.427911e-08, -1.484535e-08, -1.248164e-08, -1.095129e-08, -9.754746e-09, 
    -9.074378e-09, -8.682497e-09, -8.782535e-09, -9.105843e-09, 
    -9.730084e-09, -1.103554e-08, -1.220219e-08, -1.3275e-08, -1.317645e-08, 
    -1.302513e-08,
  -1.271288e-08, -1.202112e-08, -1.031199e-08, -9.281595e-09, -8.428712e-09, 
    -7.640933e-09, -7.358994e-09, -7.22429e-09, -7.187154e-09, -7.30979e-09, 
    -7.860169e-09, -9.035263e-09, -1.048428e-08, -1.188013e-08, -1.209176e-08,
  -1.126471e-08, -9.720808e-09, -9.37187e-09, -8.029725e-09, -6.85625e-09, 
    -5.704806e-09, -5.483571e-09, -5.342013e-09, -5.265507e-09, 
    -5.269964e-09, -5.50795e-09, -6.036489e-09, -7.24904e-09, -8.807103e-09, 
    -1.052029e-08,
  -8.763368e-09, -8.559788e-09, -7.870099e-09, -5.801726e-09, -4.415594e-09, 
    -3.253648e-09, -2.8186e-09, -2.698672e-09, -2.602939e-09, -2.812801e-09, 
    -3.261741e-09, -3.978625e-09, -4.729215e-09, -5.970527e-09, -7.568929e-09,
  -7.447404e-09, -7.55479e-09, -5.768433e-09, -3.878792e-09, -2.759521e-09, 
    -1.674893e-09, -1.255321e-09, -1.222435e-09, -1.069741e-09, 
    -1.139758e-09, -1.442064e-09, -1.917165e-09, -2.653592e-09, 
    -3.513021e-09, -4.684846e-09,
  -1.572096e-08, -1.555733e-08, -1.459976e-08, -1.381906e-08, -1.404925e-08, 
    -1.411604e-08, -1.37573e-08, -1.333402e-08, -1.338816e-08, -1.37221e-08, 
    -1.408164e-08, -1.453707e-08, -1.48822e-08, -1.520427e-08, -1.536558e-08,
  -1.486287e-08, -1.439686e-08, -1.25583e-08, -1.256986e-08, -1.251098e-08, 
    -1.234476e-08, -1.171953e-08, -1.130181e-08, -1.123436e-08, 
    -1.142648e-08, -1.183341e-08, -1.240569e-08, -1.308999e-08, 
    -1.372536e-08, -1.438615e-08,
  -1.418775e-08, -1.185108e-08, -1.127557e-08, -1.133805e-08, -1.079686e-08, 
    -9.566818e-09, -8.768152e-09, -8.287103e-09, -8.005894e-09, -7.87185e-09, 
    -7.783938e-09, -7.989046e-09, -8.601913e-09, -9.579268e-09, -1.075393e-08,
  -1.172757e-08, -1.01353e-08, -1.006521e-08, -9.753004e-09, -8.503827e-09, 
    -7.552323e-09, -6.977358e-09, -6.642343e-09, -6.366867e-09, 
    -6.083992e-09, -5.860838e-09, -5.868601e-09, -6.002946e-09, 
    -6.335853e-09, -7.052231e-09,
  -9.844774e-09, -9.419193e-09, -9.180093e-09, -8.307289e-09, -7.283448e-09, 
    -6.764608e-09, -6.43842e-09, -6.142984e-09, -5.777514e-09, -5.779333e-09, 
    -5.928321e-09, -6.101311e-09, -6.10387e-09, -6.075869e-09, -6.13593e-09,
  -8.568108e-09, -8.465402e-09, -7.884043e-09, -7.252876e-09, -6.402863e-09, 
    -6.237237e-09, -5.558209e-09, -4.988039e-09, -4.569093e-09, 
    -4.780177e-09, -5.345366e-09, -5.723225e-09, -6.037088e-09, 
    -6.154622e-09, -6.182049e-09,
  -7.456316e-09, -7.64632e-09, -7.272609e-09, -6.120382e-09, -5.875019e-09, 
    -5.591607e-09, -4.455478e-09, -3.622195e-09, -3.273648e-09, 
    -4.329881e-09, -5.269091e-09, -5.770445e-09, -5.822453e-09, -5.76376e-09, 
    -5.707995e-09,
  -6.539315e-09, -6.847912e-09, -6.079203e-09, -5.365539e-09, -5.610729e-09, 
    -5.216589e-09, -2.990422e-09, -2.684883e-09, -3.618595e-09, 
    -4.981878e-09, -5.47015e-09, -5.567099e-09, -5.225388e-09, -4.86677e-09, 
    -4.553042e-09,
  -5.84427e-09, -6.171161e-09, -5.375548e-09, -5.073405e-09, -4.721409e-09, 
    -3.91518e-09, -2.270223e-09, -2.751527e-09, -3.960357e-09, -4.867448e-09, 
    -5.036501e-09, -4.805024e-09, -4.446101e-09, -4.133616e-09, -3.978501e-09,
  -5.114581e-09, -5.415784e-09, -4.955193e-09, -4.486863e-09, -3.872934e-09, 
    -3.214689e-09, -2.656871e-09, -3.188563e-09, -2.959545e-09, -2.98261e-09, 
    -2.961856e-09, -3.011228e-09, -3.119523e-09, -3.175739e-09, -3.320646e-09,
  -1.136288e-08, -1.0195e-08, -8.661062e-09, -7.021917e-09, -5.62639e-09, 
    -4.715581e-09, -4.109456e-09, -3.729369e-09, -3.384667e-09, 
    -3.211992e-09, -3.138091e-09, -3.19612e-09, -3.393951e-09, -3.733332e-09, 
    -4.269934e-09,
  -9.793895e-09, -7.642367e-09, -6.047635e-09, -4.712758e-09, -3.501029e-09, 
    -2.67989e-09, -2.643569e-09, -2.712866e-09, -2.63389e-09, -2.420169e-09, 
    -2.227275e-09, -2.210971e-09, -2.244601e-09, -2.424729e-09, -2.645058e-09,
  -8.078402e-09, -5.857775e-09, -4.314324e-09, -2.950649e-09, -2.208819e-09, 
    -1.481917e-09, -1.846346e-09, -1.851765e-09, -1.629803e-09, 
    -1.408967e-09, -1.371219e-09, -1.446508e-09, -1.574647e-09, 
    -1.714964e-09, -1.710242e-09,
  -7.449294e-09, -5.089006e-09, -3.624411e-09, -2.600772e-09, -2.523074e-09, 
    -2.641996e-09, -3.00359e-09, -1.74356e-09, -8.634807e-10, -6.870017e-10, 
    -8.154182e-10, -1.148525e-09, -1.488654e-09, -1.790876e-09, -1.983914e-09,
  -7.884649e-09, -4.97049e-09, -4.339737e-09, -3.429647e-09, -2.874175e-09, 
    -2.976649e-09, -2.224547e-09, -1.243441e-09, -6.958056e-10, 
    -5.818674e-10, -6.424583e-10, -7.974439e-10, -1.052724e-09, -1.36814e-09, 
    -1.788232e-09,
  -8.095037e-09, -5.390531e-09, -4.196124e-09, -3.508704e-09, -2.205195e-09, 
    -1.400543e-09, -1.072651e-09, -7.582516e-10, -6.314624e-10, 
    -7.619514e-10, -9.191435e-10, -1.062091e-09, -9.607318e-10, 
    -8.243079e-10, -8.478227e-10,
  -8.638709e-09, -5.779119e-09, -3.84007e-09, -2.890107e-09, -1.81258e-09, 
    -7.777126e-10, -7.419859e-10, -9.9261e-10, -1.461691e-09, -2.348561e-09, 
    -2.839425e-09, -3.250411e-09, -3.134035e-09, -2.690712e-09, -1.943224e-09,
  -9.208961e-09, -6.427634e-09, -3.833619e-09, -2.777991e-09, -1.595187e-09, 
    -1.49131e-09, -1.431937e-09, -1.240261e-09, -2.036571e-09, -3.103434e-09, 
    -3.973963e-09, -4.307472e-09, -4.502033e-09, -4.607803e-09, -4.629759e-09,
  -9.655598e-09, -7.067301e-09, -4.484947e-09, -3.495044e-09, -2.164564e-09, 
    -2.233707e-09, -1.909891e-09, -2.003008e-09, -2.469454e-09, 
    -2.817504e-09, -2.75087e-09, -2.684188e-09, -2.743099e-09, -2.808264e-09, 
    -2.928331e-09,
  -9.685585e-09, -7.547293e-09, -5.156371e-09, -4.006418e-09, -3.513535e-09, 
    -2.396626e-09, -2.438332e-09, -2.675531e-09, -2.512383e-09, 
    -2.046868e-09, -1.916573e-09, -2.05709e-09, -2.051596e-09, -2.117103e-09, 
    -2.0508e-09,
  -5.815392e-09, -4.903367e-09, -4.850742e-09, -5.001666e-09, -5.188558e-09, 
    -5.157399e-09, -5.902275e-09, -5.135979e-09, -4.127466e-09, 
    -3.489815e-09, -3.03079e-09, -2.767198e-09, -2.555234e-09, -2.437256e-09, 
    -2.342223e-09,
  -7.653163e-09, -6.287805e-09, -6.472627e-09, -6.640949e-09, -6.171786e-09, 
    -6.283893e-09, -6.436339e-09, -5.21692e-09, -4.269419e-09, -3.52437e-09, 
    -2.998706e-09, -2.75943e-09, -2.572339e-09, -2.418899e-09, -2.316625e-09,
  -9.371746e-09, -8.927494e-09, -8.6268e-09, -7.556695e-09, -7.686956e-09, 
    -6.96665e-09, -6.616859e-09, -4.986423e-09, -3.734955e-09, -3.041239e-09, 
    -2.714728e-09, -2.606172e-09, -2.50624e-09, -2.345306e-09, -2.160122e-09,
  -1.024248e-08, -1.017692e-08, -1.006358e-08, -8.816556e-09, -7.926435e-09, 
    -6.750532e-09, -5.745148e-09, -4.379474e-09, -3.465515e-09, 
    -2.898811e-09, -2.670381e-09, -2.569551e-09, -2.440672e-09, 
    -2.329622e-09, -2.22241e-09,
  -1.014627e-08, -9.908863e-09, -9.735549e-09, -8.833818e-09, -7.493701e-09, 
    -6.544512e-09, -5.312754e-09, -4.006564e-09, -3.119265e-09, 
    -2.676215e-09, -2.58304e-09, -2.564865e-09, -2.569607e-09, -2.535994e-09, 
    -2.436789e-09,
  -9.871568e-09, -9.369815e-09, -8.976468e-09, -8.636829e-09, -7.98955e-09, 
    -6.938638e-09, -5.412362e-09, -3.897835e-09, -2.998569e-09, 
    -2.766622e-09, -2.707397e-09, -2.71032e-09, -2.670242e-09, -2.56584e-09, 
    -2.484457e-09,
  -8.561386e-09, -8.558642e-09, -8.662409e-09, -8.918313e-09, -8.346759e-09, 
    -7.035351e-09, -5.338177e-09, -3.695935e-09, -2.857924e-09, 
    -2.812493e-09, -2.916963e-09, -3.043041e-09, -3.023613e-09, -2.79003e-09, 
    -2.57754e-09,
  -7.627048e-09, -8.305417e-09, -8.945719e-09, -9.17917e-09, -8.504019e-09, 
    -7.083381e-09, -5.27832e-09, -3.477534e-09, -2.71806e-09, -2.807827e-09, 
    -3.092598e-09, -3.304056e-09, -3.183664e-09, -2.90873e-09, -2.741875e-09,
  -7.834e-09, -8.922016e-09, -9.098313e-09, -9.024455e-09, -8.231685e-09, 
    -6.829869e-09, -5.00405e-09, -3.19447e-09, -2.598486e-09, -2.808312e-09, 
    -3.169611e-09, -3.140198e-09, -2.749167e-09, -2.55717e-09, -2.712465e-09,
  -8.792383e-09, -9.284206e-09, -9.185588e-09, -8.839694e-09, -8.017249e-09, 
    -6.552635e-09, -4.631579e-09, -2.902229e-09, -2.532901e-09, 
    -3.040313e-09, -3.13021e-09, -2.929964e-09, -2.478407e-09, -2.411129e-09, 
    -2.603446e-09,
  -3.22893e-10, -4.743129e-10, -6.595105e-10, -8.967158e-10, -1.167132e-09, 
    -1.563073e-09, -2.009418e-09, -2.54981e-09, -3.059506e-09, -3.441652e-09, 
    -3.710087e-09, -3.810944e-09, -3.829895e-09, -3.828275e-09, -3.806695e-09,
  -4.42086e-10, -5.459309e-10, -7.159679e-10, -9.80668e-10, -1.431193e-09, 
    -1.939783e-09, -2.526107e-09, -3.119695e-09, -3.660238e-09, 
    -4.071301e-09, -4.300605e-09, -4.352006e-09, -4.350282e-09, 
    -4.314085e-09, -4.31481e-09,
  -6.073702e-10, -7.69893e-10, -9.628641e-10, -1.34921e-09, -1.910846e-09, 
    -2.527467e-09, -3.158652e-09, -3.823989e-09, -4.408186e-09, 
    -4.808774e-09, -4.965649e-09, -4.998897e-09, -4.96623e-09, -4.897666e-09, 
    -4.804491e-09,
  -8.103096e-10, -1.087664e-09, -1.421408e-09, -2.06136e-09, -2.777633e-09, 
    -3.431945e-09, -4.067799e-09, -4.676498e-09, -5.143278e-09, 
    -5.504125e-09, -5.570583e-09, -5.505778e-09, -5.40354e-09, -5.294371e-09, 
    -5.148721e-09,
  -1.057541e-09, -1.493922e-09, -2.105252e-09, -2.881124e-09, -3.654809e-09, 
    -4.399145e-09, -5.048621e-09, -5.713104e-09, -6.114219e-09, -6.30501e-09, 
    -6.207445e-09, -6.007579e-09, -5.727603e-09, -5.501522e-09, -5.250888e-09,
  -1.281437e-09, -2.012778e-09, -2.803642e-09, -3.658226e-09, -4.458251e-09, 
    -5.325821e-09, -5.998522e-09, -6.619488e-09, -6.844672e-09, 
    -6.703895e-09, -6.32443e-09, -5.965566e-09, -5.665884e-09, -5.441971e-09, 
    -5.258368e-09,
  -1.609358e-09, -2.652276e-09, -3.574655e-09, -4.421853e-09, -5.233896e-09, 
    -6.132157e-09, -6.751455e-09, -7.229526e-09, -7.168841e-09, 
    -6.761164e-09, -6.205253e-09, -5.778367e-09, -5.48314e-09, -5.329073e-09, 
    -5.206377e-09,
  -2.09987e-09, -3.467663e-09, -4.368032e-09, -5.095891e-09, -5.912119e-09, 
    -6.634287e-09, -7.158331e-09, -7.472578e-09, -7.110394e-09, 
    -6.502798e-09, -5.820999e-09, -5.464597e-09, -5.288481e-09, 
    -5.122313e-09, -4.822241e-09,
  -2.782286e-09, -4.343137e-09, -5.242605e-09, -5.719257e-09, -6.497988e-09, 
    -7.026626e-09, -7.52759e-09, -7.74804e-09, -6.993515e-09, -5.99461e-09, 
    -5.427293e-09, -5.14176e-09, -4.797145e-09, -4.282852e-09, -3.953547e-09,
  -3.522544e-09, -5.165478e-09, -6.124822e-09, -6.457332e-09, -7.232256e-09, 
    -7.466934e-09, -8.276328e-09, -7.722917e-09, -6.21142e-09, -5.231517e-09, 
    -4.853077e-09, -4.416926e-09, -3.992517e-09, -3.535968e-09, -3.26182e-09,
  -1.512486e-09, -2.096628e-09, -2.473529e-09, -2.541998e-09, -2.538348e-09, 
    -2.657039e-09, -2.898273e-09, -3.60687e-09, -4.759324e-09, -6.480534e-09, 
    -8.750022e-09, -1.169198e-08, -1.435867e-08, -1.519328e-08, -1.531889e-08,
  -8.675068e-10, -1.20385e-09, -1.74484e-09, -2.317101e-09, -2.530565e-09, 
    -2.62814e-09, -2.795777e-09, -3.128634e-09, -3.543584e-09, -4.115901e-09, 
    -4.925797e-09, -6.040203e-09, -7.89717e-09, -1.035505e-08, -1.25242e-08,
  -6.934218e-10, -6.691113e-10, -1.035426e-09, -1.498051e-09, -1.960143e-09, 
    -2.315002e-09, -2.557962e-09, -2.646564e-09, -2.808986e-09, 
    -3.251562e-09, -3.779075e-09, -4.34762e-09, -4.88665e-09, -5.871315e-09, 
    -7.300518e-09,
  -5.357008e-10, -4.026406e-10, -4.752642e-10, -7.5465e-10, -1.158284e-09, 
    -1.437809e-09, -1.785967e-09, -2.095509e-09, -2.300468e-09, 
    -2.479937e-09, -2.737946e-09, -3.137417e-09, -3.585306e-09, -4.2163e-09, 
    -4.953331e-09,
  -6.039634e-10, -4.637573e-10, -3.827995e-10, -3.993082e-10, -5.853316e-10, 
    -8.071782e-10, -9.700013e-10, -1.18795e-09, -1.474784e-09, -1.834403e-09, 
    -2.106355e-09, -2.285865e-09, -2.578148e-09, -3.02812e-09, -3.594221e-09,
  -6.230755e-10, -5.375493e-10, -4.276023e-10, -3.399058e-10, -3.402383e-10, 
    -4.248288e-10, -5.511533e-10, -6.597795e-10, -8.381426e-10, 
    -1.039994e-09, -1.287449e-09, -1.52691e-09, -1.711081e-09, -1.960468e-09, 
    -2.308999e-09,
  -6.561172e-10, -5.534293e-10, -4.778959e-10, -4.162138e-10, -3.466806e-10, 
    -3.193513e-10, -3.453472e-10, -3.866927e-10, -4.696064e-10, 
    -5.767027e-10, -6.971952e-10, -8.707293e-10, -1.089289e-09, 
    -1.274854e-09, -1.488064e-09,
  -7.347967e-10, -6.639397e-10, -5.645202e-10, -5.014703e-10, -4.486355e-10, 
    -3.89107e-10, -3.682712e-10, -3.535763e-10, -3.746142e-10, -4.185853e-10, 
    -4.893308e-10, -5.850735e-10, -7.264648e-10, -9.305831e-10, -1.223014e-09,
  -8.490667e-10, -7.920176e-10, -7.057489e-10, -6.000344e-10, -5.366057e-10, 
    -4.740804e-10, -4.366817e-10, -4.160942e-10, -4.302262e-10, 
    -4.702363e-10, -5.717114e-10, -7.891761e-10, -1.078425e-09, 
    -1.410599e-09, -1.715028e-09,
  -9.852561e-10, -8.823356e-10, -7.86449e-10, -6.749808e-10, -6.035213e-10, 
    -5.498443e-10, -5.36257e-10, -5.663737e-10, -7.098402e-10, -1.014571e-09, 
    -1.356568e-09, -1.600517e-09, -1.796513e-09, -1.991544e-09, -2.149137e-09,
  -4.518257e-09, -6.233349e-09, -7.518103e-09, -8.019904e-09, -7.872136e-09, 
    -7.599703e-09, -7.799779e-09, -8.156293e-09, -8.789444e-09, 
    -9.431258e-09, -9.777044e-09, -1.039968e-08, -1.092894e-08, 
    -1.127121e-08, -1.19277e-08,
  -3.437808e-09, -4.671779e-09, -6.362963e-09, -7.553287e-09, -8.015687e-09, 
    -7.908181e-09, -7.71549e-09, -7.667968e-09, -7.423075e-09, -7.802318e-09, 
    -8.665957e-09, -9.212251e-09, -1.015592e-08, -1.162478e-08, -1.280994e-08,
  -2.472174e-09, -3.584977e-09, -5.109905e-09, -6.666699e-09, -7.635909e-09, 
    -8.078099e-09, -8.051624e-09, -7.899024e-09, -7.743868e-09, 
    -7.346657e-09, -7.367154e-09, -7.726698e-09, -8.38573e-09, -9.39867e-09, 
    -1.114816e-08,
  -1.699927e-09, -2.49392e-09, -3.86858e-09, -5.503579e-09, -6.903568e-09, 
    -7.704696e-09, -8.093902e-09, -8.118782e-09, -8.257355e-09, 
    -7.963552e-09, -7.575402e-09, -7.32109e-09, -7.541098e-09, -8.001214e-09, 
    -8.917312e-09,
  -1.213688e-09, -1.790922e-09, -2.717262e-09, -4.218258e-09, -5.722948e-09, 
    -6.948029e-09, -7.622925e-09, -7.926309e-09, -8.03303e-09, -8.372007e-09, 
    -8.528968e-09, -8.037403e-09, -7.615069e-09, -7.876874e-09, -8.401167e-09,
  -9.488824e-10, -1.39773e-09, -2.04823e-09, -3.185773e-09, -4.683045e-09, 
    -5.956446e-09, -6.999608e-09, -7.434267e-09, -7.616966e-09, 
    -7.813828e-09, -8.241418e-09, -8.443063e-09, -8.472954e-09, 
    -8.350169e-09, -8.712417e-09,
  -8.785093e-10, -1.131225e-09, -1.504489e-09, -2.374301e-09, -3.651361e-09, 
    -4.995919e-09, -6.12959e-09, -6.90865e-09, -7.110601e-09, -7.232867e-09, 
    -7.503837e-09, -7.805349e-09, -8.091676e-09, -8.401856e-09, -8.882712e-09,
  -8.035298e-10, -9.671058e-10, -1.164226e-09, -1.737258e-09, -2.814961e-09, 
    -4.060873e-09, -5.20607e-09, -6.139053e-09, -6.621372e-09, -6.711262e-09, 
    -6.854278e-09, -7.082435e-09, -7.44909e-09, -7.870696e-09, -8.392351e-09,
  -7.138801e-10, -8.367007e-10, -9.610419e-10, -1.384289e-09, -2.22603e-09, 
    -3.336464e-09, -4.477931e-09, -5.331036e-09, -5.978325e-09, 
    -6.212031e-09, -6.192047e-09, -6.375878e-09, -6.785197e-09, 
    -7.142906e-09, -7.6921e-09,
  -6.999023e-10, -7.97542e-10, -8.863068e-10, -1.223379e-09, -1.915251e-09, 
    -2.886077e-09, -3.919497e-09, -4.759892e-09, -5.293329e-09, 
    -5.647191e-09, -5.677542e-09, -5.803594e-09, -6.261391e-09, 
    -6.737861e-09, -7.207905e-09,
  -2.658055e-09, -2.981434e-09, -3.399782e-09, -3.761708e-09, -4.152148e-09, 
    -4.586673e-09, -5.30457e-09, -6.181107e-09, -6.767825e-09, -7.103344e-09, 
    -7.163234e-09, -6.905324e-09, -6.463297e-09, -5.923855e-09, -5.405355e-09,
  -2.36048e-09, -2.592236e-09, -3.051249e-09, -3.47618e-09, -3.886926e-09, 
    -4.313325e-09, -4.762275e-09, -5.549611e-09, -6.5786e-09, -7.079088e-09, 
    -7.228945e-09, -7.263249e-09, -7.046972e-09, -6.593243e-09, -5.940882e-09,
  -2.141781e-09, -2.374261e-09, -2.675045e-09, -3.238026e-09, -3.647518e-09, 
    -4.035526e-09, -4.394137e-09, -4.930373e-09, -5.991981e-09, -6.89021e-09, 
    -7.277856e-09, -7.506097e-09, -7.456484e-09, -7.234849e-09, -6.599156e-09,
  -1.901605e-09, -2.202653e-09, -2.460512e-09, -2.933474e-09, -3.436813e-09, 
    -3.814331e-09, -4.162686e-09, -4.600613e-09, -5.399742e-09, -6.50922e-09, 
    -7.193221e-09, -7.594411e-09, -7.796818e-09, -7.611155e-09, -6.907653e-09,
  -1.782953e-09, -2.047477e-09, -2.320506e-09, -2.704794e-09, -3.204766e-09, 
    -3.564421e-09, -3.916558e-09, -4.282561e-09, -5.001034e-09, -6.07452e-09, 
    -7.003996e-09, -7.623764e-09, -7.846745e-09, -7.597883e-09, -6.87943e-09,
  -1.730411e-09, -1.942022e-09, -2.221343e-09, -2.553042e-09, -2.947402e-09, 
    -3.353785e-09, -3.730818e-09, -4.144515e-09, -4.661632e-09, 
    -5.651186e-09, -6.645971e-09, -7.427652e-09, -7.593401e-09, -7.42123e-09, 
    -6.834147e-09,
  -1.651897e-09, -1.842667e-09, -2.186825e-09, -2.447914e-09, -2.723785e-09, 
    -3.15732e-09, -3.536877e-09, -4.068313e-09, -4.563678e-09, -5.345353e-09, 
    -6.312983e-09, -7.207112e-09, -7.476564e-09, -7.284829e-09, -6.761034e-09,
  -1.65272e-09, -1.832289e-09, -2.117326e-09, -2.307675e-09, -2.596151e-09, 
    -3.03928e-09, -3.417638e-09, -3.983992e-09, -4.476336e-09, -5.150465e-09, 
    -6.018852e-09, -6.962909e-09, -7.26299e-09, -7.148683e-09, -6.694019e-09,
  -1.641527e-09, -1.814132e-09, -2.034511e-09, -2.238794e-09, -2.509643e-09, 
    -2.941533e-09, -3.356515e-09, -3.901951e-09, -4.368792e-09, 
    -4.891013e-09, -5.822863e-09, -6.794454e-09, -7.147905e-09, 
    -7.028881e-09, -6.603651e-09,
  -1.601731e-09, -1.74654e-09, -1.924128e-09, -2.138789e-09, -2.47772e-09, 
    -2.920133e-09, -3.2209e-09, -3.767611e-09, -4.364156e-09, -4.86527e-09, 
    -5.777165e-09, -6.850839e-09, -7.188538e-09, -7.038998e-09, -6.581383e-09,
  -4.790868e-10, -5.028017e-10, -5.17108e-10, -5.47871e-10, -5.982596e-10, 
    -6.803715e-10, -7.720471e-10, -8.748994e-10, -9.45881e-10, -1.070939e-09, 
    -1.339728e-09, -1.718629e-09, -2.067599e-09, -2.340537e-09, -2.492899e-09,
  -3.694812e-10, -3.633821e-10, -3.794529e-10, -4.276358e-10, -4.835048e-10, 
    -5.794679e-10, -6.965779e-10, -8.171117e-10, -9.550835e-10, -1.21353e-09, 
    -1.645036e-09, -2.129231e-09, -2.466883e-09, -2.827546e-09, -3.194221e-09,
  -3.195885e-10, -3.177727e-10, -3.412971e-10, -4.199897e-10, -4.620155e-10, 
    -5.808234e-10, -7.410284e-10, -8.920342e-10, -1.109111e-09, 
    -1.529663e-09, -2.1334e-09, -2.551793e-09, -3.082157e-09, -4.241116e-09, 
    -4.817224e-09,
  -3.422541e-10, -3.22097e-10, -3.313985e-10, -4.457648e-10, -5.574951e-10, 
    -6.666852e-10, -8.649261e-10, -1.093687e-09, -1.440787e-09, 
    -1.964156e-09, -2.531923e-09, -3.759695e-09, -5.460298e-09, 
    -6.372225e-09, -6.175235e-09,
  -4.0014e-10, -4.30114e-10, -4.60979e-10, -5.730733e-10, -6.973969e-10, 
    -9.37893e-10, -1.256259e-09, -1.481887e-09, -1.838092e-09, -2.699395e-09, 
    -4.272605e-09, -6.156109e-09, -6.870909e-09, -7.254591e-09, -6.98991e-09,
  -5.986562e-10, -6.232941e-10, -6.7045e-10, -8.475255e-10, -1.133484e-09, 
    -1.392451e-09, -1.623293e-09, -1.975894e-09, -2.900976e-09, 
    -4.719765e-09, -6.574794e-09, -7.663363e-09, -8.042108e-09, 
    -8.208485e-09, -7.909807e-09,
  -8.493635e-10, -8.878111e-10, -1.052379e-09, -1.330335e-09, -1.597945e-09, 
    -1.903361e-09, -2.405556e-09, -3.43847e-09, -5.064035e-09, -7.162374e-09, 
    -8.238782e-09, -8.902918e-09, -9.403001e-09, -9.740718e-09, -8.925438e-09,
  -1.302821e-09, -1.426153e-09, -1.61015e-09, -1.949214e-09, -2.268316e-09, 
    -2.813395e-09, -3.805803e-09, -5.306442e-09, -7.143945e-09, 
    -8.369895e-09, -8.774634e-09, -9.70542e-09, -1.00409e-08, -9.641586e-09, 
    -8.975666e-09,
  -1.979249e-09, -2.206088e-09, -2.518071e-09, -2.805522e-09, -3.276537e-09, 
    -4.258759e-09, -5.571563e-09, -7.2351e-09, -8.62557e-09, -9.158468e-09, 
    -9.996544e-09, -9.741103e-09, -9.222053e-09, -8.341595e-09, -8.210574e-09,
  -2.913433e-09, -3.138716e-09, -3.314319e-09, -3.671488e-09, -4.278768e-09, 
    -5.51459e-09, -6.771219e-09, -8.326173e-09, -9.356846e-09, -9.956242e-09, 
    -9.887956e-09, -9.312555e-09, -8.419145e-09, -7.721445e-09, -7.364588e-09,
  -3.051526e-09, -3.121472e-09, -3.229434e-09, -3.377023e-09, -3.57744e-09, 
    -3.77054e-09, -3.888151e-09, -3.950912e-09, -3.981785e-09, -3.955707e-09, 
    -3.902526e-09, -3.796566e-09, -3.660189e-09, -3.488121e-09, -3.295662e-09,
  -2.230603e-09, -2.319613e-09, -2.42524e-09, -2.511048e-09, -2.601735e-09, 
    -2.694877e-09, -2.780555e-09, -2.82828e-09, -2.841518e-09, -2.837393e-09, 
    -2.82786e-09, -2.788466e-09, -2.716295e-09, -2.628011e-09, -2.537403e-09,
  -1.696021e-09, -1.788622e-09, -1.895152e-09, -1.975641e-09, -2.042614e-09, 
    -2.073246e-09, -2.088882e-09, -2.095444e-09, -2.0819e-09, -2.04662e-09, 
    -2.007134e-09, -1.969924e-09, -1.937515e-09, -1.907084e-09, -1.907611e-09,
  -1.248419e-09, -1.344968e-09, -1.417459e-09, -1.494194e-09, -1.545308e-09, 
    -1.574721e-09, -1.588071e-09, -1.574374e-09, -1.55308e-09, -1.549681e-09, 
    -1.536555e-09, -1.526411e-09, -1.563652e-09, -1.727785e-09, -2.164253e-09,
  -1.030995e-09, -1.072115e-09, -1.124825e-09, -1.156888e-09, -1.176228e-09, 
    -1.189265e-09, -1.206726e-09, -1.218217e-09, -1.221737e-09, 
    -1.231052e-09, -1.248011e-09, -1.422798e-09, -1.7888e-09, -2.475324e-09, 
    -3.132593e-09,
  -9.563244e-10, -9.568094e-10, -9.498015e-10, -9.332356e-10, -9.273247e-10, 
    -9.263803e-10, -9.465355e-10, -9.672461e-10, -9.813439e-10, 
    -1.033613e-09, -1.273352e-09, -1.87799e-09, -2.601978e-09, -3.40066e-09, 
    -3.904772e-09,
  -8.580305e-10, -8.787894e-10, -8.609336e-10, -8.199045e-10, -8.288544e-10, 
    -8.126707e-10, -8.05372e-10, -8.391381e-10, -1.047212e-09, -1.542819e-09, 
    -2.248773e-09, -3.213296e-09, -3.98536e-09, -4.559034e-09, -5.016028e-09,
  -8.566937e-10, -8.402897e-10, -8.000067e-10, -7.862815e-10, -7.625854e-10, 
    -7.384789e-10, -8.016162e-10, -1.23457e-09, -2.177453e-09, -3.216656e-09, 
    -4.111895e-09, -5.035224e-09, -5.396995e-09, -5.576947e-09, -5.548111e-09,
  -7.846612e-10, -7.848531e-10, -7.545516e-10, -6.76221e-10, -6.704793e-10, 
    -8.88974e-10, -1.797564e-09, -3.415294e-09, -4.73e-09, -5.363632e-09, 
    -5.841986e-09, -5.90255e-09, -5.901148e-09, -6.051267e-09, -6.139487e-09,
  -7.159193e-10, -7.16487e-10, -7.565114e-10, -8.989211e-10, -1.594738e-09, 
    -3.108778e-09, -5.35669e-09, -6.65028e-09, -6.699951e-09, -6.816502e-09, 
    -6.929003e-09, -6.772559e-09, -6.747523e-09, -6.469933e-09, -6.248575e-09,
  -5.910977e-09, -6.285394e-09, -6.987303e-09, -8.561743e-09, -1.063386e-08, 
    -1.240247e-08, -1.345408e-08, -1.398962e-08, -1.415836e-08, 
    -1.409719e-08, -1.430199e-08, -1.475945e-08, -1.529137e-08, 
    -1.576194e-08, -1.612693e-08,
  -5.554096e-09, -5.794678e-09, -6.092494e-09, -6.501764e-09, -7.56805e-09, 
    -9.290582e-09, -1.11283e-08, -1.23306e-08, -1.307122e-08, -1.345617e-08, 
    -1.36116e-08, -1.367691e-08, -1.393304e-08, -1.420589e-08, -1.448596e-08,
  -5.112797e-09, -5.458891e-09, -5.699658e-09, -5.940945e-09, -6.236014e-09, 
    -6.870635e-09, -8.08265e-09, -9.774944e-09, -1.114486e-08, -1.198489e-08, 
    -1.24678e-08, -1.266107e-08, -1.271023e-08, -1.276379e-08, -1.28319e-08,
  -3.955637e-09, -4.615782e-09, -5.106078e-09, -5.488321e-09, -5.767334e-09, 
    -6.061055e-09, -6.471934e-09, -7.178514e-09, -8.469319e-09, 
    -9.745158e-09, -1.06221e-08, -1.117775e-08, -1.14344e-08, -1.151179e-08, 
    -1.147649e-08,
  -3.047596e-09, -3.494031e-09, -4.03578e-09, -4.621693e-09, -5.082542e-09, 
    -5.428796e-09, -5.749135e-09, -6.06184e-09, -6.472748e-09, -7.252436e-09, 
    -8.23562e-09, -9.066328e-09, -9.583839e-09, -9.830648e-09, -9.916056e-09,
  -2.531218e-09, -2.723354e-09, -3.065331e-09, -3.478588e-09, -4.027643e-09, 
    -4.56786e-09, -5.006093e-09, -5.351511e-09, -5.631429e-09, -5.933162e-09, 
    -6.370501e-09, -7.036458e-09, -7.677685e-09, -8.12294e-09, -8.303157e-09,
  -2.150292e-09, -2.338423e-09, -2.521038e-09, -2.760148e-09, -3.077834e-09, 
    -3.477124e-09, -3.964103e-09, -4.441179e-09, -4.836862e-09, 
    -5.130314e-09, -5.371466e-09, -5.644556e-09, -6.042234e-09, 
    -6.476511e-09, -6.743468e-09,
  -1.946996e-09, -2.048705e-09, -2.159262e-09, -2.318335e-09, -2.493746e-09, 
    -2.753016e-09, -3.120838e-09, -3.58309e-09, -4.055514e-09, -4.381614e-09, 
    -4.571555e-09, -4.727677e-09, -4.888819e-09, -5.097436e-09, -5.34351e-09,
  -1.829862e-09, -1.913997e-09, -1.986807e-09, -2.105604e-09, -2.24414e-09, 
    -2.412589e-09, -2.587642e-09, -2.855812e-09, -3.142566e-09, 
    -3.504065e-09, -3.779622e-09, -3.991323e-09, -4.139086e-09, 
    -4.283653e-09, -4.393566e-09,
  -1.660161e-09, -1.715694e-09, -1.780291e-09, -1.85928e-09, -1.950927e-09, 
    -2.054675e-09, -2.153057e-09, -2.2702e-09, -2.384777e-09, -2.598773e-09, 
    -2.879173e-09, -3.122189e-09, -3.289719e-09, -3.434906e-09, -3.545852e-09,
  -9.63739e-09, -1.068209e-08, -1.240581e-08, -1.413119e-08, -1.578361e-08, 
    -1.681877e-08, -1.65604e-08, -1.557672e-08, -1.30815e-08, -1.164149e-08, 
    -1.183334e-08, -1.276294e-08, -1.416885e-08, -1.624287e-08, -1.824977e-08,
  -8.742016e-09, -9.294955e-09, -1.03244e-08, -1.172462e-08, -1.333324e-08, 
    -1.550017e-08, -1.650157e-08, -1.655051e-08, -1.605362e-08, 
    -1.440374e-08, -1.23514e-08, -1.20328e-08, -1.258556e-08, -1.38488e-08, 
    -1.564255e-08,
  -7.655947e-09, -8.305564e-09, -8.95366e-09, -9.848642e-09, -1.110343e-08, 
    -1.267362e-08, -1.484167e-08, -1.636434e-08, -1.660518e-08, 
    -1.586652e-08, -1.464963e-08, -1.265948e-08, -1.214037e-08, 
    -1.248211e-08, -1.347082e-08,
  -6.205205e-09, -6.991246e-09, -7.803652e-09, -8.534038e-09, -9.348237e-09, 
    -1.04301e-08, -1.188387e-08, -1.380935e-08, -1.606358e-08, -1.692723e-08, 
    -1.633919e-08, -1.525714e-08, -1.31242e-08, -1.234902e-08, -1.239686e-08,
  -4.971126e-09, -5.482176e-09, -6.171398e-09, -7.115652e-09, -8.009703e-09, 
    -8.88923e-09, -9.811179e-09, -1.111649e-08, -1.261738e-08, -1.505023e-08, 
    -1.646694e-08, -1.656363e-08, -1.582815e-08, -1.38194e-08, -1.279974e-08,
  -4.338032e-09, -4.572194e-09, -4.897588e-09, -5.399758e-09, -6.225423e-09, 
    -7.201458e-09, -8.309983e-09, -9.340637e-09, -1.062543e-08, -1.19254e-08, 
    -1.41491e-08, -1.561439e-08, -1.640926e-08, -1.618086e-08, -1.451424e-08,
  -3.91995e-09, -4.089139e-09, -4.299704e-09, -4.565622e-09, -4.917077e-09, 
    -5.47877e-09, -6.265223e-09, -7.342368e-09, -8.572422e-09, -9.955044e-09, 
    -1.133175e-08, -1.32326e-08, -1.478497e-08, -1.597335e-08, -1.606726e-08,
  -3.588233e-09, -3.710384e-09, -3.85142e-09, -4.040607e-09, -4.297411e-09, 
    -4.599662e-09, -5.046447e-09, -5.604347e-09, -6.43062e-09, -7.689635e-09, 
    -9.073632e-09, -1.050669e-08, -1.241359e-08, -1.397585e-08, -1.5335e-08,
  -3.250569e-09, -3.419663e-09, -3.550198e-09, -3.685244e-09, -3.843215e-09, 
    -4.074289e-09, -4.332322e-09, -4.753439e-09, -5.143387e-09, 
    -5.755026e-09, -6.809996e-09, -8.006665e-09, -9.649444e-09, 
    -1.141579e-08, -1.310625e-08,
  -3.008783e-09, -3.1792e-09, -3.334705e-09, -3.462844e-09, -3.593281e-09, 
    -3.746307e-09, -3.939755e-09, -4.139826e-09, -4.493885e-09, 
    -4.803031e-09, -5.336093e-09, -6.018389e-09, -7.218854e-09, 
    -8.729321e-09, -1.039263e-08,
  -9.848045e-09, -9.993332e-09, -1.015708e-08, -1.035096e-08, -1.072972e-08, 
    -1.139582e-08, -1.275047e-08, -1.457402e-08, -1.625338e-08, 
    -1.875375e-08, -2.203093e-08, -2.348099e-08, -2.356076e-08, 
    -2.329058e-08, -2.336819e-08,
  -9.59792e-09, -9.809891e-09, -1.001077e-08, -1.021281e-08, -1.044645e-08, 
    -1.074367e-08, -1.110474e-08, -1.188382e-08, -1.331522e-08, 
    -1.484997e-08, -1.749656e-08, -2.021826e-08, -2.20078e-08, -2.304307e-08, 
    -2.325139e-08,
  -9.668454e-09, -9.766274e-09, -9.859847e-09, -1.0057e-08, -1.020233e-08, 
    -1.039699e-08, -1.066053e-08, -1.087535e-08, -1.147258e-08, 
    -1.237976e-08, -1.388994e-08, -1.612819e-08, -1.885248e-08, 
    -2.067071e-08, -2.215289e-08,
  -9.02105e-09, -9.488391e-09, -9.834333e-09, -9.999557e-09, -1.016981e-08, 
    -1.031651e-08, -1.047278e-08, -1.064028e-08, -1.086618e-08, 
    -1.122575e-08, -1.184499e-08, -1.309034e-08, -1.507705e-08, 
    -1.753217e-08, -1.931837e-08,
  -8.213868e-09, -8.720302e-09, -9.242357e-09, -9.597447e-09, -9.916378e-09, 
    -1.019949e-08, -1.047035e-08, -1.068063e-08, -1.083595e-08, 
    -1.102402e-08, -1.124216e-08, -1.156933e-08, -1.246412e-08, 
    -1.404901e-08, -1.632626e-08,
  -7.466975e-09, -7.991404e-09, -8.485398e-09, -9.018037e-09, -9.47649e-09, 
    -9.831373e-09, -1.014676e-08, -1.049181e-08, -1.083424e-08, 
    -1.115065e-08, -1.129713e-08, -1.147736e-08, -1.166959e-08, 
    -1.217941e-08, -1.317256e-08,
  -6.545948e-09, -7.106577e-09, -7.65414e-09, -8.266513e-09, -8.861807e-09, 
    -9.401275e-09, -9.828686e-09, -1.006453e-08, -1.032341e-08, 
    -1.074055e-08, -1.12943e-08, -1.161987e-08, -1.183272e-08, -1.204435e-08, 
    -1.237207e-08,
  -5.64012e-09, -6.226883e-09, -6.777904e-09, -7.361747e-09, -8.060414e-09, 
    -8.636122e-09, -9.20491e-09, -9.657311e-09, -9.932521e-09, -1.016401e-08, 
    -1.055164e-08, -1.114695e-08, -1.165126e-08, -1.20693e-08, -1.239414e-08,
  -4.683385e-09, -5.158382e-09, -5.779397e-09, -6.366252e-09, -7.022556e-09, 
    -7.706662e-09, -8.239094e-09, -8.809383e-09, -9.33246e-09, -9.833881e-09, 
    -1.020418e-08, -1.050743e-08, -1.105016e-08, -1.157605e-08, -1.223503e-08,
  -3.840447e-09, -4.289485e-09, -4.761907e-09, -5.301033e-09, -5.883763e-09, 
    -6.500537e-09, -7.187765e-09, -7.718325e-09, -8.223022e-09, 
    -8.759324e-09, -9.361214e-09, -9.901937e-09, -1.038551e-08, 
    -1.084285e-08, -1.143602e-08,
  -1.466923e-08, -1.521222e-08, -1.58469e-08, -1.644857e-08, -1.723222e-08, 
    -1.835012e-08, -1.954829e-08, -2.079892e-08, -2.147455e-08, 
    -2.178096e-08, -2.208675e-08, -2.252478e-08, -2.289409e-08, 
    -2.270343e-08, -2.227137e-08,
  -1.221567e-08, -1.299016e-08, -1.373884e-08, -1.454858e-08, -1.53404e-08, 
    -1.608359e-08, -1.7004e-08, -1.802142e-08, -1.934809e-08, -2.044911e-08, 
    -2.104707e-08, -2.16772e-08, -2.254054e-08, -2.3143e-08, -2.33356e-08,
  -1.014017e-08, -1.086934e-08, -1.146043e-08, -1.220491e-08, -1.307692e-08, 
    -1.387515e-08, -1.474197e-08, -1.550753e-08, -1.641369e-08, 
    -1.752347e-08, -1.880794e-08, -1.996188e-08, -2.118322e-08, 
    -2.226767e-08, -2.300849e-08,
  -9.173122e-09, -9.704523e-09, -1.01609e-08, -1.058124e-08, -1.109375e-08, 
    -1.184998e-08, -1.272463e-08, -1.353737e-08, -1.436472e-08, 
    -1.512335e-08, -1.59877e-08, -1.705076e-08, -1.843692e-08, -2.03046e-08, 
    -2.193014e-08,
  -8.799931e-09, -9.146916e-09, -9.231139e-09, -9.414892e-09, -9.687932e-09, 
    -1.001694e-08, -1.065442e-08, -1.149484e-08, -1.247942e-08, -1.32814e-08, 
    -1.404376e-08, -1.484612e-08, -1.574149e-08, -1.699738e-08, -1.927712e-08,
  -8.444132e-09, -8.957275e-09, -9.021559e-09, -8.981326e-09, -8.941895e-09, 
    -9.066696e-09, -9.301095e-09, -9.717413e-09, -1.042408e-08, 
    -1.134621e-08, -1.22193e-08, -1.301111e-08, -1.384417e-08, -1.472813e-08, 
    -1.58735e-08,
  -7.23136e-09, -7.718971e-09, -8.16539e-09, -8.464726e-09, -8.626204e-09, 
    -8.775102e-09, -8.872567e-09, -8.988525e-09, -9.253044e-09, 
    -9.794417e-09, -1.050407e-08, -1.132775e-08, -1.220474e-08, 
    -1.314468e-08, -1.401896e-08,
  -6.169297e-09, -6.661775e-09, -7.021979e-09, -7.478079e-09, -7.925892e-09, 
    -8.318443e-09, -8.669859e-09, -8.93546e-09, -8.91152e-09, -8.964709e-09, 
    -9.294433e-09, -9.896395e-09, -1.049879e-08, -1.135219e-08, -1.237253e-08,
  -5.370312e-09, -5.735613e-09, -6.157865e-09, -6.582677e-09, -7.040994e-09, 
    -7.559206e-09, -8.106105e-09, -8.613878e-09, -9.081591e-09, 
    -9.157105e-09, -9.095634e-09, -9.223879e-09, -9.587038e-09, 
    -1.013897e-08, -1.076079e-08,
  -4.373896e-09, -4.768825e-09, -5.170742e-09, -5.624303e-09, -5.995097e-09, 
    -6.480991e-09, -7.080295e-09, -7.682107e-09, -8.211221e-09, 
    -8.789271e-09, -9.262716e-09, -9.404072e-09, -9.398078e-09, 
    -9.496852e-09, -9.826769e-09,
  -1.950137e-08, -1.969897e-08, -1.967526e-08, -1.949355e-08, -1.934498e-08, 
    -1.911933e-08, -1.936845e-08, -2.00569e-08, -2.134612e-08, -2.270698e-08, 
    -2.34312e-08, -2.385656e-08, -2.408076e-08, -2.450809e-08, -2.46325e-08,
  -1.920514e-08, -1.954939e-08, -1.97334e-08, -1.980097e-08, -1.97177e-08, 
    -1.948845e-08, -1.917292e-08, -1.914372e-08, -1.949605e-08, 
    -2.015148e-08, -2.133276e-08, -2.260595e-08, -2.317899e-08, 
    -2.356267e-08, -2.3815e-08,
  -1.747355e-08, -1.811124e-08, -1.8516e-08, -1.89056e-08, -1.920819e-08, 
    -1.943791e-08, -1.937483e-08, -1.906761e-08, -1.878685e-08, 
    -1.869802e-08, -1.912537e-08, -1.995572e-08, -2.122122e-08, 
    -2.233851e-08, -2.311898e-08,
  -1.400825e-08, -1.486206e-08, -1.546346e-08, -1.613827e-08, -1.66346e-08, 
    -1.710318e-08, -1.778857e-08, -1.830895e-08, -1.867597e-08, 
    -1.850014e-08, -1.847492e-08, -1.857911e-08, -1.920404e-08, 
    -2.014363e-08, -2.130698e-08,
  -1.114723e-08, -1.190788e-08, -1.2596e-08, -1.335606e-08, -1.41284e-08, 
    -1.486253e-08, -1.564341e-08, -1.642571e-08, -1.712479e-08, 
    -1.773553e-08, -1.808543e-08, -1.812238e-08, -1.827427e-08, 
    -1.854069e-08, -1.910361e-08,
  -9.23847e-09, -9.792036e-09, -1.040882e-08, -1.087711e-08, -1.130966e-08, 
    -1.221885e-08, -1.334836e-08, -1.45982e-08, -1.580343e-08, -1.664547e-08, 
    -1.715504e-08, -1.763054e-08, -1.777808e-08, -1.793415e-08, -1.817116e-08,
  -7.687018e-09, -8.210374e-09, -8.864e-09, -9.453005e-09, -9.719447e-09, 
    -9.892257e-09, -1.07817e-08, -1.170538e-08, -1.269339e-08, -1.389272e-08, 
    -1.49977e-08, -1.595508e-08, -1.645666e-08, -1.694462e-08, -1.734842e-08,
  -6.091073e-09, -6.792776e-09, -7.437729e-09, -8.083972e-09, -8.633258e-09, 
    -8.621472e-09, -8.88282e-09, -9.578591e-09, -1.023338e-08, -1.098548e-08, 
    -1.197354e-08, -1.313325e-08, -1.431769e-08, -1.510048e-08, -1.567313e-08,
  -4.524704e-09, -5.048839e-09, -5.672024e-09, -6.307546e-09, -6.939565e-09, 
    -7.326386e-09, -7.515265e-09, -7.94078e-09, -8.460762e-09, -8.978472e-09, 
    -9.621807e-09, -1.034104e-08, -1.126866e-08, -1.241566e-08, -1.346515e-08,
  -3.65796e-09, -3.898223e-09, -4.363825e-09, -4.862008e-09, -5.515972e-09, 
    -5.961112e-09, -6.275857e-09, -6.591638e-09, -6.973737e-09, 
    -7.518885e-09, -8.126546e-09, -8.797269e-09, -9.404029e-09, 
    -1.016041e-08, -1.099658e-08,
  -1.991876e-08, -1.969076e-08, -1.938609e-08, -1.93125e-08, -1.928785e-08, 
    -1.931658e-08, -1.944089e-08, -1.978382e-08, -2.022707e-08, 
    -2.086934e-08, -2.122492e-08, -2.133644e-08, -2.139754e-08, 
    -2.121828e-08, -2.069814e-08,
  -2.009393e-08, -1.999722e-08, -1.975226e-08, -1.947816e-08, -1.916136e-08, 
    -1.889402e-08, -1.86742e-08, -1.854581e-08, -1.845985e-08, -1.870876e-08, 
    -1.926088e-08, -1.993936e-08, -2.058577e-08, -2.09926e-08, -2.124921e-08,
  -1.937123e-08, -1.939141e-08, -1.937103e-08, -1.916875e-08, -1.889488e-08, 
    -1.857953e-08, -1.832726e-08, -1.799484e-08, -1.786795e-08, 
    -1.763031e-08, -1.766746e-08, -1.771048e-08, -1.828782e-08, 
    -1.919213e-08, -2.007156e-08,
  -1.705066e-08, -1.713591e-08, -1.729899e-08, -1.74636e-08, -1.754261e-08, 
    -1.745924e-08, -1.725485e-08, -1.698782e-08, -1.681223e-08, 
    -1.653244e-08, -1.641469e-08, -1.632564e-08, -1.646728e-08, -1.68188e-08, 
    -1.747614e-08,
  -1.332536e-08, -1.335697e-08, -1.351017e-08, -1.376434e-08, -1.410733e-08, 
    -1.438246e-08, -1.454526e-08, -1.494409e-08, -1.51277e-08, -1.536478e-08, 
    -1.531199e-08, -1.525642e-08, -1.52778e-08, -1.549036e-08, -1.584643e-08,
  -1.056393e-08, -1.059932e-08, -1.065186e-08, -1.072393e-08, -1.082583e-08, 
    -1.10114e-08, -1.140485e-08, -1.174312e-08, -1.216783e-08, -1.275435e-08, 
    -1.32849e-08, -1.387249e-08, -1.43117e-08, -1.467169e-08, -1.490757e-08,
  -8.494846e-09, -8.545681e-09, -8.581294e-09, -8.612269e-09, -8.708207e-09, 
    -8.782782e-09, -8.894663e-09, -8.87057e-09, -9.097707e-09, -9.885662e-09, 
    -1.072352e-08, -1.174671e-08, -1.265232e-08, -1.355858e-08, -1.419009e-08,
  -7.048687e-09, -6.93201e-09, -6.943177e-09, -7.092669e-09, -7.287556e-09, 
    -7.797428e-09, -8.007337e-09, -8.159343e-09, -8.454963e-09, 
    -8.949183e-09, -9.461449e-09, -1.039129e-08, -1.129311e-08, 
    -1.204536e-08, -1.265657e-08,
  -6.134164e-09, -5.993902e-09, -5.881878e-09, -5.86754e-09, -5.985703e-09, 
    -6.330197e-09, -6.84205e-09, -7.29987e-09, -7.650714e-09, -7.826898e-09, 
    -8.002581e-09, -8.333663e-09, -8.883445e-09, -9.537132e-09, -1.036388e-08,
  -5.461049e-09, -5.298438e-09, -5.13653e-09, -4.995448e-09, -4.93788e-09, 
    -4.937074e-09, -5.040067e-09, -5.14593e-09, -5.242186e-09, -5.344817e-09, 
    -5.453557e-09, -5.618357e-09, -5.957344e-09, -6.423013e-09, -7.025814e-09,
  -1.712993e-08, -1.713909e-08, -1.720832e-08, -1.729974e-08, -1.739824e-08, 
    -1.751169e-08, -1.764785e-08, -1.786361e-08, -1.813562e-08, 
    -1.853116e-08, -1.91072e-08, -1.948473e-08, -1.987885e-08, -2.016756e-08, 
    -2.018564e-08,
  -1.809727e-08, -1.81812e-08, -1.827727e-08, -1.839861e-08, -1.855133e-08, 
    -1.872651e-08, -1.892408e-08, -1.920998e-08, -1.946743e-08, 
    -1.989375e-08, -1.996507e-08, -2.01344e-08, -2.019645e-08, -2.018853e-08, 
    -1.985996e-08,
  -1.852242e-08, -1.882652e-08, -1.903217e-08, -1.922834e-08, -1.937195e-08, 
    -1.948369e-08, -1.958775e-08, -1.962051e-08, -1.968757e-08, -1.9598e-08, 
    -1.947403e-08, -1.931966e-08, -1.90365e-08, -1.860025e-08, -1.822991e-08,
  -1.828392e-08, -1.872632e-08, -1.903058e-08, -1.932714e-08, -1.944924e-08, 
    -1.948864e-08, -1.933147e-08, -1.916772e-08, -1.873992e-08, 
    -1.825292e-08, -1.764216e-08, -1.704561e-08, -1.648002e-08, 
    -1.605528e-08, -1.589401e-08,
  -1.795098e-08, -1.814959e-08, -1.837134e-08, -1.856278e-08, -1.861346e-08, 
    -1.851632e-08, -1.822501e-08, -1.781958e-08, -1.735124e-08, 
    -1.675171e-08, -1.622116e-08, -1.574192e-08, -1.531878e-08, 
    -1.524127e-08, -1.475176e-08,
  -1.743924e-08, -1.748293e-08, -1.740528e-08, -1.738469e-08, -1.726741e-08, 
    -1.708352e-08, -1.679131e-08, -1.653146e-08, -1.60948e-08, -1.58532e-08, 
    -1.539148e-08, -1.476772e-08, -1.449747e-08, -1.390128e-08, -1.336804e-08,
  -1.625022e-08, -1.643139e-08, -1.635429e-08, -1.618665e-08, -1.59891e-08, 
    -1.573449e-08, -1.548125e-08, -1.525331e-08, -1.498536e-08, 
    -1.464868e-08, -1.410418e-08, -1.37788e-08, -1.341881e-08, -1.275979e-08, 
    -1.229429e-08,
  -1.360455e-08, -1.427171e-08, -1.463961e-08, -1.476778e-08, -1.47103e-08, 
    -1.45432e-08, -1.429305e-08, -1.400151e-08, -1.370137e-08, -1.341005e-08, 
    -1.312565e-08, -1.295183e-08, -1.227647e-08, -1.163306e-08, -1.094409e-08,
  -1.074995e-08, -1.149398e-08, -1.207758e-08, -1.246086e-08, -1.26926e-08, 
    -1.27501e-08, -1.269941e-08, -1.249993e-08, -1.225952e-08, -1.20305e-08, 
    -1.185908e-08, -1.125523e-08, -1.058732e-08, -1.003801e-08, -9.521642e-09,
  -8.585823e-09, -9.163257e-09, -9.647357e-09, -1.004719e-08, -1.035766e-08, 
    -1.054863e-08, -1.062974e-08, -1.058257e-08, -1.044503e-08, 
    -1.023479e-08, -9.953422e-09, -9.590249e-09, -9.25578e-09, -8.905255e-09, 
    -8.522529e-09,
  -1.328049e-08, -1.321459e-08, -1.365813e-08, -1.462421e-08, -1.594426e-08, 
    -1.685435e-08, -1.748508e-08, -1.774501e-08, -1.790839e-08, 
    -1.804719e-08, -1.82356e-08, -1.837982e-08, -1.873622e-08, -1.92571e-08, 
    -1.937896e-08,
  -1.456066e-08, -1.357115e-08, -1.333825e-08, -1.334153e-08, -1.379055e-08, 
    -1.469188e-08, -1.570008e-08, -1.652144e-08, -1.698689e-08, 
    -1.728483e-08, -1.74317e-08, -1.759552e-08, -1.785689e-08, -1.806251e-08, 
    -1.838604e-08,
  -1.747765e-08, -1.59183e-08, -1.459213e-08, -1.378492e-08, -1.347009e-08, 
    -1.349423e-08, -1.385173e-08, -1.464191e-08, -1.552211e-08, 
    -1.632703e-08, -1.685178e-08, -1.720676e-08, -1.739694e-08, 
    -1.755068e-08, -1.765939e-08,
  -1.782498e-08, -1.807632e-08, -1.751689e-08, -1.628215e-08, -1.511937e-08, 
    -1.431924e-08, -1.401661e-08, -1.399214e-08, -1.426665e-08, -1.47192e-08, 
    -1.530139e-08, -1.581896e-08, -1.619008e-08, -1.641843e-08, -1.656821e-08,
  -1.606544e-08, -1.67891e-08, -1.748283e-08, -1.769014e-08, -1.745865e-08, 
    -1.666288e-08, -1.571387e-08, -1.502793e-08, -1.475772e-08, 
    -1.470213e-08, -1.476344e-08, -1.491108e-08, -1.51097e-08, -1.530518e-08, 
    -1.549381e-08,
  -1.486339e-08, -1.548854e-08, -1.608063e-08, -1.659257e-08, -1.704233e-08, 
    -1.725886e-08, -1.714958e-08, -1.670309e-08, -1.61124e-08, -1.566373e-08, 
    -1.546088e-08, -1.535058e-08, -1.533138e-08, -1.538527e-08, -1.55204e-08,
  -1.296323e-08, -1.413814e-08, -1.495987e-08, -1.560255e-08, -1.608141e-08, 
    -1.642547e-08, -1.669045e-08, -1.681944e-08, -1.679912e-08, 
    -1.658489e-08, -1.627835e-08, -1.602018e-08, -1.593368e-08, 
    -1.592725e-08, -1.603569e-08,
  -9.734002e-09, -1.138931e-08, -1.297962e-08, -1.415643e-08, -1.503198e-08, 
    -1.564572e-08, -1.608318e-08, -1.630859e-08, -1.645533e-08, 
    -1.649902e-08, -1.648629e-08, -1.640604e-08, -1.630183e-08, -1.62235e-08, 
    -1.620605e-08,
  -6.984354e-09, -8.368191e-09, -9.827309e-09, -1.130204e-08, -1.290497e-08, 
    -1.425744e-08, -1.529023e-08, -1.59839e-08, -1.637967e-08, -1.656464e-08, 
    -1.665951e-08, -1.674343e-08, -1.68035e-08, -1.68346e-08, -1.678275e-08,
  -5.131445e-09, -5.879488e-09, -7.002274e-09, -8.28738e-09, -9.585142e-09, 
    -1.093557e-08, -1.236361e-08, -1.375269e-08, -1.498586e-08, 
    -1.590045e-08, -1.650508e-08, -1.687291e-08, -1.705787e-08, 
    -1.711843e-08, -1.707426e-08,
  -1.263416e-08, -1.433889e-08, -1.547193e-08, -1.696909e-08, -1.718242e-08, 
    -1.746667e-08, -1.755984e-08, -1.83261e-08, -2.0108e-08, -2.269983e-08, 
    -2.411753e-08, -2.46442e-08, -2.48687e-08, -2.56387e-08, -2.659308e-08,
  -1.191186e-08, -1.244743e-08, -1.349743e-08, -1.504571e-08, -1.658642e-08, 
    -1.732792e-08, -1.758661e-08, -1.80153e-08, -1.859069e-08, -2.042516e-08, 
    -2.291155e-08, -2.421003e-08, -2.487885e-08, -2.545691e-08, -2.622533e-08,
  -1.208302e-08, -1.199559e-08, -1.239114e-08, -1.316796e-08, -1.457346e-08, 
    -1.62861e-08, -1.757101e-08, -1.76692e-08, -1.825002e-08, -1.902899e-08, 
    -2.063614e-08, -2.290002e-08, -2.426482e-08, -2.517774e-08, -2.564395e-08,
  -1.196384e-08, -1.207385e-08, -1.196333e-08, -1.216399e-08, -1.288707e-08, 
    -1.391869e-08, -1.574424e-08, -1.741143e-08, -1.809613e-08, 
    -1.851944e-08, -1.930798e-08, -2.078935e-08, -2.254726e-08, 
    -2.435456e-08, -2.569932e-08,
  -1.071855e-08, -1.166005e-08, -1.23225e-08, -1.235691e-08, -1.23335e-08, 
    -1.269032e-08, -1.349362e-08, -1.499118e-08, -1.663012e-08, 
    -1.814962e-08, -1.88092e-08, -1.958557e-08, -2.068986e-08, -2.203581e-08, 
    -2.388672e-08,
  -8.678097e-09, -9.740644e-09, -1.077457e-08, -1.185916e-08, -1.24883e-08, 
    -1.275062e-08, -1.29038e-08, -1.346492e-08, -1.443746e-08, -1.57437e-08, 
    -1.727436e-08, -1.844499e-08, -1.936606e-08, -2.032536e-08, -2.1265e-08,
  -7.003594e-09, -7.700187e-09, -8.619875e-09, -9.689635e-09, -1.075024e-08, 
    -1.171791e-08, -1.253781e-08, -1.311127e-08, -1.366577e-08, 
    -1.432586e-08, -1.527192e-08, -1.625751e-08, -1.738166e-08, 
    -1.838448e-08, -1.910994e-08,
  -6.60127e-09, -6.678739e-09, -6.939045e-09, -7.573082e-09, -8.496312e-09, 
    -9.520379e-09, -1.057806e-08, -1.164861e-08, -1.26251e-08, -1.360335e-08, 
    -1.448842e-08, -1.529705e-08, -1.60072e-08, -1.671808e-08, -1.741252e-08,
  -6.26216e-09, -6.381635e-09, -6.452069e-09, -6.611868e-09, -6.885303e-09, 
    -7.485273e-09, -8.301418e-09, -9.350205e-09, -1.041251e-08, 
    -1.141937e-08, -1.253165e-08, -1.378939e-08, -1.490829e-08, 
    -1.598327e-08, -1.684426e-08,
  -5.512329e-09, -5.845639e-09, -6.046594e-09, -6.200983e-09, -6.382799e-09, 
    -6.57248e-09, -6.896931e-09, -7.370593e-09, -8.077165e-09, -8.987555e-09, 
    -9.899926e-09, -1.089723e-08, -1.195499e-08, -1.308393e-08, -1.424593e-08,
  -1.862401e-08, -1.832408e-08, -1.800059e-08, -1.764595e-08, -1.737617e-08, 
    -1.718366e-08, -1.725878e-08, -1.736944e-08, -1.755722e-08, 
    -1.771346e-08, -1.783011e-08, -1.781862e-08, -1.762204e-08, 
    -1.714449e-08, -1.663333e-08,
  -1.816043e-08, -1.83347e-08, -1.833022e-08, -1.805398e-08, -1.774963e-08, 
    -1.749566e-08, -1.73186e-08, -1.730264e-08, -1.744403e-08, -1.757832e-08, 
    -1.764636e-08, -1.776694e-08, -1.777698e-08, -1.767973e-08, -1.74553e-08,
  -1.684868e-08, -1.739301e-08, -1.773708e-08, -1.78954e-08, -1.773763e-08, 
    -1.751976e-08, -1.731541e-08, -1.71355e-08, -1.710522e-08, -1.724849e-08, 
    -1.736819e-08, -1.748362e-08, -1.75564e-08, -1.767389e-08, -1.771253e-08,
  -1.532718e-08, -1.61506e-08, -1.665561e-08, -1.698057e-08, -1.717948e-08, 
    -1.712391e-08, -1.702343e-08, -1.684413e-08, -1.668389e-08, 
    -1.664932e-08, -1.67679e-08, -1.695339e-08, -1.713818e-08, -1.730184e-08, 
    -1.752523e-08,
  -1.319688e-08, -1.435601e-08, -1.522869e-08, -1.580721e-08, -1.619561e-08, 
    -1.636905e-08, -1.640294e-08, -1.638775e-08, -1.622965e-08, 
    -1.614532e-08, -1.610641e-08, -1.628125e-08, -1.658929e-08, 
    -1.686485e-08, -1.713434e-08,
  -1.070519e-08, -1.182101e-08, -1.297528e-08, -1.391421e-08, -1.459915e-08, 
    -1.520412e-08, -1.544694e-08, -1.560547e-08, -1.562112e-08, 
    -1.556108e-08, -1.549497e-08, -1.547032e-08, -1.565432e-08, 
    -1.605639e-08, -1.655494e-08,
  -7.659534e-09, -9.045653e-09, -1.027446e-08, -1.147115e-08, -1.247962e-08, 
    -1.333343e-08, -1.404654e-08, -1.446294e-08, -1.480619e-08, -1.49467e-08, 
    -1.504637e-08, -1.502135e-08, -1.500997e-08, -1.510181e-08, -1.546121e-08,
  -5.105715e-09, -6.105446e-09, -7.383523e-09, -8.567655e-09, -9.759187e-09, 
    -1.087187e-08, -1.184042e-08, -1.267349e-08, -1.32981e-08, -1.38488e-08, 
    -1.417957e-08, -1.445685e-08, -1.454761e-08, -1.459072e-08, -1.467462e-08,
  -3.6274e-09, -4.222466e-09, -5.034688e-09, -6.12458e-09, -7.192248e-09, 
    -8.291003e-09, -9.334782e-09, -1.031588e-08, -1.113662e-08, 
    -1.192635e-08, -1.261188e-08, -1.320629e-08, -1.366987e-08, -1.39561e-08, 
    -1.406005e-08,
  -2.417053e-09, -2.951036e-09, -3.428296e-09, -4.115344e-09, -5.018733e-09, 
    -6.05119e-09, -7.094106e-09, -8.119514e-09, -9.013692e-09, -9.810136e-09, 
    -1.061208e-08, -1.13323e-08, -1.208053e-08, -1.266489e-08, -1.319664e-08,
  -8.081035e-09, -8.724038e-09, -9.368351e-09, -1.000892e-08, -1.059238e-08, 
    -1.10785e-08, -1.144584e-08, -1.172975e-08, -1.200635e-08, -1.246183e-08, 
    -1.303938e-08, -1.366238e-08, -1.426142e-08, -1.483272e-08, -1.53042e-08,
  -7.497447e-09, -8.122561e-09, -8.762398e-09, -9.402139e-09, -1.001062e-08, 
    -1.055181e-08, -1.104004e-08, -1.143946e-08, -1.176636e-08, 
    -1.220384e-08, -1.275902e-08, -1.336777e-08, -1.405356e-08, 
    -1.470439e-08, -1.529621e-08,
  -6.874112e-09, -7.475634e-09, -8.081432e-09, -8.746672e-09, -9.409427e-09, 
    -1.00538e-08, -1.064245e-08, -1.116315e-08, -1.158322e-08, -1.19616e-08, 
    -1.247929e-08, -1.303886e-08, -1.367249e-08, -1.427801e-08, -1.486532e-08,
  -6.175942e-09, -6.793685e-09, -7.352769e-09, -7.963392e-09, -8.620176e-09, 
    -9.301672e-09, -9.981673e-09, -1.059425e-08, -1.118726e-08, 
    -1.169602e-08, -1.222033e-08, -1.278141e-08, -1.336373e-08, 
    -1.393431e-08, -1.450139e-08,
  -5.302456e-09, -5.995347e-09, -6.695501e-09, -7.371868e-09, -8.016052e-09, 
    -8.628135e-09, -9.321495e-09, -9.970662e-09, -1.058814e-08, 
    -1.119475e-08, -1.180938e-08, -1.242604e-08, -1.306803e-08, 
    -1.367239e-08, -1.427767e-08,
  -4.233111e-09, -4.973048e-09, -5.675233e-09, -6.410515e-09, -7.146852e-09, 
    -7.859793e-09, -8.579768e-09, -9.300106e-09, -9.99554e-09, -1.063205e-08, 
    -1.12572e-08, -1.190702e-08, -1.256566e-08, -1.323423e-08, -1.386316e-08,
  -3.217123e-09, -3.901346e-09, -4.62764e-09, -5.38314e-09, -6.159958e-09, 
    -6.88659e-09, -7.662424e-09, -8.437576e-09, -9.237627e-09, -1.000887e-08, 
    -1.070956e-08, -1.138334e-08, -1.206229e-08, -1.271038e-08, -1.334795e-08,
  -2.44178e-09, -2.939937e-09, -3.566602e-09, -4.258028e-09, -5.050204e-09, 
    -5.862208e-09, -6.634263e-09, -7.430321e-09, -8.242025e-09, 
    -9.098803e-09, -9.958639e-09, -1.07193e-08, -1.147897e-08, -1.216915e-08, 
    -1.283719e-08,
  -1.679481e-09, -2.155331e-09, -2.643759e-09, -3.261313e-09, -3.939196e-09, 
    -4.719685e-09, -5.533526e-09, -6.35469e-09, -7.198881e-09, -8.06475e-09, 
    -8.920657e-09, -9.838764e-09, -1.070058e-08, -1.15094e-08, -1.226028e-08,
  -1.162989e-09, -1.485116e-09, -1.86302e-09, -2.32297e-09, -2.917938e-09, 
    -3.609003e-09, -4.410871e-09, -5.249254e-09, -6.061129e-09, 
    -6.961287e-09, -7.870069e-09, -8.746339e-09, -9.742172e-09, 
    -1.069584e-08, -1.153054e-08,
  -3.021443e-09, -3.351009e-09, -4.053324e-09, -5.188523e-09, -6.740756e-09, 
    -8.609523e-09, -1.041351e-08, -1.198392e-08, -1.328315e-08, 
    -1.438371e-08, -1.529106e-08, -1.605882e-08, -1.660328e-08, 
    -1.700403e-08, -1.733179e-08,
  -2.054856e-09, -2.285488e-09, -2.581716e-09, -3.000808e-09, -3.54341e-09, 
    -4.361721e-09, -5.567966e-09, -7.003258e-09, -8.616118e-09, 
    -1.015553e-08, -1.149983e-08, -1.251568e-08, -1.334419e-08, 
    -1.400477e-08, -1.456514e-08,
  -1.141373e-09, -1.288827e-09, -1.493522e-09, -1.792141e-09, -2.189503e-09, 
    -2.656569e-09, -3.207063e-09, -3.841908e-09, -4.699516e-09, 
    -5.787457e-09, -7.060258e-09, -8.419128e-09, -9.731084e-09, 
    -1.083083e-08, -1.163718e-08,
  -6.333064e-10, -6.620441e-10, -7.527853e-10, -8.899583e-10, -1.098128e-09, 
    -1.401485e-09, -1.761248e-09, -2.149951e-09, -2.563837e-09, 
    -3.062495e-09, -3.731303e-09, -4.627939e-09, -5.743393e-09, 
    -6.986592e-09, -8.110447e-09,
  -2.402489e-10, -2.606488e-10, -3.405063e-10, -3.854086e-10, -4.471767e-10, 
    -5.516814e-10, -7.11428e-10, -9.632632e-10, -1.303866e-09, -1.707658e-09, 
    -2.181223e-09, -2.70648e-09, -3.375168e-09, -4.278351e-09, -5.375016e-09,
  7.966485e-11, 9.328346e-11, 3.250418e-11, -4.242207e-11, -7.650634e-11, 
    -9.390821e-11, -1.52114e-10, -3.01384e-10, -5.493998e-10, -9.189369e-10, 
    -1.357649e-09, -1.829386e-09, -2.353399e-09, -2.972494e-09, -3.768361e-09,
  1.276624e-10, 1.298483e-10, 9.003569e-11, 3.708701e-11, -8.984292e-12, 
    -3.872432e-11, -5.509154e-11, -1.181306e-10, -2.503329e-10, 
    -4.961167e-10, -8.468499e-10, -1.245725e-09, -1.653724e-09, 
    -2.093772e-09, -2.615142e-09,
  -9.956625e-11, -1.27389e-10, -1.090312e-10, -9.662768e-11, -1.078473e-10, 
    -1.430195e-10, -1.456418e-10, -1.451647e-10, -1.827637e-10, 
    -2.620189e-10, -4.398328e-10, -7.117004e-10, -1.040003e-09, 
    -1.407155e-09, -1.814369e-09,
  -3.332087e-10, -3.753934e-10, -3.589118e-10, -2.96727e-10, -2.261105e-10, 
    -1.936981e-10, -1.814016e-10, -1.732746e-10, -1.6526e-10, -1.79384e-10, 
    -2.212018e-10, -3.504802e-10, -5.462473e-10, -8.267301e-10, -1.164886e-09,
  -4.219391e-10, -4.535068e-10, -4.986783e-10, -5.064674e-10, -4.627955e-10, 
    -3.821517e-10, -3.021204e-10, -2.489499e-10, -2.326257e-10, 
    -2.234282e-10, -2.272937e-10, -2.772776e-10, -3.770577e-10, -5.61154e-10, 
    -8.589245e-10,
  -1.052185e-08, -1.168546e-08, -1.315016e-08, -1.481225e-08, -1.642015e-08, 
    -1.807732e-08, -1.935221e-08, -2.003823e-08, -2.039293e-08, -1.93978e-08, 
    -1.820816e-08, -1.786529e-08, -1.796227e-08, -1.832932e-08, -1.897468e-08,
  -7.765284e-09, -8.915714e-09, -1.015318e-08, -1.14001e-08, -1.283841e-08, 
    -1.428017e-08, -1.602672e-08, -1.753079e-08, -1.869352e-08, 
    -1.940691e-08, -1.943054e-08, -1.861074e-08, -1.805923e-08, 
    -1.804954e-08, -1.822206e-08,
  -5.540328e-09, -6.368476e-09, -7.408508e-09, -8.540305e-09, -9.780842e-09, 
    -1.09916e-08, -1.240564e-08, -1.385173e-08, -1.546209e-08, -1.679354e-08, 
    -1.791942e-08, -1.851606e-08, -1.842557e-08, -1.794823e-08, -1.785338e-08,
  -4.074005e-09, -4.68446e-09, -5.236431e-09, -5.890708e-09, -6.90441e-09, 
    -8.093082e-09, -9.339445e-09, -1.062393e-08, -1.205989e-08, 
    -1.345245e-08, -1.492023e-08, -1.601189e-08, -1.690445e-08, 
    -1.735287e-08, -1.723257e-08,
  -2.293352e-09, -2.931245e-09, -3.681198e-09, -4.3842e-09, -5.040544e-09, 
    -5.719961e-09, -6.619633e-09, -7.75204e-09, -8.924671e-09, -1.012385e-08, 
    -1.133376e-08, -1.258031e-08, -1.371317e-08, -1.463798e-08, -1.539753e-08,
  -1.154975e-09, -1.461901e-09, -1.943709e-09, -2.625513e-09, -3.40375e-09, 
    -4.131103e-09, -4.785262e-09, -5.439808e-09, -6.267567e-09, 
    -7.224367e-09, -8.30363e-09, -9.439376e-09, -1.051349e-08, -1.158528e-08, 
    -1.251191e-08,
  -4.916675e-10, -6.963761e-10, -9.818077e-10, -1.334222e-09, -1.724051e-09, 
    -2.311201e-09, -3.008927e-09, -3.67558e-09, -4.230715e-09, -4.820773e-09, 
    -5.528269e-09, -6.441502e-09, -7.515463e-09, -8.687218e-09, -9.787823e-09,
  -1.004913e-10, -1.811928e-10, -3.38592e-10, -5.351399e-10, -7.321495e-10, 
    -9.686877e-10, -1.25182e-09, -1.740959e-09, -2.385156e-09, -3.119283e-09, 
    -3.789071e-09, -4.449593e-09, -5.142018e-09, -5.949901e-09, -6.868119e-09,
  2.069243e-10, 2.112175e-10, 1.852527e-10, 1.399096e-10, 4.779458e-11, 
    -8.544451e-11, -2.83618e-10, -6.057631e-10, -1.084998e-09, -1.680544e-09, 
    -2.366925e-09, -3.053529e-09, -3.681189e-09, -4.272709e-09, -4.884636e-09,
  5.491117e-10, 5.142793e-10, 4.562402e-10, 4.507845e-10, 3.481928e-10, 
    1.646316e-10, -4.511494e-11, -2.606822e-10, -5.214251e-10, -8.50245e-10, 
    -1.2765e-09, -1.816387e-09, -2.48576e-09, -3.145072e-09, -3.714079e-09,
  -1.220909e-08, -1.286287e-08, -1.359213e-08, -1.428496e-08, -1.49492e-08, 
    -1.554158e-08, -1.598604e-08, -1.66102e-08, -1.717914e-08, -1.790284e-08, 
    -1.646099e-08, -1.61248e-08, -1.723287e-08, -1.844156e-08, -1.927551e-08,
  -1.06895e-08, -1.137686e-08, -1.209157e-08, -1.299016e-08, -1.376773e-08, 
    -1.453027e-08, -1.514068e-08, -1.579002e-08, -1.63999e-08, -1.713175e-08, 
    -1.796744e-08, -1.713758e-08, -1.658036e-08, -1.724646e-08, -1.812765e-08,
  -9.162505e-09, -9.66409e-09, -1.033737e-08, -1.106056e-08, -1.181702e-08, 
    -1.252325e-08, -1.323958e-08, -1.386311e-08, -1.460404e-08, 
    -1.530386e-08, -1.631667e-08, -1.719661e-08, -1.694989e-08, 
    -1.637833e-08, -1.698583e-08,
  -7.258627e-09, -7.627388e-09, -8.152891e-09, -8.733922e-09, -9.406783e-09, 
    -1.021e-08, -1.098064e-08, -1.171812e-08, -1.23937e-08, -1.308812e-08, 
    -1.405598e-08, -1.523969e-08, -1.643022e-08, -1.664236e-08, -1.611165e-08,
  -5.777507e-09, -6.102846e-09, -6.473261e-09, -6.799112e-09, -7.241463e-09, 
    -7.905714e-09, -8.72362e-09, -9.48158e-09, -1.027058e-08, -1.104883e-08, 
    -1.183327e-08, -1.303666e-08, -1.438458e-08, -1.58591e-08, -1.657816e-08,
  -4.497008e-09, -4.915532e-09, -5.228533e-09, -5.393787e-09, -5.699944e-09, 
    -6.217938e-09, -6.897686e-09, -7.627844e-09, -8.245626e-09, 
    -8.979881e-09, -9.752507e-09, -1.070016e-08, -1.199815e-08, 
    -1.343063e-08, -1.511674e-08,
  -3.429608e-09, -3.866409e-09, -4.19283e-09, -4.404543e-09, -4.425385e-09, 
    -4.652317e-09, -5.067445e-09, -5.756017e-09, -6.508458e-09, 
    -7.220784e-09, -7.914116e-09, -8.682466e-09, -9.751186e-09, 
    -1.099127e-08, -1.278417e-08,
  -2.475265e-09, -2.784381e-09, -3.053187e-09, -3.242119e-09, -3.520055e-09, 
    -3.700034e-09, -3.633458e-09, -3.669965e-09, -4.275326e-09, 
    -5.299044e-09, -6.318749e-09, -7.176395e-09, -8.112996e-09, 
    -9.068279e-09, -1.034456e-08,
  -1.744746e-09, -1.944833e-09, -2.157317e-09, -2.292271e-09, -2.299252e-09, 
    -2.328024e-09, -2.465497e-09, -2.599022e-09, -2.753151e-09, 
    -3.196161e-09, -4.257747e-09, -5.465934e-09, -6.539904e-09, 
    -7.595057e-09, -8.641954e-09,
  -1.230932e-09, -1.503511e-09, -1.970399e-09, -2.341357e-09, -2.455297e-09, 
    -2.220153e-09, -2.003239e-09, -1.9742e-09, -2.108029e-09, -2.289492e-09, 
    -2.643583e-09, -3.584324e-09, -4.74067e-09, -5.911673e-09, -6.959997e-09,
  -9.415461e-09, -9.666835e-09, -9.953875e-09, -1.028261e-08, -1.058652e-08, 
    -1.084696e-08, -1.106042e-08, -1.123726e-08, -1.139393e-08, -1.15159e-08, 
    -1.162044e-08, -1.17113e-08, -1.182098e-08, -1.192149e-08, -1.195413e-08,
  -8.750043e-09, -9.113818e-09, -9.460085e-09, -9.776619e-09, -1.010727e-08, 
    -1.039755e-08, -1.069114e-08, -1.098566e-08, -1.128457e-08, 
    -1.151386e-08, -1.172567e-08, -1.186955e-08, -1.201068e-08, 
    -1.219099e-08, -1.231986e-08,
  -7.826715e-09, -8.261173e-09, -8.697728e-09, -9.116751e-09, -9.505754e-09, 
    -9.892484e-09, -1.025421e-08, -1.059176e-08, -1.097848e-08, 
    -1.135177e-08, -1.171707e-08, -1.203899e-08, -1.218403e-08, 
    -1.238309e-08, -1.254168e-08,
  -6.815318e-09, -7.350171e-09, -7.831971e-09, -8.317572e-09, -8.779973e-09, 
    -9.236989e-09, -9.71824e-09, -1.018063e-08, -1.06167e-08, -1.106218e-08, 
    -1.141872e-08, -1.185253e-08, -1.215286e-08, -1.230862e-08, -1.249991e-08,
  -5.581756e-09, -6.235284e-09, -6.875604e-09, -7.472638e-09, -8.015879e-09, 
    -8.541696e-09, -9.079461e-09, -9.654323e-09, -1.01806e-08, -1.068309e-08, 
    -1.108867e-08, -1.142367e-08, -1.183982e-08, -1.211534e-08, -1.229303e-08,
  -4.384716e-09, -5.040275e-09, -5.715071e-09, -6.43114e-09, -7.091827e-09, 
    -7.671391e-09, -8.241514e-09, -8.887814e-09, -9.556397e-09, 
    -1.011085e-08, -1.059993e-08, -1.097151e-08, -1.131223e-08, 
    -1.164681e-08, -1.189758e-08,
  -3.349607e-09, -3.968623e-09, -4.614561e-09, -5.293439e-09, -5.98304e-09, 
    -6.653758e-09, -7.301776e-09, -7.978864e-09, -8.678889e-09, 
    -9.333628e-09, -9.800419e-09, -1.03394e-08, -1.06999e-08, -1.105301e-08, 
    -1.131381e-08,
  -2.559208e-09, -3.1237e-09, -3.704207e-09, -4.308353e-09, -4.91263e-09, 
    -5.5449e-09, -6.227988e-09, -6.94164e-09, -7.646745e-09, -8.30714e-09, 
    -8.955976e-09, -9.379515e-09, -9.95999e-09, -1.036154e-08, -1.073136e-08,
  -1.804307e-09, -2.376237e-09, -2.958337e-09, -3.568393e-09, -4.169146e-09, 
    -4.743814e-09, -5.361748e-09, -5.99463e-09, -6.658884e-09, -7.312579e-09, 
    -7.917938e-09, -8.534646e-09, -8.995691e-09, -9.661099e-09, -1.009791e-08,
  -1.233505e-09, -1.692751e-09, -2.221053e-09, -2.760091e-09, -3.41247e-09, 
    -4.025718e-09, -4.642305e-09, -5.208223e-09, -5.786671e-09, 
    -6.443681e-09, -7.028793e-09, -7.626221e-09, -8.180362e-09, 
    -8.662666e-09, -9.234229e-09,
  -7.92163e-09, -8.121246e-09, -8.402666e-09, -8.695751e-09, -8.976316e-09, 
    -9.224466e-09, -9.440217e-09, -9.65538e-09, -9.800051e-09, -9.948416e-09, 
    -1.005201e-08, -1.008638e-08, -1.000929e-08, -9.893729e-09, -9.88816e-09,
  -7.580555e-09, -7.693904e-09, -7.864185e-09, -8.102132e-09, -8.31292e-09, 
    -8.540234e-09, -8.716078e-09, -8.904127e-09, -8.983707e-09, 
    -9.102731e-09, -9.192486e-09, -9.19155e-09, -9.10824e-09, -9.024914e-09, 
    -9.055222e-09,
  -7.717508e-09, -7.995366e-09, -8.063759e-09, -8.165595e-09, -8.247312e-09, 
    -8.351096e-09, -8.472395e-09, -8.575378e-09, -8.735807e-09, 
    -8.948183e-09, -9.160343e-09, -8.990292e-09, -8.728759e-09, 
    -8.715857e-09, -8.761702e-09,
  -6.705196e-09, -7.295036e-09, -7.771319e-09, -8.155081e-09, -8.474336e-09, 
    -8.621984e-09, -8.769943e-09, -8.808371e-09, -8.94136e-09, -9.140637e-09, 
    -9.324776e-09, -9.180697e-09, -8.723999e-09, -8.819036e-09, -9.238477e-09,
  -5.057389e-09, -5.724815e-09, -6.414034e-09, -6.998797e-09, -7.551241e-09, 
    -7.980801e-09, -8.342218e-09, -8.662104e-09, -8.825033e-09, 
    -9.005279e-09, -9.281076e-09, -9.694449e-09, -9.721392e-09, 
    -9.434078e-09, -9.493633e-09,
  -3.318572e-09, -3.971624e-09, -4.666247e-09, -5.348329e-09, -6.004762e-09, 
    -6.612139e-09, -7.109279e-09, -7.634014e-09, -8.061368e-09, 
    -8.417754e-09, -8.745154e-09, -9.087182e-09, -9.419621e-09, -9.59934e-09, 
    -9.678088e-09,
  -1.522153e-09, -2.064317e-09, -2.679756e-09, -3.34809e-09, -4.026425e-09, 
    -4.704006e-09, -5.36173e-09, -6.017794e-09, -6.646263e-09, -7.185411e-09, 
    -7.681281e-09, -8.156334e-09, -8.589617e-09, -9.0755e-09, -9.458828e-09,
  -4.696955e-10, -7.044038e-10, -1.067034e-09, -1.52706e-09, -2.093549e-09, 
    -2.732411e-09, -3.467117e-09, -4.222488e-09, -4.997362e-09, 
    -5.728098e-09, -6.412683e-09, -7.006268e-09, -7.52384e-09, -7.975767e-09, 
    -8.486169e-09,
  2.642573e-11, -1.222397e-10, -3.320213e-10, -6.378859e-10, -9.660654e-10, 
    -1.409962e-09, -1.969197e-09, -2.63564e-09, -3.394307e-09, -4.25181e-09, 
    -5.121476e-09, -5.930124e-09, -6.558852e-09, -7.10523e-09, -7.580565e-09,
  2.586887e-10, 7.257443e-11, -8.732495e-11, -3.296922e-10, -5.824171e-10, 
    -8.86872e-10, -1.277353e-09, -1.770134e-09, -2.377349e-09, -3.066824e-09, 
    -3.812749e-09, -4.598359e-09, -5.323114e-09, -5.980079e-09, -6.555713e-09,
  -8.618636e-09, -8.718786e-09, -8.898179e-09, -9.119292e-09, -9.394959e-09, 
    -9.695256e-09, -1.002084e-08, -1.036881e-08, -1.075537e-08, 
    -1.115093e-08, -1.155422e-08, -1.198512e-08, -1.241717e-08, 
    -1.288058e-08, -1.334846e-08,
  -7.710164e-09, -7.813477e-09, -7.975933e-09, -8.187412e-09, -8.430835e-09, 
    -8.696791e-09, -8.969736e-09, -9.254046e-09, -9.537179e-09, 
    -9.806515e-09, -1.008233e-08, -1.036494e-08, -1.066276e-08, 
    -1.098893e-08, -1.130495e-08,
  -7.142137e-09, -7.223791e-09, -7.31729e-09, -7.422481e-09, -7.546669e-09, 
    -7.688852e-09, -7.850969e-09, -8.041249e-09, -8.252993e-09, 
    -8.476559e-09, -8.721714e-09, -8.969676e-09, -9.251751e-09, 
    -9.537891e-09, -9.802754e-09,
  -6.274054e-09, -6.284794e-09, -6.277298e-09, -6.240056e-09, -6.237789e-09, 
    -6.254721e-09, -6.301671e-09, -6.379554e-09, -6.500757e-09, 
    -6.674159e-09, -6.908341e-09, -7.192328e-09, -7.505083e-09, 
    -7.815986e-09, -8.106757e-09,
  -5.154004e-09, -5.077939e-09, -4.984847e-09, -4.921598e-09, -4.915117e-09, 
    -4.940768e-09, -4.983535e-09, -5.054268e-09, -5.159864e-09, 
    -5.291739e-09, -5.466701e-09, -5.671304e-09, -5.94282e-09, -6.294455e-09, 
    -6.709969e-09,
  -3.904927e-09, -3.812923e-09, -3.705056e-09, -3.660373e-09, -3.657342e-09, 
    -3.654551e-09, -3.665566e-09, -3.7127e-09, -3.814e-09, -3.95459e-09, 
    -4.132648e-09, -4.335812e-09, -4.567847e-09, -4.831569e-09, -5.091427e-09,
  -2.617057e-09, -2.524541e-09, -2.428561e-09, -2.376696e-09, -2.343153e-09, 
    -2.290539e-09, -2.235991e-09, -2.206413e-09, -2.229984e-09, 
    -2.327112e-09, -2.500279e-09, -2.658883e-09, -2.873854e-09, 
    -3.040887e-09, -3.212857e-09,
  -1.474093e-09, -1.37874e-09, -1.306119e-09, -1.270214e-09, -1.231957e-09, 
    -1.16627e-09, -1.07908e-09, -1.024995e-09, -1.020891e-09, -1.10323e-09, 
    -1.247113e-09, -1.425985e-09, -1.604078e-09, -1.783099e-09, -1.982803e-09,
  -7.731847e-10, -6.85814e-10, -6.142271e-10, -5.681742e-10, -4.927125e-10, 
    -3.867461e-10, -2.486527e-10, -2.005811e-10, -2.749812e-10, 
    -4.620451e-10, -6.903869e-10, -9.790304e-10, -1.344243e-09, 
    -1.705471e-09, -2.091994e-09,
  -3.266428e-10, -2.267816e-10, -1.734187e-10, -1.117594e-10, -2.8483e-11, 
    1.299011e-11, 5.273949e-11, 1.484676e-11, -1.518081e-10, -4.475035e-10, 
    -7.985388e-10, -1.16866e-09, -1.556188e-09, -1.945194e-09, -2.343318e-09,
  -2.014439e-08, -1.981871e-08, -1.956483e-08, -1.913757e-08, -1.849701e-08, 
    -1.757679e-08, -1.629058e-08, -1.467405e-08, -1.291455e-08, 
    -1.104198e-08, -9.318715e-09, -7.946393e-09, -7.135741e-09, 
    -6.884533e-09, -6.908005e-09,
  -1.686477e-08, -1.653581e-08, -1.614577e-08, -1.560378e-08, -1.49064e-08, 
    -1.391714e-08, -1.268299e-08, -1.128052e-08, -9.728466e-09, 
    -8.288081e-09, -7.235451e-09, -6.590195e-09, -6.421981e-09, 
    -6.565158e-09, -6.762149e-09,
  -1.419786e-08, -1.413324e-08, -1.380736e-08, -1.315672e-08, -1.233333e-08, 
    -1.132466e-08, -1.025032e-08, -9.012822e-09, -7.881961e-09, -7.10521e-09, 
    -6.671201e-09, -6.675866e-09, -6.982355e-09, -7.25765e-09, -7.486286e-09,
  -1.169538e-08, -1.17201e-08, -1.154052e-08, -1.106093e-08, -1.036537e-08, 
    -9.514582e-09, -8.477567e-09, -7.524304e-09, -6.913802e-09, 
    -6.685405e-09, -6.859078e-09, -7.168181e-09, -7.363519e-09, 
    -7.460283e-09, -7.50189e-09,
  -1.042716e-08, -1.025913e-08, -1.002285e-08, -9.638232e-09, -9.072411e-09, 
    -8.223943e-09, -7.460433e-09, -7.0346e-09, -6.959322e-09, -7.15417e-09, 
    -7.351024e-09, -7.363193e-09, -7.299076e-09, -7.118813e-09, -6.706551e-09,
  -9.373013e-09, -9.162926e-09, -8.89624e-09, -8.497294e-09, -7.899734e-09, 
    -7.353001e-09, -7.08595e-09, -7.01542e-09, -7.059497e-09, -6.93039e-09, 
    -6.70603e-09, -6.383343e-09, -5.946016e-09, -5.319135e-09, -4.832557e-09,
  -8.140983e-09, -7.967023e-09, -7.700614e-09, -7.333638e-09, -6.981035e-09, 
    -6.72899e-09, -6.572273e-09, -6.338403e-09, -6.071469e-09, -5.702783e-09, 
    -5.195991e-09, -4.563051e-09, -3.847894e-09, -3.383898e-09, -3.154233e-09,
  -6.654536e-09, -6.541429e-09, -6.344266e-09, -6.121284e-09, -5.886205e-09, 
    -5.586843e-09, -5.241479e-09, -4.829123e-09, -4.282675e-09, 
    -3.622941e-09, -2.883626e-09, -2.249977e-09, -1.926742e-09, 
    -1.790385e-09, -1.724288e-09,
  -5.116549e-09, -5.031798e-09, -4.854845e-09, -4.604025e-09, -4.27268e-09, 
    -3.851022e-09, -3.361829e-09, -2.763434e-09, -2.103185e-09, 
    -1.497669e-09, -1.129658e-09, -9.948454e-10, -9.896717e-10, 
    -1.009402e-09, -1.023216e-09,
  -3.635135e-09, -3.478349e-09, -3.235742e-09, -2.9222e-09, -2.546125e-09, 
    -2.153042e-09, -1.671109e-09, -1.188154e-09, -8.262862e-10, 
    -6.519207e-10, -6.175105e-10, -6.249568e-10, -6.412114e-10, 
    -6.510926e-10, -7.089575e-10,
  -7.803772e-09, -8.402537e-09, -9.231197e-09, -1.036363e-08, -1.156585e-08, 
    -1.276655e-08, -1.407666e-08, -1.537742e-08, -1.651516e-08, 
    -1.777135e-08, -1.898104e-08, -2.009668e-08, -2.1172e-08, -2.169111e-08, 
    -2.188838e-08,
  -7.933657e-09, -8.424599e-09, -9.08797e-09, -1.004367e-08, -1.119619e-08, 
    -1.244203e-08, -1.366696e-08, -1.479952e-08, -1.598212e-08, -1.70541e-08, 
    -1.805944e-08, -1.881708e-08, -1.947751e-08, -1.988131e-08, -2.007097e-08,
  -8.00203e-09, -8.424392e-09, -8.999193e-09, -9.76453e-09, -1.084864e-08, 
    -1.206511e-08, -1.325291e-08, -1.447408e-08, -1.557407e-08, 
    -1.645163e-08, -1.709313e-08, -1.75617e-08, -1.781244e-08, -1.814046e-08, 
    -1.828e-08,
  -7.895203e-09, -8.429034e-09, -9.030708e-09, -9.705353e-09, -1.065216e-08, 
    -1.176789e-08, -1.311763e-08, -1.439037e-08, -1.530453e-08, 
    -1.595735e-08, -1.630235e-08, -1.649235e-08, -1.651952e-08, 
    -1.669248e-08, -1.67551e-08,
  -7.796882e-09, -8.346602e-09, -8.920036e-09, -9.551063e-09, -1.043425e-08, 
    -1.170494e-08, -1.295265e-08, -1.396614e-08, -1.467967e-08, 
    -1.511546e-08, -1.530757e-08, -1.54077e-08, -1.548426e-08, -1.554106e-08, 
    -1.544375e-08,
  -7.718659e-09, -8.391589e-09, -8.859661e-09, -9.480447e-09, -1.043999e-08, 
    -1.151095e-08, -1.243737e-08, -1.315664e-08, -1.364704e-08, 
    -1.399143e-08, -1.417468e-08, -1.430022e-08, -1.436323e-08, 
    -1.432938e-08, -1.414872e-08,
  -7.511797e-09, -8.37854e-09, -9.061004e-09, -9.672975e-09, -1.026044e-08, 
    -1.085786e-08, -1.143195e-08, -1.188017e-08, -1.22311e-08, -1.256269e-08, 
    -1.285107e-08, -1.309338e-08, -1.306385e-08, -1.284194e-08, -1.252798e-08,
  -7.275026e-09, -8.04003e-09, -8.724665e-09, -9.317975e-09, -9.657604e-09, 
    -9.887302e-09, -1.016639e-08, -1.05494e-08, -1.095359e-08, -1.130815e-08, 
    -1.161731e-08, -1.161116e-08, -1.152354e-08, -1.134862e-08, -1.096931e-08,
  -6.412265e-09, -7.020247e-09, -7.511432e-09, -7.932726e-09, -8.248538e-09, 
    -8.519632e-09, -8.817248e-09, -9.080965e-09, -9.485565e-09, 
    -9.727097e-09, -9.891918e-09, -9.853252e-09, -9.681053e-09, 
    -9.417992e-09, -9.131085e-09,
  -5.391299e-09, -5.853596e-09, -6.282236e-09, -6.686158e-09, -7.017638e-09, 
    -7.258489e-09, -7.536413e-09, -7.709741e-09, -7.855367e-09, 
    -7.940412e-09, -7.961366e-09, -7.940778e-09, -7.852268e-09, 
    -7.588947e-09, -7.250335e-09,
  -5.534847e-09, -4.676381e-09, -4.095564e-09, -3.847555e-09, -3.730462e-09, 
    -3.826496e-09, -4.043089e-09, -4.154763e-09, -4.329921e-09, 
    -4.573992e-09, -4.65053e-09, -4.793009e-09, -5.119117e-09, -5.586107e-09, 
    -6.367415e-09,
  -6.096139e-09, -5.347499e-09, -4.441385e-09, -3.938287e-09, -3.781182e-09, 
    -3.765886e-09, -3.949176e-09, -4.153577e-09, -4.223954e-09, 
    -4.421244e-09, -4.60341e-09, -4.70711e-09, -4.942688e-09, -5.345223e-09, 
    -5.871228e-09,
  -6.447824e-09, -5.931683e-09, -5.100533e-09, -4.245283e-09, -3.85439e-09, 
    -3.748466e-09, -3.847494e-09, -4.039261e-09, -4.186405e-09, 
    -4.338371e-09, -4.465302e-09, -4.609537e-09, -4.748004e-09, 
    -5.104404e-09, -5.550812e-09,
  -6.722521e-09, -6.345921e-09, -5.670401e-09, -4.760171e-09, -4.090622e-09, 
    -3.824447e-09, -3.782607e-09, -3.99154e-09, -4.139668e-09, -4.238745e-09, 
    -4.378376e-09, -4.487188e-09, -4.608647e-09, -4.785977e-09, -5.229079e-09,
  -6.918652e-09, -6.763767e-09, -6.221263e-09, -5.401902e-09, -4.467328e-09, 
    -3.979311e-09, -3.810023e-09, -3.898764e-09, -4.136959e-09, 
    -4.256485e-09, -4.304738e-09, -4.382274e-09, -4.506009e-09, 
    -4.627334e-09, -4.88763e-09,
  -6.709191e-09, -6.749132e-09, -6.529841e-09, -5.931962e-09, -5.054073e-09, 
    -4.301104e-09, -3.916894e-09, -3.871995e-09, -4.027463e-09, 
    -4.266109e-09, -4.340933e-09, -4.32534e-09, -4.370134e-09, -4.525937e-09, 
    -4.745726e-09,
  -6.475947e-09, -6.679562e-09, -6.55948e-09, -6.317055e-09, -5.527942e-09, 
    -4.728467e-09, -4.114685e-09, -3.953529e-09, -3.98558e-09, -4.202003e-09, 
    -4.379078e-09, -4.441207e-09, -4.416793e-09, -4.49883e-09, -4.621993e-09,
  -6.049512e-09, -6.353406e-09, -6.513838e-09, -6.509025e-09, -6.035367e-09, 
    -5.213669e-09, -4.435079e-09, -4.082186e-09, -4.014884e-09, 
    -4.126949e-09, -4.345821e-09, -4.52697e-09, -4.615798e-09, -4.705321e-09, 
    -4.777474e-09,
  -5.706795e-09, -6.11419e-09, -6.304089e-09, -6.611074e-09, -6.351324e-09, 
    -5.563554e-09, -4.839976e-09, -4.374831e-09, -4.118729e-09, 
    -4.089988e-09, -4.245103e-09, -4.494678e-09, -4.680953e-09, 
    -4.774098e-09, -4.807383e-09,
  -5.181489e-09, -5.786122e-09, -6.13531e-09, -6.481915e-09, -6.650306e-09, 
    -6.136889e-09, -5.254126e-09, -4.616949e-09, -4.284271e-09, 
    -4.182238e-09, -4.326009e-09, -4.613327e-09, -4.866771e-09, 
    -5.019964e-09, -5.094697e-09,
  -4.875754e-09, -5.031632e-09, -5.107384e-09, -5.140041e-09, -5.043538e-09, 
    -4.916985e-09, -4.770105e-09, -4.67858e-09, -4.610988e-09, -4.626696e-09, 
    -4.696708e-09, -4.697652e-09, -4.668446e-09, -4.61826e-09, -4.620098e-09,
  -5.042618e-09, -5.169386e-09, -5.20465e-09, -5.196732e-09, -5.118887e-09, 
    -5.006555e-09, -4.779913e-09, -4.632717e-09, -4.534346e-09, 
    -4.562371e-09, -4.643711e-09, -4.669793e-09, -4.633177e-09, 
    -4.562827e-09, -4.59295e-09,
  -5.014563e-09, -5.32175e-09, -5.480437e-09, -5.407097e-09, -5.134163e-09, 
    -4.91853e-09, -4.715917e-09, -4.50271e-09, -4.397355e-09, -4.405109e-09, 
    -4.545001e-09, -4.580759e-09, -4.614012e-09, -4.547837e-09, -4.54409e-09,
  -5.177491e-09, -5.613831e-09, -5.791645e-09, -5.501796e-09, -5.046466e-09, 
    -4.553846e-09, -4.374172e-09, -4.347079e-09, -4.286897e-09, 
    -4.321885e-09, -4.522723e-09, -4.663889e-09, -4.678399e-09, 
    -4.683543e-09, -4.654996e-09,
  -5.64465e-09, -6.158521e-09, -5.979059e-09, -5.437031e-09, -4.853038e-09, 
    -4.269952e-09, -4.115634e-09, -4.263122e-09, -4.402851e-09, -4.36293e-09, 
    -4.522028e-09, -4.828256e-09, -4.853708e-09, -4.82301e-09, -4.805778e-09,
  -6.288165e-09, -6.326165e-09, -5.950494e-09, -5.400507e-09, -4.687345e-09, 
    -4.179575e-09, -4.007008e-09, -4.141008e-09, -4.448957e-09, 
    -4.555385e-09, -4.756855e-09, -4.994301e-09, -5.117418e-09, 
    -5.165576e-09, -5.04548e-09,
  -6.566743e-09, -6.334423e-09, -5.80275e-09, -5.21778e-09, -4.477182e-09, 
    -4.045361e-09, -3.950764e-09, -4.064449e-09, -4.41386e-09, -4.672498e-09, 
    -4.843432e-09, -4.990408e-09, -5.045622e-09, -5.241154e-09, -5.395119e-09,
  -6.828114e-09, -6.29022e-09, -5.720996e-09, -5.179418e-09, -4.576063e-09, 
    -4.058877e-09, -3.88076e-09, -3.897694e-09, -4.246294e-09, -4.613023e-09, 
    -4.786112e-09, -4.894701e-09, -4.904324e-09, -5.026179e-09, -5.061371e-09,
  -6.720486e-09, -6.331624e-09, -5.806544e-09, -5.208295e-09, -4.61938e-09, 
    -4.164124e-09, -3.925341e-09, -3.898726e-09, -4.121988e-09, 
    -4.473385e-09, -4.754449e-09, -4.875262e-09, -4.798799e-09, 
    -4.771864e-09, -4.782946e-09,
  -6.901729e-09, -6.585139e-09, -5.869401e-09, -5.270936e-09, -4.747183e-09, 
    -4.291827e-09, -3.944573e-09, -3.814773e-09, -3.845594e-09, 
    -4.142292e-09, -4.443554e-09, -4.61423e-09, -4.655901e-09, -4.640345e-09, 
    -4.632965e-09,
  -5.400428e-09, -5.202383e-09, -5.013896e-09, -4.853033e-09, -4.71243e-09, 
    -4.57089e-09, -4.454612e-09, -4.353596e-09, -4.299816e-09, -4.289831e-09, 
    -4.325966e-09, -4.404402e-09, -4.514333e-09, -4.663135e-09, -4.821999e-09,
  -4.67811e-09, -4.612509e-09, -4.552266e-09, -4.474866e-09, -4.392416e-09, 
    -4.328728e-09, -4.29417e-09, -4.285044e-09, -4.313831e-09, -4.381023e-09, 
    -4.491736e-09, -4.641169e-09, -4.819929e-09, -4.982544e-09, -5.122161e-09,
  -4.400894e-09, -4.411035e-09, -4.392247e-09, -4.361522e-09, -4.348894e-09, 
    -4.356277e-09, -4.379127e-09, -4.425683e-09, -4.488912e-09, 
    -4.588209e-09, -4.727241e-09, -4.903883e-09, -5.02459e-09, -5.10664e-09, 
    -5.109718e-09,
  -4.11674e-09, -4.150718e-09, -4.188584e-09, -4.23536e-09, -4.2998e-09, 
    -4.365461e-09, -4.420471e-09, -4.470593e-09, -4.535193e-09, 
    -4.696791e-09, -4.829833e-09, -4.888685e-09, -4.901161e-09, 
    -4.840517e-09, -4.789682e-09,
  -3.942464e-09, -4.006929e-09, -4.112858e-09, -4.245271e-09, -4.336842e-09, 
    -4.423744e-09, -4.468893e-09, -4.538516e-09, -4.674147e-09, 
    -4.818416e-09, -4.832275e-09, -4.844404e-09, -4.839687e-09, 
    -4.835601e-09, -4.825455e-09,
  -3.740247e-09, -3.920218e-09, -4.104146e-09, -4.280898e-09, -4.377459e-09, 
    -4.44895e-09, -4.510469e-09, -4.641383e-09, -4.803922e-09, -4.852308e-09, 
    -4.913293e-09, -4.997371e-09, -5.00055e-09, -5.046365e-09, -5.045105e-09,
  -3.631855e-09, -3.889124e-09, -4.131941e-09, -4.295654e-09, -4.424106e-09, 
    -4.457135e-09, -4.57072e-09, -4.699962e-09, -4.830255e-09, -5.014994e-09, 
    -5.224395e-09, -5.076144e-09, -5.000423e-09, -5.14332e-09, -5.706049e-09,
  -3.641498e-09, -3.955696e-09, -4.162641e-09, -4.372275e-09, -4.461401e-09, 
    -4.494829e-09, -4.497674e-09, -4.575752e-09, -4.891329e-09, 
    -5.274629e-09, -5.313854e-09, -4.877179e-09, -4.878121e-09, 
    -5.342403e-09, -5.950774e-09,
  -3.709443e-09, -4.020364e-09, -4.258346e-09, -4.429413e-09, -4.48929e-09, 
    -4.526854e-09, -4.401277e-09, -4.436892e-09, -4.950957e-09, 
    -5.578348e-09, -5.493991e-09, -5.023138e-09, -5.054432e-09, 
    -5.423808e-09, -5.910616e-09,
  -3.756694e-09, -4.149272e-09, -4.377218e-09, -4.543147e-09, -4.415306e-09, 
    -4.345635e-09, -4.209402e-09, -4.223697e-09, -4.751155e-09, 
    -5.861119e-09, -5.928972e-09, -5.636609e-09, -5.530687e-09, 
    -5.628791e-09, -5.617192e-09,
  -1.800671e-08, -1.77372e-08, -1.740722e-08, -1.71336e-08, -1.672078e-08, 
    -1.627197e-08, -1.560337e-08, -1.482969e-08, -1.395475e-08, 
    -1.307451e-08, -1.215994e-08, -1.121786e-08, -1.027868e-08, 
    -9.359953e-09, -8.515935e-09,
  -1.664773e-08, -1.648446e-08, -1.63243e-08, -1.608118e-08, -1.57326e-08, 
    -1.52009e-08, -1.450972e-08, -1.368498e-08, -1.2783e-08, -1.18333e-08, 
    -1.085181e-08, -9.846095e-09, -8.859469e-09, -7.96032e-09, -7.16653e-09,
  -1.489911e-08, -1.488803e-08, -1.483368e-08, -1.470903e-08, -1.43921e-08, 
    -1.38771e-08, -1.321013e-08, -1.242296e-08, -1.153071e-08, -1.054595e-08, 
    -9.56425e-09, -8.576011e-09, -7.664749e-09, -6.88818e-09, -6.235148e-09,
  -1.289026e-08, -1.318449e-08, -1.323102e-08, -1.319319e-08, -1.29735e-08, 
    -1.254452e-08, -1.199631e-08, -1.129119e-08, -1.044702e-08, 
    -9.501283e-09, -8.561727e-09, -7.640993e-09, -6.837616e-09, 
    -6.178054e-09, -5.616419e-09,
  -1.084804e-08, -1.139033e-08, -1.161586e-08, -1.168542e-08, -1.157077e-08, 
    -1.12473e-08, -1.08135e-08, -1.01951e-08, -9.404951e-09, -8.557004e-09, 
    -7.695513e-09, -6.889789e-09, -6.204858e-09, -5.626034e-09, -5.202627e-09,
  -8.795564e-09, -9.552381e-09, -9.983797e-09, -1.018945e-08, -1.019493e-08, 
    -1.007008e-08, -9.727676e-09, -9.204077e-09, -8.505441e-09, 
    -7.743066e-09, -6.960348e-09, -6.262679e-09, -5.652057e-09, 
    -5.212611e-09, -4.929062e-09,
  -7.221625e-09, -7.866589e-09, -8.366237e-09, -8.696259e-09, -8.855985e-09, 
    -8.831454e-09, -8.603755e-09, -8.139442e-09, -7.577992e-09, 
    -6.935312e-09, -6.292967e-09, -5.705427e-09, -5.258694e-09, 
    -4.968389e-09, -4.849414e-09,
  -6.262263e-09, -6.696027e-09, -7.113158e-09, -7.444616e-09, -7.658486e-09, 
    -7.706099e-09, -7.547972e-09, -7.216423e-09, -6.748721e-09, 
    -6.241066e-09, -5.735968e-09, -5.316036e-09, -5.012297e-09, 
    -4.878021e-09, -4.875303e-09,
  -5.343096e-09, -5.851555e-09, -6.258702e-09, -6.563344e-09, -6.764145e-09, 
    -6.775436e-09, -6.643943e-09, -6.389656e-09, -6.072788e-09, 
    -5.699126e-09, -5.333406e-09, -5.053979e-09, -4.868433e-09, 
    -4.822104e-09, -4.898278e-09,
  -4.772018e-09, -5.184348e-09, -5.553848e-09, -5.852693e-09, -6.09002e-09, 
    -6.093178e-09, -5.936248e-09, -5.78244e-09, -5.560099e-09, -5.341112e-09, 
    -5.10152e-09, -4.985584e-09, -4.971083e-09, -5.034199e-09, -5.196632e-09,
  -2.329845e-08, -2.357518e-08, -2.385149e-08, -2.41552e-08, -2.431524e-08, 
    -2.44652e-08, -2.420679e-08, -2.381604e-08, -2.324498e-08, -2.24518e-08, 
    -2.188972e-08, -2.130114e-08, -2.0875e-08, -2.053849e-08, -2.013234e-08,
  -2.168289e-08, -2.2506e-08, -2.306765e-08, -2.315932e-08, -2.346708e-08, 
    -2.347442e-08, -2.319516e-08, -2.307028e-08, -2.244767e-08, 
    -2.200835e-08, -2.154089e-08, -2.109526e-08, -2.072295e-08, 
    -2.024256e-08, -1.967152e-08,
  -1.905117e-08, -2.07039e-08, -2.177554e-08, -2.21557e-08, -2.241565e-08, 
    -2.260361e-08, -2.253964e-08, -2.255275e-08, -2.205485e-08, 
    -2.171158e-08, -2.109731e-08, -2.065859e-08, -2.010921e-08, 
    -1.951425e-08, -1.880952e-08,
  -1.608235e-08, -1.810185e-08, -1.970854e-08, -2.076472e-08, -2.140592e-08, 
    -2.175468e-08, -2.184914e-08, -2.189287e-08, -2.142115e-08, 
    -2.115583e-08, -2.043222e-08, -2.0017e-08, -1.94612e-08, -1.871821e-08, 
    -1.784886e-08,
  -1.315341e-08, -1.50451e-08, -1.67672e-08, -1.832606e-08, -1.934961e-08, 
    -2.019131e-08, -2.054235e-08, -2.074039e-08, -2.043526e-08, 
    -2.010863e-08, -1.955031e-08, -1.912167e-08, -1.846385e-08, 
    -1.764959e-08, -1.662752e-08,
  -1.043311e-08, -1.264784e-08, -1.430337e-08, -1.5886e-08, -1.714843e-08, 
    -1.820436e-08, -1.877188e-08, -1.920115e-08, -1.924738e-08, -1.89947e-08, 
    -1.865317e-08, -1.821176e-08, -1.752582e-08, -1.672252e-08, -1.566394e-08,
  -7.333117e-09, -9.628024e-09, -1.183696e-08, -1.351477e-08, -1.493968e-08, 
    -1.617152e-08, -1.696609e-08, -1.751147e-08, -1.776126e-08, 
    -1.771628e-08, -1.753133e-08, -1.711037e-08, -1.652091e-08, 
    -1.569578e-08, -1.46498e-08,
  -5.554102e-09, -7.085414e-09, -9.111713e-09, -1.118585e-08, -1.274299e-08, 
    -1.41355e-08, -1.517212e-08, -1.582135e-08, -1.629514e-08, -1.640908e-08, 
    -1.634847e-08, -1.601251e-08, -1.550483e-08, -1.46736e-08, -1.378112e-08,
  -4.166742e-09, -5.373273e-09, -6.906089e-09, -8.790659e-09, -1.065059e-08, 
    -1.208523e-08, -1.334105e-08, -1.415915e-08, -1.472837e-08, 
    -1.506463e-08, -1.507904e-08, -1.494714e-08, -1.441875e-08, 
    -1.373751e-08, -1.276906e-08,
  -3.123563e-09, -4.155317e-09, -5.374878e-09, -6.817524e-09, -8.523664e-09, 
    -1.018428e-08, -1.148838e-08, -1.253449e-08, -1.319151e-08, 
    -1.366003e-08, -1.378805e-08, -1.371859e-08, -1.332638e-08, 
    -1.266949e-08, -1.187845e-08,
  -1.954704e-08, -2.078692e-08, -2.222209e-08, -2.29246e-08, -2.371625e-08, 
    -2.456083e-08, -2.591447e-08, -2.581635e-08, -2.626611e-08, 
    -2.579893e-08, -2.550428e-08, -2.521116e-08, -2.455631e-08, 
    -2.370117e-08, -2.320476e-08,
  -1.818855e-08, -1.93909e-08, -2.059045e-08, -2.204693e-08, -2.287722e-08, 
    -2.34434e-08, -2.467965e-08, -2.573542e-08, -2.641608e-08, -2.604892e-08, 
    -2.587116e-08, -2.544798e-08, -2.500416e-08, -2.466435e-08, -2.364723e-08,
  -1.626874e-08, -1.808602e-08, -1.929e-08, -2.052425e-08, -2.200649e-08, 
    -2.280014e-08, -2.361534e-08, -2.447932e-08, -2.547983e-08, 
    -2.554155e-08, -2.531554e-08, -2.536953e-08, -2.484667e-08, 
    -2.422701e-08, -2.333488e-08,
  -1.34306e-08, -1.56475e-08, -1.779838e-08, -1.926749e-08, -2.078322e-08, 
    -2.20023e-08, -2.300053e-08, -2.381518e-08, -2.457634e-08, -2.510749e-08, 
    -2.501332e-08, -2.46367e-08, -2.451278e-08, -2.438539e-08, -2.377698e-08,
  -1.042091e-08, -1.278106e-08, -1.513503e-08, -1.735227e-08, -1.902762e-08, 
    -2.074838e-08, -2.193882e-08, -2.304045e-08, -2.398015e-08, 
    -2.454466e-08, -2.475494e-08, -2.444381e-08, -2.439058e-08, 
    -2.393109e-08, -2.340685e-08,
  -7.69746e-09, -9.934776e-09, -1.231762e-08, -1.477076e-08, -1.693504e-08, 
    -1.880186e-08, -2.046796e-08, -2.177282e-08, -2.280628e-08, 
    -2.390144e-08, -2.436571e-08, -2.412506e-08, -2.404637e-08, 
    -2.385925e-08, -2.332978e-08,
  -5.210207e-09, -7.061117e-09, -9.31334e-09, -1.195954e-08, -1.435297e-08, 
    -1.657072e-08, -1.841152e-08, -2.005142e-08, -2.137995e-08, 
    -2.242139e-08, -2.342013e-08, -2.358954e-08, -2.33841e-08, -2.332406e-08, 
    -2.281882e-08,
  -3.616563e-09, -4.951017e-09, -6.617736e-09, -8.870227e-09, -1.155924e-08, 
    -1.382251e-08, -1.606621e-08, -1.781415e-08, -1.943421e-08, 
    -2.099477e-08, -2.186041e-08, -2.258277e-08, -2.249486e-08, 
    -2.240444e-08, -2.210286e-08,
  -2.54743e-09, -3.447782e-09, -4.715101e-09, -6.290669e-09, -8.626379e-09, 
    -1.105459e-08, -1.325335e-08, -1.54201e-08, -1.692555e-08, -1.862469e-08, 
    -2.010318e-08, -2.109082e-08, -2.156462e-08, -2.139994e-08, -2.122388e-08,
  -1.811269e-09, -2.360116e-09, -3.289095e-09, -4.455033e-09, -6.052938e-09, 
    -8.407408e-09, -1.054869e-08, -1.274953e-08, -1.467012e-08, 
    -1.613629e-08, -1.766354e-08, -1.902483e-08, -2.01744e-08, -2.049353e-08, 
    -2.033685e-08,
  -1.343928e-08, -1.431559e-08, -1.495796e-08, -1.543095e-08, -1.635604e-08, 
    -1.762996e-08, -1.961878e-08, -2.164795e-08, -2.402337e-08, 
    -2.498081e-08, -2.565477e-08, -2.573367e-08, -2.538964e-08, 
    -2.517655e-08, -2.539845e-08,
  -1.304518e-08, -1.336582e-08, -1.415449e-08, -1.463081e-08, -1.53233e-08, 
    -1.601471e-08, -1.728127e-08, -1.871941e-08, -2.083908e-08, 
    -2.313173e-08, -2.465827e-08, -2.588418e-08, -2.627064e-08, 
    -2.602925e-08, -2.553384e-08,
  -1.302943e-08, -1.317002e-08, -1.351439e-08, -1.396635e-08, -1.439965e-08, 
    -1.500009e-08, -1.562503e-08, -1.691278e-08, -1.809791e-08, 
    -2.019374e-08, -2.191523e-08, -2.347051e-08, -2.487409e-08, 
    -2.565576e-08, -2.617313e-08,
  -1.214855e-08, -1.272019e-08, -1.312186e-08, -1.364194e-08, -1.397625e-08, 
    -1.433751e-08, -1.469437e-08, -1.53953e-08, -1.644937e-08, -1.775122e-08, 
    -1.930914e-08, -2.05753e-08, -2.231619e-08, -2.375446e-08, -2.477142e-08,
  -1.00332e-08, -1.139315e-08, -1.22119e-08, -1.282981e-08, -1.345516e-08, 
    -1.394e-08, -1.426374e-08, -1.466241e-08, -1.526538e-08, -1.637369e-08, 
    -1.744198e-08, -1.861591e-08, -1.975255e-08, -2.123025e-08, -2.273576e-08,
  -6.615619e-09, -8.725833e-09, -1.036186e-08, -1.160978e-08, -1.242112e-08, 
    -1.315133e-08, -1.368121e-08, -1.415275e-08, -1.461265e-08, 
    -1.519109e-08, -1.626565e-08, -1.706551e-08, -1.797837e-08, 
    -1.893674e-08, -2.019776e-08,
  -3.786411e-09, -5.309321e-09, -7.19933e-09, -9.073058e-09, -1.064812e-08, 
    -1.187307e-08, -1.280943e-08, -1.340639e-08, -1.396276e-08, 
    -1.459905e-08, -1.515689e-08, -1.607609e-08, -1.678577e-08, 
    -1.757419e-08, -1.828086e-08,
  -2.539094e-09, -3.123817e-09, -4.160997e-09, -5.735924e-09, -7.508779e-09, 
    -9.291507e-09, -1.084407e-08, -1.218523e-08, -1.304789e-08, 
    -1.371539e-08, -1.445357e-08, -1.500604e-08, -1.586842e-08, 
    -1.653425e-08, -1.720716e-08,
  -2.188367e-09, -2.369256e-09, -2.755426e-09, -3.462874e-09, -4.57402e-09, 
    -6.076484e-09, -7.76866e-09, -9.433982e-09, -1.106224e-08, -1.229913e-08, 
    -1.33934e-08, -1.421917e-08, -1.490476e-08, -1.576125e-08, -1.642556e-08,
  -1.799714e-09, -2.017187e-09, -2.229306e-09, -2.512566e-09, -2.988445e-09, 
    -3.742297e-09, -4.902791e-09, -6.363485e-09, -7.978995e-09, 
    -9.605415e-09, -1.110123e-08, -1.251824e-08, -1.377137e-08, 
    -1.466345e-08, -1.551559e-08,
  -1.37081e-08, -1.32244e-08, -1.302158e-08, -1.344873e-08, -1.432092e-08, 
    -1.511184e-08, -1.614787e-08, -1.722229e-08, -1.808692e-08, 
    -1.869205e-08, -1.992387e-08, -2.262187e-08, -2.595859e-08, 
    -2.701913e-08, -2.595416e-08,
  -1.428105e-08, -1.38076e-08, -1.334292e-08, -1.305693e-08, -1.333495e-08, 
    -1.391318e-08, -1.473187e-08, -1.578777e-08, -1.709335e-08, 
    -1.795017e-08, -1.85828e-08, -2.000195e-08, -2.277442e-08, -2.618561e-08, 
    -2.802209e-08,
  -1.418423e-08, -1.431958e-08, -1.393414e-08, -1.346537e-08, -1.3107e-08, 
    -1.315406e-08, -1.359793e-08, -1.436045e-08, -1.550408e-08, 
    -1.686812e-08, -1.774931e-08, -1.840776e-08, -1.959618e-08, 
    -2.210773e-08, -2.497976e-08,
  -1.282068e-08, -1.385335e-08, -1.427285e-08, -1.404226e-08, -1.359344e-08, 
    -1.318046e-08, -1.304556e-08, -1.324138e-08, -1.394581e-08, 
    -1.518879e-08, -1.65524e-08, -1.751759e-08, -1.799486e-08, -1.896972e-08, 
    -2.070336e-08,
  -1.075689e-08, -1.231563e-08, -1.349646e-08, -1.407414e-08, -1.404313e-08, 
    -1.369059e-08, -1.330181e-08, -1.29793e-08, -1.296125e-08, -1.34857e-08, 
    -1.467308e-08, -1.612482e-08, -1.711854e-08, -1.762394e-08, -1.818818e-08,
  -8.801149e-09, -1.040401e-08, -1.184362e-08, -1.30864e-08, -1.378579e-08, 
    -1.389355e-08, -1.36574e-08, -1.3319e-08, -1.294586e-08, -1.275826e-08, 
    -1.299009e-08, -1.396612e-08, -1.53103e-08, -1.646007e-08, -1.702614e-08,
  -6.772708e-09, -8.35157e-09, -9.918745e-09, -1.131585e-08, -1.258187e-08, 
    -1.343256e-08, -1.366486e-08, -1.357479e-08, -1.327659e-08, 
    -1.297356e-08, -1.266591e-08, -1.268095e-08, -1.312286e-08, 
    -1.415219e-08, -1.52615e-08,
  -5.026849e-09, -6.292534e-09, -7.886966e-09, -9.37095e-09, -1.068441e-08, 
    -1.196697e-08, -1.292166e-08, -1.337722e-08, -1.337807e-08, 
    -1.322131e-08, -1.29255e-08, -1.25994e-08, -1.250553e-08, -1.252689e-08, 
    -1.304842e-08,
  -3.498316e-09, -4.585075e-09, -5.807901e-09, -7.368424e-09, -8.776054e-09, 
    -1.000925e-08, -1.126215e-08, -1.229952e-08, -1.296459e-08, 
    -1.313859e-08, -1.311974e-08, -1.285751e-08, -1.260141e-08, 
    -1.240769e-08, -1.224143e-08,
  -2.450779e-09, -3.185999e-09, -4.182273e-09, -5.375986e-09, -6.862532e-09, 
    -8.154451e-09, -9.283931e-09, -1.040899e-08, -1.148859e-08, 
    -1.232404e-08, -1.273042e-08, -1.289027e-08, -1.275096e-08, 
    -1.266174e-08, -1.248164e-08,
  -4.473533e-09, -5.892151e-09, -7.299712e-09, -8.869582e-09, -1.033856e-08, 
    -1.177888e-08, -1.321146e-08, -1.493399e-08, -1.638709e-08, 
    -1.806777e-08, -1.909669e-08, -1.994184e-08, -2.005863e-08, 
    -2.070361e-08, -2.145762e-08,
  -3.589181e-09, -4.839465e-09, -6.321313e-09, -7.79366e-09, -9.436831e-09, 
    -1.092541e-08, -1.226854e-08, -1.381707e-08, -1.542092e-08, 
    -1.683822e-08, -1.838723e-08, -1.945715e-08, -1.989221e-08, 
    -2.009769e-08, -2.126368e-08,
  -2.731501e-09, -3.869347e-09, -5.228538e-09, -6.763984e-09, -8.343789e-09, 
    -1.000596e-08, -1.13938e-08, -1.281608e-08, -1.439337e-08, -1.590134e-08, 
    -1.725341e-08, -1.864191e-08, -1.960525e-08, -1.986768e-08, -2.049961e-08,
  -1.993559e-09, -2.941585e-09, -4.189806e-09, -5.647662e-09, -7.262834e-09, 
    -8.920265e-09, -1.045988e-08, -1.189159e-08, -1.344122e-08, 
    -1.494277e-08, -1.635976e-08, -1.758318e-08, -1.875095e-08, 
    -1.950333e-08, -2.010731e-08,
  -1.470663e-09, -2.160245e-09, -3.185181e-09, -4.544081e-09, -6.075198e-09, 
    -7.801515e-09, -9.445352e-09, -1.093731e-08, -1.253944e-08, 
    -1.411223e-08, -1.561118e-08, -1.671943e-08, -1.771125e-08, 
    -1.861211e-08, -1.939289e-08,
  -1.08432e-09, -1.592249e-09, -2.342233e-09, -3.499048e-09, -4.927684e-09, 
    -6.542366e-09, -8.315497e-09, -9.920379e-09, -1.153237e-08, 
    -1.324275e-08, -1.482434e-08, -1.617366e-08, -1.69344e-08, -1.757884e-08, 
    -1.849339e-08,
  -9.110396e-10, -1.124456e-09, -1.696114e-09, -2.565413e-09, -3.854264e-09, 
    -5.349964e-09, -7.083814e-09, -8.797586e-09, -1.048796e-08, 
    -1.222951e-08, -1.394849e-08, -1.545211e-08, -1.654118e-08, 
    -1.680027e-08, -1.725236e-08,
  -8.872424e-10, -8.980132e-10, -1.178541e-09, -1.854646e-09, -2.833519e-09, 
    -4.189149e-09, -5.818844e-09, -7.62261e-09, -9.363372e-09, -1.114616e-08, 
    -1.299083e-08, -1.463768e-08, -1.598355e-08, -1.66004e-08, -1.652675e-08,
  -9.624473e-10, -8.900085e-10, -9.350595e-10, -1.283587e-09, -2.05189e-09, 
    -3.124128e-09, -4.547197e-09, -6.313801e-09, -8.161376e-09, 
    -1.002052e-08, -1.191044e-08, -1.376032e-08, -1.528728e-08, -1.6326e-08, 
    -1.644628e-08,
  -1.037755e-09, -9.543304e-10, -9.164179e-10, -9.965048e-10, -1.411327e-09, 
    -2.262359e-09, -3.406619e-09, -4.947375e-09, -6.803742e-09, 
    -8.741831e-09, -1.074383e-08, -1.272318e-08, -1.449418e-08, 
    -1.579727e-08, -1.635377e-08,
  -2.630125e-09, -2.516469e-09, -2.648931e-09, -2.913986e-09, -3.307894e-09, 
    -3.83882e-09, -4.387355e-09, -5.327414e-09, -7.110442e-09, -9.01237e-09, 
    -1.149961e-08, -1.383803e-08, -1.575866e-08, -1.710075e-08, -1.813436e-08,
  -1.784827e-09, -1.679447e-09, -1.697197e-09, -1.873832e-09, -2.168718e-09, 
    -2.45058e-09, -2.97591e-09, -3.762255e-09, -4.987313e-09, -6.80104e-09, 
    -9.317001e-09, -1.213628e-08, -1.476298e-08, -1.636478e-08, -1.775511e-08,
  -1.456585e-09, -1.362824e-09, -1.193863e-09, -1.216686e-09, -1.367642e-09, 
    -1.559376e-09, -1.793516e-09, -2.391989e-09, -3.437961e-09, 
    -4.954316e-09, -7.154612e-09, -9.797004e-09, -1.286056e-08, 
    -1.546047e-08, -1.697641e-08,
  -1.132774e-09, -1.175507e-09, -1.108011e-09, -9.844503e-10, -9.337402e-10, 
    -1.003756e-09, -1.141925e-09, -1.433314e-09, -2.057371e-09, 
    -3.184192e-09, -5.118499e-09, -7.714799e-09, -1.067779e-08, 
    -1.374841e-08, -1.600153e-08,
  -9.635136e-10, -9.986947e-10, -1.043205e-09, -1.034846e-09, -9.123978e-10, 
    -8.481046e-10, -8.709609e-10, -1.023166e-09, -1.402228e-09, 
    -2.031678e-09, -3.275465e-09, -5.498075e-09, -8.484626e-09, 
    -1.179034e-08, -1.436833e-08,
  -7.994509e-10, -8.204155e-10, -8.724879e-10, -9.823233e-10, -9.702515e-10, 
    -8.969061e-10, -8.603997e-10, -8.576052e-10, -1.094891e-09, -1.50968e-09, 
    -2.186539e-09, -3.699348e-09, -6.174522e-09, -9.551428e-09, -1.267053e-08,
  -6.407828e-10, -6.286103e-10, -6.937308e-10, -8.309842e-10, -9.615211e-10, 
    -9.638017e-10, -9.474276e-10, -9.171064e-10, -9.615748e-10, -1.25182e-09, 
    -1.675966e-09, -2.529632e-09, -4.415078e-09, -7.246955e-09, -1.058391e-08,
  -5.454447e-10, -5.068272e-10, -5.374891e-10, -6.245761e-10, -8.078871e-10, 
    -9.113378e-10, -9.593186e-10, -9.960279e-10, -9.78465e-10, -1.104011e-09, 
    -1.436963e-09, -1.888364e-09, -3.106572e-09, -5.484416e-09, -8.452514e-09,
  -5.901138e-10, -5.527565e-10, -5.429173e-10, -5.679901e-10, -6.491147e-10, 
    -7.811979e-10, -8.859118e-10, -9.631883e-10, -1.029987e-09, 
    -1.065075e-09, -1.296768e-09, -1.614444e-09, -2.254003e-09, 
    -4.000515e-09, -6.666583e-09,
  -5.938893e-10, -5.249501e-10, -5.005933e-10, -5.052248e-10, -5.472728e-10, 
    -6.432586e-10, -7.3374e-10, -8.94449e-10, -1.007121e-09, -1.082451e-09, 
    -1.213836e-09, -1.467098e-09, -1.852043e-09, -2.885827e-09, -5.117693e-09,
  -1.937113e-08, -1.957631e-08, -2.00319e-08, -2.059189e-08, -2.104612e-08, 
    -2.129923e-08, -2.167275e-08, -2.210091e-08, -2.258759e-08, 
    -2.296687e-08, -2.294701e-08, -2.25449e-08, -2.211248e-08, -2.169955e-08, 
    -2.104766e-08,
  -1.870408e-08, -1.853547e-08, -1.857223e-08, -1.886642e-08, -1.942232e-08, 
    -1.992597e-08, -2.024729e-08, -2.05758e-08, -2.093751e-08, -2.143134e-08, 
    -2.169629e-08, -2.149805e-08, -2.124719e-08, -2.084497e-08, -2.029893e-08,
  -1.615795e-08, -1.746576e-08, -1.775918e-08, -1.746221e-08, -1.743976e-08, 
    -1.794525e-08, -1.855017e-08, -1.905326e-08, -1.944172e-08, 
    -1.983622e-08, -2.02641e-08, -2.023854e-08, -1.993825e-08, -1.963265e-08, 
    -1.933251e-08,
  -1.249562e-08, -1.395818e-08, -1.553e-08, -1.659437e-08, -1.645986e-08, 
    -1.640521e-08, -1.66661e-08, -1.72865e-08, -1.788271e-08, -1.841716e-08, 
    -1.88516e-08, -1.896397e-08, -1.869362e-08, -1.849941e-08, -1.813422e-08,
  -7.563056e-09, -1.025341e-08, -1.180119e-08, -1.319822e-08, -1.47209e-08, 
    -1.549825e-08, -1.545149e-08, -1.562489e-08, -1.602343e-08, 
    -1.656538e-08, -1.710408e-08, -1.759493e-08, -1.753683e-08, 
    -1.742115e-08, -1.718519e-08,
  -3.728302e-09, -5.471136e-09, -7.528466e-09, -9.617231e-09, -1.089011e-08, 
    -1.233493e-08, -1.36004e-08, -1.414771e-08, -1.433373e-08, -1.469849e-08, 
    -1.503366e-08, -1.562672e-08, -1.58371e-08, -1.608355e-08, -1.631759e-08,
  -2.412591e-09, -2.6624e-09, -3.691054e-09, -5.393555e-09, -7.452299e-09, 
    -8.853733e-09, -1.002268e-08, -1.125639e-08, -1.210361e-08, 
    -1.268041e-08, -1.297676e-08, -1.349353e-08, -1.390435e-08, 
    -1.427653e-08, -1.473111e-08,
  -2.16195e-09, -2.124555e-09, -2.137394e-09, -2.574192e-09, -3.721655e-09, 
    -5.418059e-09, -6.961651e-09, -7.968827e-09, -8.953981e-09, 
    -9.906157e-09, -1.056626e-08, -1.107823e-08, -1.161748e-08, 
    -1.215912e-08, -1.269488e-08,
  -1.482021e-09, -1.700525e-09, -1.721065e-09, -1.717157e-09, -1.833756e-09, 
    -2.436384e-09, -3.698098e-09, -5.244475e-09, -6.150995e-09, 
    -6.972181e-09, -7.815087e-09, -8.407627e-09, -8.902749e-09, 
    -9.543445e-09, -1.008799e-08,
  -5.300217e-10, -9.242079e-10, -1.193735e-09, -1.264231e-09, -1.266126e-09, 
    -1.347274e-09, -1.635343e-09, -2.472912e-09, -3.630972e-09, -4.54025e-09, 
    -5.095588e-09, -5.845932e-09, -6.46649e-09, -7.009105e-09, -7.641781e-09,
  -1.877979e-08, -1.744036e-08, -1.572496e-08, -1.474778e-08, -1.379862e-08, 
    -1.354279e-08, -1.267824e-08, -1.194175e-08, -1.165389e-08, 
    -1.183458e-08, -1.184714e-08, -1.202822e-08, -1.282391e-08, 
    -1.457893e-08, -1.651489e-08,
  -1.999472e-08, -1.891548e-08, -1.755792e-08, -1.605231e-08, -1.492275e-08, 
    -1.410187e-08, -1.37432e-08, -1.289277e-08, -1.244781e-08, -1.237145e-08, 
    -1.23711e-08, -1.249817e-08, -1.320689e-08, -1.506009e-08, -1.721617e-08,
  -1.861443e-08, -1.960636e-08, -1.893779e-08, -1.755869e-08, -1.612037e-08, 
    -1.515139e-08, -1.431151e-08, -1.379731e-08, -1.30533e-08, -1.28537e-08, 
    -1.299739e-08, -1.329223e-08, -1.386277e-08, -1.535713e-08, -1.757095e-08,
  -1.547508e-08, -1.720942e-08, -1.896767e-08, -1.933815e-08, -1.77563e-08, 
    -1.633779e-08, -1.541619e-08, -1.460479e-08, -1.394735e-08, -1.34492e-08, 
    -1.343732e-08, -1.379003e-08, -1.455831e-08, -1.571871e-08, -1.783831e-08,
  -1.291504e-08, -1.413852e-08, -1.585565e-08, -1.794116e-08, -1.942684e-08, 
    -1.797619e-08, -1.653422e-08, -1.564733e-08, -1.482374e-08, 
    -1.422001e-08, -1.419476e-08, -1.449629e-08, -1.488459e-08, 
    -1.601288e-08, -1.801716e-08,
  -9.741336e-09, -1.138848e-08, -1.299126e-08, -1.46371e-08, -1.6973e-08, 
    -1.928643e-08, -1.868122e-08, -1.681253e-08, -1.59408e-08, -1.509177e-08, 
    -1.466784e-08, -1.507841e-08, -1.563913e-08, -1.642606e-08, -1.788318e-08,
  -7.029826e-09, -7.837277e-09, -9.794911e-09, -1.176172e-08, -1.367502e-08, 
    -1.606861e-08, -1.867059e-08, -1.92313e-08, -1.732992e-08, -1.624694e-08, 
    -1.540495e-08, -1.539272e-08, -1.578308e-08, -1.683932e-08, -1.797602e-08,
  -5.711774e-09, -5.854096e-09, -6.555297e-09, -8.367603e-09, -1.046296e-08, 
    -1.277121e-08, -1.523734e-08, -1.792129e-08, -1.940571e-08, 
    -1.790723e-08, -1.655406e-08, -1.581846e-08, -1.590494e-08, 
    -1.656589e-08, -1.797528e-08,
  -5.211628e-09, -5.062333e-09, -5.177055e-09, -5.836721e-09, -7.35376e-09, 
    -9.452406e-09, -1.188717e-08, -1.465822e-08, -1.714006e-08, 
    -1.927073e-08, -1.848567e-08, -1.689282e-08, -1.616976e-08, 
    -1.621072e-08, -1.750892e-08,
  -4.889222e-09, -4.667369e-09, -4.570772e-09, -4.610505e-09, -5.270378e-09, 
    -6.514793e-09, -8.340514e-09, -1.084301e-08, -1.377935e-08, 
    -1.625445e-08, -1.877827e-08, -1.884621e-08, -1.722577e-08, 
    -1.638112e-08, -1.67745e-08,
  -1.819753e-08, -1.874272e-08, -1.922194e-08, -1.955225e-08, -2.002673e-08, 
    -2.03279e-08, -2.000899e-08, -1.916744e-08, -1.805029e-08, -1.645646e-08, 
    -1.500603e-08, -1.380337e-08, -1.278992e-08, -1.19267e-08, -1.122605e-08,
  -1.826653e-08, -1.87681e-08, -1.91442e-08, -1.961918e-08, -1.990232e-08, 
    -2.027582e-08, -2.038824e-08, -1.979563e-08, -1.884708e-08, 
    -1.709662e-08, -1.563314e-08, -1.445366e-08, -1.346933e-08, 
    -1.254871e-08, -1.155231e-08,
  -1.853445e-08, -1.897347e-08, -1.937023e-08, -1.971173e-08, -2.00931e-08, 
    -2.038291e-08, -2.057095e-08, -2.038901e-08, -1.952948e-08, 
    -1.826053e-08, -1.670565e-08, -1.540007e-08, -1.428327e-08, 
    -1.301023e-08, -1.197324e-08,
  -1.869808e-08, -1.903292e-08, -1.944177e-08, -1.986075e-08, -2.001219e-08, 
    -2.041671e-08, -2.05207e-08, -2.061913e-08, -2.013098e-08, -1.923592e-08, 
    -1.765488e-08, -1.634194e-08, -1.49402e-08, -1.358748e-08, -1.246132e-08,
  -1.876716e-08, -1.915249e-08, -1.947443e-08, -1.986168e-08, -2.008884e-08, 
    -2.024226e-08, -2.021238e-08, -2.0145e-08, -2.012455e-08, -1.972642e-08, 
    -1.863831e-08, -1.725283e-08, -1.591097e-08, -1.456607e-08, -1.324512e-08,
  -1.808301e-08, -1.870903e-08, -1.921276e-08, -1.956437e-08, -1.986793e-08, 
    -2.002703e-08, -1.998051e-08, -1.968833e-08, -1.959833e-08, 
    -1.962227e-08, -1.906435e-08, -1.803895e-08, -1.674596e-08, 
    -1.555111e-08, -1.427712e-08,
  -1.678407e-08, -1.754646e-08, -1.815597e-08, -1.868893e-08, -1.90884e-08, 
    -1.93856e-08, -1.930944e-08, -1.90659e-08, -1.880757e-08, -1.876739e-08, 
    -1.87867e-08, -1.823691e-08, -1.726016e-08, -1.614887e-08, -1.51008e-08,
  -1.52961e-08, -1.60682e-08, -1.668204e-08, -1.723154e-08, -1.772887e-08, 
    -1.826763e-08, -1.842158e-08, -1.82223e-08, -1.801918e-08, -1.771788e-08, 
    -1.781366e-08, -1.773573e-08, -1.737891e-08, -1.646052e-08, -1.54832e-08,
  -1.339422e-08, -1.419511e-08, -1.489718e-08, -1.550799e-08, -1.597865e-08, 
    -1.65402e-08, -1.699689e-08, -1.715383e-08, -1.699601e-08, -1.680745e-08, 
    -1.660542e-08, -1.679104e-08, -1.68654e-08, -1.655914e-08, -1.587446e-08,
  -1.266863e-08, -1.277191e-08, -1.302984e-08, -1.344192e-08, -1.39869e-08, 
    -1.450587e-08, -1.512838e-08, -1.551573e-08, -1.56512e-08, -1.555865e-08, 
    -1.550178e-08, -1.54066e-08, -1.5725e-08, -1.601257e-08, -1.595891e-08,
  -1.43031e-08, -1.522147e-08, -1.552716e-08, -1.546927e-08, -1.514627e-08, 
    -1.500655e-08, -1.499672e-08, -1.608207e-08, -1.710154e-08, 
    -1.793851e-08, -1.837856e-08, -1.857209e-08, -1.866901e-08, 
    -1.849525e-08, -1.791449e-08,
  -1.367795e-08, -1.451983e-08, -1.508384e-08, -1.54205e-08, -1.532962e-08, 
    -1.491987e-08, -1.466706e-08, -1.501633e-08, -1.605883e-08, 
    -1.702051e-08, -1.784574e-08, -1.827511e-08, -1.853424e-08, 
    -1.816732e-08, -1.761847e-08,
  -1.337794e-08, -1.391688e-08, -1.456694e-08, -1.503607e-08, -1.500042e-08, 
    -1.493098e-08, -1.457327e-08, -1.457348e-08, -1.513112e-08, 
    -1.577778e-08, -1.671132e-08, -1.751434e-08, -1.802346e-08, 
    -1.782545e-08, -1.759551e-08,
  -1.294414e-08, -1.346512e-08, -1.399474e-08, -1.439114e-08, -1.455656e-08, 
    -1.470206e-08, -1.459818e-08, -1.446338e-08, -1.462458e-08, 
    -1.501816e-08, -1.573055e-08, -1.685552e-08, -1.765146e-08, 
    -1.782986e-08, -1.792295e-08,
  -1.270971e-08, -1.308747e-08, -1.356135e-08, -1.390961e-08, -1.40246e-08, 
    -1.414613e-08, -1.424515e-08, -1.424462e-08, -1.42929e-08, -1.458004e-08, 
    -1.541205e-08, -1.652219e-08, -1.73147e-08, -1.770128e-08, -1.815063e-08,
  -1.188144e-08, -1.257383e-08, -1.305925e-08, -1.331488e-08, -1.343666e-08, 
    -1.348035e-08, -1.376872e-08, -1.402683e-08, -1.417017e-08, 
    -1.472632e-08, -1.548523e-08, -1.647738e-08, -1.726597e-08, 
    -1.776492e-08, -1.817666e-08,
  -1.12302e-08, -1.173596e-08, -1.228966e-08, -1.278717e-08, -1.311544e-08, 
    -1.309609e-08, -1.31999e-08, -1.343375e-08, -1.404425e-08, -1.491713e-08, 
    -1.585128e-08, -1.667695e-08, -1.730958e-08, -1.770235e-08, -1.806932e-08,
  -1.108183e-08, -1.130057e-08, -1.171317e-08, -1.223362e-08, -1.24111e-08, 
    -1.230768e-08, -1.231124e-08, -1.289504e-08, -1.382974e-08, 
    -1.479256e-08, -1.577704e-08, -1.658311e-08, -1.714421e-08, -1.76299e-08, 
    -1.80026e-08,
  -1.036627e-08, -1.074072e-08, -1.119536e-08, -1.166562e-08, -1.181269e-08, 
    -1.178849e-08, -1.193933e-08, -1.263873e-08, -1.368931e-08, 
    -1.464659e-08, -1.536627e-08, -1.603436e-08, -1.677561e-08, 
    -1.744645e-08, -1.786977e-08,
  -9.811882e-09, -1.022186e-08, -1.081697e-08, -1.14729e-08, -1.195346e-08, 
    -1.207692e-08, -1.213053e-08, -1.24413e-08, -1.324898e-08, -1.410164e-08, 
    -1.484778e-08, -1.564056e-08, -1.632776e-08, -1.6888e-08, -1.73524e-08,
  -1.021984e-08, -1.081445e-08, -1.148717e-08, -1.227528e-08, -1.339787e-08, 
    -1.497998e-08, -1.614025e-08, -1.703275e-08, -1.795251e-08, 
    -1.884897e-08, -1.951392e-08, -1.994146e-08, -2.02617e-08, -2.074055e-08, 
    -2.123333e-08,
  -8.71534e-09, -9.767512e-09, -1.06563e-08, -1.14603e-08, -1.207048e-08, 
    -1.309918e-08, -1.456976e-08, -1.562876e-08, -1.647112e-08, 
    -1.719078e-08, -1.790099e-08, -1.843946e-08, -1.88361e-08, -1.940096e-08, 
    -1.981159e-08,
  -7.746703e-09, -8.672211e-09, -9.624176e-09, -1.049077e-08, -1.122941e-08, 
    -1.182104e-08, -1.279211e-08, -1.406174e-08, -1.501727e-08, 
    -1.576757e-08, -1.646686e-08, -1.710073e-08, -1.77e-08, -1.835415e-08, 
    -1.862402e-08,
  -7.102433e-09, -7.83056e-09, -8.723378e-09, -9.568058e-09, -1.031389e-08, 
    -1.088139e-08, -1.153419e-08, -1.247283e-08, -1.355951e-08, 
    -1.453231e-08, -1.525187e-08, -1.572196e-08, -1.630176e-08, -1.69197e-08, 
    -1.710635e-08,
  -6.16503e-09, -7.167651e-09, -7.835878e-09, -8.707062e-09, -9.499312e-09, 
    -1.013526e-08, -1.069674e-08, -1.14122e-08, -1.225774e-08, -1.310011e-08, 
    -1.378817e-08, -1.429934e-08, -1.495561e-08, -1.554058e-08, -1.58012e-08,
  -5.416063e-09, -6.427752e-09, -7.310406e-09, -7.982333e-09, -8.761192e-09, 
    -9.534817e-09, -1.02438e-08, -1.10041e-08, -1.167081e-08, -1.210904e-08, 
    -1.243252e-08, -1.27753e-08, -1.333626e-08, -1.392928e-08, -1.442352e-08,
  -5.003024e-09, -5.568734e-09, -6.431891e-09, -7.240239e-09, -7.901575e-09, 
    -8.833238e-09, -9.900917e-09, -1.083504e-08, -1.131215e-08, 
    -1.146732e-08, -1.152073e-08, -1.172424e-08, -1.214887e-08, -1.25709e-08, 
    -1.30263e-08,
  -4.843306e-09, -5.41026e-09, -6.016418e-09, -6.781099e-09, -7.706026e-09, 
    -8.625239e-09, -9.57011e-09, -1.022578e-08, -1.051903e-08, -1.064332e-08, 
    -1.080085e-08, -1.107116e-08, -1.14698e-08, -1.178956e-08, -1.21194e-08,
  -4.562766e-09, -5.03299e-09, -5.625915e-09, -6.310364e-09, -7.200436e-09, 
    -7.996475e-09, -8.642494e-09, -9.157138e-09, -9.551191e-09, 
    -9.891774e-09, -1.033637e-08, -1.078756e-08, -1.115643e-08, 
    -1.147698e-08, -1.178712e-08,
  -4.773225e-09, -4.930951e-09, -5.269156e-09, -5.708958e-09, -6.331632e-09, 
    -6.937983e-09, -7.387027e-09, -7.836927e-09, -8.401761e-09, 
    -9.096217e-09, -9.757445e-09, -1.021669e-08, -1.069407e-08, 
    -1.109758e-08, -1.148416e-08,
  -5.809216e-09, -6.530687e-09, -7.335999e-09, -8.394766e-09, -9.578002e-09, 
    -1.089899e-08, -1.193504e-08, -1.307074e-08, -1.422383e-08, 
    -1.580797e-08, -1.718319e-08, -1.842301e-08, -1.915145e-08, 
    -1.963988e-08, -2.014036e-08,
  -4.255667e-09, -5.16852e-09, -5.908094e-09, -6.721375e-09, -7.65603e-09, 
    -8.629085e-09, -9.588739e-09, -1.073547e-08, -1.200866e-08, 
    -1.331054e-08, -1.453779e-08, -1.584632e-08, -1.699653e-08, 
    -1.785008e-08, -1.844782e-08,
  -3.489935e-09, -3.823965e-09, -4.633792e-09, -5.372863e-09, -6.10507e-09, 
    -6.949823e-09, -7.673467e-09, -8.562623e-09, -9.679063e-09, 
    -1.087705e-08, -1.20207e-08, -1.306874e-08, -1.421322e-08, -1.526794e-08, 
    -1.627198e-08,
  -3.572558e-09, -3.429186e-09, -3.533301e-09, -4.129548e-09, -4.831122e-09, 
    -5.542101e-09, -6.208382e-09, -6.817043e-09, -7.610173e-09, 
    -8.594976e-09, -9.618766e-09, -1.060244e-08, -1.166508e-08, 
    -1.263431e-08, -1.362869e-08,
  -3.826671e-09, -3.658864e-09, -3.458398e-09, -3.446236e-09, -3.738644e-09, 
    -4.295152e-09, -4.982084e-09, -5.553875e-09, -6.128931e-09, 
    -6.819606e-09, -7.639374e-09, -8.494657e-09, -9.385689e-09, -1.03168e-08, 
    -1.125582e-08,
  -3.867041e-09, -3.81597e-09, -3.712321e-09, -3.555983e-09, -3.509538e-09, 
    -3.639442e-09, -4.033351e-09, -4.549571e-09, -5.089482e-09, 
    -5.657383e-09, -6.177645e-09, -6.846148e-09, -7.592923e-09, 
    -8.394413e-09, -9.181267e-09,
  -3.431315e-09, -3.534874e-09, -3.645686e-09, -3.646936e-09, -3.602149e-09, 
    -3.62608e-09, -3.76652e-09, -4.04187e-09, -4.398545e-09, -4.864205e-09, 
    -5.364562e-09, -5.820129e-09, -6.363486e-09, -6.972852e-09, -7.649588e-09,
  -2.983236e-09, -3.021763e-09, -3.129276e-09, -3.316831e-09, -3.45124e-09, 
    -3.516473e-09, -3.660977e-09, -3.873951e-09, -4.139501e-09, -4.42861e-09, 
    -4.82106e-09, -5.240021e-09, -5.679696e-09, -6.135862e-09, -6.64456e-09,
  -2.452345e-09, -2.485204e-09, -2.555576e-09, -2.704519e-09, -2.900845e-09, 
    -3.106719e-09, -3.321807e-09, -3.555807e-09, -3.835016e-09, 
    -4.128057e-09, -4.423852e-09, -4.739949e-09, -5.128671e-09, 
    -5.582604e-09, -6.037081e-09,
  -2.106449e-09, -2.090579e-09, -2.137593e-09, -2.259899e-09, -2.429859e-09, 
    -2.651585e-09, -2.858707e-09, -3.050711e-09, -3.299946e-09, 
    -3.644546e-09, -4.001828e-09, -4.325069e-09, -4.653333e-09, 
    -5.060909e-09, -5.523924e-09,
  -1.5263e-08, -1.632145e-08, -1.705046e-08, -1.755773e-08, -1.83768e-08, 
    -1.845037e-08, -1.879662e-08, -1.932969e-08, -1.98872e-08, -2.044605e-08, 
    -2.102917e-08, -2.155841e-08, -2.173917e-08, -2.18421e-08, -2.218032e-08,
  -1.360504e-08, -1.501609e-08, -1.634e-08, -1.717127e-08, -1.780384e-08, 
    -1.858568e-08, -1.910064e-08, -1.961831e-08, -2.002229e-08, 
    -2.028059e-08, -2.03692e-08, -2.061985e-08, -2.111432e-08, -2.156679e-08, 
    -2.181561e-08,
  -1.132523e-08, -1.304275e-08, -1.470238e-08, -1.617102e-08, -1.707958e-08, 
    -1.753038e-08, -1.807699e-08, -1.868999e-08, -1.92716e-08, -1.985195e-08, 
    -2.01855e-08, -2.018284e-08, -1.998256e-08, -1.999839e-08, -2.032018e-08,
  -9.016103e-09, -1.048141e-08, -1.215361e-08, -1.399599e-08, -1.570308e-08, 
    -1.68886e-08, -1.715905e-08, -1.750963e-08, -1.797802e-08, -1.85707e-08, 
    -1.924175e-08, -1.977496e-08, -1.988965e-08, -1.950623e-08, -1.932396e-08,
  -7.55278e-09, -8.524225e-09, -9.63861e-09, -1.107923e-08, -1.279224e-08, 
    -1.474118e-08, -1.618555e-08, -1.678306e-08, -1.700364e-08, 
    -1.727547e-08, -1.772545e-08, -1.835113e-08, -1.905237e-08, 
    -1.938922e-08, -1.898456e-08,
  -6.638772e-09, -7.196472e-09, -7.968088e-09, -8.899879e-09, -9.988248e-09, 
    -1.147178e-08, -1.321302e-08, -1.479504e-08, -1.572022e-08, 
    -1.622654e-08, -1.646585e-08, -1.676487e-08, -1.725857e-08, 
    -1.792217e-08, -1.828578e-08,
  -5.981158e-09, -6.397274e-09, -6.838012e-09, -7.452254e-09, -8.077308e-09, 
    -8.865745e-09, -1.003635e-08, -1.156169e-08, -1.303164e-08, -1.41557e-08, 
    -1.482155e-08, -1.515973e-08, -1.539214e-08, -1.58084e-08, -1.641347e-08,
  -5.499755e-09, -5.839736e-09, -6.225107e-09, -6.606014e-09, -7.063073e-09, 
    -7.473844e-09, -7.98237e-09, -8.845058e-09, -1.001145e-08, -1.130887e-08, 
    -1.247159e-08, -1.315577e-08, -1.352423e-08, -1.374245e-08, -1.401426e-08,
  -5.263703e-09, -5.451263e-09, -5.733118e-09, -6.050618e-09, -6.399537e-09, 
    -6.726088e-09, -6.99526e-09, -7.351612e-09, -7.89113e-09, -8.617538e-09, 
    -9.617658e-09, -1.060368e-08, -1.131049e-08, -1.172397e-08, -1.198789e-08,
  -4.965786e-09, -5.131996e-09, -5.314942e-09, -5.553455e-09, -5.819034e-09, 
    -6.080238e-09, -6.301053e-09, -6.527539e-09, -6.783652e-09, 
    -7.101666e-09, -7.526366e-09, -8.195371e-09, -8.880067e-09, 
    -9.481602e-09, -9.84207e-09,
  -4.921008e-09, -5.795869e-09, -7.620245e-09, -8.732003e-09, -9.841622e-09, 
    -1.113118e-08, -1.247839e-08, -1.353516e-08, -1.474303e-08, 
    -1.570079e-08, -1.645492e-08, -1.756703e-08, -1.866353e-08, -1.94409e-08, 
    -2.004901e-08,
  -4.501955e-09, -5.141448e-09, -6.40103e-09, -7.919321e-09, -9.072187e-09, 
    -1.021023e-08, -1.152199e-08, -1.272506e-08, -1.38498e-08, -1.507098e-08, 
    -1.606094e-08, -1.695201e-08, -1.789618e-08, -1.871689e-08, -1.942083e-08,
  -4.088749e-09, -4.651972e-09, -5.406227e-09, -6.883647e-09, -8.319859e-09, 
    -9.417072e-09, -1.062681e-08, -1.181004e-08, -1.299384e-08, 
    -1.415281e-08, -1.531998e-08, -1.639621e-08, -1.742988e-08, 
    -1.821137e-08, -1.882725e-08,
  -3.746795e-09, -4.300758e-09, -4.845079e-09, -5.763702e-09, -7.316976e-09, 
    -8.647014e-09, -9.778602e-09, -1.098796e-08, -1.208324e-08, 
    -1.332703e-08, -1.443671e-08, -1.550604e-08, -1.672736e-08, 
    -1.783219e-08, -1.856168e-08,
  -3.428088e-09, -3.959698e-09, -4.526799e-09, -5.086414e-09, -6.185853e-09, 
    -7.76423e-09, -9.005921e-09, -1.016447e-08, -1.130143e-08, -1.238512e-08, 
    -1.368053e-08, -1.468136e-08, -1.569944e-08, -1.702468e-08, -1.805623e-08,
  -3.198656e-09, -3.636178e-09, -4.164904e-09, -4.705639e-09, -5.354711e-09, 
    -6.624906e-09, -8.191917e-09, -9.416195e-09, -1.057859e-08, 
    -1.162544e-08, -1.276143e-08, -1.395729e-08, -1.487782e-08, 
    -1.590924e-08, -1.721368e-08,
  -3.131167e-09, -3.352628e-09, -3.864783e-09, -4.40629e-09, -4.940619e-09, 
    -5.730975e-09, -7.065712e-09, -8.570984e-09, -9.846115e-09, 
    -1.093771e-08, -1.199006e-08, -1.31466e-08, -1.415127e-08, -1.508655e-08, 
    -1.605448e-08,
  -3.179066e-09, -3.306922e-09, -3.557878e-09, -4.059111e-09, -4.611346e-09, 
    -5.241395e-09, -6.157619e-09, -7.528154e-09, -9.022404e-09, 
    -1.029086e-08, -1.125893e-08, -1.239342e-08, -1.344421e-08, 
    -1.441184e-08, -1.535029e-08,
  -3.162442e-09, -3.302886e-09, -3.513422e-09, -3.838351e-09, -4.296316e-09, 
    -4.843141e-09, -5.510021e-09, -6.556172e-09, -7.952695e-09, 
    -9.443846e-09, -1.069326e-08, -1.168139e-08, -1.275614e-08, 
    -1.366682e-08, -1.466492e-08,
  -3.604727e-09, -3.471285e-09, -3.405408e-09, -3.710701e-09, -4.117465e-09, 
    -4.576945e-09, -5.12455e-09, -5.795219e-09, -6.951188e-09, -8.374207e-09, 
    -9.756099e-09, -1.097816e-08, -1.200332e-08, -1.295765e-08, -1.387448e-08,
  -1.008333e-09, -1.128308e-09, -1.340079e-09, -1.591752e-09, -1.854463e-09, 
    -2.216912e-09, -2.689991e-09, -3.15334e-09, -3.739639e-09, -4.550551e-09, 
    -5.335538e-09, -6.162525e-09, -7.327766e-09, -8.45447e-09, -9.629507e-09,
  -9.999888e-10, -1.055103e-09, -1.14989e-09, -1.342942e-09, -1.615524e-09, 
    -1.9077e-09, -2.294829e-09, -2.768942e-09, -3.230603e-09, -3.904238e-09, 
    -4.730242e-09, -5.505379e-09, -6.435202e-09, -7.673781e-09, -8.786735e-09,
  -1.191274e-09, -1.079422e-09, -1.077794e-09, -1.147555e-09, -1.315762e-09, 
    -1.613594e-09, -1.943858e-09, -2.423893e-09, -2.864053e-09, -3.35883e-09, 
    -4.171734e-09, -4.984318e-09, -5.719746e-09, -6.74962e-09, -7.973538e-09,
  -1.595234e-09, -1.391101e-09, -1.219551e-09, -1.169782e-09, -1.194275e-09, 
    -1.361427e-09, -1.626652e-09, -2.022958e-09, -2.515158e-09, 
    -2.871497e-09, -3.476545e-09, -4.370749e-09, -5.159642e-09, 
    -5.910319e-09, -7.022403e-09,
  -2.01431e-09, -1.792113e-09, -1.56948e-09, -1.380228e-09, -1.266878e-09, 
    -1.273977e-09, -1.429163e-09, -1.664771e-09, -2.165124e-09, 
    -2.612179e-09, -2.967276e-09, -3.688531e-09, -4.598774e-09, 
    -5.358717e-09, -6.201033e-09,
  -2.350766e-09, -2.103566e-09, -1.8322e-09, -1.630781e-09, -1.446981e-09, 
    -1.332699e-09, -1.332451e-09, -1.446995e-09, -1.700166e-09, 
    -2.253446e-09, -2.635196e-09, -3.146388e-09, -3.941027e-09, 
    -4.841631e-09, -5.575698e-09,
  -2.586124e-09, -2.363996e-09, -2.085773e-09, -1.826451e-09, -1.619699e-09, 
    -1.441062e-09, -1.357413e-09, -1.347015e-09, -1.440714e-09, 
    -1.757244e-09, -2.306169e-09, -2.714976e-09, -3.429965e-09, 
    -4.255608e-09, -5.071319e-09,
  -2.715995e-09, -2.580082e-09, -2.336381e-09, -2.037551e-09, -1.782714e-09, 
    -1.564843e-09, -1.420513e-09, -1.346553e-09, -1.352939e-09, 
    -1.473512e-09, -1.878682e-09, -2.399789e-09, -2.933688e-09, -3.78207e-09, 
    -4.586413e-09,
  -2.898739e-09, -2.658448e-09, -2.521886e-09, -2.254174e-09, -1.956956e-09, 
    -1.691118e-09, -1.511373e-09, -1.412908e-09, -1.37063e-09, -1.410616e-09, 
    -1.581546e-09, -2.091242e-09, -2.613544e-09, -3.328958e-09, -4.188023e-09,
  -2.902821e-09, -2.609723e-09, -2.464659e-09, -2.362723e-09, -2.140991e-09, 
    -1.869938e-09, -1.639678e-09, -1.497986e-09, -1.419525e-09, 
    -1.420889e-09, -1.488545e-09, -1.749869e-09, -2.345397e-09, 
    -2.955061e-09, -3.774731e-09,
  -1.614745e-09, -1.648367e-09, -1.702043e-09, -1.797224e-09, -1.884487e-09, 
    -1.997476e-09, -2.141018e-09, -2.321846e-09, -2.497668e-09, 
    -2.708295e-09, -2.882074e-09, -3.126798e-09, -3.464642e-09, 
    -3.919206e-09, -4.54855e-09,
  -1.381457e-09, -1.410912e-09, -1.457676e-09, -1.525977e-09, -1.60986e-09, 
    -1.687847e-09, -1.773165e-09, -1.913654e-09, -2.086411e-09, 
    -2.298461e-09, -2.516397e-09, -2.722735e-09, -2.970266e-09, 
    -3.242251e-09, -3.603275e-09,
  -1.268913e-09, -1.286755e-09, -1.30438e-09, -1.341528e-09, -1.403386e-09, 
    -1.482068e-09, -1.563809e-09, -1.656353e-09, -1.768824e-09, 
    -1.926329e-09, -2.112894e-09, -2.334928e-09, -2.560174e-09, 
    -2.800888e-09, -3.084296e-09,
  -1.223599e-09, -1.218072e-09, -1.223748e-09, -1.239128e-09, -1.265221e-09, 
    -1.316139e-09, -1.380603e-09, -1.460329e-09, -1.558652e-09, 
    -1.681135e-09, -1.834069e-09, -2.014923e-09, -2.231418e-09, 
    -2.452341e-09, -2.690726e-09,
  -1.439298e-09, -1.409657e-09, -1.364316e-09, -1.319749e-09, -1.29053e-09, 
    -1.27437e-09, -1.285708e-09, -1.319821e-09, -1.367497e-09, -1.441906e-09, 
    -1.560417e-09, -1.723539e-09, -1.919462e-09, -2.145203e-09, -2.38298e-09,
  -1.772951e-09, -1.776925e-09, -1.743924e-09, -1.660456e-09, -1.5575e-09, 
    -1.454874e-09, -1.368714e-09, -1.297888e-09, -1.282179e-09, 
    -1.297891e-09, -1.338342e-09, -1.431019e-09, -1.578777e-09, -1.78975e-09, 
    -2.05569e-09,
  -2.166414e-09, -2.193349e-09, -2.203647e-09, -2.182085e-09, -2.089352e-09, 
    -1.925919e-09, -1.725279e-09, -1.544492e-09, -1.367562e-09, 
    -1.262192e-09, -1.231933e-09, -1.244477e-09, -1.313339e-09, 
    -1.440011e-09, -1.662082e-09,
  -2.494491e-09, -2.587815e-09, -2.639144e-09, -2.687063e-09, -2.661486e-09, 
    -2.586204e-09, -2.426973e-09, -2.141402e-09, -1.83997e-09, -1.523723e-09, 
    -1.307367e-09, -1.207366e-09, -1.18696e-09, -1.228409e-09, -1.326447e-09,
  -2.745331e-09, -2.881188e-09, -2.988629e-09, -3.048909e-09, -3.105485e-09, 
    -3.120989e-09, -3.081834e-09, -2.990885e-09, -2.768786e-09, 
    -2.432466e-09, -1.955678e-09, -1.526386e-09, -1.277327e-09, 
    -1.186411e-09, -1.188102e-09,
  -3.155286e-09, -3.298553e-09, -3.356582e-09, -3.351211e-09, -3.329574e-09, 
    -3.370638e-09, -3.383e-09, -3.378148e-09, -3.285484e-09, -3.14925e-09, 
    -2.954454e-09, -2.555261e-09, -2.047112e-09, -1.54996e-09, -1.277163e-09,
  -7.250362e-09, -7.602225e-09, -7.795323e-09, -7.933942e-09, -8.020026e-09, 
    -8.074775e-09, -8.143027e-09, -8.236862e-09, -8.364099e-09, -8.53548e-09, 
    -8.722703e-09, -8.959846e-09, -9.218549e-09, -9.524548e-09, -9.925778e-09,
  -4.925489e-09, -5.276196e-09, -5.768324e-09, -6.04465e-09, -6.193272e-09, 
    -6.25061e-09, -6.282098e-09, -6.255937e-09, -6.275993e-09, -6.306302e-09, 
    -6.363355e-09, -6.439187e-09, -6.579016e-09, -6.767635e-09, -7.011253e-09,
  -3.682455e-09, -3.834212e-09, -4.052305e-09, -4.357721e-09, -4.583465e-09, 
    -4.738783e-09, -4.826119e-09, -4.85075e-09, -4.839354e-09, -4.808263e-09, 
    -4.775826e-09, -4.753059e-09, -4.758428e-09, -4.78922e-09, -4.8515e-09,
  -2.685431e-09, -2.783876e-09, -2.878968e-09, -3.018923e-09, -3.189151e-09, 
    -3.349764e-09, -3.494114e-09, -3.574932e-09, -3.61678e-09, -3.61654e-09, 
    -3.598764e-09, -3.573395e-09, -3.553911e-09, -3.554015e-09, -3.57268e-09,
  -2.003143e-09, -2.089134e-09, -2.18145e-09, -2.266973e-09, -2.360302e-09, 
    -2.463255e-09, -2.558993e-09, -2.638293e-09, -2.684008e-09, 
    -2.708293e-09, -2.72412e-09, -2.728753e-09, -2.73376e-09, -2.733595e-09, 
    -2.73978e-09,
  -1.528686e-09, -1.611324e-09, -1.700167e-09, -1.784847e-09, -1.853811e-09, 
    -1.914795e-09, -1.973095e-09, -2.026189e-09, -2.064282e-09, 
    -2.097611e-09, -2.124982e-09, -2.144994e-09, -2.158006e-09, 
    -2.161262e-09, -2.159143e-09,
  -1.172365e-09, -1.261714e-09, -1.362161e-09, -1.454189e-09, -1.528835e-09, 
    -1.583709e-09, -1.628146e-09, -1.664442e-09, -1.703609e-09, 
    -1.738779e-09, -1.774463e-09, -1.802675e-09, -1.822337e-09, 
    -1.833822e-09, -1.830407e-09,
  -9.471753e-10, -1.021706e-09, -1.108083e-09, -1.186647e-09, -1.254986e-09, 
    -1.304531e-09, -1.346322e-09, -1.389108e-09, -1.436056e-09, 
    -1.484204e-09, -1.524805e-09, -1.558121e-09, -1.584637e-09, 
    -1.608526e-09, -1.624081e-09,
  -7.661678e-10, -8.357574e-10, -9.122521e-10, -9.844834e-10, -1.04652e-09, 
    -1.097214e-09, -1.149163e-09, -1.20248e-09, -1.254062e-09, -1.30659e-09, 
    -1.350008e-09, -1.38804e-09, -1.418005e-09, -1.43994e-09, -1.458545e-09,
  -6.277062e-10, -6.940595e-10, -7.746727e-10, -8.595004e-10, -9.395793e-10, 
    -1.010991e-09, -1.082818e-09, -1.161819e-09, -1.236743e-09, 
    -1.299148e-09, -1.339059e-09, -1.362532e-09, -1.369847e-09, 
    -1.369178e-09, -1.367202e-09,
  -1.535545e-08, -1.756053e-08, -1.915667e-08, -2.054528e-08, -2.198501e-08, 
    -2.318536e-08, -2.37626e-08, -2.388783e-08, -2.411942e-08, -2.487968e-08, 
    -2.558366e-08, -2.603675e-08, -2.627686e-08, -2.600886e-08, -2.553753e-08,
  -1.046926e-08, -1.391563e-08, -1.663757e-08, -1.838332e-08, -1.988441e-08, 
    -2.136749e-08, -2.248562e-08, -2.307455e-08, -2.315995e-08, 
    -2.316708e-08, -2.380041e-08, -2.439057e-08, -2.490897e-08, 
    -2.538309e-08, -2.562901e-08,
  -7.630777e-09, -9.440869e-09, -1.258709e-08, -1.554207e-08, -1.733548e-08, 
    -1.895284e-08, -2.051747e-08, -2.159771e-08, -2.225568e-08, 
    -2.223691e-08, -2.222492e-08, -2.262435e-08, -2.310523e-08, 
    -2.361233e-08, -2.405683e-08,
  -5.802045e-09, -6.776987e-09, -8.431886e-09, -1.125513e-08, -1.443249e-08, 
    -1.623319e-08, -1.78535e-08, -1.939839e-08, -2.056601e-08, -2.12036e-08, 
    -2.12597e-08, -2.112955e-08, -2.123659e-08, -2.161261e-08, -2.20135e-08,
  -4.537163e-09, -5.16782e-09, -6.203853e-09, -7.41651e-09, -9.779616e-09, 
    -1.295658e-08, -1.497568e-08, -1.641297e-08, -1.807952e-08, -1.93408e-08, 
    -2.001138e-08, -2.02999e-08, -2.001679e-08, -1.989474e-08, -2.004822e-08,
  -3.628164e-09, -4.215892e-09, -4.858873e-09, -5.733971e-09, -6.715283e-09, 
    -8.390402e-09, -1.132372e-08, -1.352843e-08, -1.48556e-08, -1.65009e-08, 
    -1.776773e-08, -1.851633e-08, -1.891046e-08, -1.877827e-08, -1.858471e-08,
  -3.052664e-09, -3.392099e-09, -3.863689e-09, -4.500167e-09, -5.20546e-09, 
    -6.003617e-09, -7.400273e-09, -9.900147e-09, -1.204412e-08, 
    -1.340305e-08, -1.474382e-08, -1.599067e-08, -1.680697e-08, 
    -1.724654e-08, -1.733737e-08,
  -2.358066e-09, -2.669907e-09, -3.087336e-09, -3.612358e-09, -4.068213e-09, 
    -4.568105e-09, -5.26907e-09, -6.481335e-09, -8.601399e-09, -1.051451e-08, 
    -1.193762e-08, -1.303308e-08, -1.411186e-08, -1.484578e-08, -1.536699e-08,
  -1.733952e-09, -1.952346e-09, -2.263525e-09, -2.705721e-09, -3.236503e-09, 
    -3.700684e-09, -4.032662e-09, -4.585301e-09, -5.581149e-09, 
    -7.292274e-09, -8.936128e-09, -1.034334e-08, -1.135162e-08, 
    -1.217013e-08, -1.28189e-08,
  -1.401593e-09, -1.474531e-09, -1.663804e-09, -1.943213e-09, -2.30895e-09, 
    -2.792234e-09, -3.215231e-09, -3.578798e-09, -3.986273e-09, 
    -4.734467e-09, -6.052456e-09, -7.428247e-09, -8.725388e-09, 
    -9.635806e-09, -1.022784e-08,
  -1.15894e-08, -1.249793e-08, -1.454171e-08, -1.68238e-08, -1.91553e-08, 
    -2.095734e-08, -2.26767e-08, -2.466663e-08, -2.535448e-08, -2.573073e-08, 
    -2.595825e-08, -2.678513e-08, -2.651872e-08, -2.497547e-08, -2.379799e-08,
  -1.103119e-08, -1.107675e-08, -1.1776e-08, -1.353484e-08, -1.606324e-08, 
    -1.889691e-08, -2.052475e-08, -2.207871e-08, -2.408565e-08, 
    -2.533937e-08, -2.595809e-08, -2.611858e-08, -2.670051e-08, 
    -2.682117e-08, -2.54545e-08,
  -1.166589e-08, -1.097719e-08, -1.108192e-08, -1.171043e-08, -1.287609e-08, 
    -1.526241e-08, -1.83213e-08, -2.007365e-08, -2.162593e-08, -2.351153e-08, 
    -2.507752e-08, -2.594596e-08, -2.608974e-08, -2.659177e-08, -2.658014e-08,
  -1.095868e-08, -1.124041e-08, -1.061779e-08, -1.088111e-08, -1.174575e-08, 
    -1.258842e-08, -1.453195e-08, -1.757906e-08, -1.98618e-08, -2.170643e-08, 
    -2.352256e-08, -2.504118e-08, -2.586666e-08, -2.628301e-08, -2.662899e-08,
  -9.33402e-09, -1.056629e-08, -1.119394e-08, -1.09224e-08, -1.083149e-08, 
    -1.168756e-08, -1.248947e-08, -1.413104e-08, -1.706634e-08, 
    -1.964337e-08, -2.192717e-08, -2.370919e-08, -2.502488e-08, 
    -2.571707e-08, -2.641386e-08,
  -7.685534e-09, -8.686173e-09, -9.6359e-09, -1.07432e-08, -1.126795e-08, 
    -1.109098e-08, -1.132434e-08, -1.23218e-08, -1.407405e-08, -1.686725e-08, 
    -1.962793e-08, -2.207325e-08, -2.403203e-08, -2.501897e-08, -2.556502e-08,
  -6.027068e-09, -6.798733e-09, -7.669625e-09, -8.772429e-09, -9.880654e-09, 
    -1.100647e-08, -1.196748e-08, -1.158763e-08, -1.238136e-08, 
    -1.416868e-08, -1.673942e-08, -1.953215e-08, -2.206235e-08, 
    -2.409935e-08, -2.500517e-08,
  -4.391346e-09, -5.133376e-09, -5.876596e-09, -6.740189e-09, -7.906327e-09, 
    -8.869367e-09, -1.00835e-08, -1.16717e-08, -1.23787e-08, -1.323283e-08, 
    -1.447359e-08, -1.676015e-08, -1.937443e-08, -2.197772e-08, -2.405643e-08,
  -2.923924e-09, -3.636085e-09, -4.43959e-09, -5.099825e-09, -6.018633e-09, 
    -7.21235e-09, -8.264974e-09, -9.262942e-09, -1.06882e-08, -1.221691e-08, 
    -1.392878e-08, -1.52865e-08, -1.683849e-08, -1.922237e-08, -2.162035e-08,
  -1.768873e-09, -2.341455e-09, -3.022974e-09, -3.836429e-09, -4.496309e-09, 
    -5.36976e-09, -6.654212e-09, -7.791713e-09, -8.617853e-09, -9.621352e-09, 
    -1.120075e-08, -1.325552e-08, -1.510643e-08, -1.717796e-08, -1.9064e-08,
  -1.487506e-08, -1.490308e-08, -1.513801e-08, -1.534315e-08, -1.578196e-08, 
    -1.660166e-08, -1.701224e-08, -1.732825e-08, -1.768682e-08, 
    -1.792766e-08, -1.846576e-08, -1.89644e-08, -1.834866e-08, -1.65659e-08, 
    -1.436015e-08,
  -1.465655e-08, -1.443487e-08, -1.42916e-08, -1.439997e-08, -1.470988e-08, 
    -1.511755e-08, -1.594207e-08, -1.684604e-08, -1.756769e-08, 
    -1.813782e-08, -1.839168e-08, -1.871173e-08, -1.921398e-08, 
    -1.912416e-08, -1.749021e-08,
  -1.403354e-08, -1.386372e-08, -1.37208e-08, -1.364454e-08, -1.364509e-08, 
    -1.412313e-08, -1.464875e-08, -1.527187e-08, -1.609276e-08, -1.70418e-08, 
    -1.790785e-08, -1.874487e-08, -1.942772e-08, -2.011644e-08, -1.980663e-08,
  -1.318113e-08, -1.32546e-08, -1.315499e-08, -1.316078e-08, -1.316224e-08, 
    -1.328518e-08, -1.371139e-08, -1.439572e-08, -1.506693e-08, 
    -1.580429e-08, -1.634898e-08, -1.718693e-08, -1.84471e-08, -1.975547e-08, 
    -2.103903e-08,
  -1.222048e-08, -1.21418e-08, -1.214929e-08, -1.222771e-08, -1.242419e-08, 
    -1.263349e-08, -1.28302e-08, -1.318577e-08, -1.387166e-08, -1.456941e-08, 
    -1.566844e-08, -1.618765e-08, -1.671087e-08, -1.820556e-08, -2.020985e-08,
  -1.103155e-08, -1.13408e-08, -1.156006e-08, -1.15658e-08, -1.174225e-08, 
    -1.204679e-08, -1.237694e-08, -1.245966e-08, -1.285822e-08, 
    -1.348303e-08, -1.40744e-08, -1.504324e-08, -1.591475e-08, -1.650255e-08, 
    -1.813773e-08,
  -9.539274e-09, -9.921266e-09, -1.029225e-08, -1.079123e-08, -1.109971e-08, 
    -1.143034e-08, -1.154738e-08, -1.181605e-08, -1.191101e-08, 
    -1.241492e-08, -1.317228e-08, -1.376607e-08, -1.456028e-08, -1.56473e-08, 
    -1.65099e-08,
  -8.289242e-09, -8.58592e-09, -8.881086e-09, -9.129399e-09, -9.662172e-09, 
    -1.012877e-08, -1.077344e-08, -1.107604e-08, -1.131315e-08, 
    -1.152595e-08, -1.206402e-08, -1.286254e-08, -1.347712e-08, 
    -1.412846e-08, -1.541368e-08,
  -7.134739e-09, -7.426243e-09, -7.751455e-09, -8.015148e-09, -8.102972e-09, 
    -8.546316e-09, -8.976217e-09, -9.761223e-09, -1.035905e-08, 
    -1.088439e-08, -1.144738e-08, -1.191913e-08, -1.264333e-08, 
    -1.311106e-08, -1.387552e-08,
  -6.049075e-09, -6.291716e-09, -6.640986e-09, -7.075494e-09, -7.323219e-09, 
    -7.390796e-09, -7.641495e-09, -7.969616e-09, -8.79064e-09, -9.610686e-09, 
    -1.049079e-08, -1.128595e-08, -1.177801e-08, -1.237339e-08, -1.268864e-08,
  -9.581353e-09, -1.024691e-08, -1.092203e-08, -1.142243e-08, -1.189372e-08, 
    -1.246531e-08, -1.290789e-08, -1.329036e-08, -1.374313e-08, 
    -1.437005e-08, -1.515357e-08, -1.621392e-08, -1.674702e-08, 
    -1.622149e-08, -1.579161e-08,
  -1.008952e-08, -1.073623e-08, -1.135823e-08, -1.206507e-08, -1.252723e-08, 
    -1.292983e-08, -1.335172e-08, -1.372633e-08, -1.428084e-08, 
    -1.463709e-08, -1.532098e-08, -1.587096e-08, -1.664621e-08, -1.67415e-08, 
    -1.629328e-08,
  -1.03847e-08, -1.095642e-08, -1.140876e-08, -1.194203e-08, -1.251785e-08, 
    -1.293884e-08, -1.340811e-08, -1.370382e-08, -1.426957e-08, 
    -1.470334e-08, -1.536471e-08, -1.579019e-08, -1.67061e-08, -1.718296e-08, 
    -1.713951e-08,
  -1.020148e-08, -1.082621e-08, -1.140783e-08, -1.190636e-08, -1.229219e-08, 
    -1.285755e-08, -1.328514e-08, -1.365478e-08, -1.404899e-08, -1.46717e-08, 
    -1.533259e-08, -1.580044e-08, -1.647547e-08, -1.6688e-08, -1.715916e-08,
  -9.604455e-09, -1.022235e-08, -1.077544e-08, -1.131983e-08, -1.174279e-08, 
    -1.217173e-08, -1.264225e-08, -1.306989e-08, -1.345992e-08, 
    -1.381346e-08, -1.45642e-08, -1.546365e-08, -1.587545e-08, -1.617047e-08, 
    -1.560213e-08,
  -8.776695e-09, -9.292162e-09, -9.822855e-09, -1.038008e-08, -1.082545e-08, 
    -1.117662e-08, -1.15223e-08, -1.186239e-08, -1.232829e-08, -1.253119e-08, 
    -1.315337e-08, -1.425619e-08, -1.484248e-08, -1.557019e-08, -1.517064e-08,
  -8.240079e-09, -8.579674e-09, -8.932941e-09, -9.341006e-09, -9.727639e-09, 
    -1.005095e-08, -1.030759e-08, -1.047009e-08, -1.080134e-08, 
    -1.123048e-08, -1.150799e-08, -1.244742e-08, -1.344731e-08, 
    -1.395901e-08, -1.471223e-08,
  -7.648374e-09, -8.054627e-09, -8.357116e-09, -8.660285e-09, -8.952533e-09, 
    -9.164304e-09, -9.319415e-09, -9.396461e-09, -9.455198e-09, 
    -9.721025e-09, -1.001823e-08, -1.050105e-08, -1.164464e-08, -1.2358e-08, 
    -1.313684e-08,
  -6.999252e-09, -7.401131e-09, -7.798499e-09, -8.081663e-09, -8.31212e-09, 
    -8.528726e-09, -8.609478e-09, -8.68336e-09, -8.686746e-09, -8.645505e-09, 
    -8.787028e-09, -8.953015e-09, -9.589041e-09, -1.047693e-08, -1.117752e-08,
  -6.500811e-09, -6.764219e-09, -7.053077e-09, -7.392232e-09, -7.662231e-09, 
    -7.846139e-09, -8.03432e-09, -8.075825e-09, -8.174104e-09, -8.13656e-09, 
    -8.133198e-09, -8.258609e-09, -8.413267e-09, -8.947973e-09, -9.70947e-09,
  -1.496255e-08, -1.598385e-08, -1.680592e-08, -1.680351e-08, -1.654914e-08, 
    -1.627513e-08, -1.6018e-08, -1.570068e-08, -1.53105e-08, -1.472435e-08, 
    -1.395614e-08, -1.300859e-08, -1.191651e-08, -1.090461e-08, -1.017701e-08,
  -1.264978e-08, -1.414515e-08, -1.50757e-08, -1.556832e-08, -1.559559e-08, 
    -1.53169e-08, -1.513729e-08, -1.48617e-08, -1.450406e-08, -1.391916e-08, 
    -1.316277e-08, -1.219999e-08, -1.128833e-08, -1.037872e-08, -9.844405e-09,
  -1.04284e-08, -1.191471e-08, -1.323695e-08, -1.402453e-08, -1.446575e-08, 
    -1.438993e-08, -1.426688e-08, -1.40623e-08, -1.376067e-08, -1.322244e-08, 
    -1.254802e-08, -1.162577e-08, -1.079338e-08, -1.001834e-08, -9.712977e-09,
  -8.475342e-09, -9.937764e-09, -1.12131e-08, -1.238431e-08, -1.300933e-08, 
    -1.322761e-08, -1.323784e-08, -1.312335e-08, -1.292436e-08, 
    -1.248129e-08, -1.18513e-08, -1.095135e-08, -1.016614e-08, -9.602527e-09, 
    -9.474135e-09,
  -7.260557e-09, -8.17685e-09, -9.331434e-09, -1.040713e-08, -1.1405e-08, 
    -1.185156e-08, -1.205888e-08, -1.207344e-08, -1.195469e-08, 
    -1.162484e-08, -1.106843e-08, -1.028627e-08, -9.591377e-09, 
    -9.210239e-09, -9.354565e-09,
  -6.861954e-09, -7.235139e-09, -7.906457e-09, -8.705128e-09, -9.503291e-09, 
    -1.02406e-08, -1.061304e-08, -1.079269e-08, -1.082925e-08, -1.070747e-08, 
    -1.030966e-08, -9.687192e-09, -9.038327e-09, -8.864981e-09, -9.075824e-09,
  -6.666439e-09, -6.929035e-09, -7.218508e-09, -7.691987e-09, -8.201386e-09, 
    -8.743467e-09, -9.211218e-09, -9.481357e-09, -9.624245e-09, 
    -9.654431e-09, -9.48968e-09, -9.08882e-09, -8.628421e-09, -8.523578e-09, 
    -8.72634e-09,
  -6.584357e-09, -6.722144e-09, -6.885661e-09, -7.121941e-09, -7.444914e-09, 
    -7.795856e-09, -8.16099e-09, -8.499969e-09, -8.734409e-09, -8.880163e-09, 
    -8.92198e-09, -8.713989e-09, -8.428728e-09, -8.346202e-09, -8.465266e-09,
  -6.660759e-09, -6.709055e-09, -6.769878e-09, -6.849789e-09, -6.991596e-09, 
    -7.202738e-09, -7.444541e-09, -7.71009e-09, -7.985571e-09, -8.230752e-09, 
    -8.469894e-09, -8.497512e-09, -8.367581e-09, -8.259887e-09, -8.291259e-09,
  -6.743326e-09, -6.803491e-09, -6.827829e-09, -6.873656e-09, -6.912395e-09, 
    -6.992814e-09, -7.109072e-09, -7.259283e-09, -7.466085e-09, 
    -7.661419e-09, -7.953847e-09, -8.193133e-09, -8.273363e-09, 
    -8.254184e-09, -8.215681e-09,
  -1.639427e-08, -1.923804e-08, -2.187613e-08, -2.385473e-08, -2.526608e-08, 
    -2.735367e-08, -2.85162e-08, -2.861147e-08, -2.884117e-08, -2.827968e-08, 
    -2.768919e-08, -2.754976e-08, -2.676746e-08, -2.61718e-08, -2.566923e-08,
  -1.564828e-08, -1.859598e-08, -2.154848e-08, -2.411556e-08, -2.549962e-08, 
    -2.697688e-08, -2.819425e-08, -2.845937e-08, -2.838607e-08, -2.80617e-08, 
    -2.801791e-08, -2.806256e-08, -2.704435e-08, -2.629016e-08, -2.582144e-08,
  -1.415214e-08, -1.73682e-08, -2.028611e-08, -2.343584e-08, -2.562772e-08, 
    -2.695156e-08, -2.782946e-08, -2.803307e-08, -2.814801e-08, 
    -2.773791e-08, -2.791639e-08, -2.819069e-08, -2.734023e-08, 
    -2.634935e-08, -2.559009e-08,
  -1.237035e-08, -1.583691e-08, -1.884889e-08, -2.209666e-08, -2.494616e-08, 
    -2.7072e-08, -2.778229e-08, -2.781487e-08, -2.758221e-08, -2.71786e-08, 
    -2.73851e-08, -2.772058e-08, -2.721584e-08, -2.612258e-08, -2.517636e-08,
  -1.048001e-08, -1.377558e-08, -1.704645e-08, -2.032475e-08, -2.353042e-08, 
    -2.632444e-08, -2.749698e-08, -2.748248e-08, -2.759541e-08, 
    -2.689139e-08, -2.66923e-08, -2.688042e-08, -2.654924e-08, -2.569064e-08, 
    -2.48933e-08,
  -8.657557e-09, -1.15285e-08, -1.461858e-08, -1.803177e-08, -2.135845e-08, 
    -2.487559e-08, -2.662098e-08, -2.692657e-08, -2.714027e-08, 
    -2.687984e-08, -2.632474e-08, -2.61944e-08, -2.585899e-08, -2.52372e-08, 
    -2.447962e-08,
  -7.12243e-09, -9.425062e-09, -1.210869e-08, -1.527136e-08, -1.826084e-08, 
    -2.197853e-08, -2.470279e-08, -2.561755e-08, -2.611116e-08, 
    -2.615939e-08, -2.589991e-08, -2.558848e-08, -2.516145e-08, 
    -2.451071e-08, -2.359251e-08,
  -5.955086e-09, -7.650199e-09, -9.837787e-09, -1.267923e-08, -1.519609e-08, 
    -1.837981e-08, -2.163944e-08, -2.324238e-08, -2.409276e-08, 
    -2.448595e-08, -2.443965e-08, -2.417318e-08, -2.372543e-08, 
    -2.300447e-08, -2.198713e-08,
  -5.06684e-09, -6.185924e-09, -7.847447e-09, -1.024607e-08, -1.254357e-08, 
    -1.481723e-08, -1.77988e-08, -2.004063e-08, -2.126948e-08, -2.189403e-08, 
    -2.217559e-08, -2.198464e-08, -2.163171e-08, -2.085841e-08, -1.983098e-08,
  -4.612084e-09, -5.214476e-09, -6.204123e-09, -8.002952e-09, -1.010513e-08, 
    -1.197147e-08, -1.400932e-08, -1.625452e-08, -1.785915e-08, 
    -1.875832e-08, -1.919514e-08, -1.920176e-08, -1.892895e-08, -1.8241e-08, 
    -1.725286e-08,
  -5.5011e-09, -6.333327e-09, -7.278061e-09, -8.433704e-09, -9.826241e-09, 
    -1.151381e-08, -1.345379e-08, -1.571185e-08, -1.778817e-08, 
    -1.955197e-08, -2.097227e-08, -2.239954e-08, -2.355284e-08, 
    -2.465551e-08, -2.574899e-08,
  -4.350063e-09, -5.23727e-09, -6.250188e-09, -7.505109e-09, -8.935866e-09, 
    -1.070036e-08, -1.282618e-08, -1.521068e-08, -1.743093e-08, 
    -1.922706e-08, -2.066429e-08, -2.218004e-08, -2.341994e-08, 
    -2.471353e-08, -2.5592e-08,
  -3.793401e-09, -4.34749e-09, -5.21907e-09, -6.526208e-09, -8.038948e-09, 
    -9.878291e-09, -1.209301e-08, -1.466997e-08, -1.699246e-08, 
    -1.882149e-08, -2.024667e-08, -2.184897e-08, -2.318603e-08, 
    -2.444137e-08, -2.514606e-08,
  -3.210396e-09, -3.615493e-09, -4.32981e-09, -5.514029e-09, -7.120884e-09, 
    -9.047655e-09, -1.136144e-08, -1.400156e-08, -1.63786e-08, -1.839855e-08, 
    -1.984021e-08, -2.150634e-08, -2.293163e-08, -2.410727e-08, -2.484049e-08,
  -2.933016e-09, -3.148887e-09, -3.621903e-09, -4.635381e-09, -6.144627e-09, 
    -8.133918e-09, -1.055798e-08, -1.33435e-08, -1.576261e-08, -1.791003e-08, 
    -1.944424e-08, -2.118964e-08, -2.272017e-08, -2.390594e-08, -2.465029e-08,
  -2.751598e-09, -2.921458e-09, -3.185701e-09, -3.936311e-09, -5.273944e-09, 
    -7.144459e-09, -9.662062e-09, -1.254641e-08, -1.50323e-08, -1.739335e-08, 
    -1.893517e-08, -2.062928e-08, -2.226811e-08, -2.357838e-08, -2.448414e-08,
  -2.628733e-09, -2.794293e-09, -2.989882e-09, -3.482346e-09, -4.55473e-09, 
    -6.200187e-09, -8.665336e-09, -1.161279e-08, -1.427936e-08, -1.6736e-08, 
    -1.836954e-08, -1.997052e-08, -2.15784e-08, -2.309879e-08, -2.42805e-08,
  -2.52301e-09, -2.68306e-09, -2.881688e-09, -3.239552e-09, -4.033319e-09, 
    -5.399141e-09, -7.708844e-09, -1.050305e-08, -1.327933e-08, 
    -1.594825e-08, -1.794559e-08, -1.942557e-08, -2.092328e-08, 
    -2.238095e-08, -2.376977e-08,
  -2.45337e-09, -2.581771e-09, -2.786725e-09, -3.056796e-09, -3.657099e-09, 
    -4.710775e-09, -6.718562e-09, -9.421052e-09, -1.214866e-08, 
    -1.479922e-08, -1.72087e-08, -1.895587e-08, -2.037047e-08, -2.174217e-08, 
    -2.296207e-08,
  -2.38354e-09, -2.49116e-09, -2.697343e-09, -2.917325e-09, -3.364686e-09, 
    -4.129672e-09, -5.680738e-09, -8.19711e-09, -1.094203e-08, -1.363741e-08, 
    -1.611019e-08, -1.823132e-08, -1.98578e-08, -2.13301e-08, -2.258492e-08,
  -1.056904e-08, -1.122497e-08, -1.205e-08, -1.30629e-08, -1.434279e-08, 
    -1.632185e-08, -1.799989e-08, -1.911758e-08, -1.9695e-08, -1.989692e-08, 
    -2.002046e-08, -2.051629e-08, -2.109188e-08, -2.17417e-08, -2.213086e-08,
  -9.963569e-09, -1.018241e-08, -1.073895e-08, -1.167896e-08, -1.272641e-08, 
    -1.397791e-08, -1.572441e-08, -1.712674e-08, -1.840024e-08, 
    -1.905769e-08, -1.938214e-08, -1.951054e-08, -2.024747e-08, 
    -2.096279e-08, -2.150441e-08,
  -9.932034e-09, -9.804928e-09, -9.863436e-09, -1.028093e-08, -1.112844e-08, 
    -1.216166e-08, -1.343379e-08, -1.507803e-08, -1.64029e-08, -1.74431e-08, 
    -1.815998e-08, -1.86307e-08, -1.899127e-08, -1.993235e-08, -2.058521e-08,
  -1.018631e-08, -9.859021e-09, -9.583813e-09, -9.567303e-09, -9.826867e-09, 
    -1.053541e-08, -1.147934e-08, -1.268038e-08, -1.431829e-08, 
    -1.554372e-08, -1.643567e-08, -1.71192e-08, -1.766518e-08, -1.824627e-08, 
    -1.923775e-08,
  -1.022927e-08, -1.003426e-08, -9.729557e-09, -9.413779e-09, -9.319806e-09, 
    -9.484919e-09, -9.988977e-09, -1.082511e-08, -1.192511e-08, 
    -1.340834e-08, -1.45136e-08, -1.540134e-08, -1.612866e-08, -1.67507e-08, 
    -1.75219e-08,
  -8.822128e-09, -9.703812e-09, -9.938194e-09, -9.522783e-09, -9.149815e-09, 
    -8.977256e-09, -9.149073e-09, -9.515638e-09, -1.019721e-08, 
    -1.123267e-08, -1.241995e-08, -1.340348e-08, -1.427611e-08, 
    -1.505395e-08, -1.586817e-08,
  -6.728558e-09, -8.017651e-09, -9.156865e-09, -9.768277e-09, -9.485239e-09, 
    -8.904509e-09, -8.699543e-09, -8.87144e-09, -9.237032e-09, -9.759773e-09, 
    -1.066461e-08, -1.163748e-08, -1.248502e-08, -1.320622e-08, -1.40439e-08,
  -4.579284e-09, -5.876659e-09, -7.033e-09, -8.254319e-09, -9.197692e-09, 
    -9.374248e-09, -8.854967e-09, -8.470567e-09, -8.613896e-09, 
    -8.939529e-09, -9.387448e-09, -1.005295e-08, -1.101942e-08, 
    -1.167886e-08, -1.23732e-08,
  -2.676277e-09, -3.90747e-09, -5.092118e-09, -6.128888e-09, -7.22906e-09, 
    -8.301174e-09, -8.978714e-09, -8.88133e-09, -8.483476e-09, -8.439595e-09, 
    -8.730844e-09, -9.114959e-09, -9.689365e-09, -1.038331e-08, -1.105699e-08,
  -1.404135e-09, -2.093848e-09, -3.149454e-09, -4.234094e-09, -5.283316e-09, 
    -6.195301e-09, -7.211375e-09, -8.128939e-09, -8.540761e-09, -8.42954e-09, 
    -8.289172e-09, -8.447573e-09, -8.866835e-09, -9.391705e-09, -9.933968e-09,
  -5.134952e-09, -5.58327e-09, -5.872431e-09, -6.097773e-09, -6.290411e-09, 
    -6.573849e-09, -7.026738e-09, -7.628993e-09, -8.389053e-09, 
    -9.331901e-09, -1.034271e-08, -1.134488e-08, -1.224641e-08, 
    -1.318674e-08, -1.408324e-08,
  -4.008272e-09, -4.643712e-09, -5.125039e-09, -5.41577e-09, -5.634147e-09, 
    -5.873637e-09, -6.222071e-09, -6.727634e-09, -7.405808e-09, 
    -8.341721e-09, -9.381242e-09, -1.045085e-08, -1.144159e-08, 
    -1.242003e-08, -1.339774e-08,
  -3.266224e-09, -3.882513e-09, -4.480526e-09, -4.897618e-09, -5.158836e-09, 
    -5.375536e-09, -5.61778e-09, -5.968518e-09, -6.566195e-09, -7.441724e-09, 
    -8.476158e-09, -9.578806e-09, -1.06285e-08, -1.164286e-08, -1.270925e-08,
  -2.579021e-09, -3.19138e-09, -3.850926e-09, -4.469558e-09, -4.800512e-09, 
    -5.007811e-09, -5.233313e-09, -5.466203e-09, -5.828677e-09, 
    -6.613414e-09, -7.667746e-09, -8.764281e-09, -9.900987e-09, 
    -1.095825e-08, -1.202798e-08,
  -2.18646e-09, -2.652324e-09, -3.256609e-09, -3.971823e-09, -4.615134e-09, 
    -4.860415e-09, -5.019043e-09, -5.21498e-09, -5.436213e-09, -5.859833e-09, 
    -6.833281e-09, -7.997882e-09, -9.188619e-09, -1.034785e-08, -1.141544e-08,
  -1.848365e-09, -2.233896e-09, -2.704934e-09, -3.326959e-09, -4.100234e-09, 
    -4.788253e-09, -5.024998e-09, -5.122136e-09, -5.270303e-09, 
    -5.464544e-09, -5.99358e-09, -7.075855e-09, -8.255891e-09, -9.602099e-09, 
    -1.079721e-08,
  -1.471435e-09, -1.87691e-09, -2.323036e-09, -2.803156e-09, -3.461602e-09, 
    -4.262047e-09, -4.999812e-09, -5.267911e-09, -5.327121e-09, 
    -5.404416e-09, -5.549607e-09, -6.09916e-09, -7.225755e-09, -8.444722e-09, 
    -9.834222e-09,
  -1.134072e-09, -1.440325e-09, -1.883913e-09, -2.392366e-09, -2.919034e-09, 
    -3.638212e-09, -4.480151e-09, -5.223498e-09, -5.510825e-09, 
    -5.568793e-09, -5.587103e-09, -5.649193e-09, -6.141465e-09, 
    -7.205658e-09, -8.517901e-09,
  -9.817797e-10, -1.135264e-09, -1.447839e-09, -1.906074e-09, -2.465939e-09, 
    -3.075547e-09, -3.858115e-09, -4.765775e-09, -5.527981e-09, 
    -5.793845e-09, -5.789576e-09, -5.779443e-09, -5.750505e-09, 
    -6.115553e-09, -7.055389e-09,
  -8.921215e-10, -9.644642e-10, -1.138988e-09, -1.470083e-09, -1.933259e-09, 
    -2.544049e-09, -3.225402e-09, -4.065851e-09, -5.062113e-09, 
    -5.877612e-09, -6.206461e-09, -6.010323e-09, -5.977003e-09, 
    -5.910172e-09, -6.157125e-09,
  -9.977844e-09, -1.031859e-08, -1.073611e-08, -1.130942e-08, -1.184587e-08, 
    -1.227881e-08, -1.256634e-08, -1.284527e-08, -1.313137e-08, 
    -1.362043e-08, -1.443381e-08, -1.538204e-08, -1.61922e-08, -1.665142e-08, 
    -1.68885e-08,
  -9.679636e-09, -1.000963e-08, -1.039311e-08, -1.096416e-08, -1.152843e-08, 
    -1.199502e-08, -1.232154e-08, -1.25876e-08, -1.292031e-08, -1.353202e-08, 
    -1.414462e-08, -1.470719e-08, -1.50452e-08, -1.541431e-08, -1.55501e-08,
  -9.018416e-09, -9.437989e-09, -9.879948e-09, -1.042423e-08, -1.098721e-08, 
    -1.14692e-08, -1.186514e-08, -1.227602e-08, -1.266285e-08, -1.300499e-08, 
    -1.320263e-08, -1.322036e-08, -1.328852e-08, -1.345383e-08, -1.38434e-08,
  -8.194611e-09, -8.614557e-09, -8.973981e-09, -9.511566e-09, -1.009071e-08, 
    -1.061377e-08, -1.11191e-08, -1.171521e-08, -1.209193e-08, -1.217492e-08, 
    -1.19256e-08, -1.184028e-08, -1.207488e-08, -1.274842e-08, -1.342772e-08,
  -7.217549e-09, -7.848611e-09, -8.24898e-09, -8.518669e-09, -9.041362e-09, 
    -9.694624e-09, -1.034391e-08, -1.093083e-08, -1.132439e-08, 
    -1.153975e-08, -1.167852e-08, -1.174123e-08, -1.184787e-08, 
    -1.232523e-08, -1.280555e-08,
  -6.355049e-09, -6.78106e-09, -7.338204e-09, -7.758802e-09, -8.11728e-09, 
    -8.637439e-09, -9.39435e-09, -1.021888e-08, -1.078604e-08, -1.117778e-08, 
    -1.157243e-08, -1.190148e-08, -1.237557e-08, -1.309247e-08, -1.388995e-08,
  -5.67272e-09, -5.945627e-09, -6.348674e-09, -6.827836e-09, -7.324215e-09, 
    -7.802232e-09, -8.251162e-09, -8.815173e-09, -9.408683e-09, 
    -9.961665e-09, -1.056697e-08, -1.129844e-08, -1.206186e-08, 
    -1.291017e-08, -1.376745e-08,
  -4.828399e-09, -5.381511e-09, -5.602005e-09, -5.890864e-09, -6.296281e-09, 
    -6.75812e-09, -7.238407e-09, -7.662893e-09, -8.153337e-09, -8.614298e-09, 
    -9.079734e-09, -9.667334e-09, -1.044245e-08, -1.118462e-08, -1.212624e-08,
  -3.436605e-09, -4.323732e-09, -5.075921e-09, -5.350967e-09, -5.486625e-09, 
    -5.780513e-09, -6.078688e-09, -6.431934e-09, -6.830441e-09, 
    -7.458261e-09, -8.181738e-09, -8.620016e-09, -9.253378e-09, 
    -9.859587e-09, -1.038717e-08,
  -1.964649e-09, -2.974383e-09, -3.844504e-09, -4.699725e-09, -5.117258e-09, 
    -5.096535e-09, -5.212517e-09, -5.371582e-09, -5.625004e-09, 
    -6.083235e-09, -6.883593e-09, -7.699162e-09, -8.339401e-09, 
    -8.907446e-09, -9.314291e-09,
  -8.515962e-09, -9.191466e-09, -1.027765e-08, -1.179779e-08, -1.296419e-08, 
    -1.371947e-08, -1.397064e-08, -1.389692e-08, -1.384101e-08, 
    -1.365634e-08, -1.350855e-08, -1.32948e-08, -1.301157e-08, -1.268022e-08, 
    -1.235361e-08,
  -7.573129e-09, -8.126959e-09, -8.75534e-09, -9.668391e-09, -1.08018e-08, 
    -1.158759e-08, -1.219414e-08, -1.250815e-08, -1.269564e-08, 
    -1.273686e-08, -1.266692e-08, -1.247097e-08, -1.216241e-08, 
    -1.184345e-08, -1.149934e-08,
  -6.777895e-09, -7.145097e-09, -7.614394e-09, -8.160258e-09, -9.011127e-09, 
    -9.919258e-09, -1.059421e-08, -1.11944e-08, -1.15751e-08, -1.172203e-08, 
    -1.170905e-08, -1.147353e-08, -1.121443e-08, -1.085446e-08, -1.056548e-08,
  -5.950386e-09, -6.246991e-09, -6.576014e-09, -7.02435e-09, -7.561884e-09, 
    -8.380449e-09, -9.264122e-09, -1.007209e-08, -1.063831e-08, 
    -1.085982e-08, -1.077475e-08, -1.056297e-08, -1.025384e-08, 
    -9.976297e-09, -9.657452e-09,
  -5.16883e-09, -5.476379e-09, -5.715914e-09, -6.061731e-09, -6.488836e-09, 
    -7.093965e-09, -7.867158e-09, -8.795533e-09, -9.560319e-09, 
    -9.990463e-09, -1.000739e-08, -9.817985e-09, -9.504377e-09, 
    -9.258747e-09, -8.970121e-09,
  -4.216834e-09, -4.569399e-09, -4.903481e-09, -5.283526e-09, -5.685986e-09, 
    -6.177903e-09, -6.784662e-09, -7.518675e-09, -8.362808e-09, 
    -8.919327e-09, -9.195195e-09, -9.185118e-09, -9.044423e-09, 
    -8.842895e-09, -8.561512e-09,
  -3.312384e-09, -3.673324e-09, -4.032168e-09, -4.462957e-09, -4.912199e-09, 
    -5.392954e-09, -5.939084e-09, -6.55516e-09, -7.222857e-09, -7.87371e-09, 
    -8.228199e-09, -8.413697e-09, -8.403537e-09, -8.328129e-09, -8.119285e-09,
  -2.617202e-09, -2.88998e-09, -3.229456e-09, -3.649522e-09, -4.057982e-09, 
    -4.508394e-09, -5.050487e-09, -5.68609e-09, -6.314687e-09, -6.908373e-09, 
    -7.337663e-09, -7.592105e-09, -7.69966e-09, -7.680823e-09, -7.56212e-09,
  -2.089572e-09, -2.294243e-09, -2.555447e-09, -2.902525e-09, -3.272891e-09, 
    -3.697419e-09, -4.216396e-09, -4.839158e-09, -5.482522e-09, 
    -6.018746e-09, -6.487e-09, -6.779972e-09, -7.005364e-09, -7.10976e-09, 
    -7.133023e-09,
  -1.709259e-09, -1.833018e-09, -2.027569e-09, -2.276645e-09, -2.57497e-09, 
    -2.916414e-09, -3.398998e-09, -3.99273e-09, -4.63878e-09, -5.135711e-09, 
    -5.544371e-09, -5.938881e-09, -6.245567e-09, -6.447303e-09, -6.656089e-09,
  -8.633041e-09, -8.714268e-09, -8.938255e-09, -9.418518e-09, -1.003335e-08, 
    -1.049139e-08, -1.120988e-08, -1.194561e-08, -1.32559e-08, -1.486536e-08, 
    -1.636214e-08, -1.790571e-08, -1.936334e-08, -2.100698e-08, -2.235097e-08,
  -8.717068e-09, -8.710941e-09, -8.690957e-09, -8.977982e-09, -9.513986e-09, 
    -1.006562e-08, -1.050822e-08, -1.10463e-08, -1.179208e-08, -1.294076e-08, 
    -1.441525e-08, -1.590637e-08, -1.767656e-08, -1.941346e-08, -2.103453e-08,
  -8.691356e-09, -8.774093e-09, -8.738831e-09, -8.683644e-09, -8.987448e-09, 
    -9.502228e-09, -1.006013e-08, -1.03631e-08, -1.088085e-08, -1.155791e-08, 
    -1.268716e-08, -1.416177e-08, -1.579488e-08, -1.773023e-08, -1.965224e-08,
  -8.189705e-09, -8.661247e-09, -8.818686e-09, -8.822466e-09, -8.761553e-09, 
    -9.002446e-09, -9.464978e-09, -9.96489e-09, -1.028195e-08, -1.070585e-08, 
    -1.128578e-08, -1.236547e-08, -1.389662e-08, -1.567744e-08, -1.755156e-08,
  -7.779219e-09, -8.148832e-09, -8.584427e-09, -8.842592e-09, -8.886722e-09, 
    -8.805198e-09, -8.98754e-09, -9.41349e-09, -9.825709e-09, -1.011177e-08, 
    -1.029742e-08, -1.082993e-08, -1.174789e-08, -1.316887e-08, -1.499664e-08,
  -7.519001e-09, -7.807168e-09, -8.18634e-09, -8.644102e-09, -9.001136e-09, 
    -9.030221e-09, -8.896415e-09, -9.007767e-09, -9.39431e-09, -9.79109e-09, 
    -9.927975e-09, -9.92625e-09, -1.030668e-08, -1.090998e-08, -1.221571e-08,
  -7.149051e-09, -7.511441e-09, -7.824276e-09, -8.264666e-09, -8.769183e-09, 
    -9.10534e-09, -9.161968e-09, -9.018355e-09, -9.045611e-09, -9.332796e-09, 
    -9.675206e-09, -9.798951e-09, -9.756976e-09, -9.913512e-09, -1.025044e-08,
  -6.739285e-09, -7.147178e-09, -7.477529e-09, -7.863015e-09, -8.381362e-09, 
    -8.837715e-09, -9.109074e-09, -9.204029e-09, -9.14e-09, -9.102594e-09, 
    -9.298613e-09, -9.633892e-09, -9.780052e-09, -9.933999e-09, -1.000471e-08,
  -6.230709e-09, -6.718201e-09, -7.09072e-09, -7.406001e-09, -7.889707e-09, 
    -8.44128e-09, -8.848988e-09, -9.083164e-09, -9.202563e-09, -9.173613e-09, 
    -9.159666e-09, -9.377238e-09, -9.697271e-09, -9.906989e-09, -1.004056e-08,
  -5.446759e-09, -6.117213e-09, -6.609759e-09, -7.020367e-09, -7.382812e-09, 
    -7.897173e-09, -8.47386e-09, -8.882228e-09, -9.102202e-09, -9.132433e-09, 
    -9.111739e-09, -9.183787e-09, -9.430163e-09, -9.720357e-09, -9.907818e-09,
  -8.257719e-09, -8.483844e-09, -8.785412e-09, -8.961196e-09, -9.098664e-09, 
    -9.259328e-09, -9.471688e-09, -9.691663e-09, -9.889497e-09, -1.00861e-08, 
    -1.023926e-08, -1.033835e-08, -1.037805e-08, -1.038772e-08, -1.038393e-08,
  -7.0924e-09, -7.329171e-09, -7.706995e-09, -8.024416e-09, -8.30023e-09, 
    -8.555885e-09, -8.767585e-09, -9.012352e-09, -9.314051e-09, 
    -9.588498e-09, -9.96282e-09, -1.026227e-08, -1.043852e-08, -1.050168e-08, 
    -1.047619e-08,
  -6.459736e-09, -6.602298e-09, -6.866224e-09, -7.193329e-09, -7.505933e-09, 
    -7.852555e-09, -8.180999e-09, -8.52881e-09, -8.926961e-09, -9.362156e-09, 
    -9.864023e-09, -1.029431e-08, -1.058516e-08, -1.059986e-08, -1.04727e-08,
  -6.390066e-09, -6.423824e-09, -6.592721e-09, -6.807319e-09, -7.078301e-09, 
    -7.453646e-09, -7.905935e-09, -8.281772e-09, -8.644187e-09, 
    -9.145858e-09, -9.705844e-09, -1.022328e-08, -1.057463e-08, 
    -1.055918e-08, -1.03869e-08,
  -6.429715e-09, -6.492177e-09, -6.486876e-09, -6.614832e-09, -6.845435e-09, 
    -7.220975e-09, -7.659396e-09, -8.136166e-09, -8.574022e-09, 
    -9.029391e-09, -9.439137e-09, -9.933969e-09, -1.016617e-08, 
    -1.026744e-08, -1.025639e-08,
  -6.056822e-09, -6.248888e-09, -6.333952e-09, -6.48678e-09, -6.63636e-09, 
    -6.915883e-09, -7.321413e-09, -7.78529e-09, -8.332375e-09, -8.825982e-09, 
    -9.225845e-09, -9.577742e-09, -9.698274e-09, -9.84049e-09, -9.956127e-09,
  -5.395974e-09, -5.964728e-09, -6.225144e-09, -6.384127e-09, -6.563802e-09, 
    -6.783409e-09, -7.087333e-09, -7.480944e-09, -7.983721e-09, 
    -8.536911e-09, -9.005369e-09, -9.195288e-09, -9.33424e-09, -9.527518e-09, 
    -9.727416e-09,
  -4.301836e-09, -5.001055e-09, -5.606869e-09, -6.08462e-09, -6.380838e-09, 
    -6.610477e-09, -6.927907e-09, -7.26263e-09, -7.668027e-09, -8.142853e-09, 
    -8.702195e-09, -8.917928e-09, -9.068341e-09, -9.316524e-09, -9.64707e-09,
  -3.601912e-09, -4.056939e-09, -4.642876e-09, -5.227494e-09, -5.7428e-09, 
    -6.205045e-09, -6.584828e-09, -6.973609e-09, -7.374027e-09, -7.81391e-09, 
    -8.349125e-09, -8.684001e-09, -8.883564e-09, -9.133428e-09, -9.47789e-09,
  -3.149973e-09, -3.507626e-09, -3.943593e-09, -4.490672e-09, -4.94847e-09, 
    -5.463104e-09, -5.993662e-09, -6.468347e-09, -6.991316e-09, 
    -7.495495e-09, -8.051302e-09, -8.400339e-09, -8.649188e-09, 
    -8.913137e-09, -9.266757e-09,
  -1.826834e-08, -1.824265e-08, -1.817717e-08, -1.833017e-08, -1.858844e-08, 
    -1.890999e-08, -1.919395e-08, -1.956234e-08, -1.99532e-08, -2.044207e-08, 
    -2.087423e-08, -2.105011e-08, -2.094136e-08, -2.050181e-08, -1.974246e-08,
  -1.733164e-08, -1.743867e-08, -1.744897e-08, -1.754079e-08, -1.761025e-08, 
    -1.766554e-08, -1.77198e-08, -1.775953e-08, -1.778579e-08, -1.787582e-08, 
    -1.789473e-08, -1.789131e-08, -1.795584e-08, -1.797084e-08, -1.772668e-08,
  -1.625267e-08, -1.643108e-08, -1.651537e-08, -1.656782e-08, -1.648067e-08, 
    -1.634836e-08, -1.620291e-08, -1.601209e-08, -1.569477e-08, 
    -1.530375e-08, -1.482185e-08, -1.444484e-08, -1.396443e-08, 
    -1.374564e-08, -1.373778e-08,
  -1.496611e-08, -1.51695e-08, -1.532022e-08, -1.535686e-08, -1.530482e-08, 
    -1.509595e-08, -1.490204e-08, -1.462288e-08, -1.441251e-08, 
    -1.408054e-08, -1.367306e-08, -1.334389e-08, -1.308725e-08, 
    -1.310998e-08, -1.32367e-08,
  -1.350393e-08, -1.382917e-08, -1.405488e-08, -1.421554e-08, -1.428183e-08, 
    -1.419922e-08, -1.408299e-08, -1.386164e-08, -1.374911e-08, 
    -1.349461e-08, -1.345724e-08, -1.329314e-08, -1.34959e-08, -1.373165e-08, 
    -1.401258e-08,
  -1.219783e-08, -1.249745e-08, -1.275901e-08, -1.299614e-08, -1.315635e-08, 
    -1.322515e-08, -1.316075e-08, -1.309721e-08, -1.304937e-08, 
    -1.298364e-08, -1.303285e-08, -1.310343e-08, -1.348894e-08, 
    -1.372305e-08, -1.393318e-08,
  -1.107333e-08, -1.128299e-08, -1.156522e-08, -1.177352e-08, -1.195481e-08, 
    -1.216628e-08, -1.220861e-08, -1.226447e-08, -1.22954e-08, -1.235068e-08, 
    -1.239706e-08, -1.256383e-08, -1.282481e-08, -1.299472e-08, -1.293916e-08,
  -1.003228e-08, -1.037884e-08, -1.063557e-08, -1.086588e-08, -1.1024e-08, 
    -1.116515e-08, -1.130292e-08, -1.144361e-08, -1.167031e-08, 
    -1.188481e-08, -1.200987e-08, -1.226418e-08, -1.24999e-08, -1.257395e-08, 
    -1.244591e-08,
  -8.862933e-09, -9.284761e-09, -9.612019e-09, -9.952067e-09, -1.019929e-08, 
    -1.030561e-08, -1.032834e-08, -1.038712e-08, -1.050575e-08, 
    -1.072759e-08, -1.089284e-08, -1.120536e-08, -1.141344e-08, 
    -1.149651e-08, -1.142327e-08,
  -7.501728e-09, -8.011228e-09, -8.320585e-09, -8.682854e-09, -9.078976e-09, 
    -9.390012e-09, -9.56504e-09, -9.654016e-09, -9.706485e-09, -9.76244e-09, 
    -9.870421e-09, -1.004874e-08, -1.016392e-08, -1.019488e-08, -1.021085e-08,
  -2.165169e-08, -2.191694e-08, -2.181333e-08, -2.145038e-08, -2.143498e-08, 
    -2.149227e-08, -2.145405e-08, -2.137315e-08, -2.143528e-08, 
    -2.150004e-08, -2.165062e-08, -2.181654e-08, -2.199751e-08, -2.22171e-08, 
    -2.243154e-08,
  -2.182756e-08, -2.178863e-08, -2.192472e-08, -2.186198e-08, -2.166482e-08, 
    -2.156271e-08, -2.169425e-08, -2.185548e-08, -2.196284e-08, 
    -2.209376e-08, -2.215166e-08, -2.227286e-08, -2.238886e-08, -2.25306e-08, 
    -2.260212e-08,
  -2.205343e-08, -2.185883e-08, -2.195491e-08, -2.212673e-08, -2.220232e-08, 
    -2.203356e-08, -2.199939e-08, -2.202746e-08, -2.212521e-08, -2.21381e-08, 
    -2.212747e-08, -2.210081e-08, -2.212922e-08, -2.216085e-08, -2.217126e-08,
  -2.222149e-08, -2.214225e-08, -2.201327e-08, -2.197622e-08, -2.194266e-08, 
    -2.19476e-08, -2.192965e-08, -2.198822e-08, -2.200183e-08, -2.198151e-08, 
    -2.196334e-08, -2.193165e-08, -2.189478e-08, -2.181399e-08, -2.172592e-08,
  -2.18301e-08, -2.219568e-08, -2.212827e-08, -2.204876e-08, -2.197376e-08, 
    -2.200032e-08, -2.182074e-08, -2.183601e-08, -2.17016e-08, -2.171379e-08, 
    -2.169696e-08, -2.166353e-08, -2.160415e-08, -2.147276e-08, -2.133975e-08,
  -2.049643e-08, -2.152744e-08, -2.170764e-08, -2.18128e-08, -2.174592e-08, 
    -2.193385e-08, -2.195604e-08, -2.180037e-08, -2.168333e-08, 
    -2.150956e-08, -2.145889e-08, -2.135785e-08, -2.120648e-08, 
    -2.108127e-08, -2.09152e-08,
  -1.79573e-08, -1.988363e-08, -2.102236e-08, -2.150424e-08, -2.152341e-08, 
    -2.168717e-08, -2.192562e-08, -2.186967e-08, -2.179861e-08, 
    -2.165171e-08, -2.143718e-08, -2.11679e-08, -2.093808e-08, -2.072185e-08, 
    -2.049285e-08,
  -1.399178e-08, -1.635391e-08, -1.826219e-08, -1.962581e-08, -2.051046e-08, 
    -2.097544e-08, -2.138223e-08, -2.160263e-08, -2.165946e-08, 
    -2.155548e-08, -2.1239e-08, -2.091811e-08, -2.076387e-08, -2.051059e-08, 
    -2.026891e-08,
  -1.203545e-08, -1.329847e-08, -1.498338e-08, -1.660585e-08, -1.805223e-08, 
    -1.898474e-08, -1.963405e-08, -2.011728e-08, -2.048379e-08, 
    -2.031054e-08, -1.993919e-08, -1.952663e-08, -1.936583e-08, 
    -1.938049e-08, -1.917046e-08,
  -1.032285e-08, -1.098725e-08, -1.220616e-08, -1.357275e-08, -1.515531e-08, 
    -1.638169e-08, -1.717421e-08, -1.795941e-08, -1.832954e-08, 
    -1.819783e-08, -1.791926e-08, -1.808243e-08, -1.827722e-08, -1.78428e-08, 
    -1.752788e-08,
  -2.133829e-08, -2.189781e-08, -2.23089e-08, -2.268246e-08, -2.269874e-08, 
    -2.27179e-08, -2.264664e-08, -2.242075e-08, -2.21095e-08, -2.174846e-08, 
    -2.155837e-08, -2.143632e-08, -2.124786e-08, -2.110421e-08, -2.104949e-08,
  -2.053592e-08, -2.098654e-08, -2.134108e-08, -2.184296e-08, -2.208628e-08, 
    -2.209757e-08, -2.202719e-08, -2.194136e-08, -2.185762e-08, 
    -2.180787e-08, -2.171004e-08, -2.141091e-08, -2.119143e-08, 
    -2.097105e-08, -2.089939e-08,
  -1.926845e-08, -1.994431e-08, -2.044181e-08, -2.103616e-08, -2.156082e-08, 
    -2.18653e-08, -2.177346e-08, -2.16649e-08, -2.15334e-08, -2.151152e-08, 
    -2.123582e-08, -2.089124e-08, -2.070266e-08, -2.067153e-08, -2.069305e-08,
  -1.770419e-08, -1.852202e-08, -1.922134e-08, -2.003325e-08, -2.078744e-08, 
    -2.143448e-08, -2.164231e-08, -2.145249e-08, -2.115649e-08, 
    -2.102473e-08, -2.070582e-08, -2.057683e-08, -2.059353e-08, -2.06853e-08, 
    -2.079554e-08,
  -1.600408e-08, -1.70939e-08, -1.801353e-08, -1.872904e-08, -1.94578e-08, 
    -2.01461e-08, -2.088525e-08, -2.107385e-08, -2.09937e-08, -2.06998e-08, 
    -2.059424e-08, -2.045815e-08, -2.035533e-08, -2.020264e-08, -2.034638e-08,
  -1.448867e-08, -1.544409e-08, -1.666482e-08, -1.777537e-08, -1.838376e-08, 
    -1.901024e-08, -1.96721e-08, -2.042631e-08, -2.082118e-08, -2.07696e-08, 
    -2.067013e-08, -2.043473e-08, -2.021958e-08, -2.000233e-08, -1.992834e-08,
  -1.414022e-08, -1.43226e-08, -1.517923e-08, -1.662644e-08, -1.783306e-08, 
    -1.819003e-08, -1.856764e-08, -1.938863e-08, -1.992828e-08, 
    -2.067502e-08, -2.025558e-08, -2.029868e-08, -1.994291e-08, 
    -1.986598e-08, -1.971496e-08,
  -1.419021e-08, -1.436662e-08, -1.439409e-08, -1.54116e-08, -1.66338e-08, 
    -1.770065e-08, -1.825295e-08, -1.898295e-08, -1.950124e-08, 
    -2.030979e-08, -2.033785e-08, -2.053718e-08, -2.021535e-08, 
    -1.992008e-08, -1.971618e-08,
  -1.358421e-08, -1.400063e-08, -1.426008e-08, -1.444319e-08, -1.524461e-08, 
    -1.628569e-08, -1.728123e-08, -1.805554e-08, -1.883774e-08, 
    -1.968686e-08, -2.002401e-08, -2.019434e-08, -1.999652e-08, 
    -2.000593e-08, -1.999164e-08,
  -1.222271e-08, -1.301641e-08, -1.365797e-08, -1.423938e-08, -1.468669e-08, 
    -1.561461e-08, -1.640911e-08, -1.707364e-08, -1.768978e-08, 
    -1.846022e-08, -1.894202e-08, -1.943188e-08, -2.049707e-08, 
    -2.125612e-08, -2.133572e-08,
  -1.709571e-08, -1.759479e-08, -1.809382e-08, -1.853335e-08, -1.859166e-08, 
    -1.851943e-08, -1.861725e-08, -1.885172e-08, -1.927817e-08, 
    -1.983009e-08, -2.021151e-08, -2.043762e-08, -2.061306e-08, 
    -2.071887e-08, -2.075718e-08,
  -1.671096e-08, -1.72382e-08, -1.778421e-08, -1.842543e-08, -1.908943e-08, 
    -1.951551e-08, -1.970339e-08, -1.958356e-08, -1.926731e-08, 
    -1.907459e-08, -1.913045e-08, -1.933574e-08, -1.963976e-08, 
    -2.003454e-08, -2.025808e-08,
  -1.600552e-08, -1.64799e-08, -1.693421e-08, -1.746878e-08, -1.814645e-08, 
    -1.900054e-08, -1.982949e-08, -2.032773e-08, -2.024895e-08, 
    -2.000637e-08, -1.977988e-08, -1.961633e-08, -1.949517e-08, 
    -1.954195e-08, -1.970683e-08,
  -1.540318e-08, -1.573117e-08, -1.611847e-08, -1.652472e-08, -1.696156e-08, 
    -1.750375e-08, -1.830113e-08, -1.927646e-08, -2.0021e-08, -2.02336e-08, 
    -2.029247e-08, -2.018616e-08, -2.005403e-08, -1.996241e-08, -2.005974e-08,
  -1.496859e-08, -1.490702e-08, -1.517471e-08, -1.571605e-08, -1.627925e-08, 
    -1.690076e-08, -1.758554e-08, -1.839339e-08, -1.927229e-08, 
    -1.996434e-08, -2.035575e-08, -2.032055e-08, -2.023217e-08, 
    -2.024323e-08, -2.023446e-08,
  -1.546739e-08, -1.535572e-08, -1.502028e-08, -1.46917e-08, -1.507315e-08, 
    -1.55437e-08, -1.62514e-08, -1.719532e-08, -1.816724e-08, -1.925042e-08, 
    -1.99942e-08, -2.032787e-08, -2.035996e-08, -2.038039e-08, -2.03727e-08,
  -1.647587e-08, -1.662107e-08, -1.681457e-08, -1.683378e-08, -1.669151e-08, 
    -1.635838e-08, -1.596306e-08, -1.603314e-08, -1.650155e-08, 
    -1.737459e-08, -1.835091e-08, -1.933646e-08, -2.000372e-08, 
    -2.030422e-08, -2.03491e-08,
  -1.664934e-08, -1.662038e-08, -1.671247e-08, -1.738765e-08, -1.797337e-08, 
    -1.802323e-08, -1.787948e-08, -1.738957e-08, -1.701727e-08, 
    -1.704059e-08, -1.731314e-08, -1.785573e-08, -1.843383e-08, 
    -1.910483e-08, -1.957234e-08,
  -1.628753e-08, -1.641732e-08, -1.642311e-08, -1.669514e-08, -1.693663e-08, 
    -1.734438e-08, -1.790427e-08, -1.828531e-08, -1.828075e-08, -1.78447e-08, 
    -1.755409e-08, -1.744085e-08, -1.750129e-08, -1.786743e-08, -1.820387e-08,
  -1.613542e-08, -1.585271e-08, -1.579663e-08, -1.578548e-08, -1.609243e-08, 
    -1.627234e-08, -1.650349e-08, -1.69095e-08, -1.747476e-08, -1.772062e-08, 
    -1.776063e-08, -1.740266e-08, -1.700878e-08, -1.707749e-08, -1.721276e-08,
  -1.487158e-08, -1.499559e-08, -1.518141e-08, -1.534639e-08, -1.553177e-08, 
    -1.563509e-08, -1.574764e-08, -1.577286e-08, -1.582687e-08, 
    -1.584093e-08, -1.586955e-08, -1.58909e-08, -1.598384e-08, -1.611403e-08, 
    -1.623355e-08,
  -1.473488e-08, -1.491542e-08, -1.511201e-08, -1.523617e-08, -1.533492e-08, 
    -1.542887e-08, -1.553758e-08, -1.563339e-08, -1.571953e-08, 
    -1.580731e-08, -1.58384e-08, -1.588921e-08, -1.594155e-08, -1.608408e-08, 
    -1.62561e-08,
  -1.449262e-08, -1.478613e-08, -1.510505e-08, -1.536719e-08, -1.557532e-08, 
    -1.571194e-08, -1.582548e-08, -1.589201e-08, -1.590507e-08, 
    -1.589487e-08, -1.592598e-08, -1.603e-08, -1.621643e-08, -1.641254e-08, 
    -1.663499e-08,
  -1.443272e-08, -1.47085e-08, -1.494005e-08, -1.516838e-08, -1.530263e-08, 
    -1.541702e-08, -1.553367e-08, -1.560833e-08, -1.565666e-08, 
    -1.576367e-08, -1.591709e-08, -1.619781e-08, -1.647322e-08, 
    -1.667065e-08, -1.677983e-08,
  -1.453221e-08, -1.484015e-08, -1.512228e-08, -1.540439e-08, -1.559266e-08, 
    -1.575415e-08, -1.585609e-08, -1.593138e-08, -1.605091e-08, 
    -1.618396e-08, -1.641346e-08, -1.648396e-08, -1.65799e-08, -1.662941e-08, 
    -1.669826e-08,
  -1.45477e-08, -1.498243e-08, -1.525223e-08, -1.560135e-08, -1.593547e-08, 
    -1.625261e-08, -1.644448e-08, -1.67566e-08, -1.704584e-08, -1.728086e-08, 
    -1.741191e-08, -1.742428e-08, -1.734765e-08, -1.718729e-08, -1.693984e-08,
  -1.470425e-08, -1.524933e-08, -1.562541e-08, -1.586613e-08, -1.624119e-08, 
    -1.650567e-08, -1.674242e-08, -1.688027e-08, -1.718383e-08, 
    -1.751123e-08, -1.774848e-08, -1.780546e-08, -1.767663e-08, 
    -1.745239e-08, -1.707849e-08,
  -1.459222e-08, -1.498028e-08, -1.558869e-08, -1.592271e-08, -1.626358e-08, 
    -1.629548e-08, -1.646794e-08, -1.650488e-08, -1.68583e-08, -1.714098e-08, 
    -1.733821e-08, -1.722717e-08, -1.707833e-08, -1.67619e-08, -1.650969e-08,
  -1.456346e-08, -1.500023e-08, -1.541605e-08, -1.593249e-08, -1.620013e-08, 
    -1.62462e-08, -1.622367e-08, -1.647336e-08, -1.680537e-08, -1.697195e-08, 
    -1.682671e-08, -1.650761e-08, -1.619907e-08, -1.607552e-08, -1.614186e-08,
  -1.414829e-08, -1.450574e-08, -1.491355e-08, -1.550103e-08, -1.556488e-08, 
    -1.548588e-08, -1.566587e-08, -1.592172e-08, -1.570635e-08, 
    -1.528099e-08, -1.453219e-08, -1.403249e-08, -1.373581e-08, 
    -1.380775e-08, -1.404927e-08,
  -1.689516e-08, -1.709531e-08, -1.730561e-08, -1.748168e-08, -1.763365e-08, 
    -1.784509e-08, -1.809702e-08, -1.835766e-08, -1.853959e-08, 
    -1.865964e-08, -1.877921e-08, -1.889702e-08, -1.896924e-08, 
    -1.900499e-08, -1.902207e-08,
  -1.659712e-08, -1.675939e-08, -1.69281e-08, -1.710977e-08, -1.721705e-08, 
    -1.734722e-08, -1.752401e-08, -1.768917e-08, -1.785904e-08, 
    -1.799013e-08, -1.805945e-08, -1.81155e-08, -1.809246e-08, -1.804533e-08, 
    -1.795074e-08,
  -1.651551e-08, -1.661613e-08, -1.672315e-08, -1.68271e-08, -1.692521e-08, 
    -1.701686e-08, -1.713862e-08, -1.729427e-08, -1.747197e-08, 
    -1.764498e-08, -1.775909e-08, -1.777403e-08, -1.768623e-08, 
    -1.756192e-08, -1.740342e-08,
  -1.613473e-08, -1.634231e-08, -1.650871e-08, -1.664593e-08, -1.675422e-08, 
    -1.685502e-08, -1.696883e-08, -1.710323e-08, -1.728499e-08, 
    -1.747453e-08, -1.759387e-08, -1.760408e-08, -1.756725e-08, 
    -1.748835e-08, -1.74786e-08,
  -1.551085e-08, -1.574983e-08, -1.598505e-08, -1.624163e-08, -1.646027e-08, 
    -1.665887e-08, -1.677559e-08, -1.69519e-08, -1.71447e-08, -1.733082e-08, 
    -1.743245e-08, -1.753097e-08, -1.754842e-08, -1.754774e-08, -1.75232e-08,
  -1.482082e-08, -1.499655e-08, -1.524164e-08, -1.558608e-08, -1.589926e-08, 
    -1.618464e-08, -1.644057e-08, -1.66686e-08, -1.687822e-08, -1.706845e-08, 
    -1.716734e-08, -1.729232e-08, -1.730318e-08, -1.725846e-08, -1.721542e-08,
  -1.437987e-08, -1.43589e-08, -1.444993e-08, -1.470013e-08, -1.501135e-08, 
    -1.535332e-08, -1.570047e-08, -1.59829e-08, -1.619939e-08, -1.634164e-08, 
    -1.646386e-08, -1.652256e-08, -1.653809e-08, -1.653654e-08, -1.652988e-08,
  -1.414332e-08, -1.41085e-08, -1.411197e-08, -1.417488e-08, -1.430499e-08, 
    -1.450565e-08, -1.481989e-08, -1.5085e-08, -1.529915e-08, -1.539792e-08, 
    -1.54379e-08, -1.544812e-08, -1.543133e-08, -1.542498e-08, -1.538563e-08,
  -1.393223e-08, -1.385624e-08, -1.379335e-08, -1.379168e-08, -1.384045e-08, 
    -1.397763e-08, -1.422244e-08, -1.44464e-08, -1.462052e-08, -1.463191e-08, 
    -1.463849e-08, -1.457393e-08, -1.44907e-08, -1.440559e-08, -1.427854e-08,
  -1.376215e-08, -1.361609e-08, -1.350068e-08, -1.342254e-08, -1.335822e-08, 
    -1.343606e-08, -1.362135e-08, -1.384377e-08, -1.399191e-08, 
    -1.401235e-08, -1.399916e-08, -1.384688e-08, -1.365579e-08, 
    -1.341527e-08, -1.315353e-08,
  -1.971721e-08, -1.973511e-08, -1.974221e-08, -1.97282e-08, -1.975099e-08, 
    -1.971902e-08, -1.97396e-08, -1.982226e-08, -1.994987e-08, -2.007628e-08, 
    -2.019068e-08, -2.025266e-08, -2.03244e-08, -2.03881e-08, -2.058995e-08,
  -1.8391e-08, -1.830346e-08, -1.835934e-08, -1.844895e-08, -1.852043e-08, 
    -1.855773e-08, -1.859219e-08, -1.862173e-08, -1.867093e-08, 
    -1.873111e-08, -1.879561e-08, -1.888587e-08, -1.894257e-08, 
    -1.901609e-08, -1.900804e-08,
  -1.73494e-08, -1.706016e-08, -1.699535e-08, -1.690345e-08, -1.691359e-08, 
    -1.693746e-08, -1.70164e-08, -1.705343e-08, -1.710841e-08, -1.715659e-08, 
    -1.720597e-08, -1.725638e-08, -1.730387e-08, -1.737206e-08, -1.739979e-08,
  -1.650064e-08, -1.621678e-08, -1.596652e-08, -1.580963e-08, -1.568314e-08, 
    -1.55908e-08, -1.552511e-08, -1.551901e-08, -1.558418e-08, -1.565946e-08, 
    -1.573532e-08, -1.582198e-08, -1.591623e-08, -1.602502e-08, -1.612232e-08,
  -1.626807e-08, -1.590476e-08, -1.564199e-08, -1.532952e-08, -1.507886e-08, 
    -1.482394e-08, -1.463652e-08, -1.454333e-08, -1.447223e-08, 
    -1.446051e-08, -1.445775e-08, -1.449935e-08, -1.459056e-08, 
    -1.472766e-08, -1.488406e-08,
  -1.600241e-08, -1.568159e-08, -1.534737e-08, -1.498369e-08, -1.456327e-08, 
    -1.420335e-08, -1.394429e-08, -1.37886e-08, -1.367032e-08, -1.35974e-08, 
    -1.355337e-08, -1.356903e-08, -1.368021e-08, -1.387945e-08, -1.411728e-08,
  -1.52855e-08, -1.49594e-08, -1.462932e-08, -1.41651e-08, -1.371391e-08, 
    -1.333099e-08, -1.305231e-08, -1.287495e-08, -1.279279e-08, 
    -1.274763e-08, -1.276357e-08, -1.288904e-08, -1.306936e-08, 
    -1.332306e-08, -1.360634e-08,
  -1.454762e-08, -1.418235e-08, -1.381202e-08, -1.334984e-08, -1.295362e-08, 
    -1.265856e-08, -1.245899e-08, -1.236333e-08, -1.235794e-08, 
    -1.240242e-08, -1.253517e-08, -1.274101e-08, -1.294885e-08, 
    -1.320833e-08, -1.346694e-08,
  -1.416338e-08, -1.379751e-08, -1.342123e-08, -1.303968e-08, -1.275785e-08, 
    -1.253256e-08, -1.240045e-08, -1.234901e-08, -1.239372e-08, 
    -1.251556e-08, -1.272311e-08, -1.296481e-08, -1.327565e-08, 
    -1.359936e-08, -1.390204e-08,
  -1.404712e-08, -1.377924e-08, -1.355143e-08, -1.329577e-08, -1.314057e-08, 
    -1.299537e-08, -1.287547e-08, -1.280883e-08, -1.283483e-08, 
    -1.294457e-08, -1.31372e-08, -1.344105e-08, -1.380278e-08, -1.419432e-08, 
    -1.455889e-08,
  -1.779614e-08, -1.758746e-08, -1.745919e-08, -1.748448e-08, -1.74421e-08, 
    -1.749069e-08, -1.754898e-08, -1.758783e-08, -1.784637e-08, 
    -1.832055e-08, -1.899719e-08, -2.021956e-08, -2.175301e-08, 
    -2.267205e-08, -2.321264e-08,
  -1.848074e-08, -1.819546e-08, -1.799981e-08, -1.788073e-08, -1.767599e-08, 
    -1.76523e-08, -1.774435e-08, -1.789501e-08, -1.798411e-08, -1.822782e-08, 
    -1.854147e-08, -1.910859e-08, -2.014441e-08, -2.12079e-08, -2.211795e-08,
  -1.931246e-08, -1.907941e-08, -1.884247e-08, -1.867448e-08, -1.849939e-08, 
    -1.830232e-08, -1.817278e-08, -1.81798e-08, -1.830491e-08, -1.842345e-08, 
    -1.864144e-08, -1.886674e-08, -1.926345e-08, -2.009103e-08, -2.080062e-08,
  -1.965044e-08, -1.96953e-08, -1.966331e-08, -1.952398e-08, -1.93274e-08, 
    -1.917916e-08, -1.886593e-08, -1.879824e-08, -1.870303e-08, 
    -1.883406e-08, -1.88704e-08, -1.911715e-08, -1.912339e-08, -1.94907e-08, 
    -1.981639e-08,
  -1.955056e-08, -1.98546e-08, -1.991806e-08, -1.995263e-08, -1.981113e-08, 
    -1.971734e-08, -1.948409e-08, -1.941161e-08, -1.925684e-08, 
    -1.926207e-08, -1.928466e-08, -1.948318e-08, -1.963864e-08, 
    -1.971453e-08, -1.980864e-08,
  -1.943391e-08, -1.978784e-08, -1.999275e-08, -2.016601e-08, -2.01892e-08, 
    -2.025832e-08, -2.025884e-08, -2.032355e-08, -2.032785e-08, 
    -2.028309e-08, -2.015808e-08, -2.001887e-08, -1.987915e-08, 
    -1.982795e-08, -1.980031e-08,
  -1.944377e-08, -1.963422e-08, -1.99167e-08, -1.997312e-08, -2.002729e-08, 
    -2.008513e-08, -2.01812e-08, -2.032124e-08, -2.042414e-08, -2.044426e-08, 
    -2.032606e-08, -2.013757e-08, -1.988349e-08, -1.959123e-08, -1.933824e-08,
  -1.943813e-08, -1.958576e-08, -1.984887e-08, -1.972938e-08, -1.969151e-08, 
    -1.950742e-08, -1.961894e-08, -1.969278e-08, -1.958975e-08, -1.94373e-08, 
    -1.919204e-08, -1.894279e-08, -1.868341e-08, -1.843391e-08, -1.820607e-08,
  -1.898491e-08, -1.926836e-08, -1.946375e-08, -1.934499e-08, -1.878074e-08, 
    -1.88104e-08, -1.876503e-08, -1.864004e-08, -1.840198e-08, -1.805896e-08, 
    -1.766364e-08, -1.732178e-08, -1.699642e-08, -1.668386e-08, -1.644909e-08,
  -1.814869e-08, -1.849099e-08, -1.878864e-08, -1.829566e-08, -1.778288e-08, 
    -1.770419e-08, -1.757037e-08, -1.726325e-08, -1.678066e-08, 
    -1.634124e-08, -1.582643e-08, -1.54674e-08, -1.509404e-08, -1.482856e-08, 
    -1.459165e-08,
  -2.185252e-08, -2.127887e-08, -2.059758e-08, -1.98567e-08, -1.93551e-08, 
    -1.922976e-08, -1.93174e-08, -1.956772e-08, -2.034169e-08, -2.077751e-08, 
    -2.046459e-08, -1.989739e-08, -1.999123e-08, -2.128936e-08, -2.383706e-08,
  -2.164065e-08, -2.141868e-08, -2.072665e-08, -1.997076e-08, -1.934153e-08, 
    -1.896803e-08, -1.913502e-08, -1.935179e-08, -1.997448e-08, 
    -2.079385e-08, -2.102702e-08, -2.003508e-08, -1.936029e-08, 
    -2.009778e-08, -2.122355e-08,
  -2.147388e-08, -2.133359e-08, -2.085627e-08, -2.012075e-08, -1.941776e-08, 
    -1.896424e-08, -1.880874e-08, -1.903031e-08, -1.936664e-08, 
    -2.002572e-08, -2.064114e-08, -2.081616e-08, -1.960906e-08, -1.93734e-08, 
    -1.973401e-08,
  -2.113922e-08, -2.115842e-08, -2.091683e-08, -2.031675e-08, -1.957385e-08, 
    -1.896992e-08, -1.866802e-08, -1.874876e-08, -1.90786e-08, -1.94852e-08, 
    -1.987872e-08, -2.043924e-08, -2.009287e-08, -1.954844e-08, -1.899428e-08,
  -2.076646e-08, -2.074915e-08, -2.073597e-08, -2.028377e-08, -1.961983e-08, 
    -1.901594e-08, -1.852084e-08, -1.837348e-08, -1.848308e-08, 
    -1.881361e-08, -1.925602e-08, -1.97242e-08, -2.00438e-08, -1.984278e-08, 
    -1.961629e-08,
  -2.010074e-08, -2.008964e-08, -2.013011e-08, -1.989833e-08, -1.938348e-08, 
    -1.882771e-08, -1.832993e-08, -1.807392e-08, -1.797044e-08, 
    -1.803711e-08, -1.824954e-08, -1.872437e-08, -1.8968e-08, -1.950173e-08, 
    -1.921518e-08,
  -1.934884e-08, -1.93766e-08, -1.942743e-08, -1.934884e-08, -1.915125e-08, 
    -1.870823e-08, -1.819383e-08, -1.78184e-08, -1.75255e-08, -1.754648e-08, 
    -1.752626e-08, -1.769571e-08, -1.787237e-08, -1.812036e-08, -1.848334e-08,
  -1.848139e-08, -1.844659e-08, -1.857669e-08, -1.864803e-08, -1.856289e-08, 
    -1.842212e-08, -1.798653e-08, -1.770007e-08, -1.738655e-08, 
    -1.735005e-08, -1.735078e-08, -1.744623e-08, -1.752267e-08, 
    -1.762843e-08, -1.778098e-08,
  -1.764345e-08, -1.770291e-08, -1.772652e-08, -1.782294e-08, -1.787507e-08, 
    -1.781357e-08, -1.762011e-08, -1.719207e-08, -1.697688e-08, 
    -1.680664e-08, -1.694854e-08, -1.709369e-08, -1.722397e-08, 
    -1.735609e-08, -1.749996e-08,
  -1.683173e-08, -1.693688e-08, -1.71573e-08, -1.712794e-08, -1.716626e-08, 
    -1.722533e-08, -1.725037e-08, -1.697106e-08, -1.664242e-08, 
    -1.636695e-08, -1.638145e-08, -1.638129e-08, -1.648901e-08, 
    -1.654532e-08, -1.668224e-08,
  -2.01912e-08, -2.140944e-08, -2.281207e-08, -2.365667e-08, -2.377034e-08, 
    -2.370004e-08, -2.335089e-08, -2.303961e-08, -2.283819e-08, 
    -2.315373e-08, -2.335878e-08, -2.344989e-08, -2.345704e-08, 
    -2.325383e-08, -2.301707e-08,
  -1.975701e-08, -2.076662e-08, -2.224596e-08, -2.363358e-08, -2.411539e-08, 
    -2.395948e-08, -2.349494e-08, -2.323353e-08, -2.28742e-08, -2.290582e-08, 
    -2.339155e-08, -2.346997e-08, -2.321874e-08, -2.3502e-08, -2.332204e-08,
  -1.932353e-08, -2.019634e-08, -2.145914e-08, -2.311084e-08, -2.436244e-08, 
    -2.44726e-08, -2.377748e-08, -2.329489e-08, -2.286076e-08, -2.268852e-08, 
    -2.290806e-08, -2.362929e-08, -2.326407e-08, -2.296997e-08, -2.387182e-08,
  -1.86576e-08, -1.96736e-08, -2.078754e-08, -2.22385e-08, -2.398413e-08, 
    -2.475812e-08, -2.44836e-08, -2.374089e-08, -2.302271e-08, -2.254598e-08, 
    -2.255339e-08, -2.287566e-08, -2.38888e-08, -2.320195e-08, -2.334058e-08,
  -1.792323e-08, -1.898679e-08, -2.017416e-08, -2.150823e-08, -2.328157e-08, 
    -2.466434e-08, -2.485909e-08, -2.449119e-08, -2.371956e-08, 
    -2.274389e-08, -2.2401e-08, -2.238097e-08, -2.301292e-08, -2.420122e-08, 
    -2.366884e-08,
  -1.718284e-08, -1.817748e-08, -1.935369e-08, -2.064378e-08, -2.230609e-08, 
    -2.425325e-08, -2.505158e-08, -2.508912e-08, -2.446565e-08, 
    -2.372921e-08, -2.269561e-08, -2.225007e-08, -2.221715e-08, 
    -2.274768e-08, -2.375863e-08,
  -1.633441e-08, -1.745932e-08, -1.855294e-08, -1.977102e-08, -2.115076e-08, 
    -2.312542e-08, -2.449359e-08, -2.521276e-08, -2.533451e-08, 
    -2.477901e-08, -2.402355e-08, -2.306956e-08, -2.268466e-08, 
    -2.225643e-08, -2.228144e-08,
  -1.531444e-08, -1.661027e-08, -1.771081e-08, -1.883109e-08, -2.010517e-08, 
    -2.177869e-08, -2.345084e-08, -2.438781e-08, -2.49531e-08, -2.504465e-08, 
    -2.469879e-08, -2.411649e-08, -2.345819e-08, -2.302381e-08, -2.214737e-08,
  -1.435691e-08, -1.569237e-08, -1.675952e-08, -1.784544e-08, -1.892515e-08, 
    -2.030871e-08, -2.210001e-08, -2.331557e-08, -2.41203e-08, -2.46392e-08, 
    -2.478216e-08, -2.453192e-08, -2.400342e-08, -2.341133e-08, -2.270141e-08,
  -1.345452e-08, -1.466153e-08, -1.589373e-08, -1.69705e-08, -1.795766e-08, 
    -1.900365e-08, -2.039302e-08, -2.189666e-08, -2.272162e-08, -2.32862e-08, 
    -2.356545e-08, -2.371378e-08, -2.363848e-08, -2.310099e-08, -2.256258e-08,
  -1.803891e-08, -1.77716e-08, -1.748978e-08, -1.751223e-08, -1.775822e-08, 
    -1.810513e-08, -1.876801e-08, -1.969397e-08, -1.989468e-08, -2.01849e-08, 
    -2.073339e-08, -2.183572e-08, -2.338951e-08, -2.461704e-08, -2.506083e-08,
  -1.821725e-08, -1.782659e-08, -1.735097e-08, -1.725745e-08, -1.747549e-08, 
    -1.799846e-08, -1.881197e-08, -1.960622e-08, -2.012807e-08, 
    -2.042312e-08, -2.09991e-08, -2.194352e-08, -2.27551e-08, -2.365006e-08, 
    -2.377461e-08,
  -1.813108e-08, -1.77209e-08, -1.72848e-08, -1.695149e-08, -1.717184e-08, 
    -1.745804e-08, -1.857008e-08, -1.941165e-08, -2.007248e-08, -2.06548e-08, 
    -2.105724e-08, -2.19659e-08, -2.283966e-08, -2.347651e-08, -2.347926e-08,
  -1.810741e-08, -1.768673e-08, -1.724393e-08, -1.683377e-08, -1.67779e-08, 
    -1.721867e-08, -1.796731e-08, -1.930261e-08, -2.001176e-08, 
    -2.065019e-08, -2.115545e-08, -2.199427e-08, -2.271843e-08, 
    -2.347815e-08, -2.351549e-08,
  -1.787785e-08, -1.772388e-08, -1.728567e-08, -1.673369e-08, -1.649443e-08, 
    -1.673919e-08, -1.746612e-08, -1.869609e-08, -1.992201e-08, 
    -2.056926e-08, -2.119228e-08, -2.21303e-08, -2.30547e-08, -2.356619e-08, 
    -2.348066e-08,
  -1.757827e-08, -1.751073e-08, -1.735204e-08, -1.685201e-08, -1.640929e-08, 
    -1.630575e-08, -1.698407e-08, -1.803167e-08, -1.944695e-08, -2.06824e-08, 
    -2.112156e-08, -2.196354e-08, -2.293189e-08, -2.370685e-08, -2.378999e-08,
  -1.761141e-08, -1.736933e-08, -1.712859e-08, -1.686027e-08, -1.635721e-08, 
    -1.613527e-08, -1.624898e-08, -1.738216e-08, -1.854589e-08, 
    -2.025684e-08, -2.139689e-08, -2.207022e-08, -2.290583e-08, 
    -2.378731e-08, -2.371332e-08,
  -1.759209e-08, -1.748631e-08, -1.719025e-08, -1.694793e-08, -1.635022e-08, 
    -1.611328e-08, -1.592254e-08, -1.658092e-08, -1.773367e-08, 
    -1.913279e-08, -2.102007e-08, -2.208368e-08, -2.269249e-08, 
    -2.385218e-08, -2.432717e-08,
  -1.742136e-08, -1.72959e-08, -1.717954e-08, -1.697285e-08, -1.648543e-08, 
    -1.598424e-08, -1.584985e-08, -1.591433e-08, -1.695804e-08, 
    -1.803006e-08, -1.9674e-08, -2.190401e-08, -2.264821e-08, -2.344137e-08, 
    -2.392548e-08,
  -1.714515e-08, -1.72235e-08, -1.713764e-08, -1.70449e-08, -1.684459e-08, 
    -1.621475e-08, -1.579946e-08, -1.566172e-08, -1.611554e-08, 
    -1.733979e-08, -1.823335e-08, -2.035338e-08, -2.253572e-08, 
    -2.355742e-08, -2.425623e-08,
  -1.982536e-08, -2.003144e-08, -2.004381e-08, -2.021072e-08, -2.038345e-08, 
    -2.059867e-08, -2.060726e-08, -2.031959e-08, -2.020457e-08, -1.98901e-08, 
    -1.977991e-08, -1.965146e-08, -2.003061e-08, -2.016078e-08, -2.04528e-08,
  -1.975782e-08, -2.006231e-08, -2.026181e-08, -2.040165e-08, -2.04638e-08, 
    -2.074077e-08, -2.054402e-08, -2.05427e-08, -2.01572e-08, -1.997257e-08, 
    -1.986681e-08, -1.9753e-08, -1.978965e-08, -2.031567e-08, -2.081487e-08,
  -1.960815e-08, -1.986377e-08, -2.010243e-08, -2.051336e-08, -2.054689e-08, 
    -2.077362e-08, -2.069067e-08, -2.035243e-08, -2.026531e-08, 
    -1.996898e-08, -1.957111e-08, -1.953454e-08, -1.976204e-08, -2.02006e-08, 
    -2.092212e-08,
  -1.941451e-08, -1.975095e-08, -1.992789e-08, -2.0385e-08, -2.044678e-08, 
    -2.070066e-08, -2.069852e-08, -2.06002e-08, -2.021457e-08, -2.010939e-08, 
    -1.959658e-08, -1.934715e-08, -1.952866e-08, -2.022191e-08, -2.081202e-08,
  -1.916573e-08, -1.966218e-08, -1.981953e-08, -2.01487e-08, -2.03036e-08, 
    -2.040498e-08, -2.060613e-08, -2.05541e-08, -2.039401e-08, -2.002798e-08, 
    -1.950088e-08, -1.935522e-08, -1.939098e-08, -2.015015e-08, -2.069003e-08,
  -1.899199e-08, -1.947074e-08, -1.975518e-08, -2.000287e-08, -2.024939e-08, 
    -2.014813e-08, -2.037901e-08, -2.056147e-08, -2.032665e-08, 
    -2.016371e-08, -1.967391e-08, -1.920252e-08, -1.922857e-08, 
    -2.004332e-08, -2.052068e-08,
  -1.881857e-08, -1.923598e-08, -1.954941e-08, -1.972903e-08, -2.006165e-08, 
    -2.011241e-08, -2.006703e-08, -2.048583e-08, -2.035586e-08, 
    -2.011249e-08, -1.973036e-08, -1.953341e-08, -1.910045e-08, 
    -1.991255e-08, -2.030694e-08,
  -1.904544e-08, -1.907939e-08, -1.938138e-08, -1.949534e-08, -1.968906e-08, 
    -2.00044e-08, -1.996091e-08, -2.01074e-08, -2.040983e-08, -2.015277e-08, 
    -1.977399e-08, -1.930111e-08, -1.927796e-08, -1.94666e-08, -2.036293e-08,
  -1.897117e-08, -1.915899e-08, -1.926268e-08, -1.936517e-08, -1.933518e-08, 
    -1.961731e-08, -1.987323e-08, -2.009256e-08, -2.017324e-08, 
    -2.031081e-08, -1.999977e-08, -1.962724e-08, -1.899543e-08, 
    -1.918409e-08, -1.932728e-08,
  -1.869948e-08, -1.90435e-08, -1.91634e-08, -1.940397e-08, -1.923852e-08, 
    -1.930709e-08, -1.945684e-08, -2.001311e-08, -1.99666e-08, -2.007325e-08, 
    -2.009517e-08, -1.988174e-08, -1.946032e-08, -1.899096e-08, -1.913672e-08,
  -1.996254e-08, -2.008871e-08, -2.027302e-08, -2.028903e-08, -2.039259e-08, 
    -2.029438e-08, -2.041788e-08, -2.071993e-08, -2.096505e-08, -2.13881e-08, 
    -2.108931e-08, -2.101145e-08, -2.101086e-08, -2.097114e-08, -2.069799e-08,
  -1.912735e-08, -1.95001e-08, -1.965324e-08, -1.989971e-08, -2.012751e-08, 
    -2.024749e-08, -2.016628e-08, -2.059638e-08, -2.076808e-08, 
    -2.104479e-08, -2.109892e-08, -2.087507e-08, -2.072642e-08, 
    -2.081242e-08, -2.076576e-08,
  -1.826717e-08, -1.87996e-08, -1.900113e-08, -1.926089e-08, -1.962109e-08, 
    -2.005054e-08, -2.012502e-08, -2.049828e-08, -2.058316e-08, 
    -2.075301e-08, -2.088707e-08, -2.073375e-08, -2.064369e-08, 
    -2.050483e-08, -2.046221e-08,
  -1.748524e-08, -1.799975e-08, -1.837829e-08, -1.867111e-08, -1.907188e-08, 
    -1.955082e-08, -1.988862e-08, -2.01996e-08, -2.03799e-08, -2.056817e-08, 
    -2.060562e-08, -2.058872e-08, -2.04403e-08, -2.036098e-08, -2.036151e-08,
  -1.670652e-08, -1.719393e-08, -1.776381e-08, -1.808903e-08, -1.857238e-08, 
    -1.906341e-08, -1.953235e-08, -1.987544e-08, -2.020621e-08, 
    -2.034469e-08, -2.036268e-08, -2.043686e-08, -2.039669e-08, 
    -2.043803e-08, -2.037151e-08,
  -1.607113e-08, -1.670262e-08, -1.70987e-08, -1.763465e-08, -1.806819e-08, 
    -1.854681e-08, -1.904252e-08, -1.93988e-08, -1.984216e-08, -2.013923e-08, 
    -2.023202e-08, -2.026055e-08, -2.03504e-08, -2.044042e-08, -2.053705e-08,
  -1.50523e-08, -1.579525e-08, -1.645301e-08, -1.701991e-08, -1.770735e-08, 
    -1.821189e-08, -1.859732e-08, -1.89864e-08, -1.942018e-08, -1.982624e-08, 
    -2.014035e-08, -2.034743e-08, -2.041102e-08, -2.054128e-08, -2.048009e-08,
  -1.450135e-08, -1.511067e-08, -1.573477e-08, -1.636094e-08, -1.707585e-08, 
    -1.775872e-08, -1.821274e-08, -1.85872e-08, -1.907712e-08, -1.95324e-08, 
    -1.983875e-08, -2.019661e-08, -2.043007e-08, -2.061985e-08, -2.069068e-08,
  -1.389536e-08, -1.452927e-08, -1.515101e-08, -1.581097e-08, -1.644858e-08, 
    -1.721598e-08, -1.779618e-08, -1.822549e-08, -1.875948e-08, 
    -1.929008e-08, -1.970154e-08, -2.00043e-08, -2.028659e-08, -2.062498e-08, 
    -2.073906e-08,
  -1.319221e-08, -1.398997e-08, -1.46389e-08, -1.527387e-08, -1.591e-08, 
    -1.656393e-08, -1.724784e-08, -1.784181e-08, -1.838406e-08, 
    -1.898425e-08, -1.944657e-08, -1.987986e-08, -2.013825e-08, 
    -2.050179e-08, -2.065702e-08,
  -2.173339e-08, -2.162566e-08, -2.163962e-08, -2.188797e-08, -2.265901e-08, 
    -2.371948e-08, -2.437662e-08, -2.462544e-08, -2.429952e-08, 
    -2.458627e-08, -2.514157e-08, -2.623271e-08, -2.681974e-08, 
    -2.707559e-08, -2.645542e-08,
  -2.21363e-08, -2.194514e-08, -2.181015e-08, -2.17842e-08, -2.179194e-08, 
    -2.190176e-08, -2.227263e-08, -2.256616e-08, -2.303873e-08, -2.32066e-08, 
    -2.390625e-08, -2.45864e-08, -2.473599e-08, -2.50524e-08, -2.479962e-08,
  -2.217023e-08, -2.233208e-08, -2.230373e-08, -2.216287e-08, -2.191115e-08, 
    -2.181862e-08, -2.183752e-08, -2.16969e-08, -2.179288e-08, -2.171603e-08, 
    -2.213282e-08, -2.2694e-08, -2.298466e-08, -2.337004e-08, -2.373528e-08,
  -2.124497e-08, -2.184118e-08, -2.209159e-08, -2.221889e-08, -2.22101e-08, 
    -2.207625e-08, -2.189154e-08, -2.165151e-08, -2.166333e-08, 
    -2.158226e-08, -2.189066e-08, -2.202712e-08, -2.242022e-08, 
    -2.274099e-08, -2.300195e-08,
  -2.019616e-08, -2.084458e-08, -2.157227e-08, -2.194842e-08, -2.215345e-08, 
    -2.221687e-08, -2.213909e-08, -2.206353e-08, -2.190844e-08, 
    -2.186229e-08, -2.196174e-08, -2.20997e-08, -2.215967e-08, -2.226255e-08, 
    -2.233317e-08,
  -1.842544e-08, -1.917287e-08, -1.99413e-08, -2.062264e-08, -2.11683e-08, 
    -2.149135e-08, -2.17899e-08, -2.184963e-08, -2.206487e-08, -2.229583e-08, 
    -2.248435e-08, -2.26611e-08, -2.25949e-08, -2.247421e-08, -2.232603e-08,
  -1.758852e-08, -1.778182e-08, -1.836489e-08, -1.89359e-08, -1.967001e-08, 
    -2.017599e-08, -2.057793e-08, -2.082143e-08, -2.116253e-08, 
    -2.160388e-08, -2.202393e-08, -2.237477e-08, -2.266354e-08, 
    -2.277564e-08, -2.272729e-08,
  -1.717463e-08, -1.724196e-08, -1.727669e-08, -1.756799e-08, -1.790113e-08, 
    -1.843783e-08, -1.89194e-08, -1.929781e-08, -1.96207e-08, -2.001452e-08, 
    -2.048797e-08, -2.095404e-08, -2.127927e-08, -2.165759e-08, -2.18376e-08,
  -1.616898e-08, -1.653416e-08, -1.663172e-08, -1.680567e-08, -1.691022e-08, 
    -1.719175e-08, -1.743439e-08, -1.780885e-08, -1.799359e-08, 
    -1.821813e-08, -1.839001e-08, -1.881249e-08, -1.921739e-08, 
    -1.979868e-08, -2.025675e-08,
  -1.557622e-08, -1.559294e-08, -1.573423e-08, -1.574042e-08, -1.598356e-08, 
    -1.614856e-08, -1.635552e-08, -1.652291e-08, -1.679371e-08, 
    -1.693916e-08, -1.712832e-08, -1.722688e-08, -1.739457e-08, 
    -1.778706e-08, -1.826758e-08,
  -1.587758e-08, -1.713462e-08, -1.930409e-08, -2.161326e-08, -2.348619e-08, 
    -2.534173e-08, -2.751662e-08, -2.838176e-08, -2.911166e-08, 
    -2.913248e-08, -2.892121e-08, -2.865025e-08, -2.86581e-08, -2.922136e-08, 
    -2.936648e-08,
  -1.654326e-08, -1.678919e-08, -1.74992e-08, -1.900797e-08, -2.148469e-08, 
    -2.322275e-08, -2.476576e-08, -2.622208e-08, -2.704193e-08, 
    -2.757049e-08, -2.776443e-08, -2.811788e-08, -2.83545e-08, -2.825174e-08, 
    -2.799424e-08,
  -1.662752e-08, -1.679532e-08, -1.733271e-08, -1.784897e-08, -1.890705e-08, 
    -2.07359e-08, -2.235818e-08, -2.36428e-08, -2.478392e-08, -2.539827e-08, 
    -2.594232e-08, -2.632334e-08, -2.646409e-08, -2.630873e-08, -2.570866e-08,
  -1.757723e-08, -1.728374e-08, -1.722417e-08, -1.763009e-08, -1.820243e-08, 
    -1.873691e-08, -1.994101e-08, -2.113827e-08, -2.256316e-08, 
    -2.343678e-08, -2.427966e-08, -2.453887e-08, -2.471356e-08, 
    -2.460231e-08, -2.436006e-08,
  -1.889441e-08, -1.846608e-08, -1.825859e-08, -1.793782e-08, -1.813679e-08, 
    -1.845601e-08, -1.885409e-08, -1.93059e-08, -2.006614e-08, -2.101592e-08, 
    -2.181165e-08, -2.245368e-08, -2.275891e-08, -2.284115e-08, -2.280144e-08,
  -1.989148e-08, -1.972256e-08, -1.967011e-08, -1.947812e-08, -1.904913e-08, 
    -1.89945e-08, -1.916797e-08, -1.941463e-08, -1.957724e-08, -1.986147e-08, 
    -2.008963e-08, -2.045233e-08, -2.06725e-08, -2.088892e-08, -2.099424e-08,
  -1.996327e-08, -1.992911e-08, -1.985858e-08, -1.980742e-08, -1.979648e-08, 
    -1.972341e-08, -1.964936e-08, -1.971161e-08, -1.983043e-08, 
    -2.003983e-08, -2.026615e-08, -2.04481e-08, -2.068083e-08, -2.081257e-08, 
    -2.094793e-08,
  -1.983252e-08, -1.975402e-08, -1.970295e-08, -1.956656e-08, -1.948217e-08, 
    -1.938649e-08, -1.938258e-08, -1.942776e-08, -1.949338e-08, 
    -1.962537e-08, -1.9756e-08, -1.989744e-08, -2.009241e-08, -2.024458e-08, 
    -2.038555e-08,
  -1.920551e-08, -1.938153e-08, -1.950422e-08, -1.93895e-08, -1.928057e-08, 
    -1.92272e-08, -1.911794e-08, -1.90634e-08, -1.908408e-08, -1.912835e-08, 
    -1.923259e-08, -1.931279e-08, -1.946171e-08, -1.957306e-08, -1.971708e-08,
  -1.767347e-08, -1.830818e-08, -1.855129e-08, -1.868856e-08, -1.87192e-08, 
    -1.877689e-08, -1.873163e-08, -1.877564e-08, -1.869911e-08, -1.87199e-08, 
    -1.872032e-08, -1.877487e-08, -1.88262e-08, -1.890009e-08, -1.894709e-08,
  -1.51892e-08, -1.524188e-08, -1.533223e-08, -1.556388e-08, -1.60585e-08, 
    -1.675119e-08, -1.777802e-08, -1.930272e-08, -2.067683e-08, 
    -2.195937e-08, -2.329208e-08, -2.422541e-08, -2.509318e-08, -2.57824e-08, 
    -2.649412e-08,
  -1.482469e-08, -1.488252e-08, -1.505903e-08, -1.523016e-08, -1.55088e-08, 
    -1.594512e-08, -1.653145e-08, -1.736258e-08, -1.861337e-08, 
    -1.977404e-08, -2.104338e-08, -2.211786e-08, -2.321261e-08, 
    -2.407132e-08, -2.490547e-08,
  -1.463767e-08, -1.463043e-08, -1.469053e-08, -1.487048e-08, -1.504877e-08, 
    -1.530456e-08, -1.577221e-08, -1.625399e-08, -1.688628e-08, 
    -1.781699e-08, -1.889916e-08, -1.990444e-08, -2.101846e-08, -2.20522e-08, 
    -2.299916e-08,
  -1.444155e-08, -1.445586e-08, -1.452983e-08, -1.464327e-08, -1.482682e-08, 
    -1.501544e-08, -1.525477e-08, -1.557139e-08, -1.591308e-08, 
    -1.643591e-08, -1.701175e-08, -1.79181e-08, -1.866089e-08, -1.957185e-08, 
    -2.03623e-08,
  -1.432067e-08, -1.432749e-08, -1.43281e-08, -1.440278e-08, -1.448549e-08, 
    -1.468591e-08, -1.48727e-08, -1.512293e-08, -1.52945e-08, -1.556997e-08, 
    -1.593046e-08, -1.641915e-08, -1.702031e-08, -1.762423e-08, -1.820425e-08,
  -1.41222e-08, -1.423394e-08, -1.428145e-08, -1.42986e-08, -1.430021e-08, 
    -1.433458e-08, -1.439645e-08, -1.453679e-08, -1.466794e-08, 
    -1.481092e-08, -1.499896e-08, -1.519253e-08, -1.552442e-08, 
    -1.590681e-08, -1.634372e-08,
  -1.394579e-08, -1.409363e-08, -1.433542e-08, -1.442524e-08, -1.453086e-08, 
    -1.452698e-08, -1.444396e-08, -1.430325e-08, -1.4201e-08, -1.410743e-08, 
    -1.412627e-08, -1.413441e-08, -1.421997e-08, -1.432191e-08, -1.450707e-08,
  -1.446796e-08, -1.467849e-08, -1.485335e-08, -1.489279e-08, -1.494525e-08, 
    -1.496201e-08, -1.499778e-08, -1.497294e-08, -1.487945e-08, 
    -1.468141e-08, -1.450769e-08, -1.43774e-08, -1.427733e-08, -1.421723e-08, 
    -1.422779e-08,
  -1.360602e-08, -1.462573e-08, -1.54796e-08, -1.602355e-08, -1.634364e-08, 
    -1.644432e-08, -1.646446e-08, -1.644276e-08, -1.644301e-08, 
    -1.646501e-08, -1.646488e-08, -1.642156e-08, -1.636402e-08, 
    -1.628479e-08, -1.622972e-08,
  -1.284453e-08, -1.377544e-08, -1.454275e-08, -1.539567e-08, -1.605264e-08, 
    -1.660277e-08, -1.7011e-08, -1.736871e-08, -1.76071e-08, -1.777952e-08, 
    -1.788921e-08, -1.80131e-08, -1.81083e-08, -1.822624e-08, -1.831583e-08,
  -2.118721e-08, -2.116053e-08, -2.096571e-08, -2.086678e-08, -2.069889e-08, 
    -2.063388e-08, -2.071952e-08, -2.073192e-08, -2.12074e-08, -2.143738e-08, 
    -2.076166e-08, -1.993102e-08, -1.96093e-08, -1.978859e-08, -2.063451e-08,
  -2.144239e-08, -2.140684e-08, -2.140828e-08, -2.130566e-08, -2.119111e-08, 
    -2.102474e-08, -2.084216e-08, -2.065154e-08, -2.052213e-08, 
    -2.041128e-08, -1.971559e-08, -1.905261e-08, -1.878257e-08, 
    -1.910759e-08, -1.96277e-08,
  -2.12321e-08, -2.133073e-08, -2.131804e-08, -2.126972e-08, -2.112937e-08, 
    -2.095728e-08, -2.075623e-08, -2.054576e-08, -2.008079e-08, 
    -1.937469e-08, -1.872691e-08, -1.835846e-08, -1.832796e-08, 
    -1.854323e-08, -1.888598e-08,
  -2.040042e-08, -2.076701e-08, -2.101335e-08, -2.116639e-08, -2.114541e-08, 
    -2.09614e-08, -2.045355e-08, -1.970969e-08, -1.902093e-08, -1.845855e-08, 
    -1.814739e-08, -1.811221e-08, -1.816593e-08, -1.81826e-08, -1.832457e-08,
  -1.921618e-08, -1.94173e-08, -1.970489e-08, -1.989487e-08, -1.983059e-08, 
    -1.947813e-08, -1.90385e-08, -1.863291e-08, -1.821303e-08, -1.79548e-08, 
    -1.788932e-08, -1.783759e-08, -1.782971e-08, -1.783931e-08, -1.783503e-08,
  -1.847964e-08, -1.851709e-08, -1.858748e-08, -1.863757e-08, -1.85154e-08, 
    -1.832637e-08, -1.798697e-08, -1.777867e-08, -1.768443e-08, 
    -1.762964e-08, -1.758477e-08, -1.750654e-08, -1.742035e-08, 
    -1.732136e-08, -1.724692e-08,
  -1.801736e-08, -1.799183e-08, -1.79801e-08, -1.794625e-08, -1.781467e-08, 
    -1.770516e-08, -1.75783e-08, -1.751705e-08, -1.745162e-08, -1.739394e-08, 
    -1.730066e-08, -1.720328e-08, -1.708457e-08, -1.700183e-08, -1.689535e-08,
  -1.751513e-08, -1.751095e-08, -1.751888e-08, -1.751831e-08, -1.749458e-08, 
    -1.746637e-08, -1.736591e-08, -1.73093e-08, -1.725825e-08, -1.723798e-08, 
    -1.714806e-08, -1.703595e-08, -1.688938e-08, -1.678964e-08, -1.668773e-08,
  -1.678478e-08, -1.681673e-08, -1.685027e-08, -1.691077e-08, -1.697074e-08, 
    -1.701613e-08, -1.701476e-08, -1.698608e-08, -1.695167e-08, -1.6897e-08, 
    -1.682954e-08, -1.674576e-08, -1.66453e-08, -1.655302e-08, -1.645559e-08,
  -1.574281e-08, -1.580808e-08, -1.587029e-08, -1.596735e-08, -1.608734e-08, 
    -1.622445e-08, -1.633425e-08, -1.638199e-08, -1.640888e-08, 
    -1.643451e-08, -1.643477e-08, -1.637448e-08, -1.628672e-08, 
    -1.616126e-08, -1.606867e-08,
  -1.591809e-08, -1.588172e-08, -1.641111e-08, -1.738737e-08, -1.777066e-08, 
    -1.763039e-08, -1.752873e-08, -1.780363e-08, -1.826841e-08, -1.91558e-08, 
    -2.124171e-08, -2.324786e-08, -2.465228e-08, -2.493351e-08, -2.432312e-08,
  -1.604669e-08, -1.599981e-08, -1.595974e-08, -1.630646e-08, -1.698331e-08, 
    -1.749224e-08, -1.76726e-08, -1.789517e-08, -1.822199e-08, -1.901981e-08, 
    -2.077959e-08, -2.245131e-08, -2.386811e-08, -2.455423e-08, -2.442669e-08,
  -1.619898e-08, -1.619872e-08, -1.623012e-08, -1.632826e-08, -1.658432e-08, 
    -1.71413e-08, -1.751783e-08, -1.777068e-08, -1.822845e-08, -1.910606e-08, 
    -2.027836e-08, -2.146781e-08, -2.229434e-08, -2.289543e-08, -2.320612e-08,
  -1.665869e-08, -1.645708e-08, -1.645415e-08, -1.648286e-08, -1.674759e-08, 
    -1.702458e-08, -1.764529e-08, -1.838388e-08, -1.904523e-08, 
    -1.961812e-08, -2.011194e-08, -2.054853e-08, -2.118995e-08, 
    -2.176063e-08, -2.229515e-08,
  -1.698239e-08, -1.684618e-08, -1.681287e-08, -1.693393e-08, -1.725133e-08, 
    -1.782343e-08, -1.824885e-08, -1.87123e-08, -1.90253e-08, -1.945793e-08, 
    -1.964166e-08, -1.989793e-08, -2.028016e-08, -2.07867e-08, -2.141725e-08,
  -1.71423e-08, -1.730704e-08, -1.724204e-08, -1.722135e-08, -1.741502e-08, 
    -1.778596e-08, -1.822217e-08, -1.856347e-08, -1.871896e-08, 
    -1.886844e-08, -1.914977e-08, -1.944535e-08, -1.985665e-08, 
    -2.023951e-08, -2.072163e-08,
  -1.655517e-08, -1.698082e-08, -1.707829e-08, -1.71932e-08, -1.714626e-08, 
    -1.739361e-08, -1.753147e-08, -1.771303e-08, -1.79523e-08, -1.827962e-08, 
    -1.861942e-08, -1.904185e-08, -1.943234e-08, -1.984915e-08, -2.029362e-08,
  -1.604904e-08, -1.611718e-08, -1.657706e-08, -1.684685e-08, -1.706005e-08, 
    -1.709417e-08, -1.730957e-08, -1.730019e-08, -1.733821e-08, 
    -1.748844e-08, -1.789394e-08, -1.839076e-08, -1.90278e-08, -1.952951e-08, 
    -1.998347e-08,
  -1.682139e-08, -1.623195e-08, -1.590288e-08, -1.620652e-08, -1.652887e-08, 
    -1.688309e-08, -1.710821e-08, -1.754661e-08, -1.771894e-08, 
    -1.774418e-08, -1.771761e-08, -1.787463e-08, -1.818402e-08, 
    -1.862321e-08, -1.900582e-08,
  -1.811499e-08, -1.765118e-08, -1.705739e-08, -1.646463e-08, -1.649211e-08, 
    -1.665057e-08, -1.683652e-08, -1.729424e-08, -1.762971e-08, 
    -1.811987e-08, -1.836111e-08, -1.849605e-08, -1.851012e-08, 
    -1.849349e-08, -1.851194e-08,
  -1.68359e-08, -1.696736e-08, -1.70755e-08, -1.709699e-08, -1.709906e-08, 
    -1.711073e-08, -1.704029e-08, -1.708706e-08, -1.731622e-08, 
    -1.762857e-08, -1.823518e-08, -1.89149e-08, -1.970444e-08, -2.036465e-08, 
    -2.057247e-08,
  -1.696294e-08, -1.702916e-08, -1.706533e-08, -1.708401e-08, -1.706466e-08, 
    -1.704239e-08, -1.70332e-08, -1.693688e-08, -1.694598e-08, -1.712431e-08, 
    -1.747447e-08, -1.79874e-08, -1.880673e-08, -1.967055e-08, -2.023695e-08,
  -1.709767e-08, -1.711898e-08, -1.71496e-08, -1.714582e-08, -1.711022e-08, 
    -1.70607e-08, -1.7019e-08, -1.695985e-08, -1.684209e-08, -1.683592e-08, 
    -1.696515e-08, -1.72476e-08, -1.764615e-08, -1.852411e-08, -1.94891e-08,
  -1.720415e-08, -1.723942e-08, -1.725348e-08, -1.723272e-08, -1.719238e-08, 
    -1.707809e-08, -1.700499e-08, -1.690766e-08, -1.686556e-08, 
    -1.671823e-08, -1.672125e-08, -1.684111e-08, -1.700044e-08, 
    -1.734466e-08, -1.813422e-08,
  -1.700952e-08, -1.727598e-08, -1.741993e-08, -1.742054e-08, -1.735945e-08, 
    -1.722181e-08, -1.711311e-08, -1.696312e-08, -1.686464e-08, 
    -1.676177e-08, -1.65779e-08, -1.659693e-08, -1.671318e-08, -1.679246e-08, 
    -1.711562e-08,
  -1.670787e-08, -1.700758e-08, -1.733165e-08, -1.750132e-08, -1.747292e-08, 
    -1.742811e-08, -1.723007e-08, -1.716837e-08, -1.695732e-08, 
    -1.684391e-08, -1.666718e-08, -1.649118e-08, -1.654714e-08, 
    -1.659645e-08, -1.669647e-08,
  -1.65492e-08, -1.672346e-08, -1.703032e-08, -1.738709e-08, -1.750055e-08, 
    -1.754127e-08, -1.73934e-08, -1.728796e-08, -1.71285e-08, -1.689558e-08, 
    -1.669234e-08, -1.65337e-08, -1.639552e-08, -1.644396e-08, -1.649002e-08,
  -1.63737e-08, -1.649958e-08, -1.673055e-08, -1.708238e-08, -1.739716e-08, 
    -1.748168e-08, -1.748374e-08, -1.738795e-08, -1.728981e-08, 
    -1.710564e-08, -1.676546e-08, -1.6508e-08, -1.625421e-08, -1.618788e-08, 
    -1.624882e-08,
  -1.613183e-08, -1.63026e-08, -1.653307e-08, -1.68345e-08, -1.720594e-08, 
    -1.744433e-08, -1.748533e-08, -1.743909e-08, -1.739484e-08, 
    -1.734548e-08, -1.72592e-08, -1.694537e-08, -1.664462e-08, -1.630366e-08, 
    -1.616234e-08,
  -1.59033e-08, -1.598253e-08, -1.62179e-08, -1.649133e-08, -1.690948e-08, 
    -1.722746e-08, -1.740321e-08, -1.737969e-08, -1.732751e-08, 
    -1.722587e-08, -1.722352e-08, -1.715827e-08, -1.710879e-08, 
    -1.702122e-08, -1.692426e-08,
  -1.975599e-08, -1.984472e-08, -1.990098e-08, -2.062595e-08, -2.015e-08, 
    -1.927924e-08, -1.822117e-08, -1.76583e-08, -1.734726e-08, -1.72442e-08, 
    -1.723399e-08, -1.722274e-08, -1.730741e-08, -1.740508e-08, -1.754336e-08,
  -1.928917e-08, -1.955267e-08, -1.94401e-08, -1.950576e-08, -1.988311e-08, 
    -1.918592e-08, -1.849057e-08, -1.77613e-08, -1.739063e-08, -1.715836e-08, 
    -1.716099e-08, -1.708015e-08, -1.707302e-08, -1.710467e-08, -1.724064e-08,
  -1.886554e-08, -1.900047e-08, -1.909113e-08, -1.896445e-08, -1.929389e-08, 
    -1.92661e-08, -1.867136e-08, -1.801891e-08, -1.755099e-08, -1.718165e-08, 
    -1.710084e-08, -1.703277e-08, -1.697457e-08, -1.695535e-08, -1.697477e-08,
  -1.90331e-08, -1.877998e-08, -1.879311e-08, -1.882297e-08, -1.865842e-08, 
    -1.901581e-08, -1.877688e-08, -1.82425e-08, -1.775681e-08, -1.734762e-08, 
    -1.718088e-08, -1.70752e-08, -1.700885e-08, -1.694191e-08, -1.690979e-08,
  -1.93001e-08, -1.888785e-08, -1.867892e-08, -1.863244e-08, -1.858302e-08, 
    -1.858842e-08, -1.871357e-08, -1.843804e-08, -1.799798e-08, -1.76356e-08, 
    -1.736117e-08, -1.72579e-08, -1.711234e-08, -1.700435e-08, -1.690858e-08,
  -1.955884e-08, -1.90853e-08, -1.871485e-08, -1.846596e-08, -1.829207e-08, 
    -1.820312e-08, -1.828699e-08, -1.831878e-08, -1.806473e-08, 
    -1.778332e-08, -1.752909e-08, -1.744751e-08, -1.736004e-08, 
    -1.721144e-08, -1.707876e-08,
  -1.945936e-08, -1.926544e-08, -1.882658e-08, -1.845035e-08, -1.79838e-08, 
    -1.7875e-08, -1.781186e-08, -1.796501e-08, -1.799833e-08, -1.780169e-08, 
    -1.766822e-08, -1.761469e-08, -1.755957e-08, -1.744283e-08, -1.727951e-08,
  -1.947457e-08, -1.931232e-08, -1.90434e-08, -1.858148e-08, -1.805649e-08, 
    -1.765206e-08, -1.748055e-08, -1.747683e-08, -1.755724e-08, 
    -1.753566e-08, -1.763627e-08, -1.772306e-08, -1.772766e-08, 
    -1.764593e-08, -1.748031e-08,
  -1.932928e-08, -1.944195e-08, -1.922318e-08, -1.889029e-08, -1.835553e-08, 
    -1.780286e-08, -1.738148e-08, -1.714256e-08, -1.708397e-08, 
    -1.722153e-08, -1.741938e-08, -1.761855e-08, -1.774609e-08, 
    -1.776294e-08, -1.764353e-08,
  -1.869586e-08, -1.909916e-08, -1.920722e-08, -1.916041e-08, -1.895573e-08, 
    -1.837503e-08, -1.787695e-08, -1.727022e-08, -1.702663e-08, 
    -1.698651e-08, -1.718251e-08, -1.741367e-08, -1.764756e-08, 
    -1.773727e-08, -1.771395e-08,
  -2.358854e-08, -2.35494e-08, -2.352007e-08, -2.332707e-08, -2.411791e-08, 
    -2.516055e-08, -2.56953e-08, -2.594943e-08, -2.550841e-08, -2.471834e-08, 
    -2.371145e-08, -2.265009e-08, -2.206112e-08, -2.156705e-08, -2.113832e-08,
  -2.307577e-08, -2.341378e-08, -2.332832e-08, -2.310353e-08, -2.354494e-08, 
    -2.448686e-08, -2.534537e-08, -2.570265e-08, -2.565196e-08, 
    -2.458632e-08, -2.362611e-08, -2.261701e-08, -2.180119e-08, 
    -2.088534e-08, -2.045705e-08,
  -2.299921e-08, -2.314135e-08, -2.293214e-08, -2.334878e-08, -2.351593e-08, 
    -2.390693e-08, -2.434188e-08, -2.471885e-08, -2.463359e-08, 
    -2.387049e-08, -2.283418e-08, -2.195844e-08, -2.130461e-08, -2.0671e-08, 
    -2.027674e-08,
  -2.332436e-08, -2.360421e-08, -2.355355e-08, -2.348565e-08, -2.355513e-08, 
    -2.383106e-08, -2.3923e-08, -2.408438e-08, -2.361048e-08, -2.272208e-08, 
    -2.181684e-08, -2.124354e-08, -2.08198e-08, -2.0547e-08, -2.026775e-08,
  -2.458638e-08, -2.438688e-08, -2.411875e-08, -2.420849e-08, -2.438933e-08, 
    -2.459882e-08, -2.459317e-08, -2.430276e-08, -2.372773e-08, -2.2938e-08, 
    -2.198845e-08, -2.133069e-08, -2.089648e-08, -2.067141e-08, -2.040519e-08,
  -2.469667e-08, -2.464574e-08, -2.44605e-08, -2.377761e-08, -2.365932e-08, 
    -2.345709e-08, -2.372017e-08, -2.386197e-08, -2.35896e-08, -2.280771e-08, 
    -2.16858e-08, -2.089949e-08, -2.044199e-08, -2.027398e-08, -2.013547e-08,
  -2.448169e-08, -2.421713e-08, -2.370741e-08, -2.327823e-08, -2.307079e-08, 
    -2.345318e-08, -2.337046e-08, -2.301371e-08, -2.302507e-08, 
    -2.242082e-08, -2.130069e-08, -2.045181e-08, -2.007496e-08, 
    -1.987835e-08, -1.9779e-08,
  -2.482502e-08, -2.437485e-08, -2.402803e-08, -2.376581e-08, -2.333265e-08, 
    -2.285967e-08, -2.274185e-08, -2.287371e-08, -2.244979e-08, 
    -2.189589e-08, -2.104557e-08, -2.041308e-08, -1.995601e-08, -1.98108e-08, 
    -1.966753e-08,
  -2.516156e-08, -2.478799e-08, -2.416964e-08, -2.35218e-08, -2.291462e-08, 
    -2.267485e-08, -2.259514e-08, -2.285456e-08, -2.245215e-08, 
    -2.163171e-08, -2.099866e-08, -2.015234e-08, -1.979822e-08, 
    -1.946363e-08, -1.935175e-08,
  -2.519242e-08, -2.48707e-08, -2.381898e-08, -2.295952e-08, -2.215135e-08, 
    -2.217143e-08, -2.208254e-08, -2.208347e-08, -2.195858e-08, 
    -2.151429e-08, -2.093795e-08, -2.034916e-08, -1.981277e-08, 
    -1.949228e-08, -1.923609e-08,
  -1.92186e-08, -1.955478e-08, -1.974485e-08, -2.022981e-08, -2.065135e-08, 
    -2.105163e-08, -2.133238e-08, -2.17385e-08, -2.233625e-08, -2.304355e-08, 
    -2.352331e-08, -2.407833e-08, -2.436698e-08, -2.454314e-08, -2.454931e-08,
  -1.950787e-08, -1.998368e-08, -2.046458e-08, -2.067797e-08, -2.127679e-08, 
    -2.170629e-08, -2.190149e-08, -2.218685e-08, -2.262557e-08, 
    -2.317919e-08, -2.375224e-08, -2.428496e-08, -2.463096e-08, 
    -2.470775e-08, -2.455305e-08,
  -1.985567e-08, -2.021211e-08, -2.09147e-08, -2.124608e-08, -2.183923e-08, 
    -2.239756e-08, -2.248553e-08, -2.260169e-08, -2.263088e-08, 
    -2.326957e-08, -2.424655e-08, -2.472902e-08, -2.46588e-08, -2.438889e-08, 
    -2.414492e-08,
  -2.037936e-08, -2.071213e-08, -2.129618e-08, -2.190881e-08, -2.26005e-08, 
    -2.288455e-08, -2.299564e-08, -2.325221e-08, -2.362366e-08, 
    -2.428575e-08, -2.475024e-08, -2.488524e-08, -2.477644e-08, 
    -2.422763e-08, -2.367598e-08,
  -2.089748e-08, -2.138334e-08, -2.235746e-08, -2.27236e-08, -2.293425e-08, 
    -2.345595e-08, -2.384479e-08, -2.428091e-08, -2.446695e-08, 
    -2.450224e-08, -2.466625e-08, -2.43367e-08, -2.386439e-08, -2.326464e-08, 
    -2.282308e-08,
  -2.177795e-08, -2.296283e-08, -2.368785e-08, -2.343129e-08, -2.39248e-08, 
    -2.45289e-08, -2.491935e-08, -2.550819e-08, -2.584178e-08, -2.60487e-08, 
    -2.560262e-08, -2.470154e-08, -2.379736e-08, -2.327049e-08, -2.290131e-08,
  -2.313744e-08, -2.461421e-08, -2.462922e-08, -2.44773e-08, -2.518251e-08, 
    -2.587065e-08, -2.623581e-08, -2.638568e-08, -2.634026e-08, 
    -2.578439e-08, -2.610999e-08, -2.638074e-08, -2.571293e-08, 
    -2.503507e-08, -2.437427e-08,
  -2.410691e-08, -2.569173e-08, -2.604927e-08, -2.596775e-08, -2.657981e-08, 
    -2.6698e-08, -2.580097e-08, -2.643438e-08, -2.639059e-08, -2.725629e-08, 
    -2.69467e-08, -2.672189e-08, -2.596839e-08, -2.498221e-08, -2.430124e-08,
  -2.564198e-08, -2.715677e-08, -2.743436e-08, -2.7064e-08, -2.697208e-08, 
    -2.686206e-08, -2.593343e-08, -2.556066e-08, -2.537209e-08, 
    -2.520552e-08, -2.493689e-08, -2.473865e-08, -2.418329e-08, 
    -2.348625e-08, -2.283922e-08,
  -2.619562e-08, -2.746143e-08, -2.788882e-08, -2.756427e-08, -2.724801e-08, 
    -2.702089e-08, -2.705406e-08, -2.684012e-08, -2.608533e-08, 
    -2.557563e-08, -2.508967e-08, -2.414311e-08, -2.329377e-08, 
    -2.292503e-08, -2.231388e-08,
  -8.152685e-09, -8.402323e-09, -9.104325e-09, -9.876412e-09, -1.068815e-08, 
    -1.171556e-08, -1.234436e-08, -1.280306e-08, -1.38646e-08, -1.457988e-08, 
    -1.55192e-08, -1.720828e-08, -1.800713e-08, -1.819284e-08, -1.870602e-08,
  -8.206281e-09, -8.392566e-09, -8.805733e-09, -9.629744e-09, -1.036386e-08, 
    -1.128166e-08, -1.198143e-08, -1.233209e-08, -1.280468e-08, 
    -1.363886e-08, -1.432139e-08, -1.541691e-08, -1.670805e-08, 
    -1.747662e-08, -1.809729e-08,
  -8.394387e-09, -8.572486e-09, -8.860265e-09, -9.504787e-09, -1.013575e-08, 
    -1.088496e-08, -1.184792e-08, -1.225351e-08, -1.259798e-08, 
    -1.305559e-08, -1.370071e-08, -1.446169e-08, -1.557701e-08, 
    -1.660976e-08, -1.735227e-08,
  -8.912393e-09, -8.950294e-09, -9.13071e-09, -9.562251e-09, -1.020687e-08, 
    -1.086222e-08, -1.1783e-08, -1.238822e-08, -1.276033e-08, -1.299272e-08, 
    -1.3516e-08, -1.415161e-08, -1.500768e-08, -1.618667e-08, -1.7214e-08,
  -9.672852e-09, -9.68075e-09, -9.703921e-09, -1.005686e-08, -1.069297e-08, 
    -1.132183e-08, -1.19931e-08, -1.249819e-08, -1.297816e-08, -1.334344e-08, 
    -1.371731e-08, -1.44959e-08, -1.548826e-08, -1.655402e-08, -1.750516e-08,
  -1.042868e-08, -1.053614e-08, -1.061033e-08, -1.07893e-08, -1.122798e-08, 
    -1.169737e-08, -1.226287e-08, -1.289358e-08, -1.350392e-08, 
    -1.412025e-08, -1.490606e-08, -1.579557e-08, -1.667441e-08, 
    -1.746538e-08, -1.810596e-08,
  -1.095927e-08, -1.121833e-08, -1.150272e-08, -1.16786e-08, -1.215969e-08, 
    -1.269503e-08, -1.317016e-08, -1.387079e-08, -1.49365e-08, -1.580627e-08, 
    -1.630282e-08, -1.680344e-08, -1.739606e-08, -1.788329e-08, -1.824516e-08,
  -1.180342e-08, -1.224972e-08, -1.269996e-08, -1.280408e-08, -1.321935e-08, 
    -1.389745e-08, -1.478717e-08, -1.56861e-08, -1.643405e-08, -1.686426e-08, 
    -1.718497e-08, -1.750258e-08, -1.78845e-08, -1.826577e-08, -1.85004e-08,
  -1.292056e-08, -1.356597e-08, -1.394711e-08, -1.45276e-08, -1.524527e-08, 
    -1.595495e-08, -1.658307e-08, -1.694745e-08, -1.735928e-08, -1.76994e-08, 
    -1.794604e-08, -1.830158e-08, -1.884333e-08, -1.927318e-08, -1.953483e-08,
  -1.43212e-08, -1.524149e-08, -1.57672e-08, -1.646794e-08, -1.703176e-08, 
    -1.738683e-08, -1.762174e-08, -1.796674e-08, -1.837036e-08, 
    -1.886922e-08, -1.943297e-08, -2.007959e-08, -2.058508e-08, 
    -2.095945e-08, -2.143447e-08,
  -1.25794e-08, -1.327578e-08, -1.385756e-08, -1.468631e-08, -1.523701e-08, 
    -1.578949e-08, -1.668196e-08, -1.782724e-08, -1.918507e-08, 
    -2.056227e-08, -2.200733e-08, -2.275445e-08, -2.370207e-08, 
    -2.492087e-08, -2.542628e-08,
  -1.136927e-08, -1.203785e-08, -1.271049e-08, -1.33851e-08, -1.417062e-08, 
    -1.464254e-08, -1.524446e-08, -1.591086e-08, -1.699922e-08, 
    -1.803305e-08, -1.952799e-08, -2.090964e-08, -2.182634e-08, 
    -2.267092e-08, -2.376485e-08,
  -1.034144e-08, -1.08507e-08, -1.147517e-08, -1.206764e-08, -1.277374e-08, 
    -1.345962e-08, -1.396462e-08, -1.448129e-08, -1.5078e-08, -1.590253e-08, 
    -1.682424e-08, -1.798936e-08, -1.931038e-08, -2.035359e-08, -2.117434e-08,
  -9.383849e-09, -9.737986e-09, -1.020744e-08, -1.076409e-08, -1.135252e-08, 
    -1.202162e-08, -1.267823e-08, -1.320951e-08, -1.372242e-08, 
    -1.428127e-08, -1.498676e-08, -1.575612e-08, -1.664963e-08, 
    -1.775953e-08, -1.877223e-08,
  -8.617343e-09, -8.812489e-09, -9.106817e-09, -9.513396e-09, -1.003591e-08, 
    -1.061909e-08, -1.124212e-08, -1.18473e-08, -1.238554e-08, -1.292706e-08, 
    -1.347783e-08, -1.412438e-08, -1.47959e-08, -1.553034e-08, -1.641369e-08,
  -8.074431e-09, -8.064887e-09, -8.180575e-09, -8.3862e-09, -8.738478e-09, 
    -9.215444e-09, -9.813768e-09, -1.041255e-08, -1.097713e-08, -1.14988e-08, 
    -1.20185e-08, -1.258518e-08, -1.31792e-08, -1.381782e-08, -1.454102e-08,
  -7.945136e-09, -7.810107e-09, -7.724471e-09, -7.737457e-09, -7.837498e-09, 
    -8.035577e-09, -8.375522e-09, -8.917453e-09, -9.549805e-09, 
    -1.010592e-08, -1.060931e-08, -1.110294e-08, -1.16315e-08, -1.217239e-08, 
    -1.27846e-08,
  -8.235388e-09, -8.038677e-09, -7.853344e-09, -7.68047e-09, -7.60092e-09, 
    -7.579654e-09, -7.606093e-09, -7.762357e-09, -8.148334e-09, 
    -8.684907e-09, -9.304046e-09, -9.820369e-09, -1.030047e-08, 
    -1.076008e-08, -1.129348e-08,
  -8.946856e-09, -8.596135e-09, -8.361162e-09, -8.134592e-09, -7.956625e-09, 
    -7.741371e-09, -7.609371e-09, -7.489575e-09, -7.527087e-09, 
    -7.698223e-09, -8.04453e-09, -8.564077e-09, -9.17762e-09, -9.651966e-09, 
    -1.009913e-08,
  -9.761093e-09, -9.336527e-09, -8.977343e-09, -8.682768e-09, -8.471146e-09, 
    -8.294324e-09, -8.05789e-09, -7.781151e-09, -7.608929e-09, -7.593269e-09, 
    -7.658235e-09, -7.827782e-09, -8.172724e-09, -8.706033e-09, -9.262982e-09,
  -1.443196e-08, -1.47839e-08, -1.511948e-08, -1.545522e-08, -1.576653e-08, 
    -1.598661e-08, -1.635131e-08, -1.67838e-08, -1.745092e-08, -1.808421e-08, 
    -1.952507e-08, -2.06886e-08, -2.16423e-08, -2.239366e-08, -2.361792e-08,
  -1.413177e-08, -1.436675e-08, -1.473518e-08, -1.509406e-08, -1.54438e-08, 
    -1.57392e-08, -1.611455e-08, -1.648994e-08, -1.702192e-08, -1.748589e-08, 
    -1.821758e-08, -1.949822e-08, -2.080096e-08, -2.158978e-08, -2.262593e-08,
  -1.385118e-08, -1.405045e-08, -1.434184e-08, -1.469056e-08, -1.508343e-08, 
    -1.540744e-08, -1.572886e-08, -1.615192e-08, -1.658668e-08, -1.71383e-08, 
    -1.760621e-08, -1.818981e-08, -1.946291e-08, -2.075735e-08, -2.15635e-08,
  -1.348623e-08, -1.370294e-08, -1.393238e-08, -1.419015e-08, -1.453786e-08, 
    -1.494378e-08, -1.531087e-08, -1.570272e-08, -1.612184e-08, 
    -1.663067e-08, -1.717734e-08, -1.768716e-08, -1.826637e-08, 
    -1.944556e-08, -2.072048e-08,
  -1.318722e-08, -1.341173e-08, -1.358968e-08, -1.379718e-08, -1.405546e-08, 
    -1.440267e-08, -1.476754e-08, -1.517755e-08, -1.557021e-08, 
    -1.603863e-08, -1.656879e-08, -1.713777e-08, -1.765163e-08, 
    -1.828593e-08, -1.93733e-08,
  -1.289476e-08, -1.30425e-08, -1.329489e-08, -1.347616e-08, -1.367546e-08, 
    -1.394474e-08, -1.426277e-08, -1.463004e-08, -1.500966e-08, 
    -1.540807e-08, -1.588618e-08, -1.642693e-08, -1.703655e-08, 
    -1.757179e-08, -1.824779e-08,
  -1.252813e-08, -1.262095e-08, -1.276361e-08, -1.299364e-08, -1.321246e-08, 
    -1.344233e-08, -1.375507e-08, -1.407732e-08, -1.444614e-08, 
    -1.480541e-08, -1.521716e-08, -1.563398e-08, -1.617389e-08, 
    -1.676832e-08, -1.739733e-08,
  -1.228518e-08, -1.226618e-08, -1.231563e-08, -1.240098e-08, -1.258727e-08, 
    -1.277232e-08, -1.30385e-08, -1.332226e-08, -1.368227e-08, -1.407512e-08, 
    -1.448812e-08, -1.49015e-08, -1.534127e-08, -1.583812e-08, -1.638238e-08,
  -1.19533e-08, -1.191805e-08, -1.190632e-08, -1.186669e-08, -1.195761e-08, 
    -1.207557e-08, -1.224872e-08, -1.245331e-08, -1.272035e-08, 
    -1.303179e-08, -1.341727e-08, -1.383524e-08, -1.428363e-08, 
    -1.477328e-08, -1.532188e-08,
  -1.17649e-08, -1.168235e-08, -1.166605e-08, -1.161904e-08, -1.161666e-08, 
    -1.163422e-08, -1.166678e-08, -1.172828e-08, -1.186284e-08, 
    -1.205068e-08, -1.226821e-08, -1.254441e-08, -1.286882e-08, 
    -1.325667e-08, -1.372445e-08,
  -1.575559e-08, -1.631815e-08, -1.689046e-08, -1.729896e-08, -1.780392e-08, 
    -1.825305e-08, -1.877983e-08, -1.930424e-08, -1.968242e-08, 
    -2.047812e-08, -2.074493e-08, -2.060386e-08, -2.134937e-08, 
    -2.310024e-08, -2.468399e-08,
  -1.528632e-08, -1.581208e-08, -1.639523e-08, -1.680492e-08, -1.720754e-08, 
    -1.767155e-08, -1.82333e-08, -1.870912e-08, -1.922834e-08, -1.963346e-08, 
    -2.035015e-08, -2.05386e-08, -2.061654e-08, -2.13173e-08, -2.286243e-08,
  -1.484164e-08, -1.535795e-08, -1.587093e-08, -1.640459e-08, -1.673293e-08, 
    -1.712033e-08, -1.758495e-08, -1.811396e-08, -1.863776e-08, 
    -1.902328e-08, -1.95132e-08, -2.005577e-08, -2.031046e-08, -2.047844e-08, 
    -2.111893e-08,
  -1.431153e-08, -1.487475e-08, -1.535656e-08, -1.592735e-08, -1.634898e-08, 
    -1.66906e-08, -1.704151e-08, -1.744777e-08, -1.795641e-08, -1.845696e-08, 
    -1.882016e-08, -1.932058e-08, -1.981589e-08, -2.007938e-08, -2.024244e-08,
  -1.377324e-08, -1.445042e-08, -1.491588e-08, -1.544512e-08, -1.593653e-08, 
    -1.629988e-08, -1.661903e-08, -1.696452e-08, -1.732064e-08, 
    -1.773957e-08, -1.817684e-08, -1.851913e-08, -1.905263e-08, 
    -1.953118e-08, -1.983472e-08,
  -1.325778e-08, -1.401254e-08, -1.453966e-08, -1.498954e-08, -1.547873e-08, 
    -1.58318e-08, -1.616847e-08, -1.649609e-08, -1.680409e-08, -1.716558e-08, 
    -1.753859e-08, -1.786888e-08, -1.819834e-08, -1.870916e-08, -1.916121e-08,
  -1.28107e-08, -1.356983e-08, -1.419831e-08, -1.4674e-08, -1.507466e-08, 
    -1.541406e-08, -1.569279e-08, -1.604045e-08, -1.634728e-08, 
    -1.659879e-08, -1.694009e-08, -1.728199e-08, -1.755998e-08, -1.78517e-08, 
    -1.828323e-08,
  -1.244817e-08, -1.314398e-08, -1.385171e-08, -1.43594e-08, -1.470265e-08, 
    -1.500305e-08, -1.525988e-08, -1.554013e-08, -1.584612e-08, 
    -1.613311e-08, -1.637603e-08, -1.664708e-08, -1.693205e-08, 
    -1.715111e-08, -1.743848e-08,
  -1.214e-08, -1.274947e-08, -1.348448e-08, -1.403036e-08, -1.434023e-08, 
    -1.45688e-08, -1.482153e-08, -1.50763e-08, -1.532548e-08, -1.554514e-08, 
    -1.580255e-08, -1.602936e-08, -1.627706e-08, -1.652209e-08, -1.673662e-08,
  -1.188828e-08, -1.245945e-08, -1.313877e-08, -1.366163e-08, -1.3911e-08, 
    -1.409165e-08, -1.435565e-08, -1.457624e-08, -1.484108e-08, 
    -1.503653e-08, -1.523245e-08, -1.540415e-08, -1.560248e-08, 
    -1.581439e-08, -1.602314e-08,
  -1.417002e-08, -1.487871e-08, -1.542844e-08, -1.59353e-08, -1.634776e-08, 
    -1.663913e-08, -1.686179e-08, -1.704308e-08, -1.732562e-08, 
    -1.755663e-08, -1.77585e-08, -1.796235e-08, -1.830558e-08, -1.883651e-08, 
    -1.927052e-08,
  -1.281906e-08, -1.379219e-08, -1.457244e-08, -1.524479e-08, -1.58259e-08, 
    -1.618541e-08, -1.653994e-08, -1.672426e-08, -1.692632e-08, -1.72207e-08, 
    -1.754693e-08, -1.779486e-08, -1.809078e-08, -1.854579e-08, -1.9019e-08,
  -1.150444e-08, -1.245702e-08, -1.336333e-08, -1.422603e-08, -1.509875e-08, 
    -1.564501e-08, -1.605112e-08, -1.644195e-08, -1.668351e-08, 
    -1.692639e-08, -1.72846e-08, -1.762831e-08, -1.790493e-08, -1.829947e-08, 
    -1.878479e-08,
  -1.00092e-08, -1.110573e-08, -1.21309e-08, -1.302142e-08, -1.403855e-08, 
    -1.495295e-08, -1.546389e-08, -1.604766e-08, -1.633868e-08, 
    -1.667452e-08, -1.697193e-08, -1.738056e-08, -1.771843e-08, 
    -1.809872e-08, -1.850704e-08,
  -8.803825e-09, -9.779806e-09, -1.093293e-08, -1.190348e-08, -1.287236e-08, 
    -1.398652e-08, -1.473629e-08, -1.551868e-08, -1.598737e-08, -1.63877e-08, 
    -1.671319e-08, -1.709652e-08, -1.752417e-08, -1.802353e-08, -1.835595e-08,
  -7.625858e-09, -8.544392e-09, -9.641059e-09, -1.076369e-08, -1.182365e-08, 
    -1.294997e-08, -1.387168e-08, -1.479559e-08, -1.553094e-08, 
    -1.603913e-08, -1.642972e-08, -1.679309e-08, -1.717708e-08, 
    -1.782203e-08, -1.831316e-08,
  -6.531353e-09, -7.382424e-09, -8.398493e-09, -9.581639e-09, -1.066515e-08, 
    -1.196295e-08, -1.297493e-08, -1.394444e-08, -1.489597e-08, 
    -1.558869e-08, -1.616514e-08, -1.660043e-08, -1.691132e-08, 
    -1.746207e-08, -1.803048e-08,
  -5.625339e-09, -6.401025e-09, -7.297231e-09, -8.448321e-09, -9.598212e-09, 
    -1.08033e-08, -1.210941e-08, -1.309165e-08, -1.413913e-08, -1.496233e-08, 
    -1.56893e-08, -1.632897e-08, -1.674496e-08, -1.71809e-08, -1.761386e-08,
  -4.951497e-09, -5.554001e-09, -6.43715e-09, -7.461976e-09, -8.585822e-09, 
    -9.776898e-09, -1.108284e-08, -1.236091e-08, -1.338832e-08, 
    -1.434734e-08, -1.51069e-08, -1.591603e-08, -1.649672e-08, -1.692092e-08, 
    -1.734886e-08,
  -4.522738e-09, -4.999195e-09, -5.73339e-09, -6.703886e-09, -7.773358e-09, 
    -8.861893e-09, -1.003191e-08, -1.136201e-08, -1.261219e-08, -1.36452e-08, 
    -1.450974e-08, -1.533295e-08, -1.616708e-08, -1.671259e-08, -1.710075e-08,
  -2.197496e-08, -2.238946e-08, -2.268417e-08, -2.261778e-08, -2.242787e-08, 
    -2.206932e-08, -2.175767e-08, -2.154017e-08, -2.136675e-08, 
    -2.117952e-08, -2.101448e-08, -2.089026e-08, -2.078642e-08, 
    -2.063128e-08, -2.04492e-08,
  -2.10586e-08, -2.137221e-08, -2.178531e-08, -2.223542e-08, -2.251321e-08, 
    -2.233801e-08, -2.194223e-08, -2.149665e-08, -2.106714e-08, -2.07601e-08, 
    -2.058411e-08, -2.051654e-08, -2.052734e-08, -2.03883e-08, -2.022615e-08,
  -1.97286e-08, -2.033635e-08, -2.07854e-08, -2.097261e-08, -2.147624e-08, 
    -2.181266e-08, -2.170349e-08, -2.145008e-08, -2.094428e-08, 
    -2.052388e-08, -2.027082e-08, -2.012741e-08, -2.003751e-08, -1.98837e-08, 
    -1.968132e-08,
  -1.847222e-08, -1.92598e-08, -1.977154e-08, -2.022525e-08, -2.050414e-08, 
    -2.097766e-08, -2.11629e-08, -2.117816e-08, -2.082887e-08, -2.052196e-08, 
    -2.018603e-08, -1.984811e-08, -1.957696e-08, -1.929391e-08, -1.903252e-08,
  -1.719045e-08, -1.768714e-08, -1.836374e-08, -1.896383e-08, -1.942876e-08, 
    -1.979536e-08, -2.016006e-08, -2.05245e-08, -2.043959e-08, -2.018805e-08, 
    -1.992244e-08, -1.959878e-08, -1.922608e-08, -1.885083e-08, -1.854151e-08,
  -1.656304e-08, -1.66263e-08, -1.704623e-08, -1.762272e-08, -1.81179e-08, 
    -1.853818e-08, -1.900261e-08, -1.925393e-08, -1.965614e-08, 
    -1.967788e-08, -1.965848e-08, -1.952074e-08, -1.91828e-08, -1.870823e-08, 
    -1.815792e-08,
  -1.604438e-08, -1.629215e-08, -1.627257e-08, -1.654271e-08, -1.695447e-08, 
    -1.718712e-08, -1.745599e-08, -1.783195e-08, -1.828639e-08, 
    -1.877001e-08, -1.886739e-08, -1.89271e-08, -1.861246e-08, -1.82756e-08, 
    -1.78501e-08,
  -1.467542e-08, -1.543475e-08, -1.591664e-08, -1.588727e-08, -1.609491e-08, 
    -1.620596e-08, -1.650687e-08, -1.660054e-08, -1.686612e-08, 
    -1.733117e-08, -1.768673e-08, -1.787217e-08, -1.785899e-08, 
    -1.775991e-08, -1.749172e-08,
  -1.198293e-08, -1.328663e-08, -1.436599e-08, -1.50011e-08, -1.524392e-08, 
    -1.545289e-08, -1.544336e-08, -1.571713e-08, -1.587697e-08, 
    -1.604775e-08, -1.628965e-08, -1.651836e-08, -1.695277e-08, 
    -1.721752e-08, -1.731563e-08,
  -1.004112e-08, -1.085298e-08, -1.185643e-08, -1.299083e-08, -1.387355e-08, 
    -1.444874e-08, -1.475445e-08, -1.492765e-08, -1.50831e-08, -1.521023e-08, 
    -1.532338e-08, -1.557004e-08, -1.601587e-08, -1.662647e-08, -1.680843e-08,
  -1.651684e-08, -1.671274e-08, -1.691235e-08, -1.727668e-08, -1.781783e-08, 
    -1.808263e-08, -1.844577e-08, -1.880083e-08, -1.917386e-08, 
    -1.954107e-08, -1.977972e-08, -1.979383e-08, -1.966633e-08, 
    -1.937291e-08, -1.948583e-08,
  -1.594942e-08, -1.637219e-08, -1.667092e-08, -1.699902e-08, -1.731382e-08, 
    -1.788869e-08, -1.836423e-08, -1.877185e-08, -1.911571e-08, 
    -1.944667e-08, -1.982058e-08, -1.998517e-08, -2.010353e-08, 
    -2.008507e-08, -1.989578e-08,
  -1.537508e-08, -1.573788e-08, -1.618228e-08, -1.664439e-08, -1.709635e-08, 
    -1.751698e-08, -1.807998e-08, -1.880382e-08, -1.917308e-08, 
    -1.935402e-08, -1.955002e-08, -1.988421e-08, -2.0157e-08, -2.036534e-08, 
    -2.05338e-08,
  -1.499204e-08, -1.529633e-08, -1.56304e-08, -1.613871e-08, -1.660568e-08, 
    -1.71754e-08, -1.778439e-08, -1.838406e-08, -1.916063e-08, -1.941376e-08, 
    -1.954922e-08, -1.973045e-08, -2.012572e-08, -2.054711e-08, -2.082093e-08,
  -1.481883e-08, -1.49939e-08, -1.517665e-08, -1.562664e-08, -1.61949e-08, 
    -1.66286e-08, -1.740412e-08, -1.801242e-08, -1.873493e-08, -1.948591e-08, 
    -1.976228e-08, -1.999117e-08, -2.025883e-08, -2.057081e-08, -2.093118e-08,
  -1.466043e-08, -1.487332e-08, -1.499801e-08, -1.518769e-08, -1.564166e-08, 
    -1.624027e-08, -1.68423e-08, -1.767645e-08, -1.827335e-08, -1.900707e-08, 
    -1.974136e-08, -2.01806e-08, -2.058874e-08, -2.0922e-08, -2.109394e-08,
  -1.40553e-08, -1.459606e-08, -1.489856e-08, -1.504274e-08, -1.5269e-08, 
    -1.57637e-08, -1.614507e-08, -1.708204e-08, -1.783704e-08, -1.843795e-08, 
    -1.933997e-08, -2.000768e-08, -2.068338e-08, -2.095327e-08, -2.128886e-08,
  -1.385292e-08, -1.404154e-08, -1.450094e-08, -1.48968e-08, -1.512308e-08, 
    -1.540922e-08, -1.58388e-08, -1.624551e-08, -1.721043e-08, -1.777488e-08, 
    -1.87139e-08, -1.95523e-08, -2.039621e-08, -2.081752e-08, -2.116407e-08,
  -1.37497e-08, -1.396336e-08, -1.41347e-08, -1.454943e-08, -1.492001e-08, 
    -1.520151e-08, -1.551479e-08, -1.576058e-08, -1.637964e-08, 
    -1.695119e-08, -1.763085e-08, -1.848779e-08, -1.938741e-08, 
    -2.015533e-08, -2.087634e-08,
  -1.337041e-08, -1.365817e-08, -1.393833e-08, -1.418127e-08, -1.463357e-08, 
    -1.492085e-08, -1.531108e-08, -1.554787e-08, -1.580565e-08, 
    -1.624608e-08, -1.676059e-08, -1.730708e-08, -1.811901e-08, 
    -1.878521e-08, -1.960051e-08,
  -1.414139e-08, -1.425829e-08, -1.447531e-08, -1.464143e-08, -1.480979e-08, 
    -1.495674e-08, -1.513269e-08, -1.536862e-08, -1.582348e-08, 
    -1.620118e-08, -1.658291e-08, -1.69668e-08, -1.72311e-08, -1.737837e-08, 
    -1.73901e-08,
  -1.387279e-08, -1.395738e-08, -1.410179e-08, -1.432332e-08, -1.442911e-08, 
    -1.460738e-08, -1.481457e-08, -1.505969e-08, -1.541885e-08, -1.58892e-08, 
    -1.632179e-08, -1.674236e-08, -1.719711e-08, -1.751407e-08, -1.775594e-08,
  -1.364503e-08, -1.367104e-08, -1.376136e-08, -1.397601e-08, -1.415073e-08, 
    -1.430259e-08, -1.448246e-08, -1.472535e-08, -1.502775e-08, 
    -1.542614e-08, -1.595632e-08, -1.643476e-08, -1.694157e-08, 
    -1.748379e-08, -1.785475e-08,
  -1.343386e-08, -1.344754e-08, -1.349356e-08, -1.357736e-08, -1.375967e-08, 
    -1.399229e-08, -1.419081e-08, -1.440452e-08, -1.467842e-08, -1.50157e-08, 
    -1.544028e-08, -1.598014e-08, -1.654432e-08, -1.720549e-08, -1.774843e-08,
  -1.309367e-08, -1.323647e-08, -1.333905e-08, -1.338806e-08, -1.3465e-08, 
    -1.361321e-08, -1.384546e-08, -1.408311e-08, -1.430557e-08, -1.4641e-08, 
    -1.500445e-08, -1.550385e-08, -1.602581e-08, -1.671717e-08, -1.738926e-08,
  -1.250189e-08, -1.279356e-08, -1.2973e-08, -1.315904e-08, -1.326355e-08, 
    -1.33786e-08, -1.349976e-08, -1.371735e-08, -1.39248e-08, -1.418605e-08, 
    -1.45351e-08, -1.501605e-08, -1.552852e-08, -1.615146e-08, -1.682732e-08,
  -1.203086e-08, -1.229351e-08, -1.252964e-08, -1.271373e-08, -1.293029e-08, 
    -1.308634e-08, -1.325948e-08, -1.337323e-08, -1.356959e-08, 
    -1.377868e-08, -1.406625e-08, -1.449615e-08, -1.500106e-08, 
    -1.558792e-08, -1.621691e-08,
  -1.150558e-08, -1.172621e-08, -1.204289e-08, -1.22745e-08, -1.247731e-08, 
    -1.270099e-08, -1.290751e-08, -1.308786e-08, -1.322158e-08, 
    -1.342078e-08, -1.363003e-08, -1.401714e-08, -1.445726e-08, 
    -1.502652e-08, -1.56112e-08,
  -1.092794e-08, -1.11987e-08, -1.14529e-08, -1.176329e-08, -1.204e-08, 
    -1.226015e-08, -1.250068e-08, -1.270755e-08, -1.288291e-08, 
    -1.306611e-08, -1.326839e-08, -1.355115e-08, -1.392243e-08, 
    -1.442928e-08, -1.498989e-08,
  -1.022276e-08, -1.057063e-08, -1.087102e-08, -1.114912e-08, -1.148168e-08, 
    -1.180307e-08, -1.206805e-08, -1.233803e-08, -1.253728e-08, 
    -1.270081e-08, -1.292081e-08, -1.317134e-08, -1.348026e-08, 
    -1.388968e-08, -1.437559e-08,
  -2.625724e-08, -2.5606e-08, -2.476865e-08, -2.449285e-08, -2.444854e-08, 
    -2.444644e-08, -2.433236e-08, -2.383847e-08, -2.251992e-08, 
    -2.138967e-08, -2.036706e-08, -1.935934e-08, -1.905112e-08, 
    -1.867109e-08, -1.838394e-08,
  -2.560177e-08, -2.557003e-08, -2.483695e-08, -2.435177e-08, -2.414674e-08, 
    -2.393343e-08, -2.364394e-08, -2.291764e-08, -2.154504e-08, -2.07222e-08, 
    -2.005936e-08, -1.923853e-08, -1.853854e-08, -1.812909e-08, -1.784843e-08,
  -2.507146e-08, -2.513359e-08, -2.469603e-08, -2.395203e-08, -2.386241e-08, 
    -2.38315e-08, -2.34597e-08, -2.235209e-08, -2.117072e-08, -2.031332e-08, 
    -1.962488e-08, -1.868919e-08, -1.802762e-08, -1.769961e-08, -1.715469e-08,
  -2.410754e-08, -2.42691e-08, -2.399416e-08, -2.343443e-08, -2.340187e-08, 
    -2.345567e-08, -2.273289e-08, -2.149305e-08, -2.05738e-08, -1.980554e-08, 
    -1.904679e-08, -1.799783e-08, -1.734366e-08, -1.675214e-08, -1.633028e-08,
  -2.340938e-08, -2.339748e-08, -2.302691e-08, -2.257344e-08, -2.260231e-08, 
    -2.248954e-08, -2.195421e-08, -2.077972e-08, -2.007945e-08, 
    -1.937576e-08, -1.849784e-08, -1.764781e-08, -1.687432e-08, -1.62748e-08, 
    -1.617067e-08,
  -2.291291e-08, -2.280768e-08, -2.241893e-08, -2.209197e-08, -2.212583e-08, 
    -2.206795e-08, -2.159895e-08, -2.040494e-08, -1.973977e-08, 
    -1.884033e-08, -1.79959e-08, -1.729924e-08, -1.651589e-08, -1.603931e-08, 
    -1.582582e-08,
  -2.225996e-08, -2.205062e-08, -2.169394e-08, -2.138894e-08, -2.15489e-08, 
    -2.155849e-08, -2.10074e-08, -1.986095e-08, -1.920459e-08, -1.832944e-08, 
    -1.763146e-08, -1.693749e-08, -1.621568e-08, -1.588662e-08, -1.559275e-08,
  -2.163206e-08, -2.156411e-08, -2.106508e-08, -2.090306e-08, -2.108259e-08, 
    -2.105392e-08, -2.04086e-08, -1.953646e-08, -1.87502e-08, -1.794449e-08, 
    -1.735697e-08, -1.664772e-08, -1.604896e-08, -1.556636e-08, -1.512033e-08,
  -2.08179e-08, -2.086283e-08, -2.069819e-08, -2.063608e-08, -2.081009e-08, 
    -2.069846e-08, -2.01566e-08, -1.935793e-08, -1.849922e-08, -1.77476e-08, 
    -1.712641e-08, -1.638733e-08, -1.5669e-08, -1.508089e-08, -1.47399e-08,
  -1.996752e-08, -1.993e-08, -2.001802e-08, -2.005445e-08, -2.013305e-08, 
    -2.002918e-08, -1.957778e-08, -1.903373e-08, -1.824271e-08, 
    -1.738627e-08, -1.660936e-08, -1.58323e-08, -1.523615e-08, -1.484078e-08, 
    -1.448863e-08,
  -2.46502e-08, -2.551925e-08, -2.638218e-08, -2.638856e-08, -2.563031e-08, 
    -2.657995e-08, -2.686565e-08, -2.734987e-08, -2.770852e-08, -2.7529e-08, 
    -2.69758e-08, -2.684603e-08, -2.647936e-08, -2.662491e-08, -2.546271e-08,
  -2.443577e-08, -2.5523e-08, -2.650682e-08, -2.669235e-08, -2.594867e-08, 
    -2.644778e-08, -2.595947e-08, -2.611479e-08, -2.646416e-08, -2.65953e-08, 
    -2.592168e-08, -2.603486e-08, -2.673168e-08, -2.76766e-08, -2.610126e-08,
  -2.395959e-08, -2.497696e-08, -2.631152e-08, -2.709366e-08, -2.586372e-08, 
    -2.636473e-08, -2.627535e-08, -2.619918e-08, -2.627915e-08, 
    -2.653571e-08, -2.644436e-08, -2.702565e-08, -2.781923e-08, 
    -2.908618e-08, -2.690732e-08,
  -2.319894e-08, -2.436455e-08, -2.608648e-08, -2.735468e-08, -2.597588e-08, 
    -2.632261e-08, -2.590558e-08, -2.557026e-08, -2.568633e-08, 
    -2.647998e-08, -2.656765e-08, -2.738797e-08, -2.765176e-08, 
    -2.884732e-08, -2.697024e-08,
  -2.224227e-08, -2.365308e-08, -2.5396e-08, -2.721522e-08, -2.617803e-08, 
    -2.611099e-08, -2.627273e-08, -2.599576e-08, -2.604726e-08, 
    -2.662258e-08, -2.738121e-08, -2.810935e-08, -2.757562e-08, 
    -2.873749e-08, -2.739369e-08,
  -2.122661e-08, -2.296027e-08, -2.468712e-08, -2.670287e-08, -2.63276e-08, 
    -2.618279e-08, -2.648775e-08, -2.609055e-08, -2.633453e-08, 
    -2.672409e-08, -2.72564e-08, -2.774111e-08, -2.6968e-08, -2.753624e-08, 
    -2.657064e-08,
  -2.018969e-08, -2.211628e-08, -2.381167e-08, -2.609981e-08, -2.619198e-08, 
    -2.616629e-08, -2.664443e-08, -2.605072e-08, -2.62461e-08, -2.664015e-08, 
    -2.709908e-08, -2.731854e-08, -2.631784e-08, -2.634441e-08, -2.561727e-08,
  -1.909879e-08, -2.113383e-08, -2.298229e-08, -2.538297e-08, -2.581204e-08, 
    -2.619146e-08, -2.675771e-08, -2.653216e-08, -2.657179e-08, -2.67992e-08, 
    -2.685292e-08, -2.651701e-08, -2.581546e-08, -2.502777e-08, -2.391506e-08,
  -1.820253e-08, -1.999011e-08, -2.201584e-08, -2.448381e-08, -2.537063e-08, 
    -2.584176e-08, -2.662988e-08, -2.648594e-08, -2.655665e-08, 
    -2.682005e-08, -2.64064e-08, -2.588794e-08, -2.535966e-08, -2.377419e-08, 
    -2.242026e-08,
  -1.748309e-08, -1.897325e-08, -2.101197e-08, -2.339806e-08, -2.500984e-08, 
    -2.532656e-08, -2.638333e-08, -2.655908e-08, -2.71532e-08, -2.66873e-08, 
    -2.604481e-08, -2.530599e-08, -2.500254e-08, -2.305305e-08, -2.138684e-08,
  -2.205131e-08, -2.219557e-08, -2.184773e-08, -2.163869e-08, -2.152511e-08, 
    -2.125699e-08, -2.177513e-08, -2.20421e-08, -2.332036e-08, -2.618543e-08, 
    -2.599302e-08, -2.604768e-08, -2.614572e-08, -2.911453e-08, -2.952018e-08,
  -2.194309e-08, -2.197428e-08, -2.165329e-08, -2.149752e-08, -2.158022e-08, 
    -2.133899e-08, -2.176576e-08, -2.178338e-08, -2.29551e-08, -2.533693e-08, 
    -2.530408e-08, -2.568162e-08, -2.620177e-08, -2.805119e-08, -2.830936e-08,
  -2.209251e-08, -2.181628e-08, -2.165015e-08, -2.110929e-08, -2.133664e-08, 
    -2.123165e-08, -2.16673e-08, -2.197125e-08, -2.314935e-08, -2.545994e-08, 
    -2.5264e-08, -2.566431e-08, -2.61189e-08, -2.776456e-08, -2.836405e-08,
  -2.137664e-08, -2.146959e-08, -2.166475e-08, -2.125975e-08, -2.126438e-08, 
    -2.13164e-08, -2.148278e-08, -2.194819e-08, -2.280207e-08, -2.459048e-08, 
    -2.493931e-08, -2.56768e-08, -2.659081e-08, -2.782054e-08, -2.80452e-08,
  -1.997605e-08, -2.046439e-08, -2.075312e-08, -2.094914e-08, -2.112863e-08, 
    -2.139256e-08, -2.154252e-08, -2.202334e-08, -2.288143e-08, 
    -2.424783e-08, -2.491143e-08, -2.576014e-08, -2.651619e-08, 
    -2.762625e-08, -2.773296e-08,
  -1.787585e-08, -1.908731e-08, -1.951766e-08, -1.996521e-08, -2.047637e-08, 
    -2.104601e-08, -2.149442e-08, -2.193225e-08, -2.270361e-08, 
    -2.369339e-08, -2.47217e-08, -2.593454e-08, -2.644155e-08, -2.727645e-08, 
    -2.68578e-08,
  -1.592153e-08, -1.72058e-08, -1.80666e-08, -1.874511e-08, -1.946116e-08, 
    -2.039517e-08, -2.105759e-08, -2.177054e-08, -2.231707e-08, 
    -2.334178e-08, -2.452327e-08, -2.611942e-08, -2.61413e-08, -2.664919e-08, 
    -2.587603e-08,
  -1.398756e-08, -1.510613e-08, -1.627405e-08, -1.707564e-08, -1.813581e-08, 
    -1.933947e-08, -2.040844e-08, -2.134467e-08, -2.207535e-08, -2.27976e-08, 
    -2.427515e-08, -2.575731e-08, -2.575107e-08, -2.585921e-08, -2.482577e-08,
  -1.215087e-08, -1.319369e-08, -1.429922e-08, -1.525995e-08, -1.631991e-08, 
    -1.780023e-08, -1.919963e-08, -2.055291e-08, -2.147191e-08, 
    -2.246205e-08, -2.38133e-08, -2.508506e-08, -2.537687e-08, -2.541371e-08, 
    -2.428725e-08,
  -1.067818e-08, -1.150381e-08, -1.252516e-08, -1.358887e-08, -1.46421e-08, 
    -1.595856e-08, -1.759349e-08, -1.916928e-08, -2.069225e-08, 
    -2.164073e-08, -2.293411e-08, -2.442757e-08, -2.476778e-08, 
    -2.497465e-08, -2.422938e-08,
  -2.348506e-08, -2.412e-08, -2.42828e-08, -2.44682e-08, -2.459709e-08, 
    -2.511017e-08, -2.542708e-08, -2.559747e-08, -2.547222e-08, 
    -2.515277e-08, -2.500571e-08, -2.464403e-08, -2.449117e-08, 
    -2.423401e-08, -2.402339e-08,
  -2.248152e-08, -2.330262e-08, -2.392542e-08, -2.425733e-08, -2.448092e-08, 
    -2.48162e-08, -2.510621e-08, -2.531207e-08, -2.526615e-08, -2.517196e-08, 
    -2.487981e-08, -2.469496e-08, -2.447459e-08, -2.427583e-08, -2.40374e-08,
  -2.180941e-08, -2.254479e-08, -2.319374e-08, -2.38314e-08, -2.41644e-08, 
    -2.451778e-08, -2.4703e-08, -2.49063e-08, -2.497825e-08, -2.489666e-08, 
    -2.472187e-08, -2.460986e-08, -2.438731e-08, -2.421332e-08, -2.403898e-08,
  -2.120553e-08, -2.20477e-08, -2.270345e-08, -2.330447e-08, -2.385647e-08, 
    -2.426405e-08, -2.465875e-08, -2.482973e-08, -2.496925e-08, -2.4933e-08, 
    -2.48871e-08, -2.46688e-08, -2.451773e-08, -2.434847e-08, -2.42492e-08,
  -2.071764e-08, -2.134536e-08, -2.20328e-08, -2.264441e-08, -2.320349e-08, 
    -2.37261e-08, -2.419647e-08, -2.458877e-08, -2.487309e-08, -2.503218e-08, 
    -2.507824e-08, -2.490057e-08, -2.470952e-08, -2.450788e-08, -2.431893e-08,
  -2.04036e-08, -2.083973e-08, -2.131856e-08, -2.194445e-08, -2.25101e-08, 
    -2.309225e-08, -2.356909e-08, -2.402524e-08, -2.42762e-08, -2.460304e-08, 
    -2.473593e-08, -2.471393e-08, -2.454454e-08, -2.433958e-08, -2.417635e-08,
  -1.992187e-08, -2.019501e-08, -2.058757e-08, -2.110371e-08, -2.167721e-08, 
    -2.218759e-08, -2.270637e-08, -2.320833e-08, -2.360982e-08, 
    -2.394201e-08, -2.427681e-08, -2.442784e-08, -2.436951e-08, 
    -2.417666e-08, -2.399335e-08,
  -1.982696e-08, -1.981862e-08, -1.997721e-08, -2.038194e-08, -2.082426e-08, 
    -2.137183e-08, -2.18246e-08, -2.229081e-08, -2.269853e-08, -2.301512e-08, 
    -2.326795e-08, -2.350345e-08, -2.363373e-08, -2.357366e-08, -2.336409e-08,
  -1.954248e-08, -1.975171e-08, -1.979209e-08, -1.984008e-08, -2.011905e-08, 
    -2.047974e-08, -2.102056e-08, -2.147567e-08, -2.200147e-08, 
    -2.239899e-08, -2.260835e-08, -2.26857e-08, -2.274011e-08, -2.278829e-08, 
    -2.266346e-08,
  -1.846674e-08, -1.92238e-08, -1.959883e-08, -1.979348e-08, -1.977834e-08, 
    -1.984917e-08, -2.006368e-08, -2.047836e-08, -2.097722e-08, 
    -2.144149e-08, -2.174825e-08, -2.190389e-08, -2.198245e-08, 
    -2.189612e-08, -2.180939e-08,
  -2.007879e-08, -2.053974e-08, -2.104762e-08, -2.150692e-08, -2.178496e-08, 
    -2.194163e-08, -2.205761e-08, -2.196702e-08, -2.19798e-08, -2.212732e-08, 
    -2.236466e-08, -2.264754e-08, -2.286052e-08, -2.298614e-08, -2.311125e-08,
  -1.946215e-08, -2.004061e-08, -2.054544e-08, -2.108413e-08, -2.14776e-08, 
    -2.174844e-08, -2.19615e-08, -2.200031e-08, -2.201451e-08, -2.205515e-08, 
    -2.224431e-08, -2.240934e-08, -2.259886e-08, -2.26769e-08, -2.281588e-08,
  -1.886087e-08, -1.941022e-08, -1.996899e-08, -2.045586e-08, -2.093737e-08, 
    -2.128879e-08, -2.154393e-08, -2.165241e-08, -2.177935e-08, 
    -2.193749e-08, -2.218975e-08, -2.241031e-08, -2.256115e-08, 
    -2.259851e-08, -2.264528e-08,
  -1.826161e-08, -1.878181e-08, -1.926978e-08, -1.986222e-08, -2.03058e-08, 
    -2.071534e-08, -2.099337e-08, -2.112514e-08, -2.118071e-08, 
    -2.137322e-08, -2.170774e-08, -2.206117e-08, -2.232909e-08, -2.24767e-08, 
    -2.251411e-08,
  -1.676613e-08, -1.804385e-08, -1.866436e-08, -1.914926e-08, -1.970575e-08, 
    -2.01227e-08, -2.049519e-08, -2.065148e-08, -2.066986e-08, -2.077553e-08, 
    -2.104736e-08, -2.145301e-08, -2.181089e-08, -2.212116e-08, -2.231692e-08,
  -1.545096e-08, -1.661884e-08, -1.778507e-08, -1.848522e-08, -1.893732e-08, 
    -1.944632e-08, -1.987714e-08, -2.020636e-08, -2.033595e-08, -2.04079e-08, 
    -2.055533e-08, -2.082127e-08, -2.117804e-08, -2.154132e-08, -2.182545e-08,
  -1.448979e-08, -1.523799e-08, -1.634946e-08, -1.754814e-08, -1.834051e-08, 
    -1.875782e-08, -1.919467e-08, -1.954206e-08, -1.980061e-08, 
    -2.001286e-08, -2.017052e-08, -2.03529e-08, -2.060781e-08, -2.095275e-08, 
    -2.132418e-08,
  -1.356649e-08, -1.428752e-08, -1.497006e-08, -1.606801e-08, -1.724809e-08, 
    -1.80726e-08, -1.860536e-08, -1.899925e-08, -1.920725e-08, -1.946894e-08, 
    -1.975578e-08, -1.995115e-08, -2.021166e-08, -2.050208e-08, -2.090816e-08,
  -1.274582e-08, -1.347656e-08, -1.416104e-08, -1.484697e-08, -1.590269e-08, 
    -1.687667e-08, -1.766347e-08, -1.827054e-08, -1.868587e-08, 
    -1.896162e-08, -1.928217e-08, -1.952238e-08, -1.984455e-08, 
    -2.017941e-08, -2.050564e-08,
  -1.207878e-08, -1.257274e-08, -1.329789e-08, -1.394778e-08, -1.473719e-08, 
    -1.575942e-08, -1.667734e-08, -1.73684e-08, -1.791974e-08, -1.844146e-08, 
    -1.88617e-08, -1.915034e-08, -1.938859e-08, -1.962889e-08, -1.991161e-08,
  -1.47672e-08, -1.50989e-08, -1.550087e-08, -1.5898e-08, -1.630741e-08, 
    -1.647157e-08, -1.678456e-08, -1.722607e-08, -1.769658e-08, 
    -1.790835e-08, -1.802669e-08, -1.810964e-08, -1.831532e-08, 
    -1.857276e-08, -1.879946e-08,
  -1.38965e-08, -1.444911e-08, -1.494702e-08, -1.530203e-08, -1.563176e-08, 
    -1.586288e-08, -1.605909e-08, -1.648155e-08, -1.688359e-08, 
    -1.710025e-08, -1.726464e-08, -1.738217e-08, -1.753085e-08, -1.77558e-08, 
    -1.805352e-08,
  -1.329209e-08, -1.38591e-08, -1.442153e-08, -1.485299e-08, -1.513289e-08, 
    -1.537855e-08, -1.557027e-08, -1.586294e-08, -1.623303e-08, 
    -1.644112e-08, -1.658056e-08, -1.670312e-08, -1.680065e-08, 
    -1.698545e-08, -1.719793e-08,
  -1.27739e-08, -1.329107e-08, -1.383442e-08, -1.427255e-08, -1.459766e-08, 
    -1.486361e-08, -1.511114e-08, -1.538849e-08, -1.573559e-08, 
    -1.600439e-08, -1.612339e-08, -1.621477e-08, -1.629671e-08, 
    -1.640221e-08, -1.651002e-08,
  -1.246471e-08, -1.28323e-08, -1.331082e-08, -1.372489e-08, -1.409929e-08, 
    -1.437059e-08, -1.462768e-08, -1.493507e-08, -1.526832e-08, 
    -1.556448e-08, -1.573982e-08, -1.584326e-08, -1.590193e-08, 
    -1.600185e-08, -1.606879e-08,
  -1.200361e-08, -1.245975e-08, -1.285462e-08, -1.326983e-08, -1.366283e-08, 
    -1.399503e-08, -1.423095e-08, -1.454192e-08, -1.487985e-08, 
    -1.516722e-08, -1.53645e-08, -1.549512e-08, -1.558578e-08, -1.56699e-08, 
    -1.579265e-08,
  -1.123548e-08, -1.184204e-08, -1.231711e-08, -1.275999e-08, -1.317868e-08, 
    -1.357093e-08, -1.389223e-08, -1.417712e-08, -1.453971e-08, 
    -1.484472e-08, -1.508812e-08, -1.521528e-08, -1.528453e-08, 
    -1.534219e-08, -1.549106e-08,
  -1.058505e-08, -1.116441e-08, -1.173389e-08, -1.22452e-08, -1.270916e-08, 
    -1.310213e-08, -1.34617e-08, -1.376731e-08, -1.406919e-08, -1.440436e-08, 
    -1.4703e-08, -1.497299e-08, -1.515091e-08, -1.523646e-08, -1.53325e-08,
  -9.788492e-09, -1.04352e-08, -1.105136e-08, -1.164317e-08, -1.22039e-08, 
    -1.269301e-08, -1.309525e-08, -1.33974e-08, -1.368603e-08, -1.394705e-08, 
    -1.420617e-08, -1.443258e-08, -1.467104e-08, -1.488558e-08, -1.508499e-08,
  -9.196153e-09, -9.683959e-09, -1.029199e-08, -1.089053e-08, -1.15029e-08, 
    -1.207704e-08, -1.261843e-08, -1.303293e-08, -1.33707e-08, -1.360918e-08, 
    -1.38092e-08, -1.406076e-08, -1.430733e-08, -1.452691e-08, -1.469581e-08,
  -1.36477e-08, -1.356484e-08, -1.353624e-08, -1.345547e-08, -1.33283e-08, 
    -1.309349e-08, -1.29044e-08, -1.263541e-08, -1.235399e-08, -1.217752e-08, 
    -1.209419e-08, -1.210876e-08, -1.227694e-08, -1.249433e-08, -1.275047e-08,
  -1.252425e-08, -1.2479e-08, -1.234491e-08, -1.209117e-08, -1.182548e-08, 
    -1.151399e-08, -1.129248e-08, -1.107755e-08, -1.105435e-08, -1.10452e-08, 
    -1.109906e-08, -1.115211e-08, -1.13188e-08, -1.147784e-08, -1.178548e-08,
  -1.165627e-08, -1.150479e-08, -1.125773e-08, -1.094049e-08, -1.063955e-08, 
    -1.038195e-08, -1.019994e-08, -1.008044e-08, -1.002809e-08, 
    -1.005403e-08, -1.013453e-08, -1.028804e-08, -1.046811e-08, -1.0674e-08, 
    -1.089631e-08,
  -1.08338e-08, -1.061249e-08, -1.037364e-08, -1.009761e-08, -9.874375e-09, 
    -9.719506e-09, -9.617668e-09, -9.563549e-09, -9.556045e-09, 
    -9.615472e-09, -9.730285e-09, -9.88655e-09, -1.006612e-08, -1.026632e-08, 
    -1.050282e-08,
  -1.033526e-08, -1.014479e-08, -9.939797e-09, -9.728899e-09, -9.540365e-09, 
    -9.411133e-09, -9.311621e-09, -9.276469e-09, -9.289679e-09, 
    -9.366184e-09, -9.492304e-09, -9.656488e-09, -9.856081e-09, 
    -1.010185e-08, -1.038025e-08,
  -9.886182e-09, -9.766578e-09, -9.620019e-09, -9.480628e-09, -9.320686e-09, 
    -9.209542e-09, -9.156243e-09, -9.139459e-09, -9.176901e-09, 
    -9.269935e-09, -9.400261e-09, -9.572317e-09, -9.822034e-09, 
    -1.011466e-08, -1.041108e-08,
  -9.558048e-09, -9.47032e-09, -9.381618e-09, -9.263748e-09, -9.130577e-09, 
    -9.057797e-09, -9.050264e-09, -9.093376e-09, -9.171901e-09, 
    -9.305557e-09, -9.466053e-09, -9.672801e-09, -9.949024e-09, 
    -1.025045e-08, -1.050596e-08,
  -9.337321e-09, -9.236405e-09, -9.15191e-09, -9.04859e-09, -8.933833e-09, 
    -8.886027e-09, -8.877675e-09, -8.95721e-09, -9.092773e-09, -9.300468e-09, 
    -9.503852e-09, -9.788229e-09, -1.010761e-08, -1.040895e-08, -1.064837e-08,
  -9.405523e-09, -9.230411e-09, -9.112441e-09, -9.007601e-09, -8.893664e-09, 
    -8.8487e-09, -8.861252e-09, -8.943374e-09, -9.092664e-09, -9.32686e-09, 
    -9.553213e-09, -9.853343e-09, -1.019771e-08, -1.049138e-08, -1.073653e-08,
  -9.59393e-09, -9.409201e-09, -9.278338e-09, -9.164217e-09, -9.045141e-09, 
    -9.012104e-09, -9.013026e-09, -9.111851e-09, -9.217084e-09, -9.40093e-09, 
    -9.610683e-09, -9.875676e-09, -1.019279e-08, -1.043635e-08, -1.066997e-08,
  -1.828308e-08, -1.848507e-08, -1.86095e-08, -1.877118e-08, -1.88577e-08, 
    -1.896092e-08, -1.894921e-08, -1.88297e-08, -1.856704e-08, -1.819183e-08, 
    -1.761941e-08, -1.69348e-08, -1.622568e-08, -1.554065e-08, -1.493078e-08,
  -1.750522e-08, -1.771857e-08, -1.7933e-08, -1.807784e-08, -1.81374e-08, 
    -1.811498e-08, -1.798851e-08, -1.777017e-08, -1.746176e-08, 
    -1.705891e-08, -1.6497e-08, -1.584788e-08, -1.518396e-08, -1.455248e-08, 
    -1.399727e-08,
  -1.670318e-08, -1.694705e-08, -1.717273e-08, -1.729279e-08, -1.732281e-08, 
    -1.723721e-08, -1.708347e-08, -1.686158e-08, -1.65465e-08, -1.611492e-08, 
    -1.553118e-08, -1.487203e-08, -1.422056e-08, -1.361116e-08, -1.307789e-08,
  -1.591091e-08, -1.613363e-08, -1.636908e-08, -1.648134e-08, -1.649105e-08, 
    -1.640411e-08, -1.626662e-08, -1.606795e-08, -1.577251e-08, 
    -1.531095e-08, -1.471366e-08, -1.40591e-08, -1.340679e-08, -1.27947e-08, 
    -1.224076e-08,
  -1.516865e-08, -1.543957e-08, -1.560928e-08, -1.573158e-08, -1.570494e-08, 
    -1.563313e-08, -1.548353e-08, -1.528076e-08, -1.498218e-08, 
    -1.452374e-08, -1.393461e-08, -1.329227e-08, -1.264693e-08, 
    -1.206693e-08, -1.155652e-08,
  -1.445871e-08, -1.472e-08, -1.489297e-08, -1.499979e-08, -1.496909e-08, 
    -1.489088e-08, -1.473555e-08, -1.455117e-08, -1.42898e-08, -1.384244e-08, 
    -1.329422e-08, -1.266996e-08, -1.205605e-08, -1.152129e-08, -1.106751e-08,
  -1.367873e-08, -1.397597e-08, -1.419133e-08, -1.432746e-08, -1.435008e-08, 
    -1.429439e-08, -1.415232e-08, -1.397478e-08, -1.369536e-08, 
    -1.324626e-08, -1.268693e-08, -1.208537e-08, -1.149928e-08, -1.10029e-08, 
    -1.057596e-08,
  -1.280975e-08, -1.310647e-08, -1.337837e-08, -1.356438e-08, -1.365402e-08, 
    -1.362824e-08, -1.355289e-08, -1.338669e-08, -1.307225e-08, 
    -1.259705e-08, -1.206134e-08, -1.149118e-08, -1.097592e-08, -1.05248e-08, 
    -1.015895e-08,
  -1.179086e-08, -1.209557e-08, -1.24161e-08, -1.263427e-08, -1.277792e-08, 
    -1.28105e-08, -1.281503e-08, -1.27042e-08, -1.24117e-08, -1.19707e-08, 
    -1.149378e-08, -1.096976e-08, -1.05082e-08, -1.008778e-08, -9.764788e-09,
  -1.065142e-08, -1.10909e-08, -1.137675e-08, -1.161918e-08, -1.175498e-08, 
    -1.180646e-08, -1.183054e-08, -1.181751e-08, -1.156347e-08, 
    -1.124035e-08, -1.080466e-08, -1.039832e-08, -9.945304e-09, 
    -9.628055e-09, -9.309941e-09,
  -2.060612e-08, -2.01778e-08, -1.979416e-08, -1.939532e-08, -1.90113e-08, 
    -1.860375e-08, -1.817539e-08, -1.77675e-08, -1.739168e-08, -1.702475e-08, 
    -1.678694e-08, -1.6626e-08, -1.639647e-08, -1.611126e-08, -1.582393e-08,
  -1.982389e-08, -1.939112e-08, -1.895874e-08, -1.849959e-08, -1.801416e-08, 
    -1.754388e-08, -1.704015e-08, -1.655141e-08, -1.607891e-08, 
    -1.572677e-08, -1.555983e-08, -1.542593e-08, -1.521661e-08, 
    -1.496276e-08, -1.465879e-08,
  -1.868111e-08, -1.830493e-08, -1.787108e-08, -1.738492e-08, -1.688333e-08, 
    -1.638754e-08, -1.586521e-08, -1.534865e-08, -1.492675e-08, 
    -1.468594e-08, -1.453039e-08, -1.446106e-08, -1.431953e-08, 
    -1.404102e-08, -1.374449e-08,
  -1.708523e-08, -1.67566e-08, -1.640842e-08, -1.597516e-08, -1.553344e-08, 
    -1.50966e-08, -1.464283e-08, -1.422867e-08, -1.388412e-08, -1.363387e-08, 
    -1.351893e-08, -1.347655e-08, -1.330634e-08, -1.307283e-08, -1.288362e-08,
  -1.554895e-08, -1.524346e-08, -1.497942e-08, -1.467156e-08, -1.430929e-08, 
    -1.394885e-08, -1.354829e-08, -1.313221e-08, -1.276921e-08, 
    -1.257554e-08, -1.251384e-08, -1.241793e-08, -1.232744e-08, 
    -1.219752e-08, -1.210277e-08,
  -1.427729e-08, -1.405178e-08, -1.383151e-08, -1.353539e-08, -1.322995e-08, 
    -1.287718e-08, -1.244865e-08, -1.200204e-08, -1.164957e-08, 
    -1.150376e-08, -1.144022e-08, -1.141885e-08, -1.139449e-08, 
    -1.136204e-08, -1.129807e-08,
  -1.292186e-08, -1.279345e-08, -1.261521e-08, -1.235207e-08, -1.203624e-08, 
    -1.166634e-08, -1.123988e-08, -1.082944e-08, -1.052235e-08, 
    -1.044203e-08, -1.045609e-08, -1.049254e-08, -1.050932e-08, 
    -1.051124e-08, -1.04932e-08,
  -1.147577e-08, -1.135397e-08, -1.117812e-08, -1.091889e-08, -1.05976e-08, 
    -1.028574e-08, -9.898828e-09, -9.533609e-09, -9.308946e-09, 
    -9.330934e-09, -9.417341e-09, -9.52082e-09, -9.636767e-09, -9.695949e-09, 
    -9.789793e-09,
  -1.013109e-08, -1.001977e-08, -9.792485e-09, -9.477027e-09, -9.140244e-09, 
    -8.803833e-09, -8.507154e-09, -8.242823e-09, -8.222099e-09, 
    -8.390833e-09, -8.533151e-09, -8.715916e-09, -8.893163e-09, 
    -9.008735e-09, -9.160633e-09,
  -9.019036e-09, -8.851708e-09, -8.584455e-09, -8.287006e-09, -7.962506e-09, 
    -7.664259e-09, -7.435198e-09, -7.284521e-09, -7.353254e-09, 
    -7.527793e-09, -7.681157e-09, -7.8998e-09, -8.120492e-09, -8.304041e-09, 
    -8.499224e-09,
  -2.496162e-08, -2.486001e-08, -2.460479e-08, -2.428387e-08, -2.406558e-08, 
    -2.40626e-08, -2.404675e-08, -2.370982e-08, -2.345533e-08, -2.342912e-08, 
    -2.343939e-08, -2.329334e-08, -2.302396e-08, -2.305308e-08, -2.294655e-08,
  -2.474322e-08, -2.450453e-08, -2.428679e-08, -2.392857e-08, -2.372459e-08, 
    -2.347957e-08, -2.327707e-08, -2.300514e-08, -2.254064e-08, 
    -2.229773e-08, -2.218496e-08, -2.204473e-08, -2.200848e-08, 
    -2.210135e-08, -2.208248e-08,
  -2.400956e-08, -2.38968e-08, -2.400695e-08, -2.378168e-08, -2.347128e-08, 
    -2.33344e-08, -2.303658e-08, -2.275379e-08, -2.237054e-08, -2.196717e-08, 
    -2.159829e-08, -2.153345e-08, -2.14515e-08, -2.140174e-08, -2.103504e-08,
  -2.363422e-08, -2.336895e-08, -2.36143e-08, -2.367873e-08, -2.315946e-08, 
    -2.292519e-08, -2.266014e-08, -2.231117e-08, -2.198591e-08, 
    -2.154196e-08, -2.128237e-08, -2.113744e-08, -2.078561e-08, 
    -2.054602e-08, -1.992613e-08,
  -2.339587e-08, -2.313625e-08, -2.342268e-08, -2.356566e-08, -2.319162e-08, 
    -2.273836e-08, -2.238511e-08, -2.203909e-08, -2.168705e-08, 
    -2.121547e-08, -2.093724e-08, -2.052785e-08, -2.013681e-08, 
    -1.955213e-08, -1.877977e-08,
  -2.264614e-08, -2.24222e-08, -2.275975e-08, -2.296508e-08, -2.274622e-08, 
    -2.23974e-08, -2.208034e-08, -2.163855e-08, -2.11858e-08, -2.068244e-08, 
    -2.012918e-08, -1.947526e-08, -1.885468e-08, -1.809847e-08, -1.731759e-08,
  -2.154349e-08, -2.147176e-08, -2.179811e-08, -2.208312e-08, -2.212369e-08, 
    -2.183552e-08, -2.148915e-08, -2.091668e-08, -2.029665e-08, -1.96617e-08, 
    -1.894633e-08, -1.821355e-08, -1.743348e-08, -1.660479e-08, -1.586181e-08,
  -2.046881e-08, -2.056325e-08, -2.073625e-08, -2.079755e-08, -2.085915e-08, 
    -2.063467e-08, -2.018591e-08, -1.964335e-08, -1.896096e-08, -1.80587e-08, 
    -1.71716e-08, -1.639095e-08, -1.556955e-08, -1.486231e-08, -1.435482e-08,
  -1.883413e-08, -1.896839e-08, -1.918714e-08, -1.914728e-08, -1.89212e-08, 
    -1.849826e-08, -1.801657e-08, -1.734935e-08, -1.662893e-08, 
    -1.594596e-08, -1.529133e-08, -1.469851e-08, -1.405069e-08, 
    -1.355732e-08, -1.299458e-08,
  -1.700262e-08, -1.72272e-08, -1.731391e-08, -1.721712e-08, -1.698209e-08, 
    -1.662309e-08, -1.617762e-08, -1.56993e-08, -1.514389e-08, -1.453437e-08, 
    -1.396212e-08, -1.345413e-08, -1.293553e-08, -1.244139e-08, -1.185456e-08,
  -1.555857e-08, -1.568078e-08, -1.653601e-08, -1.752838e-08, -1.82028e-08, 
    -1.861685e-08, -1.905481e-08, -1.981568e-08, -2.067008e-08, 
    -2.121943e-08, -2.167395e-08, -2.194315e-08, -2.218775e-08, 
    -2.219082e-08, -2.223476e-08,
  -1.471053e-08, -1.547576e-08, -1.589691e-08, -1.690173e-08, -1.758213e-08, 
    -1.839343e-08, -1.880681e-08, -1.918542e-08, -1.976389e-08, 
    -2.016762e-08, -2.047782e-08, -2.075238e-08, -2.09889e-08, -2.110827e-08, 
    -2.120708e-08,
  -1.381729e-08, -1.486654e-08, -1.555895e-08, -1.638831e-08, -1.711014e-08, 
    -1.751142e-08, -1.837033e-08, -1.885116e-08, -1.925363e-08, 
    -1.975091e-08, -2.003632e-08, -2.013526e-08, -2.021229e-08, 
    -2.038038e-08, -2.065465e-08,
  -1.270323e-08, -1.397698e-08, -1.502006e-08, -1.577702e-08, -1.650807e-08, 
    -1.694112e-08, -1.757119e-08, -1.833169e-08, -1.884644e-08, 
    -1.933952e-08, -1.960903e-08, -1.981272e-08, -2.004524e-08, 
    -2.026731e-08, -2.071425e-08,
  -1.203732e-08, -1.2964e-08, -1.42473e-08, -1.520123e-08, -1.588251e-08, 
    -1.646786e-08, -1.683629e-08, -1.738761e-08, -1.805553e-08, 
    -1.873677e-08, -1.911916e-08, -1.952236e-08, -1.981688e-08, 
    -2.015619e-08, -2.061869e-08,
  -1.164192e-08, -1.223716e-08, -1.337856e-08, -1.458638e-08, -1.544406e-08, 
    -1.611927e-08, -1.65533e-08, -1.696558e-08, -1.744284e-08, -1.804645e-08, 
    -1.86157e-08, -1.916916e-08, -1.959565e-08, -2.000466e-08, -2.03679e-08,
  -1.14462e-08, -1.202535e-08, -1.284655e-08, -1.39729e-08, -1.488646e-08, 
    -1.555403e-08, -1.601028e-08, -1.64048e-08, -1.682259e-08, -1.728622e-08, 
    -1.777043e-08, -1.829524e-08, -1.871513e-08, -1.903522e-08, -1.918169e-08,
  -1.12897e-08, -1.194389e-08, -1.272509e-08, -1.36431e-08, -1.453994e-08, 
    -1.518215e-08, -1.562107e-08, -1.60059e-08, -1.634877e-08, -1.675957e-08, 
    -1.71587e-08, -1.758749e-08, -1.804067e-08, -1.830168e-08, -1.84028e-08,
  -1.124877e-08, -1.17948e-08, -1.2445e-08, -1.323852e-08, -1.412096e-08, 
    -1.482169e-08, -1.526754e-08, -1.564749e-08, -1.602102e-08, 
    -1.633528e-08, -1.662911e-08, -1.695923e-08, -1.740535e-08, 
    -1.779284e-08, -1.817007e-08,
  -1.129047e-08, -1.178096e-08, -1.234439e-08, -1.294299e-08, -1.365374e-08, 
    -1.439821e-08, -1.499863e-08, -1.546158e-08, -1.582232e-08, 
    -1.620825e-08, -1.648973e-08, -1.674236e-08, -1.717482e-08, 
    -1.766302e-08, -1.808956e-08,
  -3.818667e-09, -4.455406e-09, -5.113836e-09, -5.816579e-09, -6.647151e-09, 
    -7.635975e-09, -8.49251e-09, -9.376464e-09, -1.041473e-08, -1.159091e-08, 
    -1.297423e-08, -1.446343e-08, -1.586805e-08, -1.707479e-08, -1.807797e-08,
  -3.489034e-09, -4.082304e-09, -4.704672e-09, -5.322333e-09, -6.027064e-09, 
    -6.854035e-09, -7.828644e-09, -8.723585e-09, -9.581476e-09, 
    -1.058655e-08, -1.168285e-08, -1.298291e-08, -1.451236e-08, -1.58992e-08, 
    -1.720013e-08,
  -3.412028e-09, -3.841274e-09, -4.37343e-09, -4.894109e-09, -5.518652e-09, 
    -6.279635e-09, -7.13485e-09, -8.1553e-09, -9.064895e-09, -1.000981e-08, 
    -1.096017e-08, -1.187084e-08, -1.308632e-08, -1.450922e-08, -1.584613e-08,
  -3.494753e-09, -3.637302e-09, -3.957612e-09, -4.389071e-09, -4.932378e-09, 
    -5.639359e-09, -6.431968e-09, -7.347449e-09, -8.329394e-09, 
    -9.344118e-09, -1.044234e-08, -1.134765e-08, -1.226895e-08, 
    -1.334907e-08, -1.451356e-08,
  -3.645785e-09, -3.586595e-09, -3.702923e-09, -3.999969e-09, -4.45316e-09, 
    -5.096607e-09, -5.860762e-09, -6.687442e-09, -7.593226e-09, 
    -8.584665e-09, -9.744962e-09, -1.086882e-08, -1.182775e-08, 
    -1.269148e-08, -1.366774e-08,
  -3.793929e-09, -3.624347e-09, -3.554593e-09, -3.737206e-09, -4.08889e-09, 
    -4.603057e-09, -5.246898e-09, -6.006229e-09, -6.869206e-09, 
    -7.794207e-09, -8.953635e-09, -1.012056e-08, -1.130984e-08, -1.23363e-08, 
    -1.319573e-08,
  -4.137305e-09, -3.937779e-09, -3.763468e-09, -3.751042e-09, -3.95057e-09, 
    -4.364878e-09, -4.896753e-09, -5.467118e-09, -6.173816e-09, -7.04076e-09, 
    -8.009856e-09, -9.275635e-09, -1.049072e-08, -1.164753e-08, -1.274762e-08,
  -4.122679e-09, -4.167226e-09, -4.055766e-09, -3.913739e-09, -3.920645e-09, 
    -4.185642e-09, -4.695568e-09, -5.243751e-09, -5.81389e-09, -6.484119e-09, 
    -7.31504e-09, -8.273674e-09, -9.561606e-09, -1.077904e-08, -1.19612e-08,
  -4.376478e-09, -4.341024e-09, -4.404864e-09, -4.319007e-09, -4.241637e-09, 
    -4.367524e-09, -4.642763e-09, -5.080703e-09, -5.600252e-09, 
    -6.136555e-09, -6.801087e-09, -7.596221e-09, -8.618969e-09, 
    -9.883202e-09, -1.112556e-08,
  -4.349515e-09, -4.430078e-09, -4.443381e-09, -4.467597e-09, -4.416386e-09, 
    -4.449149e-09, -4.792668e-09, -5.140489e-09, -5.541426e-09, -5.99694e-09, 
    -6.495231e-09, -7.078728e-09, -7.827671e-09, -8.883346e-09, -1.01457e-08,
  -3.321766e-09, -3.342449e-09, -3.492979e-09, -3.661973e-09, -3.829533e-09, 
    -4.033868e-09, -4.264762e-09, -4.481455e-09, -4.679021e-09, 
    -4.881172e-09, -5.1156e-09, -5.437995e-09, -5.901463e-09, -6.532367e-09, 
    -7.230806e-09,
  -3.162266e-09, -3.18105e-09, -3.22279e-09, -3.321786e-09, -3.460817e-09, 
    -3.619794e-09, -3.824796e-09, -4.061665e-09, -4.290325e-09, 
    -4.504012e-09, -4.713659e-09, -4.933884e-09, -5.181866e-09, 
    -5.487445e-09, -5.882232e-09,
  -3.084512e-09, -3.119626e-09, -3.168044e-09, -3.247725e-09, -3.326804e-09, 
    -3.40953e-09, -3.524703e-09, -3.660646e-09, -3.827719e-09, -4.011052e-09, 
    -4.19088e-09, -4.371929e-09, -4.555146e-09, -4.731482e-09, -4.919684e-09,
  -2.981032e-09, -3.050394e-09, -3.13188e-09, -3.207866e-09, -3.23962e-09, 
    -3.249777e-09, -3.279187e-09, -3.346633e-09, -3.434457e-09, -3.55369e-09, 
    -3.677218e-09, -3.817395e-09, -3.974173e-09, -4.118165e-09, -4.276353e-09,
  -2.901537e-09, -2.968563e-09, -3.039921e-09, -3.105258e-09, -3.133891e-09, 
    -3.150562e-09, -3.147138e-09, -3.157833e-09, -3.173176e-09, 
    -3.217252e-09, -3.300101e-09, -3.429294e-09, -3.570604e-09, 
    -3.696969e-09, -3.808829e-09,
  -2.803561e-09, -2.842085e-09, -2.884822e-09, -2.930271e-09, -2.970629e-09, 
    -3.009816e-09, -3.038932e-09, -3.051928e-09, -3.049933e-09, 
    -3.036711e-09, -3.030584e-09, -3.077052e-09, -3.182028e-09, -3.30596e-09, 
    -3.441679e-09,
  -2.769215e-09, -2.771678e-09, -2.779974e-09, -2.79022e-09, -2.813449e-09, 
    -2.84837e-09, -2.894801e-09, -2.934073e-09, -2.955058e-09, -2.950633e-09, 
    -2.929613e-09, -2.913196e-09, -2.917035e-09, -2.967441e-09, -3.075617e-09,
  -2.703149e-09, -2.702338e-09, -2.6901e-09, -2.686368e-09, -2.698491e-09, 
    -2.724793e-09, -2.762351e-09, -2.805508e-09, -2.847656e-09, 
    -2.869958e-09, -2.882699e-09, -2.87248e-09, -2.856087e-09, -2.833304e-09, 
    -2.844193e-09,
  -2.76527e-09, -2.781079e-09, -2.776936e-09, -2.770175e-09, -2.769102e-09, 
    -2.769161e-09, -2.778204e-09, -2.801326e-09, -2.842092e-09, -2.88181e-09, 
    -2.906783e-09, -2.906589e-09, -2.898325e-09, -2.879958e-09, -2.862165e-09,
  -2.828148e-09, -2.834165e-09, -2.845092e-09, -2.845166e-09, -2.860927e-09, 
    -2.885168e-09, -2.906137e-09, -2.905867e-09, -2.922091e-09, -2.94289e-09, 
    -2.963872e-09, -2.973252e-09, -2.955448e-09, -2.939455e-09, -2.921872e-09,
  -6.649428e-09, -6.898265e-09, -7.210888e-09, -7.5585e-09, -7.992514e-09, 
    -8.451425e-09, -8.937656e-09, -9.46068e-09, -9.980407e-09, -1.084037e-08, 
    -1.218483e-08, -1.388905e-08, -1.54904e-08, -1.734823e-08, -1.957019e-08,
  -5.633594e-09, -5.774623e-09, -6.003969e-09, -6.27836e-09, -6.602475e-09, 
    -6.990666e-09, -7.358711e-09, -7.805891e-09, -8.333841e-09, 
    -8.832443e-09, -9.52762e-09, -1.057822e-08, -1.190079e-08, -1.342381e-08, 
    -1.513058e-08,
  -4.898021e-09, -4.996136e-09, -5.135328e-09, -5.343447e-09, -5.591262e-09, 
    -5.846243e-09, -6.185002e-09, -6.496957e-09, -6.872767e-09, 
    -7.322625e-09, -7.763018e-09, -8.330043e-09, -9.147578e-09, 
    -1.021204e-08, -1.146137e-08,
  -4.120044e-09, -4.224288e-09, -4.328253e-09, -4.465992e-09, -4.64755e-09, 
    -4.866151e-09, -5.114526e-09, -5.397124e-09, -5.663523e-09, 
    -5.975675e-09, -6.365526e-09, -6.771984e-09, -7.272953e-09, 
    -7.982329e-09, -8.864881e-09,
  -3.571453e-09, -3.641776e-09, -3.697361e-09, -3.772645e-09, -3.881306e-09, 
    -4.037974e-09, -4.230817e-09, -4.454305e-09, -4.682216e-09, -4.89148e-09, 
    -5.169454e-09, -5.491494e-09, -5.80534e-09, -6.236174e-09, -6.827855e-09,
  -3.149043e-09, -3.200358e-09, -3.267103e-09, -3.316027e-09, -3.380427e-09, 
    -3.456933e-09, -3.577668e-09, -3.725626e-09, -3.911029e-09, -4.09979e-09, 
    -4.281495e-09, -4.53567e-09, -4.775686e-09, -5.020274e-09, -5.337929e-09,
  -2.837101e-09, -2.894385e-09, -2.968698e-09, -3.029135e-09, -3.092844e-09, 
    -3.149869e-09, -3.21693e-09, -3.289819e-09, -3.382617e-09, -3.504713e-09, 
    -3.650155e-09, -3.805702e-09, -3.993842e-09, -4.190576e-09, -4.387926e-09,
  -2.534615e-09, -2.60117e-09, -2.668445e-09, -2.722674e-09, -2.776872e-09, 
    -2.841374e-09, -2.899864e-09, -2.973796e-09, -3.035836e-09, 
    -3.094734e-09, -3.176225e-09, -3.270035e-09, -3.403222e-09, 
    -3.558902e-09, -3.714049e-09,
  -2.337723e-09, -2.398205e-09, -2.45888e-09, -2.5097e-09, -2.555004e-09, 
    -2.59664e-09, -2.671385e-09, -2.737902e-09, -2.799964e-09, -2.854965e-09, 
    -2.904222e-09, -2.952693e-09, -3.012385e-09, -3.112837e-09, -3.235912e-09,
  -2.199983e-09, -2.258465e-09, -2.324333e-09, -2.368317e-09, -2.383573e-09, 
    -2.449467e-09, -2.509957e-09, -2.572557e-09, -2.639559e-09, 
    -2.707199e-09, -2.755894e-09, -2.794686e-09, -2.838108e-09, 
    -2.895505e-09, -2.985668e-09,
  -8.539338e-09, -8.548315e-09, -8.683543e-09, -8.891524e-09, -9.116971e-09, 
    -9.293987e-09, -9.560002e-09, -9.836751e-09, -1.030042e-08, 
    -1.101943e-08, -1.182003e-08, -1.27125e-08, -1.387869e-08, -1.548097e-08, 
    -1.734044e-08,
  -7.619078e-09, -7.636768e-09, -7.730429e-09, -7.913159e-09, -8.166221e-09, 
    -8.39668e-09, -8.676142e-09, -8.992598e-09, -9.347265e-09, -9.834008e-09, 
    -1.050969e-08, -1.126028e-08, -1.215893e-08, -1.340339e-08, -1.490525e-08,
  -6.902572e-09, -6.944226e-09, -7.020942e-09, -7.130405e-09, -7.322989e-09, 
    -7.536881e-09, -7.762976e-09, -8.076251e-09, -8.441454e-09, -8.83561e-09, 
    -9.375567e-09, -9.99693e-09, -1.076542e-08, -1.161911e-08, -1.28795e-08,
  -6.177401e-09, -6.217903e-09, -6.302904e-09, -6.39035e-09, -6.543115e-09, 
    -6.761064e-09, -7.006505e-09, -7.244668e-09, -7.576702e-09, 
    -7.927522e-09, -8.371104e-09, -8.903175e-09, -9.513644e-09, 
    -1.025766e-08, -1.110441e-08,
  -5.515834e-09, -5.55522e-09, -5.631061e-09, -5.749639e-09, -5.876344e-09, 
    -6.067341e-09, -6.312048e-09, -6.568934e-09, -6.838662e-09, 
    -7.160542e-09, -7.496022e-09, -7.932582e-09, -8.478202e-09, 
    -9.049018e-09, -9.822586e-09,
  -4.826163e-09, -4.849956e-09, -4.951963e-09, -5.064426e-09, -5.206116e-09, 
    -5.387082e-09, -5.611773e-09, -5.890944e-09, -6.18622e-09, -6.488972e-09, 
    -6.815889e-09, -7.108992e-09, -7.54198e-09, -8.037927e-09, -8.605902e-09,
  -4.242693e-09, -4.234359e-09, -4.33247e-09, -4.465603e-09, -4.608129e-09, 
    -4.769861e-09, -4.937314e-09, -5.166776e-09, -5.465618e-09, 
    -5.808969e-09, -6.16536e-09, -6.511029e-09, -6.82036e-09, -7.251838e-09, 
    -7.646777e-09,
  -3.639846e-09, -3.649917e-09, -3.753999e-09, -3.892401e-09, -4.052378e-09, 
    -4.217955e-09, -4.378172e-09, -4.517307e-09, -4.729011e-09, 
    -5.033642e-09, -5.348356e-09, -5.769706e-09, -6.164976e-09, 
    -6.558088e-09, -6.996431e-09,
  -3.110962e-09, -3.106525e-09, -3.213732e-09, -3.334304e-09, -3.488024e-09, 
    -3.654126e-09, -3.844804e-09, -4.011351e-09, -4.154308e-09, 
    -4.366304e-09, -4.626433e-09, -4.926689e-09, -5.329229e-09, 
    -5.759726e-09, -6.203532e-09,
  -2.644906e-09, -2.652873e-09, -2.754746e-09, -2.850084e-09, -2.94074e-09, 
    -3.071345e-09, -3.231655e-09, -3.42512e-09, -3.604086e-09, -3.773918e-09, 
    -4.01133e-09, -4.269526e-09, -4.57892e-09, -4.946633e-09, -5.359721e-09,
  -1.14576e-08, -1.118153e-08, -1.099336e-08, -1.088923e-08, -1.083667e-08, 
    -1.08201e-08, -1.084318e-08, -1.09073e-08, -1.101213e-08, -1.113947e-08, 
    -1.128123e-08, -1.146206e-08, -1.171237e-08, -1.20427e-08, -1.23821e-08,
  -1.01093e-08, -9.855223e-09, -9.69966e-09, -9.578802e-09, -9.516403e-09, 
    -9.517297e-09, -9.604679e-09, -9.753238e-09, -9.950723e-09, -1.01239e-08, 
    -1.03051e-08, -1.048074e-08, -1.07308e-08, -1.101804e-08, -1.138439e-08,
  -9.008112e-09, -8.833903e-09, -8.729878e-09, -8.622314e-09, -8.551843e-09, 
    -8.547027e-09, -8.583982e-09, -8.684158e-09, -8.824007e-09, -9.05657e-09, 
    -9.282004e-09, -9.523053e-09, -9.791147e-09, -1.009196e-08, -1.043583e-08,
  -7.889699e-09, -7.792443e-09, -7.732063e-09, -7.664744e-09, -7.62362e-09, 
    -7.61966e-09, -7.638118e-09, -7.705825e-09, -7.813548e-09, -7.985513e-09, 
    -8.236365e-09, -8.500837e-09, -8.793109e-09, -9.088294e-09, -9.42355e-09,
  -7.130546e-09, -7.045648e-09, -6.99906e-09, -6.960015e-09, -6.942934e-09, 
    -6.949421e-09, -6.971861e-09, -7.010011e-09, -7.082009e-09, 
    -7.193556e-09, -7.368686e-09, -7.612678e-09, -7.904291e-09, 
    -8.233545e-09, -8.502432e-09,
  -6.566742e-09, -6.457848e-09, -6.411976e-09, -6.364887e-09, -6.3396e-09, 
    -6.341868e-09, -6.359398e-09, -6.399421e-09, -6.451777e-09, 
    -6.539695e-09, -6.669084e-09, -6.846122e-09, -7.083789e-09, 
    -7.388878e-09, -7.717391e-09,
  -6.03355e-09, -5.92047e-09, -5.861656e-09, -5.804571e-09, -5.76795e-09, 
    -5.761587e-09, -5.789769e-09, -5.827571e-09, -5.881837e-09, 
    -5.961486e-09, -6.073746e-09, -6.217084e-09, -6.402347e-09, 
    -6.652763e-09, -6.947008e-09,
  -5.549522e-09, -5.430458e-09, -5.362209e-09, -5.28327e-09, -5.234318e-09, 
    -5.210154e-09, -5.234871e-09, -5.274797e-09, -5.335057e-09, 
    -5.414055e-09, -5.516316e-09, -5.644691e-09, -5.797147e-09, 
    -6.008254e-09, -6.262437e-09,
  -5.020221e-09, -4.902684e-09, -4.828161e-09, -4.754289e-09, -4.690403e-09, 
    -4.659024e-09, -4.661862e-09, -4.704825e-09, -4.768676e-09, 
    -4.850246e-09, -4.965606e-09, -5.105132e-09, -5.251868e-09, 
    -5.435131e-09, -5.660931e-09,
  -4.503714e-09, -4.388109e-09, -4.317254e-09, -4.232245e-09, -4.160989e-09, 
    -4.122765e-09, -4.114361e-09, -4.144548e-09, -4.184027e-09, 
    -4.253737e-09, -4.359133e-09, -4.504115e-09, -4.64992e-09, -4.856742e-09, 
    -5.09464e-09,
  -1.589856e-08, -1.554582e-08, -1.510931e-08, -1.461077e-08, -1.414324e-08, 
    -1.374939e-08, -1.338774e-08, -1.304466e-08, -1.276556e-08, -1.25451e-08, 
    -1.240586e-08, -1.231361e-08, -1.224458e-08, -1.219434e-08, -1.220719e-08,
  -1.449535e-08, -1.415048e-08, -1.3818e-08, -1.337414e-08, -1.297264e-08, 
    -1.260964e-08, -1.225698e-08, -1.192746e-08, -1.164473e-08, 
    -1.143363e-08, -1.130557e-08, -1.120399e-08, -1.111201e-08, 
    -1.104536e-08, -1.103236e-08,
  -1.368707e-08, -1.342085e-08, -1.308127e-08, -1.260261e-08, -1.220241e-08, 
    -1.184098e-08, -1.152458e-08, -1.119333e-08, -1.088826e-08, 
    -1.066397e-08, -1.049105e-08, -1.037111e-08, -1.025697e-08, 
    -1.016852e-08, -1.014667e-08,
  -1.28434e-08, -1.255712e-08, -1.221102e-08, -1.172023e-08, -1.129038e-08, 
    -1.097069e-08, -1.066568e-08, -1.033944e-08, -1.003407e-08, 
    -9.804384e-09, -9.63143e-09, -9.529055e-09, -9.421123e-09, -9.320779e-09, 
    -9.261813e-09,
  -1.20952e-08, -1.176237e-08, -1.140646e-08, -1.088178e-08, -1.051477e-08, 
    -1.024582e-08, -9.954255e-09, -9.638113e-09, -9.344099e-09, 
    -9.114183e-09, -8.964495e-09, -8.878112e-09, -8.800195e-09, 
    -8.712816e-09, -8.644757e-09,
  -1.104319e-08, -1.065659e-08, -1.028505e-08, -9.805042e-09, -9.506952e-09, 
    -9.280567e-09, -8.992523e-09, -8.674062e-09, -8.377055e-09, 
    -8.138445e-09, -7.980534e-09, -7.909359e-09, -7.888779e-09, -7.87787e-09, 
    -7.872164e-09,
  -9.952457e-09, -9.485381e-09, -9.113006e-09, -8.779151e-09, -8.56506e-09, 
    -8.312321e-09, -7.97972e-09, -7.670629e-09, -7.409126e-09, -7.218823e-09, 
    -7.08025e-09, -7.027417e-09, -7.029804e-09, -7.06604e-09, -7.100458e-09,
  -8.777213e-09, -8.371097e-09, -8.025967e-09, -7.750098e-09, -7.516473e-09, 
    -7.235584e-09, -6.882409e-09, -6.585061e-09, -6.375752e-09, 
    -6.258699e-09, -6.16528e-09, -6.130207e-09, -6.15473e-09, -6.208275e-09, 
    -6.279266e-09,
  -7.703345e-09, -7.266602e-09, -6.963742e-09, -6.699683e-09, -6.382102e-09, 
    -6.082613e-09, -5.795413e-09, -5.571227e-09, -5.43489e-09, -5.366903e-09, 
    -5.317647e-09, -5.309916e-09, -5.348353e-09, -5.415354e-09, -5.503396e-09,
  -6.728829e-09, -6.211227e-09, -5.890261e-09, -5.604756e-09, -5.290058e-09, 
    -5.014596e-09, -4.782487e-09, -4.626349e-09, -4.537319e-09, -4.49954e-09, 
    -4.479083e-09, -4.514464e-09, -4.576703e-09, -4.661437e-09, -4.763725e-09,
  -1.981541e-08, -1.961762e-08, -1.946705e-08, -1.928622e-08, -1.916329e-08, 
    -1.902742e-08, -1.891324e-08, -1.883479e-08, -1.868855e-08, 
    -1.855692e-08, -1.841692e-08, -1.829031e-08, -1.814126e-08, 
    -1.804964e-08, -1.798669e-08,
  -1.932595e-08, -1.902174e-08, -1.889602e-08, -1.86403e-08, -1.848927e-08, 
    -1.82569e-08, -1.813565e-08, -1.795916e-08, -1.777257e-08, -1.757581e-08, 
    -1.740708e-08, -1.726299e-08, -1.715862e-08, -1.706231e-08, -1.698638e-08,
  -1.870171e-08, -1.845173e-08, -1.828125e-08, -1.806506e-08, -1.784411e-08, 
    -1.763165e-08, -1.747259e-08, -1.729908e-08, -1.710236e-08, 
    -1.688807e-08, -1.668462e-08, -1.651021e-08, -1.63416e-08, -1.620008e-08, 
    -1.607837e-08,
  -1.788739e-08, -1.762662e-08, -1.740964e-08, -1.702573e-08, -1.687704e-08, 
    -1.667228e-08, -1.654158e-08, -1.635919e-08, -1.615564e-08, 
    -1.595744e-08, -1.575031e-08, -1.549263e-08, -1.524417e-08, 
    -1.497547e-08, -1.477875e-08,
  -1.675083e-08, -1.656485e-08, -1.633449e-08, -1.594181e-08, -1.580323e-08, 
    -1.570293e-08, -1.555583e-08, -1.541406e-08, -1.523326e-08, 
    -1.504345e-08, -1.484137e-08, -1.458963e-08, -1.433899e-08, 
    -1.405957e-08, -1.381084e-08,
  -1.540648e-08, -1.525819e-08, -1.511541e-08, -1.484573e-08, -1.46772e-08, 
    -1.466281e-08, -1.453437e-08, -1.43986e-08, -1.422016e-08, -1.403228e-08, 
    -1.385345e-08, -1.367001e-08, -1.342705e-08, -1.320046e-08, -1.297229e-08,
  -1.426954e-08, -1.406379e-08, -1.399898e-08, -1.381616e-08, -1.369544e-08, 
    -1.373919e-08, -1.366653e-08, -1.352363e-08, -1.333907e-08, 
    -1.315637e-08, -1.296235e-08, -1.274479e-08, -1.250885e-08, -1.22881e-08, 
    -1.207089e-08,
  -1.319093e-08, -1.299455e-08, -1.302515e-08, -1.295099e-08, -1.298597e-08, 
    -1.290786e-08, -1.274179e-08, -1.251562e-08, -1.228823e-08, 
    -1.209851e-08, -1.182449e-08, -1.152645e-08, -1.12622e-08, -1.104107e-08, 
    -1.082007e-08,
  -1.234461e-08, -1.215225e-08, -1.218583e-08, -1.205753e-08, -1.201786e-08, 
    -1.189831e-08, -1.164105e-08, -1.142903e-08, -1.117798e-08, 
    -1.094532e-08, -1.063952e-08, -1.033069e-08, -1.00677e-08, -9.822004e-09, 
    -9.596146e-09,
  -1.117867e-08, -1.112226e-08, -1.110728e-08, -1.099424e-08, -1.094769e-08, 
    -1.084671e-08, -1.066374e-08, -1.041302e-08, -1.009678e-08, 
    -9.768003e-09, -9.407542e-09, -9.06299e-09, -8.785485e-09, -8.532681e-09, 
    -8.303091e-09,
  -2.57166e-08, -2.51952e-08, -2.518795e-08, -2.451492e-08, -2.374777e-08, 
    -2.208729e-08, -1.943182e-08, -1.67607e-08, -1.49063e-08, -1.775928e-08, 
    -1.959092e-08, -2.030095e-08, -2.072574e-08, -2.099107e-08, -2.109914e-08,
  -2.494749e-08, -2.467471e-08, -2.444317e-08, -2.389152e-08, -2.33312e-08, 
    -2.183584e-08, -1.672453e-08, -1.537799e-08, -1.48203e-08, -1.846884e-08, 
    -1.879135e-08, -1.859292e-08, -1.907977e-08, -1.942341e-08, -1.964053e-08,
  -2.421885e-08, -2.396963e-08, -2.356899e-08, -2.336165e-08, -2.273369e-08, 
    -2.097148e-08, -1.761026e-08, -1.722672e-08, -1.802233e-08, 
    -2.053884e-08, -2.005903e-08, -1.972995e-08, -2.004476e-08, 
    -2.005738e-08, -1.984028e-08,
  -2.321537e-08, -2.29547e-08, -2.264595e-08, -2.23144e-08, -2.173602e-08, 
    -1.958587e-08, -1.89723e-08, -1.887014e-08, -2.03707e-08, -2.055094e-08, 
    -1.976658e-08, -1.961918e-08, -1.922178e-08, -1.888352e-08, -1.858855e-08,
  -2.193492e-08, -2.17879e-08, -2.149137e-08, -2.1062e-08, -2.067529e-08, 
    -1.998919e-08, -2.074744e-08, -2.015621e-08, -2.0633e-08, -2.004769e-08, 
    -1.923767e-08, -1.86862e-08, -1.82856e-08, -1.794206e-08, -1.76995e-08,
  -2.073661e-08, -2.059192e-08, -2.022605e-08, -1.9693e-08, -1.916907e-08, 
    -1.89538e-08, -1.895297e-08, -1.978494e-08, -1.979141e-08, -1.929465e-08, 
    -1.872859e-08, -1.835379e-08, -1.783394e-08, -1.731854e-08, -1.693531e-08,
  -1.927525e-08, -1.904641e-08, -1.86771e-08, -1.810491e-08, -1.759801e-08, 
    -1.780588e-08, -1.815014e-08, -1.844732e-08, -1.811793e-08, 
    -1.748468e-08, -1.704996e-08, -1.679452e-08, -1.645348e-08, 
    -1.612962e-08, -1.589863e-08,
  -1.729119e-08, -1.704058e-08, -1.675164e-08, -1.642212e-08, -1.61907e-08, 
    -1.616537e-08, -1.626658e-08, -1.596333e-08, -1.547795e-08, 
    -1.474603e-08, -1.459317e-08, -1.448636e-08, -1.435052e-08, 
    -1.418723e-08, -1.406637e-08,
  -1.497552e-08, -1.494818e-08, -1.489748e-08, -1.495214e-08, -1.484401e-08, 
    -1.47557e-08, -1.455237e-08, -1.424638e-08, -1.346021e-08, -1.301433e-08, 
    -1.296563e-08, -1.296854e-08, -1.286743e-08, -1.272309e-08, -1.255664e-08,
  -1.159023e-08, -1.203453e-08, -1.245917e-08, -1.275179e-08, -1.288036e-08, 
    -1.274533e-08, -1.258266e-08, -1.224815e-08, -1.139187e-08, 
    -1.107717e-08, -1.105605e-08, -1.096724e-08, -1.091442e-08, 
    -1.081487e-08, -1.06618e-08,
  -2.532441e-08, -2.566479e-08, -2.579717e-08, -2.601526e-08, -2.619627e-08, 
    -2.623293e-08, -2.630783e-08, -2.670391e-08, -2.737909e-08, 
    -2.733383e-08, -2.784841e-08, -2.700819e-08, -2.615823e-08, 
    -2.608442e-08, -2.611998e-08,
  -2.424664e-08, -2.466415e-08, -2.488928e-08, -2.507253e-08, -2.523295e-08, 
    -2.528537e-08, -2.538579e-08, -2.580663e-08, -2.635183e-08, 
    -2.650727e-08, -2.634856e-08, -2.616495e-08, -2.51255e-08, -2.50536e-08, 
    -2.476993e-08,
  -2.248761e-08, -2.293127e-08, -2.333533e-08, -2.368168e-08, -2.392328e-08, 
    -2.415933e-08, -2.432925e-08, -2.473807e-08, -2.51399e-08, -2.535855e-08, 
    -2.494192e-08, -2.456562e-08, -2.407729e-08, -2.388483e-08, -2.357475e-08,
  -1.996125e-08, -2.066671e-08, -2.124257e-08, -2.183471e-08, -2.224685e-08, 
    -2.264229e-08, -2.292745e-08, -2.343267e-08, -2.381408e-08, 
    -2.393477e-08, -2.363979e-08, -2.297066e-08, -2.272451e-08, 
    -2.267977e-08, -2.260492e-08,
  -1.753472e-08, -1.824477e-08, -1.88298e-08, -1.946997e-08, -2.001914e-08, 
    -2.057444e-08, -2.104466e-08, -2.165589e-08, -2.208357e-08, -2.22104e-08, 
    -2.188191e-08, -2.125384e-08, -2.107088e-08, -2.125753e-08, -2.130859e-08,
  -1.546157e-08, -1.618262e-08, -1.677883e-08, -1.730107e-08, -1.78087e-08, 
    -1.827709e-08, -1.88131e-08, -1.93883e-08, -1.978678e-08, -1.996578e-08, 
    -1.959268e-08, -1.912604e-08, -1.915728e-08, -1.935586e-08, -1.952232e-08,
  -1.314364e-08, -1.402187e-08, -1.473668e-08, -1.531737e-08, -1.578366e-08, 
    -1.628665e-08, -1.671036e-08, -1.714222e-08, -1.749575e-08, 
    -1.761047e-08, -1.707259e-08, -1.690767e-08, -1.716698e-08, 
    -1.745093e-08, -1.762533e-08,
  -1.068341e-08, -1.16041e-08, -1.247169e-08, -1.323321e-08, -1.377434e-08, 
    -1.431535e-08, -1.474429e-08, -1.516343e-08, -1.546484e-08, 
    -1.535562e-08, -1.497303e-08, -1.504023e-08, -1.543998e-08, 
    -1.558006e-08, -1.561199e-08,
  -7.914449e-09, -8.824995e-09, -9.76551e-09, -1.064618e-08, -1.13538e-08, 
    -1.198603e-08, -1.255031e-08, -1.294495e-08, -1.325843e-08, 
    -1.320059e-08, -1.324566e-08, -1.356907e-08, -1.383578e-08, 
    -1.390424e-08, -1.401598e-08,
  -5.499009e-09, -6.304478e-09, -7.159784e-09, -8.041929e-09, -8.798479e-09, 
    -9.41758e-09, -9.946831e-09, -1.04047e-08, -1.078902e-08, -1.107211e-08, 
    -1.132981e-08, -1.164619e-08, -1.178573e-08, -1.201679e-08, -1.225793e-08,
  -1.930044e-08, -1.973922e-08, -2.020359e-08, -2.075006e-08, -2.145436e-08, 
    -2.215606e-08, -2.288916e-08, -2.348767e-08, -2.385751e-08, 
    -2.408976e-08, -2.437327e-08, -2.47857e-08, -2.525209e-08, -2.56676e-08, 
    -2.599019e-08,
  -1.915741e-08, -1.949847e-08, -1.986799e-08, -2.021577e-08, -2.054952e-08, 
    -2.099589e-08, -2.153154e-08, -2.20498e-08, -2.273987e-08, -2.342251e-08, 
    -2.378889e-08, -2.402866e-08, -2.433334e-08, -2.476897e-08, -2.517853e-08,
  -1.846141e-08, -1.884102e-08, -1.91708e-08, -1.953225e-08, -1.987722e-08, 
    -2.014333e-08, -2.046388e-08, -2.084281e-08, -2.126845e-08, 
    -2.178391e-08, -2.231486e-08, -2.272971e-08, -2.30377e-08, -2.329775e-08, 
    -2.361652e-08,
  -1.75778e-08, -1.800573e-08, -1.831911e-08, -1.863173e-08, -1.898148e-08, 
    -1.929914e-08, -1.957453e-08, -1.981342e-08, -2.001854e-08, 
    -2.030419e-08, -2.062496e-08, -2.106283e-08, -2.131011e-08, -2.15707e-08, 
    -2.175716e-08,
  -1.612641e-08, -1.667516e-08, -1.71101e-08, -1.748148e-08, -1.782293e-08, 
    -1.81957e-08, -1.84321e-08, -1.86934e-08, -1.890784e-08, -1.910341e-08, 
    -1.927003e-08, -1.945053e-08, -1.968399e-08, -1.988728e-08, -2.002066e-08,
  -1.425702e-08, -1.481801e-08, -1.534771e-08, -1.583104e-08, -1.624095e-08, 
    -1.656331e-08, -1.685213e-08, -1.712081e-08, -1.737002e-08, 
    -1.756761e-08, -1.780711e-08, -1.801335e-08, -1.819402e-08, 
    -1.837791e-08, -1.850126e-08,
  -1.21716e-08, -1.271296e-08, -1.323893e-08, -1.376999e-08, -1.423217e-08, 
    -1.45636e-08, -1.479771e-08, -1.497827e-08, -1.520646e-08, -1.545744e-08, 
    -1.568514e-08, -1.593233e-08, -1.614911e-08, -1.636606e-08, -1.658189e-08,
  -1.022132e-08, -1.055537e-08, -1.096417e-08, -1.14584e-08, -1.19617e-08, 
    -1.232642e-08, -1.257891e-08, -1.277995e-08, -1.298601e-08, 
    -1.317037e-08, -1.33954e-08, -1.356003e-08, -1.37515e-08, -1.391198e-08, 
    -1.408442e-08,
  -8.686122e-09, -8.801288e-09, -9.043811e-09, -9.302995e-09, -9.646976e-09, 
    -1.000181e-08, -1.030798e-08, -1.059309e-08, -1.083804e-08, 
    -1.105434e-08, -1.126827e-08, -1.147636e-08, -1.163823e-08, -1.17779e-08, 
    -1.189717e-08,
  -7.190577e-09, -7.320502e-09, -7.465291e-09, -7.640535e-09, -7.881612e-09, 
    -8.128824e-09, -8.387627e-09, -8.615653e-09, -8.83062e-09, -9.048303e-09, 
    -9.228522e-09, -9.410309e-09, -9.585838e-09, -9.756174e-09, -9.924321e-09 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
