netcdf atmos_daily.00010101-00010701.pv350K.tile3 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pv350K(time, grid_yt, grid_xt) ;
		pv350K:_FillValue = -1.e+10f ;
		pv350K:missing_value = -1.e+10f ;
		pv350K:units = "(K m**2) / (kg s)" ;
		pv350K:long_name = "350-K potential vorticity; needs x350 scaling" ;
		pv350K:cell_methods = "time: mean" ;
		pv350K:time_avg_info = "average_T1,average_T2,average_DT" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile3.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.0008770345, 0.4596241, 0.9892928, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.01035247, 0.004304647, 0.6546783, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.8534847, 0.8118016, 0.9951549, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9894952, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4452189, 0.3028796, 0.7140614, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9903189, 0.3150955, 0.0007410151, 0, 0.02645395, 
    0.9012984, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.681631, 0, 0, 0, 0.004980796, 0.7708192, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5536854, 0, 0, 0, 0.004666397, 0.9395298, 1,
  1, 1, 1, 1, 1, 1, 1, 0.9995009, 0.3626226, 0, 0, 0, 0, 0.8367797, 1,
  1, 1, 1, 1, 1, 0.8451425, 0.7016711, 0.3953246, 0, 0, 0, 0, 0.006316811, 
    0.8673657, 1 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pv350K =
  1.956544e-08, 1.929139e-08, 1.919465e-08, 1.878182e-08, 1.871692e-08, 
    1.831042e-08, 1.848399e-08, 1.917274e-08, 1.987178e-08, 2.160755e-08, 
    2.175548e-08, 2.084801e-08, 2.093063e-08, 2.1128e-08, 2.145071e-08,
  1.924618e-08, 1.861085e-08, 1.843349e-08, 1.855146e-08, 1.847449e-08, 
    1.821514e-08, 1.820239e-08, 1.875827e-08, 1.981038e-08, 2.071397e-08, 
    2.108209e-08, 1.994096e-08, 2.03695e-08, 2.105738e-08, 2.125602e-08,
  1.896625e-08, 1.810602e-08, 1.798871e-08, 1.805245e-08, 1.844115e-08, 
    1.807105e-08, 1.798877e-08, 1.854827e-08, 1.941428e-08, 2.046698e-08, 
    2.079022e-08, 1.923211e-08, 1.957046e-08, 2.050581e-08, 1.971832e-08,
  1.920405e-08, 1.867191e-08, 1.812325e-08, 1.838725e-08, 1.856698e-08, 
    1.830087e-08, 1.801886e-08, 1.840346e-08, 1.949506e-08, 2.096569e-08, 
    2.206437e-08, 2.043815e-08, 2.04335e-08, 2.051314e-08, 1.911095e-08,
  1.942533e-08, 1.846354e-08, 1.831368e-08, 1.838679e-08, 1.815388e-08, 
    1.819651e-08, 1.850711e-08, 1.884478e-08, 1.977738e-08, 2.056808e-08, 
    1.973866e-08, 1.956512e-08, 2.063411e-08, 1.937932e-08, 1.905385e-08,
  1.888121e-08, 1.82102e-08, 1.774435e-08, 1.823549e-08, 1.81034e-08, 
    1.789324e-08, 1.778577e-08, 1.84599e-08, 1.94196e-08, 1.934291e-08, 
    1.838104e-08, 1.773349e-08, 1.869901e-08, 1.872253e-08, 1.900003e-08,
  1.839111e-08, 1.789692e-08, 1.771645e-08, 1.79536e-08, 1.776288e-08, 
    1.762466e-08, 1.797826e-08, 1.862255e-08, 1.900095e-08, 1.859529e-08, 
    1.796657e-08, 1.772472e-08, 1.770177e-08, 1.816552e-08, 1.935776e-08,
  1.814538e-08, 1.789054e-08, 1.76629e-08, 1.812831e-08, 1.795586e-08, 
    1.755651e-08, 1.754161e-08, 1.816586e-08, 1.881464e-08, 1.822258e-08, 
    1.733837e-08, 1.679241e-08, 1.70251e-08, 1.78871e-08, 1.840157e-08,
  1.775092e-08, 1.778386e-08, 1.777956e-08, 1.82177e-08, 1.805073e-08, 
    1.778231e-08, 1.789656e-08, 1.873038e-08, 1.861127e-08, 1.754958e-08, 
    1.683749e-08, 1.659093e-08, 1.685156e-08, 1.742378e-08, 1.846872e-08,
  1.745179e-08, 1.758454e-08, 1.773803e-08, 1.795321e-08, 1.758535e-08, 
    1.758132e-08, 1.792253e-08, 1.82116e-08, 1.781129e-08, 1.673896e-08, 
    1.65018e-08, 1.636424e-08, 1.671453e-08, 1.780003e-08, 1.89503e-08,
  1.284792e-08, 1.337274e-08, 1.402606e-08, 1.427087e-08, 1.486801e-08, 
    1.541114e-08, 1.567895e-08, 1.606956e-08, 1.656348e-08, 1.744238e-08, 
    1.761592e-08, 1.712817e-08, 1.734801e-08, 1.702644e-08, 1.739368e-08,
  1.252309e-08, 1.296808e-08, 1.370908e-08, 1.388071e-08, 1.435606e-08, 
    1.499736e-08, 1.529603e-08, 1.578218e-08, 1.624612e-08, 1.658054e-08, 
    1.706531e-08, 1.655964e-08, 1.725105e-08, 1.707437e-08, 1.754331e-08,
  1.243465e-08, 1.253128e-08, 1.325905e-08, 1.367172e-08, 1.423599e-08, 
    1.463746e-08, 1.491136e-08, 1.55521e-08, 1.603732e-08, 1.648305e-08, 
    1.679708e-08, 1.620301e-08, 1.679161e-08, 1.641904e-08, 1.647339e-08,
  1.176321e-08, 1.219938e-08, 1.302712e-08, 1.337391e-08, 1.365925e-08, 
    1.439421e-08, 1.465397e-08, 1.523886e-08, 1.600995e-08, 1.652107e-08, 
    1.754443e-08, 1.736618e-08, 1.756589e-08, 1.707791e-08, 1.703027e-08,
  1.164646e-08, 1.196141e-08, 1.26927e-08, 1.294381e-08, 1.355718e-08, 
    1.41557e-08, 1.446652e-08, 1.518274e-08, 1.55272e-08, 1.610172e-08, 
    1.625066e-08, 1.723986e-08, 1.782862e-08, 1.735403e-08, 1.753455e-08,
  1.134944e-08, 1.183594e-08, 1.239274e-08, 1.267751e-08, 1.336807e-08, 
    1.382597e-08, 1.421159e-08, 1.469671e-08, 1.535252e-08, 1.611543e-08, 
    1.649473e-08, 1.669392e-08, 1.775549e-08, 1.823309e-08, 1.779278e-08,
  1.133091e-08, 1.18341e-08, 1.2095e-08, 1.259474e-08, 1.330295e-08, 
    1.380561e-08, 1.411691e-08, 1.472077e-08, 1.562712e-08, 1.611647e-08, 
    1.676504e-08, 1.732451e-08, 1.829287e-08, 1.878465e-08, 1.761505e-08,
  1.109911e-08, 1.173844e-08, 1.192149e-08, 1.263294e-08, 1.343114e-08, 
    1.385068e-08, 1.421764e-08, 1.447347e-08, 1.519767e-08, 1.632447e-08, 
    1.712563e-08, 1.7632e-08, 1.861812e-08, 1.87518e-08, 1.76241e-08,
  1.114344e-08, 1.163664e-08, 1.197623e-08, 1.277034e-08, 1.321191e-08, 
    1.358466e-08, 1.404774e-08, 1.451294e-08, 1.526839e-08, 1.685586e-08, 
    1.740907e-08, 1.783043e-08, 1.80845e-08, 1.825886e-08, 1.764112e-08,
  1.099663e-08, 1.132945e-08, 1.175073e-08, 1.268676e-08, 1.32745e-08, 
    1.355677e-08, 1.418207e-08, 1.521078e-08, 1.621811e-08, 1.734021e-08, 
    1.7663e-08, 1.776802e-08, 1.751608e-08, 1.738387e-08, 1.750762e-08,
  1.434228e-08, 1.37052e-08, 1.322355e-08, 1.294443e-08, 1.267345e-08, 
    1.233616e-08, 1.209791e-08, 1.189569e-08, 1.162552e-08, 1.232281e-08, 
    1.392814e-08, 1.461243e-08, 1.445987e-08, 1.39144e-08, 1.44538e-08,
  1.446241e-08, 1.38914e-08, 1.341683e-08, 1.314478e-08, 1.275475e-08, 
    1.243481e-08, 1.22812e-08, 1.213766e-08, 1.207718e-08, 1.251748e-08, 
    1.396813e-08, 1.459092e-08, 1.449721e-08, 1.429368e-08, 1.448021e-08,
  1.531562e-08, 1.409448e-08, 1.356932e-08, 1.299759e-08, 1.269091e-08, 
    1.260626e-08, 1.250521e-08, 1.27403e-08, 1.233387e-08, 1.31082e-08, 
    1.44121e-08, 1.473052e-08, 1.455648e-08, 1.449693e-08, 1.430297e-08,
  1.553789e-08, 1.407991e-08, 1.353046e-08, 1.324652e-08, 1.325761e-08, 
    1.296603e-08, 1.292018e-08, 1.298726e-08, 1.275225e-08, 1.421973e-08, 
    1.507973e-08, 1.509247e-08, 1.476088e-08, 1.419094e-08, 1.418414e-08,
  1.512831e-08, 1.442123e-08, 1.42501e-08, 1.427806e-08, 1.399087e-08, 
    1.361829e-08, 1.331335e-08, 1.339126e-08, 1.389886e-08, 1.592438e-08, 
    1.560632e-08, 1.446949e-08, 1.375401e-08, 1.331072e-08, 1.44209e-08,
  1.541847e-08, 1.524003e-08, 1.506284e-08, 1.50623e-08, 1.437972e-08, 
    1.418908e-08, 1.382348e-08, 1.370007e-08, 1.587601e-08, 1.523496e-08, 
    1.364876e-08, 1.27132e-08, 1.297123e-08, 1.286888e-08, 1.494872e-08,
  1.567795e-08, 1.557864e-08, 1.547474e-08, 1.511543e-08, 1.494558e-08, 
    1.437241e-08, 1.391807e-08, 1.371328e-08, 1.295227e-08, 1.225852e-08, 
    1.18863e-08, 1.211967e-08, 1.260769e-08, 1.3222e-08, 1.500365e-08,
  1.60476e-08, 1.573191e-08, 1.536126e-08, 1.484284e-08, 1.459517e-08, 
    1.456112e-08, 1.40002e-08, 1.379505e-08, 1.113589e-08, 1.109104e-08, 
    1.157539e-08, 1.222781e-08, 1.280272e-08, 1.345988e-08, 1.435667e-08,
  1.529957e-08, 1.540328e-08, 1.480659e-08, 1.424192e-08, 1.397385e-08, 
    1.363603e-08, 1.385409e-08, 1.324639e-08, 1.282276e-08, 1.257813e-08, 
    1.301816e-08, 1.327399e-08, 1.304933e-08, 1.367251e-08, 1.373038e-08,
  1.455544e-08, 1.448643e-08, 1.438512e-08, 1.394735e-08, 1.377711e-08, 
    1.294938e-08, 1.320711e-08, 1.348655e-08, 1.342187e-08, 1.351617e-08, 
    1.370446e-08, 1.371667e-08, 1.373534e-08, 1.371426e-08, 1.407482e-08,
  1.597086e-08, 1.646711e-08, 1.603986e-08, 1.611204e-08, 1.680495e-08, 
    1.733961e-08, 1.733333e-08, 1.716462e-08, 1.704336e-08, 1.662475e-08, 
    1.671011e-08, 1.644657e-08, 1.673056e-08, 1.618363e-08, 1.618309e-08,
  1.679242e-08, 1.625924e-08, 1.63415e-08, 1.607593e-08, 1.749012e-08, 
    1.774039e-08, 1.75045e-08, 1.742121e-08, 1.736198e-08, 1.718532e-08, 
    1.701373e-08, 1.675154e-08, 1.707584e-08, 1.684804e-08, 1.665098e-08,
  1.736957e-08, 1.721249e-08, 1.735485e-08, 1.675613e-08, 1.765031e-08, 
    1.768958e-08, 1.786834e-08, 1.762581e-08, 1.783272e-08, 1.762487e-08, 
    1.768296e-08, 1.739048e-08, 1.783779e-08, 1.770358e-08, 1.74522e-08,
  1.76179e-08, 1.807982e-08, 1.744871e-08, 1.701905e-08, 1.739876e-08, 
    1.746522e-08, 1.773099e-08, 1.753797e-08, 1.753712e-08, 1.78452e-08, 
    1.82386e-08, 1.869321e-08, 1.913822e-08, 1.917805e-08, 1.89219e-08,
  1.794586e-08, 1.818135e-08, 1.805269e-08, 1.697132e-08, 1.738021e-08, 
    1.764403e-08, 1.771509e-08, 1.741956e-08, 1.747017e-08, 1.898845e-08, 
    1.861645e-08, 2.025586e-08, 2.013082e-08, 2.013384e-08, 2.023609e-08,
  1.894417e-08, 1.951858e-08, 1.862894e-08, 1.807488e-08, 1.798707e-08, 
    1.82325e-08, 1.822835e-08, 1.836289e-08, 1.761999e-08, 1.719747e-08, 
    2.042279e-08, 2.012047e-08, 1.969305e-08, 1.849809e-08, 1.934322e-08,
  1.890232e-08, 1.879235e-08, 1.847795e-08, 1.829294e-08, 1.739728e-08, 
    1.74029e-08, 1.750522e-08, 1.770007e-08, 1.764372e-08, 1.666363e-08, 
    1.596265e-08, 1.581657e-08, 1.495532e-08, 1.55188e-08, 1.820188e-08,
  1.908773e-08, 1.895854e-08, 1.942855e-08, 1.860572e-08, 1.824747e-08, 
    1.802759e-08, 1.824684e-08, 1.783867e-08, 1.573397e-08, 1.58997e-08, 
    1.496162e-08, 1.494116e-08, 1.378691e-08, 1.326307e-08, 1.483737e-08,
  1.998015e-08, 1.99649e-08, 2.077469e-08, 2.016142e-08, 1.991666e-08, 
    1.962024e-08, 1.972844e-08, 1.939566e-08, 1.800457e-08, 1.843694e-08, 
    1.79592e-08, 1.787045e-08, 1.745594e-08, 1.517478e-08, 1.322328e-08,
  2.059929e-08, 2.065638e-08, 2.105139e-08, 2.118798e-08, 2.065985e-08, 
    2.038306e-08, 2.012409e-08, 2.012046e-08, 2.011528e-08, 2.008305e-08, 
    1.978969e-08, 1.9592e-08, 1.946109e-08, 1.761783e-08, 1.650278e-08,
  2.00482e-08, 2.066246e-08, 2.085074e-08, 2.181588e-08, 2.217927e-08, 
    2.20709e-08, 2.191909e-08, 2.247371e-08, 2.308424e-08, 2.183639e-08, 
    2.136171e-08, 2.079199e-08, 2.111717e-08, 2.05459e-08, 2.0035e-08,
  2.082227e-08, 2.103173e-08, 2.164746e-08, 2.201945e-08, 2.285928e-08, 
    2.308159e-08, 2.273528e-08, 2.296985e-08, 2.313605e-08, 2.226451e-08, 
    2.137321e-08, 2.122523e-08, 2.165821e-08, 2.109879e-08, 2.046766e-08,
  2.066629e-08, 2.175677e-08, 2.265825e-08, 2.259386e-08, 2.313923e-08, 
    2.369865e-08, 2.296616e-08, 2.277259e-08, 2.311219e-08, 2.238931e-08, 
    2.184928e-08, 2.165613e-08, 2.211404e-08, 2.128083e-08, 2.140858e-08,
  2.133394e-08, 2.294671e-08, 2.296427e-08, 2.292882e-08, 2.306173e-08, 
    2.295935e-08, 2.212351e-08, 2.229732e-08, 2.204582e-08, 2.187884e-08, 
    2.137325e-08, 2.092661e-08, 2.131937e-08, 2.08404e-08, 2.173622e-08,
  2.251778e-08, 2.390189e-08, 2.386231e-08, 2.339553e-08, 2.299808e-08, 
    2.291487e-08, 2.285863e-08, 2.234094e-08, 2.180265e-08, 2.231555e-08, 
    2.136116e-08, 2.229225e-08, 2.170213e-08, 2.181897e-08, 2.223806e-08,
  2.357166e-08, 2.429547e-08, 2.34819e-08, 2.30241e-08, 2.28912e-08, 
    2.290253e-08, 2.260383e-08, 2.221973e-08, 2.252287e-08, 2.203489e-08, 
    2.298868e-08, 2.272765e-08, 2.262097e-08, 2.177317e-08, 2.270303e-08,
  2.415856e-08, 2.394854e-08, 2.283488e-08, 2.273174e-08, 2.2724e-08, 
    2.273906e-08, 2.244961e-08, 2.244366e-08, 2.297405e-08, 2.24366e-08, 
    2.265389e-08, 2.257538e-08, 2.275076e-08, 2.201756e-08, 2.297003e-08,
  2.399557e-08, 2.353176e-08, 2.269988e-08, 2.284067e-08, 2.313336e-08, 
    2.307516e-08, 2.278114e-08, 2.282614e-08, 2.265647e-08, 2.254655e-08, 
    2.282633e-08, 2.302478e-08, 2.337409e-08, 2.287189e-08, 2.3459e-08,
  2.407936e-08, 2.386419e-08, 2.313858e-08, 2.33807e-08, 2.368185e-08, 
    2.349046e-08, 2.30017e-08, 2.305808e-08, 2.282818e-08, 2.316311e-08, 
    2.344272e-08, 2.367609e-08, 2.386356e-08, 2.368283e-08, 2.399629e-08,
  2.378631e-08, 2.348356e-08, 2.256918e-08, 2.271705e-08, 2.293576e-08, 
    2.309979e-08, 2.276254e-08, 2.297856e-08, 2.330718e-08, 2.368994e-08, 
    2.389054e-08, 2.404517e-08, 2.43177e-08, 2.455175e-08, 2.453281e-08,
  1.462342e-08, 1.636847e-08, 1.729664e-08, 1.8175e-08, 1.922526e-08, 
    2.053207e-08, 2.132608e-08, 2.251846e-08, 2.414418e-08, 2.445428e-08, 
    2.218868e-08, 2.174334e-08, 2.269211e-08, 2.177888e-08, 2.224325e-08,
  1.603879e-08, 1.711279e-08, 1.815063e-08, 1.927884e-08, 2.009905e-08, 
    2.135184e-08, 2.200994e-08, 2.361991e-08, 2.516744e-08, 2.37135e-08, 
    2.22863e-08, 2.24413e-08, 2.289645e-08, 2.20538e-08, 2.216478e-08,
  1.722479e-08, 1.775252e-08, 1.854777e-08, 1.97521e-08, 2.106483e-08, 
    2.210652e-08, 2.264697e-08, 2.432928e-08, 2.484909e-08, 2.340174e-08, 
    2.254078e-08, 2.27751e-08, 2.246563e-08, 2.22776e-08, 2.266377e-08,
  1.879536e-08, 1.87095e-08, 1.947132e-08, 2.069759e-08, 2.207339e-08, 
    2.263778e-08, 2.319818e-08, 2.440671e-08, 2.431566e-08, 2.219447e-08, 
    2.17663e-08, 2.280103e-08, 2.308173e-08, 2.343266e-08, 2.341284e-08,
  1.996846e-08, 1.979321e-08, 2.088351e-08, 2.202436e-08, 2.257839e-08, 
    2.251708e-08, 2.319848e-08, 2.355631e-08, 2.169385e-08, 1.946081e-08, 
    2.065345e-08, 2.282498e-08, 2.457756e-08, 2.377429e-08, 2.256027e-08,
  2.058249e-08, 2.099249e-08, 2.172392e-08, 2.218427e-08, 2.232604e-08, 
    2.237578e-08, 2.293842e-08, 2.200068e-08, 2.093784e-08, 1.940896e-08, 
    2.235213e-08, 2.229176e-08, 2.441571e-08, 2.428908e-08, 2.233819e-08,
  2.105864e-08, 2.185401e-08, 2.266516e-08, 2.243781e-08, 2.305296e-08, 
    2.254645e-08, 2.244321e-08, 2.137899e-08, 2.129573e-08, 2.169426e-08, 
    2.413605e-08, 2.288368e-08, 2.444008e-08, 2.445749e-08, 2.346341e-08,
  2.214026e-08, 2.286297e-08, 2.258797e-08, 2.219981e-08, 2.313835e-08, 
    2.241634e-08, 2.239703e-08, 2.215697e-08, 2.259667e-08, 2.26362e-08, 
    2.361033e-08, 2.291786e-08, 2.446516e-08, 2.416096e-08, 2.322767e-08,
  2.318019e-08, 2.310282e-08, 2.252375e-08, 2.251792e-08, 2.305423e-08, 
    2.237376e-08, 2.231729e-08, 2.173498e-08, 2.239279e-08, 2.340767e-08, 
    2.34193e-08, 2.294573e-08, 2.338417e-08, 2.356963e-08, 2.255087e-08,
  2.342488e-08, 2.297755e-08, 2.212212e-08, 2.171571e-08, 2.201176e-08, 
    2.180588e-08, 2.144553e-08, 2.270016e-08, 2.340515e-08, 2.343995e-08, 
    2.304199e-08, 2.296947e-08, 2.322495e-08, 2.270876e-08, 2.234386e-08,
  2.357694e-08, 2.340491e-08, 2.353429e-08, 2.362434e-08, 2.375948e-08, 
    2.305513e-08, 2.232741e-08, 2.235918e-08, 2.22564e-08, 2.296905e-08, 
    2.280751e-08, 2.330925e-08, 2.373586e-08, 2.319777e-08, 2.325479e-08,
  2.406349e-08, 2.315551e-08, 2.327146e-08, 2.364844e-08, 2.343616e-08, 
    2.290565e-08, 2.221744e-08, 2.224589e-08, 2.206956e-08, 2.233723e-08, 
    2.225259e-08, 2.302327e-08, 2.35526e-08, 2.382797e-08, 2.320486e-08,
  2.356197e-08, 2.1862e-08, 2.239024e-08, 2.270978e-08, 2.278397e-08, 
    2.192952e-08, 2.116488e-08, 2.15011e-08, 2.19927e-08, 2.233555e-08, 
    2.275724e-08, 2.324264e-08, 2.351111e-08, 2.384036e-08, 2.355019e-08,
  2.388964e-08, 2.271509e-08, 2.251671e-08, 2.196795e-08, 2.166453e-08, 
    2.128237e-08, 2.048182e-08, 2.060613e-08, 2.148321e-08, 2.190967e-08, 
    2.275147e-08, 2.342431e-08, 2.385299e-08, 2.493138e-08, 2.424021e-08,
  2.33598e-08, 2.210223e-08, 2.188654e-08, 2.066024e-08, 2.061032e-08, 
    2.062728e-08, 2.010302e-08, 2.007286e-08, 2.044798e-08, 2.066444e-08, 
    2.171958e-08, 2.359496e-08, 2.524429e-08, 2.506487e-08, 2.342149e-08,
  2.153972e-08, 2.13056e-08, 2.019493e-08, 1.944158e-08, 2.017724e-08, 
    2.006147e-08, 1.957059e-08, 1.935036e-08, 1.995259e-08, 2.050378e-08, 
    2.234659e-08, 2.275757e-08, 2.517305e-08, 2.579237e-08, 2.502349e-08,
  2.117407e-08, 2.13395e-08, 1.897026e-08, 1.819047e-08, 1.948299e-08, 
    1.96371e-08, 1.933253e-08, 1.967743e-08, 2.057917e-08, 2.115473e-08, 
    2.268132e-08, 2.288674e-08, 2.514406e-08, 2.668527e-08, 2.411107e-08,
  2.042411e-08, 1.86047e-08, 1.680455e-08, 1.762386e-08, 1.965897e-08, 
    1.887454e-08, 1.923252e-08, 1.942399e-08, 1.975314e-08, 2.06343e-08, 
    2.183431e-08, 2.24833e-08, 2.461308e-08, 2.559849e-08, 2.248117e-08,
  1.800854e-08, 1.759811e-08, 1.698811e-08, 1.799962e-08, 1.920801e-08, 
    1.837737e-08, 1.917863e-08, 1.906911e-08, 1.927895e-08, 2.099038e-08, 
    2.207465e-08, 2.250744e-08, 2.360487e-08, 2.32475e-08, 2.144279e-08,
  1.758838e-08, 1.864202e-08, 1.603505e-08, 1.729833e-08, 1.822265e-08, 
    1.804126e-08, 1.890316e-08, 1.998642e-08, 2.066937e-08, 2.151327e-08, 
    2.227745e-08, 2.275647e-08, 2.31232e-08, 2.122825e-08, 2.214898e-08,
  2.435388e-08, 2.455207e-08, 2.184762e-08, 2.110041e-08, 2.098672e-08, 
    2.161695e-08, 2.179102e-08, 2.358179e-08, 2.423647e-08, 2.158384e-08, 
    1.700461e-08, 1.713607e-08, 1.849121e-08, 1.634027e-08, 1.562921e-08,
  2.553496e-08, 2.349715e-08, 2.115784e-08, 2.1599e-08, 2.230891e-08, 
    2.283438e-08, 2.294034e-08, 2.457147e-08, 2.609969e-08, 2.28408e-08, 
    1.591036e-08, 1.748524e-08, 1.636961e-08, 1.534973e-08, 1.493378e-08,
  2.32046e-08, 2.107979e-08, 2.110222e-08, 2.328757e-08, 2.32905e-08, 
    2.290562e-08, 2.366324e-08, 2.410101e-08, 2.494573e-08, 2.140315e-08, 
    2.131948e-08, 2.220682e-08, 1.923936e-08, 1.714113e-08, 1.711895e-08,
  1.987023e-08, 2.080386e-08, 2.231044e-08, 2.385848e-08, 2.286768e-08, 
    2.257332e-08, 2.356847e-08, 2.261762e-08, 2.08999e-08, 2.007872e-08, 
    2.006379e-08, 2.228361e-08, 2.078087e-08, 1.833998e-08, 1.918309e-08,
  2.10055e-08, 2.07249e-08, 2.243898e-08, 2.148344e-08, 2.127827e-08, 
    2.124645e-08, 2.134938e-08, 2.125878e-08, 2.09662e-08, 1.926341e-08, 
    1.959172e-08, 1.927309e-08, 1.588115e-08, 1.547099e-08, 1.675167e-08,
  2.051659e-08, 2.139274e-08, 2.284814e-08, 2.154566e-08, 2.013774e-08, 
    2.112095e-08, 2.134541e-08, 2.136971e-08, 2.109669e-08, 1.845947e-08, 
    1.870204e-08, 1.668729e-08, 1.529341e-08, 1.621647e-08, 1.815868e-08,
  2.133015e-08, 2.278893e-08, 2.291717e-08, 2.079864e-08, 2.022084e-08, 
    2.245644e-08, 2.205345e-08, 2.15591e-08, 1.924604e-08, 1.804211e-08, 
    1.634887e-08, 1.580626e-08, 1.565505e-08, 1.640888e-08, 1.796606e-08,
  2.245069e-08, 2.313702e-08, 2.214147e-08, 2.061251e-08, 2.253221e-08, 
    2.268391e-08, 2.163271e-08, 1.867072e-08, 1.619988e-08, 1.58748e-08, 
    1.603043e-08, 1.65726e-08, 1.737626e-08, 1.80217e-08, 1.760151e-08,
  2.383023e-08, 2.338959e-08, 2.183948e-08, 2.197151e-08, 2.188315e-08, 
    2.128909e-08, 2.111907e-08, 1.903428e-08, 1.74853e-08, 1.862924e-08, 
    1.88136e-08, 1.847846e-08, 1.820472e-08, 1.751509e-08, 1.67229e-08,
  2.432887e-08, 2.443662e-08, 2.270876e-08, 2.295206e-08, 2.303247e-08, 
    2.254079e-08, 2.169526e-08, 1.961431e-08, 1.930883e-08, 1.882833e-08, 
    1.787686e-08, 1.777257e-08, 1.823439e-08, 1.669761e-08, 1.828047e-08,
  2.247859e-08, 2.323431e-08, 2.34761e-08, 2.299134e-08, 2.253119e-08, 
    2.231566e-08, 2.149216e-08, 2.207252e-08, 2.162342e-08, 2.23554e-08, 
    2.085819e-08, 2.090226e-08, 2.164299e-08, 2.16672e-08, 2.209372e-08,
  2.409909e-08, 2.376551e-08, 2.32269e-08, 2.27668e-08, 2.274028e-08, 
    2.230468e-08, 2.153496e-08, 2.211493e-08, 2.193385e-08, 2.245701e-08, 
    2.160779e-08, 2.156127e-08, 2.194667e-08, 2.192908e-08, 2.124082e-08,
  2.511022e-08, 2.333464e-08, 2.344825e-08, 2.319571e-08, 2.242511e-08, 
    2.138176e-08, 2.121389e-08, 2.128218e-08, 2.211184e-08, 2.222092e-08, 
    2.165872e-08, 2.229386e-08, 2.321901e-08, 2.402454e-08, 2.564694e-08,
  2.442488e-08, 2.298807e-08, 2.317599e-08, 2.25316e-08, 2.149544e-08, 
    2.09334e-08, 2.095829e-08, 2.125893e-08, 2.161742e-08, 2.083893e-08, 
    2.207453e-08, 2.389352e-08, 2.442802e-08, 2.661843e-08, 2.579892e-08,
  2.375822e-08, 2.311109e-08, 2.309174e-08, 2.22624e-08, 2.119779e-08, 
    2.108486e-08, 2.102676e-08, 2.134583e-08, 2.134261e-08, 2.172928e-08, 
    2.269443e-08, 2.402887e-08, 2.466697e-08, 2.50205e-08, 2.169885e-08,
  2.38384e-08, 2.327368e-08, 2.258187e-08, 2.194668e-08, 2.160082e-08, 
    2.155517e-08, 2.153455e-08, 2.178641e-08, 2.217392e-08, 2.272004e-08, 
    2.282982e-08, 2.23123e-08, 2.304e-08, 2.299145e-08, 2.099992e-08,
  2.311919e-08, 2.311815e-08, 2.264896e-08, 2.215504e-08, 2.174444e-08, 
    2.14796e-08, 2.152484e-08, 2.2198e-08, 2.261136e-08, 2.274145e-08, 
    2.259165e-08, 2.226046e-08, 2.285548e-08, 2.305861e-08, 2.02179e-08,
  2.321522e-08, 2.373117e-08, 2.26638e-08, 2.221818e-08, 2.195266e-08, 
    2.168054e-08, 2.19318e-08, 2.221399e-08, 2.262203e-08, 2.265162e-08, 
    2.21443e-08, 2.176453e-08, 2.216434e-08, 2.142037e-08, 2.011302e-08,
  2.272505e-08, 2.336743e-08, 2.256215e-08, 2.229728e-08, 2.214751e-08, 
    2.196715e-08, 2.21035e-08, 2.26805e-08, 2.299604e-08, 2.237717e-08, 
    2.215941e-08, 2.225002e-08, 2.226797e-08, 2.104585e-08, 2.040133e-08,
  2.321723e-08, 2.345653e-08, 2.259972e-08, 2.23181e-08, 2.208538e-08, 
    2.214834e-08, 2.2377e-08, 2.311707e-08, 2.261623e-08, 2.234205e-08, 
    2.27849e-08, 2.254729e-08, 2.199272e-08, 2.117275e-08, 2.033649e-08,
  2.044072e-08, 2.105591e-08, 2.086102e-08, 2.072166e-08, 2.026069e-08, 
    2.050507e-08, 2.058069e-08, 2.109019e-08, 2.079688e-08, 2.139446e-08, 
    2.152472e-08, 2.174298e-08, 2.231786e-08, 2.224299e-08, 2.202886e-08,
  2.122196e-08, 2.123155e-08, 2.006975e-08, 2.087152e-08, 2.097092e-08, 
    2.085916e-08, 2.089687e-08, 2.111395e-08, 2.062646e-08, 2.125199e-08, 
    2.133561e-08, 2.202018e-08, 2.265471e-08, 2.262968e-08, 2.264355e-08,
  2.207835e-08, 2.114978e-08, 2.030472e-08, 2.223466e-08, 2.216497e-08, 
    2.10772e-08, 2.080991e-08, 2.090331e-08, 2.084625e-08, 2.125054e-08, 
    2.153914e-08, 2.259419e-08, 2.319359e-08, 2.278177e-08, 2.331529e-08,
  1.983287e-08, 1.984849e-08, 2.09212e-08, 2.20817e-08, 2.067171e-08, 
    2.014255e-08, 2.052314e-08, 2.073826e-08, 2.121819e-08, 2.20387e-08, 
    2.363807e-08, 2.460365e-08, 2.35931e-08, 2.296907e-08, 2.41631e-08,
  1.905085e-08, 1.99788e-08, 2.077371e-08, 1.940255e-08, 1.944481e-08, 
    2.005094e-08, 2.074318e-08, 2.129516e-08, 2.251211e-08, 2.36923e-08, 
    2.429846e-08, 2.392006e-08, 2.249503e-08, 2.248001e-08, 2.427766e-08,
  1.938381e-08, 1.963049e-08, 1.929443e-08, 1.859961e-08, 1.932349e-08, 
    2.05318e-08, 2.103205e-08, 2.143513e-08, 2.21568e-08, 2.24664e-08, 
    2.255299e-08, 2.120011e-08, 2.143667e-08, 2.264973e-08, 2.183058e-08,
  1.835881e-08, 1.800184e-08, 1.808557e-08, 1.875118e-08, 2.048502e-08, 
    2.151239e-08, 2.13107e-08, 2.112908e-08, 2.177219e-08, 2.074059e-08, 
    2.070808e-08, 2.07106e-08, 2.158494e-08, 2.273515e-08, 2.116118e-08,
  1.72758e-08, 1.686706e-08, 1.814811e-08, 2.018268e-08, 2.15529e-08, 
    2.178851e-08, 2.100732e-08, 2.079291e-08, 1.999656e-08, 2.03575e-08, 
    2.08262e-08, 2.110656e-08, 2.229974e-08, 2.263052e-08, 2.174206e-08,
  1.662617e-08, 1.783893e-08, 1.945425e-08, 2.113953e-08, 2.066112e-08, 
    2.056071e-08, 2.048627e-08, 2.040409e-08, 2.002995e-08, 2.141581e-08, 
    2.171059e-08, 2.200357e-08, 2.253207e-08, 2.255255e-08, 2.236191e-08,
  1.716214e-08, 1.843326e-08, 1.989108e-08, 1.999621e-08, 1.930045e-08, 
    1.983667e-08, 2.061386e-08, 2.141078e-08, 2.171861e-08, 2.216412e-08, 
    2.2241e-08, 2.252567e-08, 2.279571e-08, 2.232995e-08, 2.277848e-08,
  2.173568e-08, 2.175221e-08, 2.141683e-08, 2.164944e-08, 2.139397e-08, 
    2.110456e-08, 2.030401e-08, 2.030844e-08, 1.985382e-08, 1.945869e-08, 
    1.942672e-08, 1.890732e-08, 1.791058e-08, 1.801743e-08, 1.878779e-08,
  2.529876e-08, 2.362892e-08, 2.253701e-08, 2.12216e-08, 2.128259e-08, 
    2.159959e-08, 2.164857e-08, 2.090743e-08, 2.013777e-08, 2.066595e-08, 
    1.993123e-08, 1.92859e-08, 1.881594e-08, 1.923113e-08, 1.912067e-08,
  2.283512e-08, 2.523607e-08, 2.315611e-08, 2.220999e-08, 2.262058e-08, 
    2.226133e-08, 2.21804e-08, 2.003454e-08, 2.040493e-08, 2.147315e-08, 
    2.116578e-08, 2.000593e-08, 2.081021e-08, 2.273586e-08, 2.206037e-08,
  2.314544e-08, 2.370889e-08, 2.320929e-08, 2.305748e-08, 2.309786e-08, 
    2.251885e-08, 2.12229e-08, 1.890657e-08, 1.99143e-08, 2.296368e-08, 
    2.471308e-08, 2.260352e-08, 2.297345e-08, 2.50363e-08, 2.345831e-08,
  2.345688e-08, 2.468763e-08, 2.428898e-08, 2.213983e-08, 2.173168e-08, 
    2.248944e-08, 2.198074e-08, 2.304032e-08, 2.178627e-08, 2.732812e-08, 
    2.530967e-08, 2.101539e-08, 2.05415e-08, 2.20846e-08, 2.257252e-08,
  2.595598e-08, 2.727175e-08, 2.746578e-08, 2.580661e-08, 2.366267e-08, 
    2.2772e-08, 2.163641e-08, 2.179239e-08, 2.385494e-08, 2.468772e-08, 
    2.00775e-08, 1.744856e-08, 1.901211e-08, 1.845451e-08, 2.277227e-08,
  2.773487e-08, 2.755859e-08, 2.818597e-08, 2.682e-08, 2.657337e-08, 
    2.537873e-08, 2.530991e-08, 2.445851e-08, 2.392313e-08, 1.96425e-08, 
    1.77753e-08, 1.922117e-08, 1.761752e-08, 1.710263e-08, 2.279037e-08,
  2.811911e-08, 2.711438e-08, 2.775498e-08, 2.706043e-08, 2.646753e-08, 
    2.604778e-08, 2.604233e-08, 2.624729e-08, 2.64765e-08, 2.463639e-08, 
    2.293901e-08, 2.151493e-08, 1.933207e-08, 2.03754e-08, 2.284808e-08,
  2.65734e-08, 2.6384e-08, 2.716603e-08, 2.677523e-08, 2.568106e-08, 
    2.652824e-08, 2.680515e-08, 2.744576e-08, 2.689779e-08, 2.579475e-08, 
    2.386747e-08, 2.394139e-08, 1.960778e-08, 1.897163e-08, 2.204669e-08,
  2.572624e-08, 2.558211e-08, 2.704431e-08, 2.612624e-08, 2.573658e-08, 
    2.554459e-08, 2.59394e-08, 2.557579e-08, 2.473395e-08, 2.517968e-08, 
    2.555132e-08, 2.46428e-08, 2.490835e-08, 2.154365e-08, 2.125105e-08,
  2.258927e-08, 2.346909e-08, 2.405786e-08, 2.428727e-08, 2.415834e-08, 
    2.394102e-08, 2.423789e-08, 2.407594e-08, 2.411028e-08, 2.317693e-08, 
    2.294853e-08, 2.269435e-08, 2.325622e-08, 2.331476e-08, 2.221701e-08,
  2.251489e-08, 2.316565e-08, 2.369274e-08, 2.329873e-08, 2.280494e-08, 
    2.254741e-08, 2.296369e-08, 2.237416e-08, 2.354715e-08, 2.363298e-08, 
    2.437578e-08, 2.402897e-08, 2.394108e-08, 2.447404e-08, 2.263296e-08,
  2.293013e-08, 2.247046e-08, 2.253312e-08, 2.184836e-08, 2.157251e-08, 
    2.225058e-08, 2.239139e-08, 2.098093e-08, 2.111398e-08, 2.163639e-08, 
    2.256417e-08, 2.30861e-08, 2.254825e-08, 2.333108e-08, 2.101886e-08,
  2.255352e-08, 2.232739e-08, 2.238704e-08, 2.284019e-08, 2.363728e-08, 
    2.430004e-08, 2.389234e-08, 2.362625e-08, 2.200538e-08, 2.19239e-08, 
    2.315962e-08, 2.310169e-08, 2.384334e-08, 2.41632e-08, 2.074677e-08,
  2.261769e-08, 2.220693e-08, 2.28541e-08, 2.370289e-08, 2.432672e-08, 
    2.477602e-08, 2.468053e-08, 2.50128e-08, 2.382634e-08, 2.597164e-08, 
    2.521166e-08, 2.361334e-08, 2.259011e-08, 2.204266e-08, 2.041712e-08,
  2.25531e-08, 2.265719e-08, 2.259816e-08, 2.3492e-08, 2.388004e-08, 
    2.441308e-08, 2.468655e-08, 2.512052e-08, 2.600939e-08, 2.699797e-08, 
    2.455066e-08, 2.417278e-08, 2.312462e-08, 2.073439e-08, 2.267639e-08,
  2.298533e-08, 2.234098e-08, 2.242205e-08, 2.332919e-08, 2.347507e-08, 
    2.376911e-08, 2.410945e-08, 2.535917e-08, 2.59152e-08, 2.558534e-08, 
    2.565904e-08, 2.572058e-08, 2.472229e-08, 2.223197e-08, 2.523157e-08,
  2.299729e-08, 2.28028e-08, 2.269986e-08, 2.320291e-08, 2.301221e-08, 
    2.3313e-08, 2.376646e-08, 2.468398e-08, 2.541513e-08, 2.530378e-08, 
    2.571205e-08, 2.558901e-08, 2.509998e-08, 2.456525e-08, 2.735811e-08,
  2.332814e-08, 2.329378e-08, 2.286078e-08, 2.322418e-08, 2.331615e-08, 
    2.389805e-08, 2.413205e-08, 2.474085e-08, 2.463338e-08, 2.471398e-08, 
    2.508902e-08, 2.555355e-08, 2.550008e-08, 2.631279e-08, 2.714527e-08,
  2.348854e-08, 2.335418e-08, 2.341668e-08, 2.339509e-08, 2.402137e-08, 
    2.471265e-08, 2.455841e-08, 2.45946e-08, 2.464315e-08, 2.473231e-08, 
    2.543988e-08, 2.520336e-08, 2.560768e-08, 2.654594e-08, 2.65687e-08,
  2.029747e-08, 2.165507e-08, 2.233156e-08, 2.258412e-08, 2.193445e-08, 
    2.197327e-08, 2.281801e-08, 2.429822e-08, 2.483254e-08, 2.588521e-08, 
    2.532985e-08, 2.387605e-08, 2.350607e-08, 2.230267e-08, 2.22495e-08,
  1.832417e-08, 2.04915e-08, 2.266282e-08, 2.365894e-08, 2.227465e-08, 
    2.242294e-08, 2.323106e-08, 2.459348e-08, 2.544421e-08, 2.549984e-08, 
    2.435585e-08, 2.372402e-08, 2.308416e-08, 2.275723e-08, 2.313766e-08,
  1.982453e-08, 2.001222e-08, 2.219817e-08, 2.367951e-08, 2.34117e-08, 
    2.243602e-08, 2.272214e-08, 2.449623e-08, 2.564002e-08, 2.48437e-08, 
    2.395423e-08, 2.406427e-08, 2.347746e-08, 2.281452e-08, 2.377887e-08,
  2.208099e-08, 2.190221e-08, 2.296514e-08, 2.336741e-08, 2.300979e-08, 
    2.314402e-08, 2.302978e-08, 2.408482e-08, 2.443502e-08, 2.327878e-08, 
    2.459849e-08, 2.57229e-08, 2.409792e-08, 2.420672e-08, 2.433554e-08,
  2.411269e-08, 2.297881e-08, 2.310989e-08, 2.371659e-08, 2.338299e-08, 
    2.340384e-08, 2.406417e-08, 2.46358e-08, 2.384963e-08, 2.247612e-08, 
    2.280875e-08, 2.411844e-08, 2.42228e-08, 2.681966e-08, 2.429847e-08,
  2.31417e-08, 2.269172e-08, 2.251459e-08, 2.33202e-08, 2.320245e-08, 
    2.35402e-08, 2.360639e-08, 2.334588e-08, 2.278006e-08, 2.221053e-08, 
    2.37747e-08, 2.382859e-08, 2.402366e-08, 2.773888e-08, 2.475525e-08,
  2.239957e-08, 2.239317e-08, 2.21372e-08, 2.291582e-08, 2.372136e-08, 
    2.396481e-08, 2.363419e-08, 2.359743e-08, 2.356482e-08, 2.40422e-08, 
    2.438291e-08, 2.360135e-08, 2.543388e-08, 2.80989e-08, 2.402037e-08,
  2.264445e-08, 2.291092e-08, 2.235641e-08, 2.351619e-08, 2.453857e-08, 
    2.529013e-08, 2.457027e-08, 2.404136e-08, 2.35476e-08, 2.407031e-08, 
    2.455962e-08, 2.483575e-08, 2.64587e-08, 2.577042e-08, 2.260885e-08,
  2.259055e-08, 2.366695e-08, 2.3016e-08, 2.365769e-08, 2.45711e-08, 
    2.489533e-08, 2.33656e-08, 2.271589e-08, 2.324235e-08, 2.508127e-08, 
    2.531796e-08, 2.525703e-08, 2.566384e-08, 2.42579e-08, 2.369999e-08,
  2.378947e-08, 2.372563e-08, 2.310689e-08, 2.28873e-08, 2.314373e-08, 
    2.319179e-08, 2.266828e-08, 2.319355e-08, 2.523531e-08, 2.541621e-08, 
    2.503308e-08, 2.51948e-08, 2.530808e-08, 2.496406e-08, 2.514039e-08,
  1.585219e-08, 1.749266e-08, 1.897334e-08, 2.005509e-08, 2.008411e-08, 
    2.084226e-08, 2.130699e-08, 2.206509e-08, 2.309542e-08, 2.215411e-08, 
    2.228048e-08, 2.217405e-08, 2.15983e-08, 1.87521e-08, 1.824185e-08,
  1.768198e-08, 1.878653e-08, 2.04366e-08, 2.108631e-08, 2.092763e-08, 
    2.167927e-08, 2.195312e-08, 2.269603e-08, 2.385075e-08, 2.336108e-08, 
    2.244253e-08, 2.248032e-08, 2.091927e-08, 1.912349e-08, 1.967834e-08,
  1.920403e-08, 2.056418e-08, 2.078964e-08, 2.205428e-08, 2.248641e-08, 
    2.215513e-08, 2.240997e-08, 2.288266e-08, 2.362304e-08, 2.31294e-08, 
    2.291929e-08, 2.338565e-08, 2.123729e-08, 1.819511e-08, 2.06538e-08,
  2.068996e-08, 2.075921e-08, 2.121608e-08, 2.216289e-08, 2.207078e-08, 
    2.148005e-08, 2.23482e-08, 2.228462e-08, 2.282053e-08, 2.183164e-08, 
    2.036324e-08, 2.037508e-08, 2.088696e-08, 2.02093e-08, 2.440447e-08,
  2.110819e-08, 2.045058e-08, 2.093077e-08, 2.165594e-08, 2.137451e-08, 
    2.16401e-08, 2.1219e-08, 2.14237e-08, 2.032501e-08, 1.669424e-08, 
    1.777878e-08, 1.989308e-08, 2.077157e-08, 2.518888e-08, 2.764935e-08,
  2.144281e-08, 2.168543e-08, 2.183304e-08, 2.158309e-08, 2.124912e-08, 
    2.064828e-08, 2.026809e-08, 1.984573e-08, 1.722844e-08, 1.790396e-08, 
    2.304606e-08, 2.373673e-08, 2.40864e-08, 2.782227e-08, 2.623623e-08,
  1.990669e-08, 2.114965e-08, 2.182602e-08, 2.099113e-08, 2.145172e-08, 
    2.139929e-08, 2.175054e-08, 2.044588e-08, 1.994756e-08, 2.223162e-08, 
    2.339702e-08, 2.307342e-08, 2.547428e-08, 2.819203e-08, 2.104114e-08,
  2.024748e-08, 2.065869e-08, 2.137176e-08, 2.179928e-08, 2.231479e-08, 
    2.358436e-08, 2.298649e-08, 2.25891e-08, 2.177376e-08, 2.287108e-08, 
    2.363015e-08, 2.440224e-08, 2.682766e-08, 2.702814e-08, 2.112723e-08,
  2.004793e-08, 2.071023e-08, 2.163032e-08, 2.210123e-08, 2.301754e-08, 
    2.309165e-08, 2.238724e-08, 2.120314e-08, 2.152117e-08, 2.381988e-08, 
    2.440898e-08, 2.462758e-08, 2.524607e-08, 2.424838e-08, 2.302132e-08,
  2.048264e-08, 2.116018e-08, 2.129782e-08, 2.150419e-08, 2.164942e-08, 
    2.110312e-08, 2.066093e-08, 2.144367e-08, 2.424641e-08, 2.490412e-08, 
    2.448776e-08, 2.457726e-08, 2.486806e-08, 2.451012e-08, 2.458018e-08,
  2.011917e-08, 1.936531e-08, 1.863661e-08, 1.867409e-08, 1.898393e-08, 
    1.885135e-08, 1.899929e-08, 1.98544e-08, 2.054788e-08, 2.145162e-08, 
    2.264986e-08, 2.456781e-08, 2.435691e-08, 2.498436e-08, 2.442687e-08,
  1.922321e-08, 1.828109e-08, 1.857985e-08, 1.906371e-08, 1.884191e-08, 
    1.892093e-08, 1.993758e-08, 2.018989e-08, 2.046895e-08, 2.06302e-08, 
    2.144712e-08, 2.16303e-08, 2.186826e-08, 2.398182e-08, 2.329755e-08,
  1.719227e-08, 1.805349e-08, 1.885348e-08, 1.916569e-08, 1.898424e-08, 
    2.007992e-08, 2.056104e-08, 2.080205e-08, 2.157945e-08, 1.995026e-08, 
    2.116336e-08, 1.993707e-08, 2.172563e-08, 2.394819e-08, 2.284914e-08,
  1.826935e-08, 1.940768e-08, 1.946778e-08, 1.932665e-08, 2.068156e-08, 
    2.082413e-08, 2.055708e-08, 2.033723e-08, 2.115261e-08, 2.225175e-08, 
    2.324193e-08, 2.061429e-08, 2.115188e-08, 2.168481e-08, 2.25826e-08,
  1.933959e-08, 2.05529e-08, 2.133512e-08, 2.150216e-08, 2.139027e-08, 
    2.165381e-08, 2.151975e-08, 2.151774e-08, 2.142065e-08, 2.204963e-08, 
    2.18136e-08, 2.057378e-08, 2.119732e-08, 2.168763e-08, 2.343139e-08,
  2.003579e-08, 2.100834e-08, 2.102729e-08, 2.099048e-08, 2.112463e-08, 
    2.170086e-08, 2.102453e-08, 1.99954e-08, 1.932486e-08, 2.003114e-08, 
    2.104577e-08, 2.01226e-08, 2.155494e-08, 2.080874e-08, 2.259326e-08,
  2.106851e-08, 2.101987e-08, 2.046789e-08, 2.083958e-08, 2.150624e-08, 
    2.111611e-08, 2.012068e-08, 1.944573e-08, 1.950056e-08, 1.890347e-08, 
    2.018828e-08, 2.056815e-08, 2.129215e-08, 2.17263e-08, 1.783485e-08,
  2.106656e-08, 2.063411e-08, 2.072135e-08, 2.126605e-08, 2.130659e-08, 
    2.060092e-08, 2.00013e-08, 1.981919e-08, 2.026527e-08, 2.002524e-08, 
    2.074335e-08, 2.055889e-08, 2.164296e-08, 2.194246e-08, 1.780181e-08,
  2.066679e-08, 2.115976e-08, 2.119567e-08, 2.163628e-08, 2.176079e-08, 
    2.111196e-08, 2.067051e-08, 2.081801e-08, 2.052299e-08, 2.04401e-08, 
    2.080853e-08, 2.094626e-08, 2.162729e-08, 2.055899e-08, 2.045914e-08,
  2.115852e-08, 2.170341e-08, 2.188442e-08, 2.228214e-08, 2.214788e-08, 
    2.167854e-08, 2.106465e-08, 2.078764e-08, 2.068853e-08, 2.048421e-08, 
    2.08351e-08, 2.073965e-08, 2.117488e-08, 2.181462e-08, 2.225539e-08,
  1.573195e-08, 1.708136e-08, 1.715985e-08, 1.753196e-08, 1.784834e-08, 
    1.830745e-08, 1.842416e-08, 1.86235e-08, 1.818438e-08, 1.891626e-08, 
    2.029356e-08, 1.997648e-08, 1.970126e-08, 1.983761e-08, 2.086208e-08,
  1.668932e-08, 1.661141e-08, 1.704717e-08, 1.726117e-08, 1.754779e-08, 
    1.767572e-08, 1.804524e-08, 1.818606e-08, 1.833429e-08, 1.909339e-08, 
    1.964861e-08, 1.948531e-08, 2.0034e-08, 2.057442e-08, 2.073412e-08,
  1.529768e-08, 1.714039e-08, 1.749337e-08, 1.756828e-08, 1.746431e-08, 
    1.82538e-08, 1.858477e-08, 1.856586e-08, 1.912443e-08, 1.945241e-08, 
    1.961745e-08, 1.946609e-08, 2.002338e-08, 2.009069e-08, 1.847943e-08,
  1.598437e-08, 1.773183e-08, 1.72007e-08, 1.724281e-08, 1.808875e-08, 
    1.820058e-08, 1.848653e-08, 1.881559e-08, 1.948873e-08, 2.01738e-08, 
    2.097517e-08, 2.146716e-08, 2.092942e-08, 1.952349e-08, 1.642401e-08,
  1.663613e-08, 1.790981e-08, 1.805404e-08, 1.83517e-08, 1.855455e-08, 
    1.868082e-08, 1.898153e-08, 1.916238e-08, 2.012865e-08, 2.143452e-08, 
    2.18429e-08, 2.052935e-08, 1.889427e-08, 1.640942e-08, 1.489373e-08,
  1.744662e-08, 1.768984e-08, 1.754186e-08, 1.752128e-08, 1.744453e-08, 
    1.804575e-08, 1.815637e-08, 1.888249e-08, 2.045571e-08, 2.07954e-08, 
    2.023266e-08, 1.766022e-08, 1.644793e-08, 1.458556e-08, 1.506911e-08,
  1.740326e-08, 1.704039e-08, 1.71917e-08, 1.70377e-08, 1.715105e-08, 
    1.802121e-08, 1.821894e-08, 1.890689e-08, 1.915473e-08, 1.808073e-08, 
    1.636555e-08, 1.546014e-08, 1.458228e-08, 1.446085e-08, 1.509296e-08,
  1.667908e-08, 1.645473e-08, 1.621102e-08, 1.60369e-08, 1.684122e-08, 
    1.763651e-08, 1.817032e-08, 1.835596e-08, 1.668251e-08, 1.605476e-08, 
    1.52386e-08, 1.49576e-08, 1.459691e-08, 1.498737e-08, 1.516196e-08,
  1.564382e-08, 1.587993e-08, 1.584369e-08, 1.643311e-08, 1.723935e-08, 
    1.729377e-08, 1.812863e-08, 1.716842e-08, 1.522983e-08, 1.579293e-08, 
    1.545387e-08, 1.517827e-08, 1.432704e-08, 1.498259e-08, 1.543859e-08,
  1.455534e-08, 1.545033e-08, 1.648285e-08, 1.632262e-08, 1.561831e-08, 
    1.608886e-08, 1.601079e-08, 1.581915e-08, 1.519739e-08, 1.53451e-08, 
    1.549433e-08, 1.521127e-08, 1.475499e-08, 1.431522e-08, 1.440362e-08,
  1.24187e-08, 1.340563e-08, 1.329027e-08, 1.386999e-08, 1.44574e-08, 
    1.505682e-08, 1.558756e-08, 1.567551e-08, 1.571493e-08, 1.596316e-08, 
    1.720098e-08, 1.632702e-08, 1.63733e-08, 1.606577e-08, 1.648097e-08,
  1.347237e-08, 1.375842e-08, 1.40278e-08, 1.443901e-08, 1.464201e-08, 
    1.513814e-08, 1.540422e-08, 1.515648e-08, 1.553525e-08, 1.572354e-08, 
    1.656831e-08, 1.586911e-08, 1.664995e-08, 1.64955e-08, 1.696532e-08,
  1.313516e-08, 1.429223e-08, 1.479135e-08, 1.479079e-08, 1.491123e-08, 
    1.563508e-08, 1.563332e-08, 1.51364e-08, 1.581353e-08, 1.54335e-08, 
    1.648825e-08, 1.599945e-08, 1.67619e-08, 1.642688e-08, 1.68031e-08,
  1.408272e-08, 1.512179e-08, 1.465194e-08, 1.483508e-08, 1.51923e-08, 
    1.544277e-08, 1.549373e-08, 1.514979e-08, 1.579968e-08, 1.534996e-08, 
    1.593012e-08, 1.650325e-08, 1.666782e-08, 1.64249e-08, 1.576413e-08,
  1.450569e-08, 1.512803e-08, 1.519488e-08, 1.511268e-08, 1.546172e-08, 
    1.58208e-08, 1.554338e-08, 1.561757e-08, 1.534553e-08, 1.460775e-08, 
    1.544256e-08, 1.609149e-08, 1.545579e-08, 1.447826e-08, 1.372109e-08,
  1.558092e-08, 1.575663e-08, 1.577762e-08, 1.56492e-08, 1.557597e-08, 
    1.5734e-08, 1.497738e-08, 1.503643e-08, 1.3377e-08, 1.401056e-08, 
    1.507227e-08, 1.513871e-08, 1.50371e-08, 1.279934e-08, 1.495239e-08,
  1.581809e-08, 1.606491e-08, 1.573773e-08, 1.581468e-08, 1.574388e-08, 
    1.572161e-08, 1.585047e-08, 1.573055e-08, 1.446201e-08, 1.485181e-08, 
    1.527098e-08, 1.573171e-08, 1.554948e-08, 1.333948e-08, 1.751988e-08,
  1.563022e-08, 1.606227e-08, 1.637919e-08, 1.610687e-08, 1.614757e-08, 
    1.635423e-08, 1.633422e-08, 1.664076e-08, 1.565634e-08, 1.6194e-08, 
    1.623616e-08, 1.670586e-08, 1.754199e-08, 1.585323e-08, 1.733601e-08,
  1.630737e-08, 1.654332e-08, 1.683097e-08, 1.672597e-08, 1.674666e-08, 
    1.671209e-08, 1.649552e-08, 1.649777e-08, 1.609775e-08, 1.668125e-08, 
    1.651193e-08, 1.713022e-08, 1.755593e-08, 1.647864e-08, 1.566538e-08,
  1.678987e-08, 1.652063e-08, 1.661844e-08, 1.670566e-08, 1.665173e-08, 
    1.645651e-08, 1.639882e-08, 1.644115e-08, 1.711284e-08, 1.700208e-08, 
    1.698263e-08, 1.708485e-08, 1.766408e-08, 1.703712e-08, 1.707038e-08,
  1.04698e-08, 1.089877e-08, 1.140526e-08, 1.180408e-08, 1.223456e-08, 
    1.26796e-08, 1.307915e-08, 1.354431e-08, 1.384504e-08, 1.405898e-08, 
    1.472398e-08, 1.497917e-08, 1.49689e-08, 1.54067e-08, 1.56277e-08,
  1.373799e-08, 1.397291e-08, 1.403231e-08, 1.406142e-08, 1.435933e-08, 
    1.431188e-08, 1.441568e-08, 1.46282e-08, 1.477957e-08, 1.500039e-08, 
    1.540864e-08, 1.556865e-08, 1.572816e-08, 1.632179e-08, 1.686245e-08,
  1.546739e-08, 1.591903e-08, 1.563439e-08, 1.594172e-08, 1.580582e-08, 
    1.579369e-08, 1.568231e-08, 1.56461e-08, 1.581877e-08, 1.604502e-08, 
    1.64757e-08, 1.637172e-08, 1.695066e-08, 1.795188e-08, 1.790806e-08,
  1.726889e-08, 1.703993e-08, 1.725849e-08, 1.748042e-08, 1.737519e-08, 
    1.72174e-08, 1.701352e-08, 1.68189e-08, 1.741301e-08, 1.780927e-08, 
    1.882306e-08, 1.850205e-08, 1.913373e-08, 1.930215e-08, 1.875847e-08,
  1.860095e-08, 1.83683e-08, 1.813789e-08, 1.795491e-08, 1.802418e-08, 
    1.817075e-08, 1.819707e-08, 1.9379e-08, 2.090727e-08, 2.095461e-08, 
    1.96582e-08, 1.899606e-08, 1.901423e-08, 1.881553e-08, 1.926358e-08,
  1.952661e-08, 2.008984e-08, 1.945292e-08, 1.938153e-08, 1.868587e-08, 
    1.849007e-08, 1.759043e-08, 1.814008e-08, 2.006446e-08, 2.066843e-08, 
    1.817337e-08, 1.857057e-08, 1.947125e-08, 1.781895e-08, 1.947461e-08,
  1.986079e-08, 1.964902e-08, 2.016314e-08, 1.974265e-08, 1.983347e-08, 
    1.962588e-08, 1.973111e-08, 2.064018e-08, 1.896393e-08, 1.716092e-08, 
    1.595306e-08, 1.82131e-08, 1.85296e-08, 1.711334e-08, 1.931963e-08,
  2.046235e-08, 2.01191e-08, 2.03494e-08, 2.014978e-08, 2.035955e-08, 
    1.977725e-08, 2.003368e-08, 2.207312e-08, 2.137141e-08, 1.958029e-08, 
    1.829163e-08, 1.904035e-08, 1.904606e-08, 1.863302e-08, 1.965046e-08,
  2.062785e-08, 2.070582e-08, 2.071223e-08, 2.041707e-08, 2.077875e-08, 
    2.058703e-08, 2.007838e-08, 2.052545e-08, 2.07593e-08, 1.875756e-08, 
    1.837932e-08, 1.911257e-08, 1.914339e-08, 1.903977e-08, 1.908498e-08,
  2.034998e-08, 2.009308e-08, 2.077359e-08, 1.984177e-08, 1.907622e-08, 
    1.960102e-08, 2.017948e-08, 1.909113e-08, 1.844236e-08, 1.788965e-08, 
    1.813087e-08, 1.819737e-08, 1.852703e-08, 1.827684e-08, 1.836498e-08,
  1.211774e-08, 1.282526e-08, 1.351429e-08, 1.43522e-08, 1.48357e-08, 
    1.520746e-08, 1.550256e-08, 1.608035e-08, 1.655176e-08, 1.601392e-08, 
    1.527855e-08, 1.590744e-08, 1.593594e-08, 1.538153e-08, 1.5357e-08,
  1.5369e-08, 1.611905e-08, 1.645661e-08, 1.680007e-08, 1.734727e-08, 
    1.715139e-08, 1.722926e-08, 1.767638e-08, 1.782026e-08, 1.748696e-08, 
    1.705575e-08, 1.724271e-08, 1.67665e-08, 1.657245e-08, 1.598183e-08,
  1.808841e-08, 1.760018e-08, 1.787802e-08, 1.84337e-08, 1.879611e-08, 
    1.8135e-08, 1.811473e-08, 1.844073e-08, 1.866886e-08, 1.846641e-08, 
    1.834361e-08, 1.776991e-08, 1.683046e-08, 1.725014e-08, 1.613111e-08,
  1.895132e-08, 1.798301e-08, 1.861283e-08, 1.902328e-08, 1.881448e-08, 
    1.866964e-08, 1.894826e-08, 1.948622e-08, 1.929629e-08, 1.953248e-08, 
    1.948801e-08, 1.766807e-08, 1.700445e-08, 1.719697e-08, 1.718753e-08,
  1.814067e-08, 1.787283e-08, 1.834694e-08, 1.849917e-08, 1.880174e-08, 
    1.910645e-08, 1.945693e-08, 1.97437e-08, 1.949316e-08, 1.846981e-08, 
    1.777152e-08, 1.692696e-08, 1.533686e-08, 1.751184e-08, 1.983214e-08,
  1.842209e-08, 1.859259e-08, 1.89128e-08, 1.924463e-08, 1.964248e-08, 
    1.976377e-08, 1.977287e-08, 1.95599e-08, 1.859501e-08, 1.907213e-08, 
    1.887092e-08, 1.733895e-08, 1.708034e-08, 1.932339e-08, 2.207136e-08,
  1.819105e-08, 1.896273e-08, 1.920748e-08, 1.947208e-08, 1.963612e-08, 
    1.990692e-08, 1.979161e-08, 1.953513e-08, 1.920164e-08, 1.906887e-08, 
    1.837432e-08, 1.863248e-08, 1.832012e-08, 1.960541e-08, 2.172931e-08,
  1.847687e-08, 1.960163e-08, 1.97252e-08, 1.977286e-08, 2.0123e-08, 
    2.0479e-08, 2.047335e-08, 2.01583e-08, 2.039605e-08, 2.081149e-08, 
    2.071685e-08, 2.007896e-08, 1.895938e-08, 1.961561e-08, 2.167452e-08,
  1.881772e-08, 1.984793e-08, 2.003809e-08, 2.040246e-08, 2.065181e-08, 
    2.071815e-08, 2.080094e-08, 2.046014e-08, 2.100094e-08, 2.185106e-08, 
    2.173151e-08, 2.175438e-08, 2.083025e-08, 2.092545e-08, 2.225902e-08,
  1.951905e-08, 2.041273e-08, 2.032203e-08, 2.074375e-08, 2.099766e-08, 
    2.10022e-08, 2.107521e-08, 2.149634e-08, 2.227925e-08, 2.273449e-08, 
    2.285978e-08, 2.269221e-08, 2.265472e-08, 2.249465e-08, 2.31064e-08,
  1.121119e-08, 1.128746e-08, 1.140444e-08, 1.170183e-08, 1.188509e-08, 
    1.196894e-08, 1.220231e-08, 1.250176e-08, 1.281223e-08, 1.301187e-08, 
    1.346035e-08, 1.408021e-08, 1.422111e-08, 1.436206e-08, 1.434897e-08,
  1.292608e-08, 1.288607e-08, 1.272585e-08, 1.266755e-08, 1.295601e-08, 
    1.311849e-08, 1.328817e-08, 1.334864e-08, 1.377459e-08, 1.414991e-08, 
    1.438363e-08, 1.49783e-08, 1.447766e-08, 1.472529e-08, 1.428379e-08,
  1.379668e-08, 1.403833e-08, 1.405731e-08, 1.402584e-08, 1.417023e-08, 
    1.444545e-08, 1.471186e-08, 1.424287e-08, 1.427294e-08, 1.485406e-08, 
    1.470555e-08, 1.522841e-08, 1.461029e-08, 1.488003e-08, 1.42259e-08,
  1.476447e-08, 1.509309e-08, 1.538644e-08, 1.5018e-08, 1.495945e-08, 
    1.469781e-08, 1.465309e-08, 1.438013e-08, 1.440569e-08, 1.469779e-08, 
    1.438447e-08, 1.339375e-08, 1.376029e-08, 1.45001e-08, 1.543861e-08,
  1.527476e-08, 1.52083e-08, 1.517958e-08, 1.43058e-08, 1.415269e-08, 
    1.4662e-08, 1.438187e-08, 1.425705e-08, 1.434669e-08, 1.458824e-08, 
    1.409484e-08, 1.391041e-08, 1.395184e-08, 1.58261e-08, 1.608364e-08,
  1.481185e-08, 1.580031e-08, 1.527614e-08, 1.493283e-08, 1.431847e-08, 
    1.426451e-08, 1.384562e-08, 1.363681e-08, 1.281075e-08, 1.340608e-08, 
    1.55218e-08, 1.50594e-08, 1.5058e-08, 1.754064e-08, 1.706887e-08,
  1.497049e-08, 1.629855e-08, 1.669812e-08, 1.605497e-08, 1.581566e-08, 
    1.537106e-08, 1.547428e-08, 1.52082e-08, 1.472198e-08, 1.551254e-08, 
    1.620569e-08, 1.550202e-08, 1.725754e-08, 1.944312e-08, 1.666389e-08,
  1.553825e-08, 1.689931e-08, 1.802032e-08, 1.784408e-08, 1.754304e-08, 
    1.743066e-08, 1.724074e-08, 1.709332e-08, 1.619711e-08, 1.723703e-08, 
    1.732281e-08, 1.756374e-08, 1.884747e-08, 1.785219e-08, 1.342101e-08,
  1.702303e-08, 1.823615e-08, 1.85468e-08, 1.932295e-08, 1.892474e-08, 
    1.87343e-08, 1.81614e-08, 1.695621e-08, 1.759459e-08, 1.911179e-08, 
    1.894708e-08, 1.891514e-08, 1.88869e-08, 1.601699e-08, 1.445902e-08,
  1.979764e-08, 1.964213e-08, 1.949596e-08, 1.994024e-08, 1.955922e-08, 
    1.887471e-08, 1.827308e-08, 1.887938e-08, 2.074421e-08, 2.085428e-08, 
    2.036714e-08, 2.01391e-08, 2.020212e-08, 1.889435e-08, 1.847898e-08,
  1.30259e-08, 1.303836e-08, 1.31724e-08, 1.356123e-08, 1.373172e-08, 
    1.388652e-08, 1.403902e-08, 1.436502e-08, 1.50589e-08, 1.435833e-08, 
    1.372998e-08, 1.433037e-08, 1.607653e-08, 1.696092e-08, 1.689243e-08,
  1.701572e-08, 1.714145e-08, 1.640927e-08, 1.616014e-08, 1.695179e-08, 
    1.687286e-08, 1.679619e-08, 1.677508e-08, 1.760977e-08, 1.674021e-08, 
    1.646679e-08, 1.714151e-08, 1.844224e-08, 1.86153e-08, 1.734076e-08,
  1.893701e-08, 1.980693e-08, 1.911115e-08, 1.895334e-08, 1.887814e-08, 
    1.871695e-08, 1.889333e-08, 1.891799e-08, 1.919578e-08, 1.795567e-08, 
    1.77425e-08, 1.918107e-08, 1.998076e-08, 1.941509e-08, 1.752799e-08,
  2.004256e-08, 2.068857e-08, 2.045912e-08, 2.043499e-08, 1.996598e-08, 
    1.994773e-08, 2.076223e-08, 2.059522e-08, 1.984321e-08, 1.889471e-08, 
    1.695602e-08, 1.815728e-08, 1.903886e-08, 1.876097e-08, 1.868592e-08,
  2.072687e-08, 2.03822e-08, 2.059087e-08, 1.970241e-08, 1.926469e-08, 
    1.951596e-08, 1.99383e-08, 1.965381e-08, 1.792011e-08, 1.582831e-08, 
    1.581088e-08, 1.770172e-08, 1.672634e-08, 1.766085e-08, 1.748482e-08,
  2.161934e-08, 2.172337e-08, 2.192099e-08, 2.105805e-08, 2.062857e-08, 
    2.013832e-08, 1.932718e-08, 1.826512e-08, 1.639394e-08, 1.61336e-08, 
    1.868332e-08, 1.840094e-08, 1.700005e-08, 1.859889e-08, 1.725198e-08,
  2.273465e-08, 2.315333e-08, 2.334484e-08, 2.294984e-08, 2.241486e-08, 
    2.196695e-08, 2.135858e-08, 2.012765e-08, 1.871741e-08, 1.981419e-08, 
    1.987801e-08, 1.854804e-08, 1.982989e-08, 2.094856e-08, 1.771565e-08,
  2.355636e-08, 2.413989e-08, 2.457266e-08, 2.424563e-08, 2.376421e-08, 
    2.354516e-08, 2.314237e-08, 2.224459e-08, 2.116851e-08, 2.125086e-08, 
    2.0729e-08, 2.051402e-08, 2.122938e-08, 2.07483e-08, 1.73303e-08,
  2.554179e-08, 2.569931e-08, 2.587504e-08, 2.573503e-08, 2.505569e-08, 
    2.470677e-08, 2.433803e-08, 2.285955e-08, 2.260364e-08, 2.284956e-08, 
    2.268591e-08, 2.197159e-08, 2.168427e-08, 2.034147e-08, 1.961398e-08,
  2.611288e-08, 2.57434e-08, 2.608312e-08, 2.614042e-08, 2.586944e-08, 
    2.553722e-08, 2.48794e-08, 2.418972e-08, 2.494747e-08, 2.432348e-08, 
    2.415596e-08, 2.299719e-08, 2.29365e-08, 2.186211e-08, 2.191321e-08,
  2.17816e-08, 2.186435e-08, 2.2063e-08, 2.212457e-08, 2.18384e-08, 
    2.161544e-08, 2.118349e-08, 2.121913e-08, 2.103843e-08, 2.057102e-08, 
    1.907648e-08, 1.852016e-08, 1.851734e-08, 1.831889e-08, 1.833027e-08,
  2.512784e-08, 2.495772e-08, 2.436186e-08, 2.394504e-08, 2.370619e-08, 
    2.325656e-08, 2.275817e-08, 2.252527e-08, 2.250727e-08, 2.170236e-08, 
    2.080491e-08, 2.023338e-08, 2.041015e-08, 2.044122e-08, 2.062237e-08,
  2.542491e-08, 2.463163e-08, 2.410004e-08, 2.419224e-08, 2.391368e-08, 
    2.353743e-08, 2.362028e-08, 2.318273e-08, 2.307554e-08, 2.257852e-08, 
    2.190908e-08, 2.195176e-08, 2.254979e-08, 2.302243e-08, 2.306862e-08,
  2.46454e-08, 2.410428e-08, 2.400287e-08, 2.456078e-08, 2.48731e-08, 
    2.479644e-08, 2.491559e-08, 2.463775e-08, 2.474571e-08, 2.38984e-08, 
    2.354865e-08, 2.331617e-08, 2.406313e-08, 2.544997e-08, 2.626891e-08,
  2.411008e-08, 2.371494e-08, 2.397195e-08, 2.422392e-08, 2.435964e-08, 
    2.459154e-08, 2.475432e-08, 2.472248e-08, 2.476021e-08, 2.513204e-08, 
    2.444969e-08, 2.374802e-08, 2.324323e-08, 2.402829e-08, 2.5314e-08,
  2.523663e-08, 2.478476e-08, 2.477015e-08, 2.489574e-08, 2.484502e-08, 
    2.471304e-08, 2.470161e-08, 2.470329e-08, 2.481149e-08, 2.494755e-08, 
    2.416458e-08, 2.471304e-08, 2.352096e-08, 2.429854e-08, 2.48848e-08,
  2.424345e-08, 2.435916e-08, 2.420771e-08, 2.440823e-08, 2.426507e-08, 
    2.428107e-08, 2.412141e-08, 2.430484e-08, 2.422387e-08, 2.454718e-08, 
    2.442124e-08, 2.425522e-08, 2.373138e-08, 2.34035e-08, 2.426243e-08,
  2.421546e-08, 2.430407e-08, 2.410938e-08, 2.423235e-08, 2.394893e-08, 
    2.399516e-08, 2.404235e-08, 2.427252e-08, 2.473131e-08, 2.43826e-08, 
    2.474708e-08, 2.426224e-08, 2.398109e-08, 2.415583e-08, 2.518094e-08,
  2.429083e-08, 2.357151e-08, 2.337617e-08, 2.325514e-08, 2.317585e-08, 
    2.369972e-08, 2.421751e-08, 2.47025e-08, 2.518914e-08, 2.492393e-08, 
    2.559044e-08, 2.530805e-08, 2.541272e-08, 2.527768e-08, 2.614681e-08,
  2.296841e-08, 2.162147e-08, 2.121315e-08, 2.131653e-08, 2.143332e-08, 
    2.193612e-08, 2.254346e-08, 2.294322e-08, 2.416863e-08, 2.464928e-08, 
    2.572773e-08, 2.552081e-08, 2.617828e-08, 2.629829e-08, 2.63495e-08,
  1.994002e-08, 2.058291e-08, 2.118754e-08, 2.224219e-08, 2.26418e-08, 
    2.251946e-08, 2.274662e-08, 2.27474e-08, 2.270703e-08, 2.180631e-08, 
    1.905673e-08, 1.971185e-08, 2.050246e-08, 2.05601e-08, 2.008626e-08,
  2.262432e-08, 2.35146e-08, 2.29809e-08, 2.32564e-08, 2.417451e-08, 
    2.303491e-08, 2.261974e-08, 2.228815e-08, 2.193367e-08, 2.106802e-08, 
    1.969153e-08, 1.937501e-08, 1.983209e-08, 1.931305e-08, 1.964184e-08,
  2.505137e-08, 2.388197e-08, 2.306433e-08, 2.262854e-08, 2.271448e-08, 
    2.172154e-08, 2.117708e-08, 2.159886e-08, 2.12694e-08, 2.031699e-08, 
    1.996052e-08, 2.017275e-08, 2.053876e-08, 1.956484e-08, 2.066115e-08,
  2.392933e-08, 2.164685e-08, 2.192088e-08, 2.207224e-08, 2.124786e-08, 
    2.110961e-08, 2.180479e-08, 2.245365e-08, 2.191007e-08, 2.098976e-08, 
    1.968526e-08, 2.031904e-08, 2.133134e-08, 2.143312e-08, 2.325492e-08,
  2.186894e-08, 2.104493e-08, 2.141881e-08, 2.135159e-08, 2.150851e-08, 
    2.18605e-08, 2.265547e-08, 2.292111e-08, 2.259609e-08, 2.095495e-08, 
    2.067796e-08, 2.220112e-08, 2.307819e-08, 2.394125e-08, 2.500323e-08,
  2.315029e-08, 2.383397e-08, 2.400355e-08, 2.449621e-08, 2.491032e-08, 
    2.484238e-08, 2.474369e-08, 2.468049e-08, 2.390223e-08, 2.342306e-08, 
    2.526068e-08, 2.489674e-08, 2.491895e-08, 2.49167e-08, 2.508049e-08,
  2.468028e-08, 2.511167e-08, 2.526232e-08, 2.548222e-08, 2.540456e-08, 
    2.550701e-08, 2.512844e-08, 2.521063e-08, 2.491383e-08, 2.512122e-08, 
    2.500889e-08, 2.443845e-08, 2.448362e-08, 2.407019e-08, 2.36003e-08,
  2.585801e-08, 2.5947e-08, 2.607823e-08, 2.589607e-08, 2.592904e-08, 
    2.581464e-08, 2.566848e-08, 2.535486e-08, 2.4609e-08, 2.370755e-08, 
    2.310874e-08, 2.210643e-08, 2.16515e-08, 2.142129e-08, 2.131879e-08,
  2.698837e-08, 2.64746e-08, 2.588222e-08, 2.492438e-08, 2.342704e-08, 
    2.231315e-08, 2.149814e-08, 2.025448e-08, 1.95214e-08, 1.918106e-08, 
    1.910671e-08, 1.887413e-08, 1.915704e-08, 1.919289e-08, 1.952356e-08,
  2.493324e-08, 2.294521e-08, 2.128482e-08, 1.97329e-08, 1.861213e-08, 
    1.831669e-08, 1.787499e-08, 1.808757e-08, 1.868376e-08, 1.885004e-08, 
    1.926442e-08, 1.947208e-08, 1.997408e-08, 2.031354e-08, 2.056488e-08,
  2.200248e-08, 2.337273e-08, 2.446432e-08, 2.522335e-08, 2.528122e-08, 
    2.572539e-08, 2.59603e-08, 2.648117e-08, 2.693719e-08, 2.652154e-08, 
    2.51582e-08, 2.560617e-08, 2.592593e-08, 2.520931e-08, 2.494592e-08,
  2.612176e-08, 2.758997e-08, 2.688481e-08, 2.664263e-08, 2.754745e-08, 
    2.743396e-08, 2.749752e-08, 2.797227e-08, 2.835975e-08, 2.833857e-08, 
    2.723303e-08, 2.729085e-08, 2.708941e-08, 2.60844e-08, 2.644431e-08,
  2.852362e-08, 2.849423e-08, 2.788495e-08, 2.844425e-08, 2.855776e-08, 
    2.923402e-08, 2.887901e-08, 2.934689e-08, 2.932122e-08, 2.926275e-08, 
    2.817403e-08, 2.793379e-08, 2.695253e-08, 2.661116e-08, 2.675052e-08,
  2.888541e-08, 2.833787e-08, 2.880458e-08, 2.931458e-08, 2.916074e-08, 
    2.956091e-08, 2.930752e-08, 2.93114e-08, 2.866289e-08, 2.784603e-08, 
    2.697458e-08, 2.776011e-08, 2.710313e-08, 2.665602e-08, 2.543665e-08,
  2.777583e-08, 2.794028e-08, 2.824008e-08, 2.82308e-08, 2.833998e-08, 
    2.761256e-08, 2.760888e-08, 2.68788e-08, 2.63451e-08, 2.545078e-08, 
    2.486436e-08, 2.462601e-08, 2.342636e-08, 2.289733e-08, 2.206305e-08,
  2.831415e-08, 2.785756e-08, 2.700211e-08, 2.654207e-08, 2.537419e-08, 
    2.463075e-08, 2.367187e-08, 2.299543e-08, 2.2049e-08, 2.127026e-08, 
    2.021205e-08, 1.982739e-08, 1.979863e-08, 1.948394e-08, 2.025697e-08,
  2.607133e-08, 2.431681e-08, 2.312871e-08, 2.156664e-08, 2.033971e-08, 
    1.93894e-08, 1.847029e-08, 1.81381e-08, 1.769097e-08, 1.755219e-08, 
    1.782835e-08, 1.811023e-08, 1.848877e-08, 1.86394e-08, 1.982288e-08,
  2.191534e-08, 2.062261e-08, 1.90168e-08, 1.776791e-08, 1.680587e-08, 
    1.642211e-08, 1.630712e-08, 1.698364e-08, 1.701371e-08, 1.730935e-08, 
    1.775729e-08, 1.826539e-08, 1.905711e-08, 1.973398e-08, 2.094918e-08,
  1.773886e-08, 1.685802e-08, 1.582447e-08, 1.597421e-08, 1.61454e-08, 
    1.683819e-08, 1.740666e-08, 1.834878e-08, 1.853248e-08, 1.897803e-08, 
    1.971272e-08, 1.98934e-08, 2.004628e-08, 2.062263e-08, 2.052765e-08,
  1.561003e-08, 1.557391e-08, 1.65421e-08, 1.775718e-08, 1.889979e-08, 
    2.026085e-08, 2.098052e-08, 2.185504e-08, 2.208413e-08, 2.205874e-08, 
    2.214041e-08, 2.186407e-08, 2.178187e-08, 2.180895e-08, 2.178844e-08,
  2.532615e-08, 2.472038e-08, 2.478026e-08, 2.497118e-08, 2.496289e-08, 
    2.457613e-08, 2.441083e-08, 2.417588e-08, 2.401856e-08, 2.358204e-08, 
    2.364964e-08, 2.346459e-08, 2.37852e-08, 2.329356e-08, 2.319819e-08,
  2.470167e-08, 2.431136e-08, 2.464216e-08, 2.425775e-08, 2.373351e-08, 
    2.308998e-08, 2.29438e-08, 2.254112e-08, 2.232343e-08, 2.169682e-08, 
    2.212425e-08, 2.158344e-08, 2.197785e-08, 2.148008e-08, 2.169362e-08,
  2.461203e-08, 2.214161e-08, 2.23573e-08, 2.13598e-08, 2.025545e-08, 
    2.04399e-08, 2.011066e-08, 1.983724e-08, 1.958987e-08, 1.939836e-08, 
    1.912272e-08, 1.916283e-08, 1.922505e-08, 1.93677e-08, 1.924884e-08,
  2.386125e-08, 2.187815e-08, 2.033366e-08, 1.965628e-08, 2.055885e-08, 
    2.022649e-08, 1.941786e-08, 1.952277e-08, 1.945467e-08, 1.934685e-08, 
    2.147735e-08, 2.194662e-08, 2.084583e-08, 2.083289e-08, 1.96384e-08,
  2.15156e-08, 2.131274e-08, 2.140057e-08, 2.097313e-08, 2.097618e-08, 
    2.103919e-08, 2.108802e-08, 2.079828e-08, 2.180845e-08, 2.338279e-08, 
    2.330653e-08, 2.257294e-08, 2.199284e-08, 2.174147e-08, 2.013275e-08,
  2.133538e-08, 2.163045e-08, 2.156396e-08, 2.177988e-08, 2.21929e-08, 
    2.26872e-08, 2.248692e-08, 2.310948e-08, 2.455975e-08, 2.437448e-08, 
    2.283476e-08, 2.252266e-08, 2.498065e-08, 2.217806e-08, 2.131568e-08,
  2.270103e-08, 2.293706e-08, 2.292693e-08, 2.30271e-08, 2.311987e-08, 
    2.392156e-08, 2.434033e-08, 2.506787e-08, 2.563585e-08, 2.446947e-08, 
    2.454661e-08, 2.455139e-08, 2.437756e-08, 2.206933e-08, 2.39916e-08,
  2.363992e-08, 2.353035e-08, 2.392948e-08, 2.402355e-08, 2.367049e-08, 
    2.428624e-08, 2.480604e-08, 2.538456e-08, 2.625379e-08, 2.539074e-08, 
    2.512641e-08, 2.479151e-08, 2.4359e-08, 2.489618e-08, 2.644871e-08,
  2.497741e-08, 2.463231e-08, 2.50466e-08, 2.52461e-08, 2.485602e-08, 
    2.518385e-08, 2.686586e-08, 2.810647e-08, 2.684675e-08, 2.481983e-08, 
    2.488943e-08, 2.474589e-08, 2.454173e-08, 2.636552e-08, 2.561627e-08,
  2.590062e-08, 2.615981e-08, 2.643693e-08, 2.640077e-08, 2.672183e-08, 
    2.685417e-08, 2.726289e-08, 2.680393e-08, 2.479424e-08, 2.521718e-08, 
    2.529234e-08, 2.477928e-08, 2.461256e-08, 2.510884e-08, 2.475316e-08,
  2.506599e-08, 2.412903e-08, 2.403062e-08, 2.26739e-08, 2.139878e-08, 
    2.218206e-08, 2.44981e-08, 2.578752e-08, 2.450821e-08, 2.357167e-08, 
    2.362221e-08, 2.415453e-08, 2.365443e-08, 2.250397e-08, 2.291172e-08,
  2.48394e-08, 2.45653e-08, 2.426426e-08, 2.214591e-08, 2.088755e-08, 
    2.278135e-08, 2.458452e-08, 2.521425e-08, 2.44954e-08, 2.315826e-08, 
    2.360667e-08, 2.348935e-08, 2.29229e-08, 2.273764e-08, 2.421995e-08,
  2.543762e-08, 2.484965e-08, 2.336521e-08, 2.122358e-08, 2.193546e-08, 
    2.332279e-08, 2.379707e-08, 2.445979e-08, 2.390996e-08, 2.406172e-08, 
    2.466036e-08, 2.281733e-08, 2.228511e-08, 2.393878e-08, 2.384304e-08,
  2.697292e-08, 2.601564e-08, 2.256575e-08, 2.073074e-08, 2.199244e-08, 
    2.343698e-08, 2.34511e-08, 2.300322e-08, 2.392087e-08, 2.475274e-08, 
    2.450165e-08, 2.333807e-08, 2.37045e-08, 2.517067e-08, 2.233275e-08,
  2.856417e-08, 2.702791e-08, 2.268719e-08, 2.065196e-08, 2.115458e-08, 
    2.302686e-08, 2.314134e-08, 2.247419e-08, 2.375821e-08, 2.196849e-08, 
    2.03435e-08, 2.245575e-08, 2.573011e-08, 2.375711e-08, 2.163044e-08,
  2.761409e-08, 2.585159e-08, 2.017453e-08, 1.970095e-08, 2.107708e-08, 
    2.216036e-08, 2.160289e-08, 2.068353e-08, 2.108272e-08, 1.956284e-08, 
    2.141378e-08, 2.236577e-08, 2.455653e-08, 2.366352e-08, 2.351486e-08,
  2.786578e-08, 2.57983e-08, 2.003651e-08, 2.037245e-08, 2.107808e-08, 
    2.216493e-08, 2.236243e-08, 2.1687e-08, 2.1609e-08, 2.084928e-08, 
    2.229809e-08, 2.225949e-08, 2.408211e-08, 2.472308e-08, 2.380182e-08,
  2.724586e-08, 2.232593e-08, 2.060206e-08, 2.079858e-08, 2.17898e-08, 
    2.302305e-08, 2.338052e-08, 2.15931e-08, 2.02408e-08, 2.083534e-08, 
    2.175985e-08, 2.23911e-08, 2.394799e-08, 2.452504e-08, 2.260354e-08,
  2.646089e-08, 2.526658e-08, 2.338785e-08, 2.156236e-08, 2.259157e-08, 
    2.456349e-08, 2.238039e-08, 2.096018e-08, 1.993542e-08, 2.201116e-08, 
    2.25531e-08, 2.249349e-08, 2.279009e-08, 2.221657e-08, 2.156031e-08,
  2.825159e-08, 2.95687e-08, 2.463408e-08, 2.115074e-08, 2.17077e-08, 
    2.329764e-08, 2.046359e-08, 2.076491e-08, 2.178454e-08, 2.247804e-08, 
    2.19278e-08, 2.220056e-08, 2.23411e-08, 2.178262e-08, 2.248464e-08,
  2.878475e-08, 3.179925e-08, 3.241272e-08, 3.293551e-08, 3.777227e-08, 
    3.715028e-08, 3.30983e-08, 3.453431e-08, 3.189934e-08, 2.633017e-08, 
    1.965348e-08, 1.668451e-08, 1.795594e-08, 1.744533e-08, 1.751845e-08,
  2.983997e-08, 3.225072e-08, 3.398625e-08, 3.51214e-08, 3.735551e-08, 
    3.491486e-08, 3.261113e-08, 3.464588e-08, 3.027972e-08, 2.495536e-08, 
    1.987009e-08, 1.986461e-08, 2.045551e-08, 1.746107e-08, 1.779971e-08,
  3.253083e-08, 3.356718e-08, 3.398226e-08, 3.568327e-08, 3.63819e-08, 
    3.251734e-08, 2.964694e-08, 2.721069e-08, 2.449106e-08, 2.323753e-08, 
    2.47023e-08, 2.279861e-08, 2.065948e-08, 1.668215e-08, 1.976215e-08,
  3.081106e-08, 3.148327e-08, 3.334498e-08, 3.284145e-08, 3.12597e-08, 
    2.831273e-08, 2.581406e-08, 2.277162e-08, 2.147735e-08, 2.154645e-08, 
    1.783689e-08, 1.726984e-08, 1.807429e-08, 1.963209e-08, 2.331348e-08,
  3.107448e-08, 3.205464e-08, 3.185741e-08, 2.954573e-08, 2.868448e-08, 
    2.473046e-08, 2.199658e-08, 1.965494e-08, 2.012348e-08, 1.760286e-08, 
    1.690665e-08, 1.903477e-08, 2.164049e-08, 2.401458e-08, 2.379605e-08,
  3.261094e-08, 3.283894e-08, 3.232404e-08, 3.009348e-08, 2.807788e-08, 
    2.39327e-08, 2.130888e-08, 2.06935e-08, 2.04953e-08, 2.044688e-08, 
    2.247954e-08, 2.25902e-08, 2.291602e-08, 2.489075e-08, 2.389427e-08,
  3.487046e-08, 3.415972e-08, 3.204877e-08, 3.051043e-08, 2.646706e-08, 
    2.218317e-08, 2.0703e-08, 2.216102e-08, 2.186503e-08, 2.189478e-08, 
    2.263053e-08, 2.22843e-08, 2.409359e-08, 2.513636e-08, 2.408918e-08,
  3.507091e-08, 3.36191e-08, 3.171234e-08, 2.887135e-08, 2.590607e-08, 
    2.329565e-08, 2.348331e-08, 2.309164e-08, 2.198955e-08, 2.24377e-08, 
    2.280006e-08, 2.298668e-08, 2.447023e-08, 2.378747e-08, 2.222751e-08,
  3.535028e-08, 3.336883e-08, 3.114055e-08, 2.769034e-08, 2.521686e-08, 
    2.425903e-08, 2.355053e-08, 2.256335e-08, 2.224741e-08, 2.284318e-08, 
    2.324115e-08, 2.32347e-08, 2.339898e-08, 2.237455e-08, 2.213257e-08,
  3.541971e-08, 3.257662e-08, 2.981181e-08, 2.60393e-08, 2.406925e-08, 
    2.455399e-08, 2.390929e-08, 2.328039e-08, 2.309344e-08, 2.333735e-08, 
    2.353004e-08, 2.349083e-08, 2.338881e-08, 2.278351e-08, 2.296536e-08,
  2.242053e-08, 2.275705e-08, 2.317621e-08, 2.328715e-08, 2.385746e-08, 
    2.559538e-08, 2.614751e-08, 2.755881e-08, 2.867329e-08, 2.697774e-08, 
    2.458547e-08, 2.569331e-08, 2.511368e-08, 2.521761e-08, 2.535264e-08,
  2.252396e-08, 2.259142e-08, 2.305685e-08, 2.357693e-08, 2.452884e-08, 
    2.541062e-08, 2.520428e-08, 2.726431e-08, 2.852464e-08, 2.623599e-08, 
    2.574232e-08, 2.647867e-08, 2.510356e-08, 2.569858e-08, 2.467381e-08,
  2.304576e-08, 2.267852e-08, 2.284174e-08, 2.342106e-08, 2.494932e-08, 
    2.491965e-08, 2.490912e-08, 2.679713e-08, 2.775252e-08, 2.649392e-08, 
    2.727023e-08, 2.597194e-08, 2.517386e-08, 2.573846e-08, 2.439765e-08,
  2.282655e-08, 2.282166e-08, 2.318532e-08, 2.365919e-08, 2.458876e-08, 
    2.479599e-08, 2.484322e-08, 2.641959e-08, 2.749837e-08, 2.59062e-08, 
    2.705185e-08, 2.489833e-08, 2.63862e-08, 2.508938e-08, 2.265454e-08,
  2.282757e-08, 2.285728e-08, 2.323481e-08, 2.380127e-08, 2.462903e-08, 
    2.49928e-08, 2.554432e-08, 2.684436e-08, 2.632649e-08, 2.452066e-08, 
    2.342043e-08, 2.481581e-08, 2.951567e-08, 2.408981e-08, 2.298985e-08,
  2.2503e-08, 2.245462e-08, 2.261513e-08, 2.332249e-08, 2.430086e-08, 
    2.481301e-08, 2.559471e-08, 2.676799e-08, 2.537946e-08, 2.344983e-08, 
    2.468563e-08, 2.593646e-08, 2.741064e-08, 2.532722e-08, 2.600351e-08,
  2.214932e-08, 2.229056e-08, 2.265938e-08, 2.320018e-08, 2.399791e-08, 
    2.425466e-08, 2.50558e-08, 2.550835e-08, 2.437928e-08, 2.426082e-08, 
    2.60512e-08, 2.523078e-08, 2.712985e-08, 2.736194e-08, 2.608749e-08,
  2.208326e-08, 2.231649e-08, 2.257618e-08, 2.311834e-08, 2.375731e-08, 
    2.414346e-08, 2.498964e-08, 2.549557e-08, 2.472822e-08, 2.461226e-08, 
    2.537844e-08, 2.541612e-08, 2.726943e-08, 2.86677e-08, 2.452086e-08,
  2.203994e-08, 2.224667e-08, 2.255155e-08, 2.31411e-08, 2.394982e-08, 
    2.417495e-08, 2.459056e-08, 2.501352e-08, 2.458602e-08, 2.475498e-08, 
    2.504162e-08, 2.478878e-08, 2.617013e-08, 2.552342e-08, 2.338441e-08,
  2.220568e-08, 2.231838e-08, 2.251727e-08, 2.293833e-08, 2.376994e-08, 
    2.400439e-08, 2.416709e-08, 2.492563e-08, 2.536275e-08, 2.5193e-08, 
    2.516535e-08, 2.496681e-08, 2.533326e-08, 2.452546e-08, 2.440701e-08,
  1.939704e-08, 2.024908e-08, 2.078011e-08, 2.124035e-08, 2.118919e-08, 
    2.125984e-08, 2.128418e-08, 2.171625e-08, 2.282371e-08, 2.409415e-08, 
    2.301097e-08, 2.369922e-08, 2.355568e-08, 2.32541e-08, 2.259097e-08,
  2.047836e-08, 2.115691e-08, 2.11827e-08, 2.138515e-08, 2.148865e-08, 
    2.189722e-08, 2.185777e-08, 2.246483e-08, 2.337364e-08, 2.364255e-08, 
    2.299197e-08, 2.283925e-08, 2.369476e-08, 2.316194e-08, 2.135027e-08,
  2.172427e-08, 2.128532e-08, 2.12479e-08, 2.18917e-08, 2.224975e-08, 
    2.239499e-08, 2.204441e-08, 2.255508e-08, 2.311996e-08, 2.343138e-08, 
    2.332287e-08, 2.290237e-08, 2.347744e-08, 2.191513e-08, 2.132536e-08,
  2.131195e-08, 2.042019e-08, 2.099743e-08, 2.209319e-08, 2.201964e-08, 
    2.221015e-08, 2.245138e-08, 2.252778e-08, 2.280306e-08, 2.244655e-08, 
    2.180859e-08, 2.16415e-08, 2.252009e-08, 2.19704e-08, 2.317923e-08,
  2.054414e-08, 2.079264e-08, 2.134858e-08, 2.139399e-08, 2.158515e-08, 
    2.162903e-08, 2.165e-08, 2.173864e-08, 2.151932e-08, 2.057828e-08, 
    2.110881e-08, 2.205753e-08, 2.289497e-08, 2.229278e-08, 2.318125e-08,
  2.147829e-08, 2.107733e-08, 2.121857e-08, 2.148014e-08, 2.146326e-08, 
    2.128287e-08, 2.111038e-08, 2.093697e-08, 2.117334e-08, 2.163604e-08, 
    2.232708e-08, 2.168536e-08, 2.220401e-08, 2.422479e-08, 2.380225e-08,
  2.105039e-08, 2.101494e-08, 2.124257e-08, 2.123606e-08, 2.118697e-08, 
    2.135654e-08, 2.125537e-08, 2.13687e-08, 2.191902e-08, 2.220768e-08, 
    2.166469e-08, 2.098649e-08, 2.248448e-08, 2.51874e-08, 2.184485e-08,
  2.035427e-08, 2.057831e-08, 2.090847e-08, 2.096961e-08, 2.139342e-08, 
    2.183475e-08, 2.163163e-08, 2.139685e-08, 2.099872e-08, 2.076172e-08, 
    2.061152e-08, 2.10423e-08, 2.30036e-08, 2.377291e-08, 2.164827e-08,
  2.055904e-08, 2.05579e-08, 2.071382e-08, 2.100481e-08, 2.138307e-08, 
    2.194382e-08, 2.140943e-08, 2.080394e-08, 2.017556e-08, 2.083654e-08, 
    2.101905e-08, 2.118085e-08, 2.199861e-08, 2.186009e-08, 2.082215e-08,
  2.031275e-08, 2.046815e-08, 2.091228e-08, 2.117377e-08, 2.13884e-08, 
    2.133712e-08, 2.017612e-08, 2.026936e-08, 2.119217e-08, 2.110413e-08, 
    2.085211e-08, 2.104197e-08, 2.156634e-08, 2.119695e-08, 2.160221e-08,
  2.177839e-08, 2.220986e-08, 2.210689e-08, 2.325279e-08, 2.345728e-08, 
    2.381634e-08, 2.321343e-08, 2.255582e-08, 2.24598e-08, 2.139941e-08, 
    2.085508e-08, 2.107113e-08, 2.205947e-08, 2.309122e-08, 2.180457e-08,
  2.256955e-08, 2.364646e-08, 2.26011e-08, 2.324701e-08, 2.444332e-08, 
    2.454144e-08, 2.306128e-08, 2.286143e-08, 2.216761e-08, 2.108054e-08, 
    2.13693e-08, 2.235316e-08, 2.27427e-08, 2.179798e-08, 1.990433e-08,
  2.321271e-08, 2.445963e-08, 2.40013e-08, 2.393723e-08, 2.478076e-08, 
    2.377441e-08, 2.204098e-08, 2.224771e-08, 2.125398e-08, 2.112547e-08, 
    2.126172e-08, 2.254466e-08, 2.153434e-08, 1.98127e-08, 2.013788e-08,
  2.297875e-08, 2.324552e-08, 2.278448e-08, 2.344673e-08, 2.253918e-08, 
    2.230112e-08, 2.234573e-08, 2.210349e-08, 2.051246e-08, 2.166015e-08, 
    1.849125e-08, 1.707042e-08, 1.895476e-08, 1.957611e-08, 2.150422e-08,
  2.31858e-08, 2.31682e-08, 2.288398e-08, 2.19166e-08, 2.24043e-08, 
    2.258401e-08, 2.290744e-08, 2.224796e-08, 2.14944e-08, 2.131082e-08, 
    2.000913e-08, 2.100582e-08, 2.248919e-08, 2.251566e-08, 2.272125e-08,
  2.396867e-08, 2.332016e-08, 2.288817e-08, 2.283529e-08, 2.305778e-08, 
    2.297934e-08, 2.282476e-08, 2.300939e-08, 2.034225e-08, 1.80268e-08, 
    2.340218e-08, 2.222406e-08, 2.122875e-08, 2.040042e-08, 2.135612e-08,
  2.407429e-08, 2.352227e-08, 2.333608e-08, 2.356372e-08, 2.347527e-08, 
    2.348794e-08, 2.300896e-08, 2.342815e-08, 2.205059e-08, 2.029726e-08, 
    2.011151e-08, 1.928979e-08, 2.0396e-08, 2.077985e-08, 2.048336e-08,
  2.399107e-08, 2.321175e-08, 2.318785e-08, 2.314509e-08, 2.306175e-08, 
    2.297716e-08, 2.275325e-08, 2.278287e-08, 2.119098e-08, 2.138308e-08, 
    2.101637e-08, 2.101692e-08, 2.158982e-08, 2.149351e-08, 2.01954e-08,
  2.442852e-08, 2.247187e-08, 2.195534e-08, 2.226844e-08, 2.219284e-08, 
    2.250046e-08, 2.240086e-08, 2.200478e-08, 2.076356e-08, 2.165973e-08, 
    2.159212e-08, 2.180601e-08, 2.194983e-08, 2.180479e-08, 2.099011e-08,
  2.546757e-08, 2.158656e-08, 2.132716e-08, 2.150971e-08, 2.136209e-08, 
    2.150033e-08, 2.128123e-08, 2.17354e-08, 2.277914e-08, 2.28547e-08, 
    2.253417e-08, 2.269891e-08, 2.278043e-08, 2.253405e-08, 2.230902e-08,
  2.404854e-08, 2.506537e-08, 2.643878e-08, 2.676202e-08, 2.63135e-08, 
    2.495924e-08, 2.437831e-08, 2.423105e-08, 2.379269e-08, 2.326645e-08, 
    2.436228e-08, 2.457515e-08, 2.482892e-08, 2.490918e-08, 2.462535e-08,
  2.422846e-08, 2.589051e-08, 2.73697e-08, 2.682656e-08, 2.566417e-08, 
    2.433703e-08, 2.350514e-08, 2.319315e-08, 2.1953e-08, 2.228795e-08, 
    2.360174e-08, 2.394992e-08, 2.443558e-08, 2.391993e-08, 2.376088e-08,
  2.55543e-08, 2.671513e-08, 2.651839e-08, 2.542639e-08, 2.393219e-08, 
    2.295027e-08, 2.177004e-08, 2.138937e-08, 2.093157e-08, 2.188136e-08, 
    2.296944e-08, 2.383948e-08, 2.43824e-08, 2.348379e-08, 2.465964e-08,
  2.609103e-08, 2.702801e-08, 2.615873e-08, 2.446919e-08, 2.296521e-08, 
    2.195297e-08, 2.075409e-08, 2.05471e-08, 2.039714e-08, 2.160587e-08, 
    2.11821e-08, 2.248734e-08, 2.348709e-08, 2.307099e-08, 2.310742e-08,
  2.773626e-08, 2.721177e-08, 2.53889e-08, 2.349329e-08, 2.205833e-08, 
    2.085255e-08, 2.03529e-08, 2.004616e-08, 2.077216e-08, 2.088858e-08, 
    2.090321e-08, 2.323293e-08, 2.302267e-08, 2.230591e-08, 2.283386e-08,
  2.77489e-08, 2.63679e-08, 2.453894e-08, 2.368658e-08, 2.191062e-08, 
    2.076671e-08, 2.002758e-08, 2.013157e-08, 2.022639e-08, 2.071948e-08, 
    2.231822e-08, 2.229702e-08, 2.275865e-08, 2.176023e-08, 2.527178e-08,
  2.800897e-08, 2.555814e-08, 2.461897e-08, 2.36469e-08, 2.093933e-08, 
    1.999953e-08, 1.941096e-08, 2.023076e-08, 1.980483e-08, 2.07032e-08, 
    2.124517e-08, 2.17977e-08, 2.225841e-08, 2.227172e-08, 2.527684e-08,
  2.782233e-08, 2.575043e-08, 2.513685e-08, 2.33553e-08, 2.020156e-08, 
    1.958531e-08, 1.913294e-08, 1.947954e-08, 1.89223e-08, 1.90133e-08, 
    1.921191e-08, 2.034802e-08, 2.093477e-08, 2.236643e-08, 2.284397e-08,
  2.739438e-08, 2.591816e-08, 2.556647e-08, 2.355522e-08, 2.004824e-08, 
    1.955148e-08, 1.87384e-08, 1.909087e-08, 1.879189e-08, 1.903301e-08, 
    1.890199e-08, 1.882959e-08, 1.99434e-08, 2.091909e-08, 2.09174e-08,
  2.717551e-08, 2.627018e-08, 2.666197e-08, 2.477804e-08, 2.091123e-08, 
    1.954239e-08, 1.838162e-08, 1.838897e-08, 1.871903e-08, 1.799781e-08, 
    1.751267e-08, 1.762981e-08, 1.929066e-08, 1.984629e-08, 2.137634e-08,
  2.017273e-08, 2.057894e-08, 2.082313e-08, 2.099038e-08, 2.224695e-08, 
    2.379834e-08, 2.469054e-08, 2.525018e-08, 2.486219e-08, 2.376855e-08, 
    2.178358e-08, 2.105591e-08, 2.083817e-08, 2.016547e-08, 2.01188e-08,
  2.062158e-08, 2.130094e-08, 2.116898e-08, 2.157901e-08, 2.326633e-08, 
    2.464501e-08, 2.506436e-08, 2.558272e-08, 2.52549e-08, 2.364149e-08, 
    2.154896e-08, 2.09059e-08, 2.0461e-08, 1.979015e-08, 2.02453e-08,
  2.085645e-08, 2.119032e-08, 2.155713e-08, 2.261839e-08, 2.410376e-08, 
    2.5099e-08, 2.507431e-08, 2.510884e-08, 2.423237e-08, 2.239741e-08, 
    2.164917e-08, 2.085975e-08, 2.032414e-08, 1.988138e-08, 2.059293e-08,
  2.084799e-08, 2.119254e-08, 2.171237e-08, 2.303132e-08, 2.410068e-08, 
    2.471436e-08, 2.504025e-08, 2.470027e-08, 2.325469e-08, 2.21043e-08, 
    2.120077e-08, 1.989197e-08, 1.991857e-08, 2.012565e-08, 1.979836e-08,
  2.117589e-08, 2.178438e-08, 2.241578e-08, 2.28496e-08, 2.433314e-08, 
    2.449705e-08, 2.420502e-08, 2.319965e-08, 2.19839e-08, 2.091768e-08, 
    1.985325e-08, 1.956836e-08, 1.974951e-08, 1.916958e-08, 1.899891e-08,
  2.222539e-08, 2.226989e-08, 2.235953e-08, 2.317952e-08, 2.47748e-08, 
    2.432826e-08, 2.377219e-08, 2.251084e-08, 2.164199e-08, 2.051878e-08, 
    2.061311e-08, 1.987543e-08, 1.877018e-08, 1.84681e-08, 1.936089e-08,
  2.168228e-08, 2.174181e-08, 2.247049e-08, 2.415912e-08, 2.498904e-08, 
    2.46691e-08, 2.337396e-08, 2.249596e-08, 2.212493e-08, 2.127203e-08, 
    2.040053e-08, 1.954828e-08, 1.82431e-08, 1.82629e-08, 1.989845e-08,
  2.183259e-08, 2.231163e-08, 2.288396e-08, 2.466818e-08, 2.482203e-08, 
    2.472322e-08, 2.328695e-08, 2.311781e-08, 2.186963e-08, 2.084036e-08, 
    2.052165e-08, 1.974409e-08, 1.829162e-08, 1.864369e-08, 1.78068e-08,
  2.103883e-08, 2.195713e-08, 2.315181e-08, 2.457163e-08, 2.439434e-08, 
    2.461952e-08, 2.322465e-08, 2.223696e-08, 2.030239e-08, 2.110483e-08, 
    2.042611e-08, 1.91698e-08, 1.761491e-08, 1.647686e-08, 1.592862e-08,
  2.111407e-08, 2.257473e-08, 2.362056e-08, 2.424426e-08, 2.402591e-08, 
    2.385735e-08, 2.293823e-08, 2.149736e-08, 2.114461e-08, 2.059216e-08, 
    2.00461e-08, 1.91064e-08, 1.808135e-08, 1.693195e-08, 1.616801e-08,
  2.087736e-08, 2.182813e-08, 2.168774e-08, 2.226204e-08, 2.25583e-08, 
    2.274901e-08, 2.301683e-08, 2.310041e-08, 2.280282e-08, 2.273628e-08, 
    2.336874e-08, 2.358267e-08, 2.38715e-08, 2.348292e-08, 2.299645e-08,
  2.121892e-08, 2.216128e-08, 2.228312e-08, 2.26653e-08, 2.273638e-08, 
    2.336626e-08, 2.341598e-08, 2.322506e-08, 2.303798e-08, 2.282381e-08, 
    2.331941e-08, 2.354124e-08, 2.337111e-08, 2.303696e-08, 2.26224e-08,
  2.069347e-08, 2.291999e-08, 2.360317e-08, 2.352717e-08, 2.319209e-08, 
    2.415634e-08, 2.368107e-08, 2.29619e-08, 2.310782e-08, 2.296322e-08, 
    2.31898e-08, 2.319877e-08, 2.258125e-08, 2.233188e-08, 2.217116e-08,
  2.119432e-08, 2.320146e-08, 2.309339e-08, 2.30805e-08, 2.327382e-08, 
    2.342675e-08, 2.320426e-08, 2.316778e-08, 2.253924e-08, 2.340796e-08, 
    2.269142e-08, 2.104568e-08, 2.165387e-08, 2.223311e-08, 2.291996e-08,
  2.224986e-08, 2.414668e-08, 2.459869e-08, 2.413596e-08, 2.465061e-08, 
    2.413929e-08, 2.397343e-08, 2.315504e-08, 2.304788e-08, 2.333591e-08, 
    2.240398e-08, 2.257906e-08, 2.234118e-08, 2.311489e-08, 2.435993e-08,
  2.382305e-08, 2.437444e-08, 2.391127e-08, 2.417186e-08, 2.346758e-08, 
    2.29436e-08, 2.220475e-08, 2.208153e-08, 2.196466e-08, 2.201133e-08, 
    2.345074e-08, 2.365905e-08, 2.217538e-08, 2.205973e-08, 2.410197e-08,
  2.368578e-08, 2.349801e-08, 2.34556e-08, 2.289864e-08, 2.231142e-08, 
    2.216773e-08, 2.184885e-08, 2.214543e-08, 2.267742e-08, 2.30372e-08, 
    2.332182e-08, 2.291986e-08, 2.171864e-08, 2.177117e-08, 2.285981e-08,
  2.382061e-08, 2.324128e-08, 2.278684e-08, 2.239202e-08, 2.206961e-08, 
    2.189737e-08, 2.207629e-08, 2.308535e-08, 2.296542e-08, 2.327104e-08, 
    2.306997e-08, 2.318813e-08, 2.212233e-08, 2.171942e-08, 2.169163e-08,
  2.25256e-08, 2.208592e-08, 2.264691e-08, 2.267954e-08, 2.193819e-08, 
    2.183444e-08, 2.259449e-08, 2.29624e-08, 2.318471e-08, 2.381348e-08, 
    2.366785e-08, 2.249362e-08, 2.124472e-08, 2.017026e-08, 1.968653e-08,
  2.208187e-08, 2.240717e-08, 2.310301e-08, 2.217538e-08, 2.20185e-08, 
    2.205213e-08, 2.248313e-08, 2.274801e-08, 2.436814e-08, 2.377398e-08, 
    2.224099e-08, 2.11186e-08, 2.091176e-08, 2.014298e-08, 1.991438e-08,
  2.157231e-08, 2.121997e-08, 2.126897e-08, 2.121493e-08, 2.15879e-08, 
    2.141188e-08, 2.1309e-08, 2.134273e-08, 2.120083e-08, 2.16663e-08, 
    2.339806e-08, 2.366781e-08, 2.351657e-08, 2.352711e-08, 2.376608e-08,
  2.14302e-08, 2.12722e-08, 2.112506e-08, 2.130116e-08, 2.133559e-08, 
    2.06292e-08, 2.096953e-08, 2.072904e-08, 2.07946e-08, 2.168625e-08, 
    2.282788e-08, 2.320592e-08, 2.328147e-08, 2.430773e-08, 2.41568e-08,
  2.056084e-08, 2.132038e-08, 2.177203e-08, 2.1517e-08, 2.072202e-08, 
    2.104073e-08, 2.109102e-08, 2.06724e-08, 2.103761e-08, 2.19957e-08, 
    2.285824e-08, 2.268786e-08, 2.314066e-08, 2.420031e-08, 2.345267e-08,
  2.080065e-08, 2.137377e-08, 2.104231e-08, 2.064922e-08, 2.072778e-08, 
    2.08567e-08, 2.071273e-08, 2.103341e-08, 2.157045e-08, 2.34475e-08, 
    2.464508e-08, 2.389662e-08, 2.380455e-08, 2.37029e-08, 2.112765e-08,
  2.057374e-08, 2.126444e-08, 2.151618e-08, 2.11954e-08, 2.125165e-08, 
    2.119074e-08, 2.178488e-08, 2.234787e-08, 2.383746e-08, 2.572936e-08, 
    2.543515e-08, 2.512046e-08, 2.483516e-08, 2.188828e-08, 2.169988e-08,
  2.110035e-08, 2.117125e-08, 2.101179e-08, 2.099662e-08, 2.062323e-08, 
    2.111217e-08, 2.154492e-08, 2.24501e-08, 2.371418e-08, 2.43404e-08, 
    2.263789e-08, 2.188936e-08, 2.178464e-08, 1.973998e-08, 2.238164e-08,
  2.095284e-08, 2.074175e-08, 2.09851e-08, 2.077167e-08, 2.089718e-08, 
    2.137687e-08, 2.178267e-08, 2.284726e-08, 2.37827e-08, 2.238101e-08, 
    2.13704e-08, 2.130171e-08, 1.997682e-08, 1.92191e-08, 2.419751e-08,
  2.089139e-08, 2.048502e-08, 2.063111e-08, 2.086333e-08, 2.094372e-08, 
    2.109741e-08, 2.153606e-08, 2.25348e-08, 2.188635e-08, 2.157594e-08, 
    2.116885e-08, 2.133066e-08, 2.067957e-08, 2.169883e-08, 2.422339e-08,
  1.970749e-08, 1.971958e-08, 2.075269e-08, 2.115291e-08, 2.086784e-08, 
    2.096548e-08, 2.197286e-08, 2.221315e-08, 2.23874e-08, 2.233678e-08, 
    2.253099e-08, 2.246118e-08, 2.191279e-08, 2.292726e-08, 2.287173e-08,
  1.971916e-08, 2.00351e-08, 2.105453e-08, 2.095614e-08, 2.120526e-08, 
    2.150019e-08, 2.241291e-08, 2.271938e-08, 2.287943e-08, 2.237191e-08, 
    2.286294e-08, 2.226915e-08, 2.257398e-08, 2.269494e-08, 2.24887e-08,
  2.392762e-08, 2.409637e-08, 2.374726e-08, 2.328595e-08, 2.32832e-08, 
    2.340265e-08, 2.430864e-08, 2.443351e-08, 2.431068e-08, 2.331282e-08, 
    2.415327e-08, 2.382092e-08, 2.285593e-08, 2.152893e-08, 2.132996e-08,
  2.385416e-08, 2.345746e-08, 2.330997e-08, 2.296903e-08, 2.288301e-08, 
    2.346159e-08, 2.369937e-08, 2.374977e-08, 2.325376e-08, 2.295117e-08, 
    2.288486e-08, 2.246016e-08, 2.163033e-08, 2.208549e-08, 2.312581e-08,
  2.170473e-08, 2.294323e-08, 2.296415e-08, 2.329496e-08, 2.29952e-08, 
    2.405077e-08, 2.396122e-08, 2.361679e-08, 2.337264e-08, 2.284367e-08, 
    2.271339e-08, 2.217736e-08, 2.178912e-08, 2.337522e-08, 2.285216e-08,
  2.231207e-08, 2.338289e-08, 2.304195e-08, 2.304441e-08, 2.341895e-08, 
    2.407171e-08, 2.37698e-08, 2.387461e-08, 2.319009e-08, 2.378845e-08, 
    2.395333e-08, 2.37745e-08, 2.325319e-08, 2.364175e-08, 2.038627e-08,
  2.278541e-08, 2.407181e-08, 2.460484e-08, 2.466559e-08, 2.543293e-08, 
    2.522889e-08, 2.539544e-08, 2.491492e-08, 2.479154e-08, 2.549612e-08, 
    2.453459e-08, 2.406459e-08, 2.279136e-08, 2.079878e-08, 1.882437e-08,
  2.38527e-08, 2.469952e-08, 2.427323e-08, 2.517113e-08, 2.482096e-08, 
    2.466429e-08, 2.411571e-08, 2.364803e-08, 2.322686e-08, 2.344767e-08, 
    2.215116e-08, 2.128384e-08, 2.110844e-08, 1.88153e-08, 2.006612e-08,
  2.401691e-08, 2.419242e-08, 2.45056e-08, 2.462882e-08, 2.434475e-08, 
    2.393709e-08, 2.351273e-08, 2.287145e-08, 2.29019e-08, 2.170496e-08, 
    2.080335e-08, 2.084107e-08, 1.965882e-08, 1.848459e-08, 2.34452e-08,
  2.460883e-08, 2.465704e-08, 2.452876e-08, 2.466944e-08, 2.397989e-08, 
    2.346954e-08, 2.256129e-08, 2.215331e-08, 2.130887e-08, 2.060422e-08, 
    2.029615e-08, 2.062835e-08, 1.969564e-08, 2.043304e-08, 2.365876e-08,
  2.344917e-08, 2.351709e-08, 2.359018e-08, 2.372403e-08, 2.231923e-08, 
    2.194952e-08, 2.119759e-08, 2.092616e-08, 2.058823e-08, 1.999043e-08, 
    2.031605e-08, 2.071826e-08, 2.055933e-08, 2.173657e-08, 2.324376e-08,
  2.346858e-08, 2.354816e-08, 2.361275e-08, 2.295839e-08, 2.176623e-08, 
    2.13309e-08, 2.072258e-08, 2.034568e-08, 2.005904e-08, 1.993153e-08, 
    2.061786e-08, 2.07562e-08, 2.114372e-08, 2.213577e-08, 2.243092e-08,
  2.311469e-08, 2.399247e-08, 2.433012e-08, 2.43552e-08, 2.398392e-08, 
    2.367519e-08, 2.257826e-08, 2.183833e-08, 2.088235e-08, 2.023531e-08, 
    2.250326e-08, 2.291144e-08, 2.394392e-08, 2.421701e-08, 2.464548e-08,
  2.434765e-08, 2.456543e-08, 2.460649e-08, 2.368014e-08, 2.29517e-08, 
    2.174403e-08, 2.074034e-08, 2.035075e-08, 1.992895e-08, 2.103068e-08, 
    2.211758e-08, 2.261162e-08, 2.40945e-08, 2.503946e-08, 2.610521e-08,
  2.376947e-08, 2.407067e-08, 2.327753e-08, 2.248824e-08, 2.087851e-08, 
    2.069666e-08, 2.018899e-08, 2.026238e-08, 2.065193e-08, 2.140297e-08, 
    2.262123e-08, 2.353569e-08, 2.556526e-08, 2.607015e-08, 2.603936e-08,
  2.284108e-08, 2.289302e-08, 2.167955e-08, 2.040138e-08, 1.999016e-08, 
    2.002906e-08, 1.98061e-08, 2.04658e-08, 2.08462e-08, 2.300787e-08, 
    2.499586e-08, 2.719099e-08, 2.711195e-08, 2.646764e-08, 2.334601e-08,
  2.136584e-08, 2.102226e-08, 2.047279e-08, 1.999757e-08, 2.019365e-08, 
    2.009976e-08, 2.090622e-08, 2.184331e-08, 2.339146e-08, 2.489279e-08, 
    2.530509e-08, 2.52816e-08, 2.447274e-08, 2.262833e-08, 2.024427e-08,
  2.044097e-08, 2.031892e-08, 1.979824e-08, 1.998397e-08, 1.966302e-08, 
    2.015269e-08, 2.086881e-08, 2.219275e-08, 2.314329e-08, 2.423162e-08, 
    2.346215e-08, 2.237056e-08, 2.192103e-08, 1.97716e-08, 2.049715e-08,
  1.977832e-08, 1.957913e-08, 1.947831e-08, 1.965805e-08, 1.975881e-08, 
    2.067615e-08, 2.164904e-08, 2.314307e-08, 2.345698e-08, 2.291459e-08, 
    2.206593e-08, 2.165245e-08, 2.061251e-08, 1.88854e-08, 2.066614e-08,
  1.922582e-08, 1.934978e-08, 1.924084e-08, 1.986867e-08, 2.01521e-08, 
    2.135207e-08, 2.210584e-08, 2.206822e-08, 2.194523e-08, 2.16002e-08, 
    2.079444e-08, 2.032541e-08, 1.933115e-08, 1.89059e-08, 2.02048e-08,
  1.849852e-08, 1.934921e-08, 1.978365e-08, 2.093389e-08, 2.085961e-08, 
    2.14846e-08, 2.153762e-08, 2.151571e-08, 2.166966e-08, 2.070366e-08, 
    2.014407e-08, 1.955027e-08, 1.88776e-08, 1.914167e-08, 1.955282e-08,
  1.898969e-08, 2.018355e-08, 2.077083e-08, 2.097049e-08, 2.125824e-08, 
    2.177555e-08, 2.129976e-08, 2.130628e-08, 2.024651e-08, 1.97115e-08, 
    1.939005e-08, 1.904857e-08, 1.895519e-08, 1.953426e-08, 1.978398e-08,
  2.163583e-08, 2.224779e-08, 2.164077e-08, 2.184012e-08, 2.176471e-08, 
    2.231631e-08, 2.214326e-08, 2.165626e-08, 1.996892e-08, 1.91766e-08, 
    2.025608e-08, 2.043119e-08, 2.027124e-08, 2.054525e-08, 2.109034e-08,
  2.280964e-08, 2.173576e-08, 2.151562e-08, 2.157731e-08, 2.098988e-08, 
    2.099746e-08, 2.022332e-08, 2.026682e-08, 1.920673e-08, 1.979616e-08, 
    2.020785e-08, 2.026426e-08, 2.039319e-08, 2.148365e-08, 2.275499e-08,
  2.035296e-08, 2.071938e-08, 2.055999e-08, 2.033909e-08, 1.98531e-08, 
    2.036775e-08, 2.048293e-08, 2.038479e-08, 1.988653e-08, 2.023576e-08, 
    2.048754e-08, 2.050497e-08, 2.146433e-08, 2.261403e-08, 2.26374e-08,
  1.978288e-08, 2.073936e-08, 2.026372e-08, 1.991204e-08, 2.058283e-08, 
    2.080999e-08, 2.06786e-08, 2.059688e-08, 2.05838e-08, 2.125775e-08, 
    2.297577e-08, 2.424667e-08, 2.361456e-08, 2.305053e-08, 2.139932e-08,
  1.979426e-08, 2.076901e-08, 2.078922e-08, 2.14267e-08, 2.191999e-08, 
    2.215025e-08, 2.208565e-08, 2.201775e-08, 2.260862e-08, 2.442892e-08, 
    2.460747e-08, 2.378563e-08, 2.217217e-08, 2.151945e-08, 2.180256e-08,
  2.031645e-08, 2.056689e-08, 2.134788e-08, 2.232401e-08, 2.198895e-08, 
    2.251923e-08, 2.201438e-08, 2.258483e-08, 2.354336e-08, 2.426715e-08, 
    2.257176e-08, 2.196878e-08, 2.25221e-08, 2.14097e-08, 2.222879e-08,
  2.03648e-08, 2.145206e-08, 2.218531e-08, 2.229049e-08, 2.265593e-08, 
    2.272478e-08, 2.261961e-08, 2.360226e-08, 2.353794e-08, 2.274617e-08, 
    2.235161e-08, 2.300027e-08, 2.238911e-08, 2.161312e-08, 2.356161e-08,
  2.21097e-08, 2.290549e-08, 2.256244e-08, 2.341041e-08, 2.288029e-08, 
    2.240809e-08, 2.238496e-08, 2.28934e-08, 2.324376e-08, 2.348079e-08, 
    2.368402e-08, 2.378217e-08, 2.340033e-08, 2.301658e-08, 2.408118e-08,
  2.266913e-08, 2.287995e-08, 2.346474e-08, 2.400482e-08, 2.276191e-08, 
    2.291355e-08, 2.341636e-08, 2.51674e-08, 2.489631e-08, 2.411872e-08, 
    2.407993e-08, 2.422964e-08, 2.403128e-08, 2.419985e-08, 2.480469e-08,
  2.299749e-08, 2.365996e-08, 2.469357e-08, 2.445818e-08, 2.456778e-08, 
    2.505579e-08, 2.531421e-08, 2.528872e-08, 2.417444e-08, 2.4403e-08, 
    2.475163e-08, 2.487183e-08, 2.484531e-08, 2.524144e-08, 2.529859e-08,
  2.381811e-08, 2.118296e-08, 2.041624e-08, 2.109703e-08, 2.238118e-08, 
    2.425216e-08, 2.504003e-08, 2.520962e-08, 2.473095e-08, 2.450318e-08, 
    2.585921e-08, 2.551742e-08, 2.425405e-08, 2.409389e-08, 2.441784e-08,
  2.134543e-08, 2.022868e-08, 2.061966e-08, 2.176123e-08, 2.31821e-08, 
    2.427453e-08, 2.491784e-08, 2.505808e-08, 2.497411e-08, 2.511819e-08, 
    2.50467e-08, 2.436859e-08, 2.432479e-08, 2.519951e-08, 2.591785e-08,
  1.967512e-08, 2.023028e-08, 2.266938e-08, 2.350315e-08, 2.352798e-08, 
    2.514123e-08, 2.55484e-08, 2.535628e-08, 2.526703e-08, 2.491403e-08, 
    2.456491e-08, 2.417364e-08, 2.575472e-08, 2.655113e-08, 2.614863e-08,
  1.996616e-08, 2.205713e-08, 2.265167e-08, 2.34895e-08, 2.485083e-08, 
    2.512678e-08, 2.517185e-08, 2.583343e-08, 2.54676e-08, 2.547389e-08, 
    2.546721e-08, 2.652032e-08, 2.727067e-08, 2.624201e-08, 2.418923e-08,
  2.201201e-08, 2.479928e-08, 2.661383e-08, 2.714616e-08, 2.67863e-08, 
    2.676307e-08, 2.690255e-08, 2.682078e-08, 2.694998e-08, 2.74137e-08, 
    2.676575e-08, 2.542577e-08, 2.381232e-08, 2.291997e-08, 2.380594e-08,
  2.411703e-08, 2.529415e-08, 2.645018e-08, 2.637849e-08, 2.577981e-08, 
    2.600044e-08, 2.596695e-08, 2.648818e-08, 2.739343e-08, 2.645871e-08, 
    2.498664e-08, 2.394094e-08, 2.332249e-08, 2.196854e-08, 2.481994e-08,
  2.562076e-08, 2.680672e-08, 2.656842e-08, 2.63023e-08, 2.616865e-08, 
    2.589117e-08, 2.591569e-08, 2.637368e-08, 2.641862e-08, 2.510884e-08, 
    2.4424e-08, 2.368587e-08, 2.236786e-08, 2.14662e-08, 2.559726e-08,
  2.691689e-08, 2.670418e-08, 2.66861e-08, 2.618756e-08, 2.546392e-08, 
    2.503746e-08, 2.506201e-08, 2.51117e-08, 2.554401e-08, 2.478015e-08, 
    2.409296e-08, 2.272483e-08, 2.233489e-08, 2.14532e-08, 2.299673e-08,
  2.721801e-08, 2.7438e-08, 2.736806e-08, 2.632594e-08, 2.599026e-08, 
    2.57742e-08, 2.552468e-08, 2.569774e-08, 2.499955e-08, 2.417937e-08, 
    2.329656e-08, 2.224317e-08, 2.225615e-08, 2.170963e-08, 2.25149e-08,
  2.856016e-08, 2.846184e-08, 2.831602e-08, 2.703631e-08, 2.69048e-08, 
    2.591682e-08, 2.485271e-08, 2.489085e-08, 2.401423e-08, 2.374482e-08, 
    2.289355e-08, 2.215991e-08, 2.245163e-08, 2.255107e-08, 2.337416e-08,
  2.072953e-08, 2.146448e-08, 2.308408e-08, 2.561855e-08, 3.027473e-08, 
    3.134188e-08, 2.97187e-08, 2.765667e-08, 2.520088e-08, 2.319809e-08, 
    2.270623e-08, 2.312374e-08, 2.350303e-08, 2.438483e-08, 2.497821e-08,
  2.192067e-08, 2.335993e-08, 2.610425e-08, 2.934329e-08, 3.258727e-08, 
    3.007035e-08, 2.747626e-08, 2.58989e-08, 2.385954e-08, 2.248203e-08, 
    2.342076e-08, 2.410012e-08, 2.4574e-08, 2.554175e-08, 2.524224e-08,
  2.350597e-08, 2.604957e-08, 2.987005e-08, 3.118495e-08, 3.056547e-08, 
    2.787563e-08, 2.480004e-08, 2.309783e-08, 2.250504e-08, 2.339235e-08, 
    2.40915e-08, 2.392852e-08, 2.47178e-08, 2.530501e-08, 2.471037e-08,
  2.409555e-08, 2.912174e-08, 3.134844e-08, 3.172971e-08, 2.962369e-08, 
    2.438012e-08, 2.245302e-08, 2.281195e-08, 2.416521e-08, 2.507428e-08, 
    2.524277e-08, 2.626129e-08, 2.584577e-08, 2.524411e-08, 2.338501e-08,
  2.707582e-08, 3.189831e-08, 3.196214e-08, 2.892164e-08, 2.48389e-08, 
    2.245385e-08, 2.27371e-08, 2.411451e-08, 2.492321e-08, 2.583338e-08, 
    2.560037e-08, 2.486908e-08, 2.38526e-08, 2.282533e-08, 2.330551e-08,
  3.047636e-08, 3.113612e-08, 2.922249e-08, 2.683087e-08, 2.439574e-08, 
    2.245218e-08, 2.345642e-08, 2.432807e-08, 2.419882e-08, 2.437027e-08, 
    2.336906e-08, 2.318788e-08, 2.375159e-08, 2.299314e-08, 2.468398e-08,
  3.221562e-08, 3.073111e-08, 2.828176e-08, 2.532783e-08, 2.23162e-08, 
    2.264818e-08, 2.370412e-08, 2.382169e-08, 2.33856e-08, 2.320809e-08, 
    2.347774e-08, 2.39187e-08, 2.377188e-08, 2.315993e-08, 2.428891e-08,
  3.315764e-08, 2.932518e-08, 2.700421e-08, 2.355975e-08, 2.196132e-08, 
    2.348748e-08, 2.446445e-08, 2.392299e-08, 2.341952e-08, 2.380952e-08, 
    2.434493e-08, 2.425042e-08, 2.39389e-08, 2.384621e-08, 2.43216e-08,
  3.249504e-08, 2.92873e-08, 2.693343e-08, 2.397915e-08, 2.290234e-08, 
    2.444148e-08, 2.544066e-08, 2.519502e-08, 2.431194e-08, 2.472801e-08, 
    2.465225e-08, 2.432989e-08, 2.37617e-08, 2.352498e-08, 2.344213e-08,
  3.201278e-08, 2.912725e-08, 2.676448e-08, 2.362018e-08, 2.370639e-08, 
    2.627042e-08, 2.629211e-08, 2.532077e-08, 2.497398e-08, 2.508882e-08, 
    2.462459e-08, 2.416698e-08, 2.374996e-08, 2.348606e-08, 2.342865e-08,
  2.36346e-08, 2.402996e-08, 2.58246e-08, 2.638746e-08, 2.662282e-08, 
    2.551559e-08, 2.523896e-08, 2.539722e-08, 2.5165e-08, 2.41791e-08, 
    2.478976e-08, 2.421751e-08, 2.412548e-08, 2.428916e-08, 2.480597e-08,
  2.112566e-08, 2.193943e-08, 2.552639e-08, 2.600805e-08, 2.532261e-08, 
    2.486759e-08, 2.505445e-08, 2.488882e-08, 2.480834e-08, 2.486163e-08, 
    2.51949e-08, 2.457224e-08, 2.444592e-08, 2.502037e-08, 2.554472e-08,
  2.065262e-08, 2.259414e-08, 2.481525e-08, 2.538937e-08, 2.557439e-08, 
    2.508277e-08, 2.475176e-08, 2.487118e-08, 2.531993e-08, 2.519575e-08, 
    2.51948e-08, 2.444379e-08, 2.466904e-08, 2.530387e-08, 2.549437e-08,
  2.288182e-08, 2.416928e-08, 2.452249e-08, 2.570921e-08, 2.753756e-08, 
    2.615877e-08, 2.478366e-08, 2.499425e-08, 2.621343e-08, 2.75717e-08, 
    2.844602e-08, 2.783787e-08, 2.63069e-08, 2.548311e-08, 2.466221e-08,
  2.316631e-08, 2.518963e-08, 2.699782e-08, 2.734673e-08, 2.597269e-08, 
    2.590078e-08, 2.619809e-08, 2.704575e-08, 2.930379e-08, 2.886848e-08, 
    2.768559e-08, 2.798472e-08, 2.619025e-08, 2.378924e-08, 2.389971e-08,
  2.281429e-08, 2.419536e-08, 2.512468e-08, 2.617474e-08, 2.680495e-08, 
    2.628805e-08, 2.603957e-08, 2.70518e-08, 2.729001e-08, 2.723064e-08, 
    2.535791e-08, 2.546903e-08, 2.537504e-08, 2.372007e-08, 2.442454e-08,
  2.281017e-08, 2.398611e-08, 2.47904e-08, 2.599097e-08, 2.602497e-08, 
    2.571469e-08, 2.559396e-08, 2.573395e-08, 2.605496e-08, 2.509012e-08, 
    2.557297e-08, 2.572308e-08, 2.440066e-08, 2.56014e-08, 2.535984e-08,
  2.199606e-08, 2.309936e-08, 2.417541e-08, 2.535603e-08, 2.597834e-08, 
    2.538073e-08, 2.46101e-08, 2.47174e-08, 2.478278e-08, 2.503496e-08, 
    2.559435e-08, 2.572862e-08, 2.628523e-08, 2.832477e-08, 2.60104e-08,
  2.109152e-08, 2.247715e-08, 2.391558e-08, 2.545868e-08, 2.678488e-08, 
    2.699125e-08, 2.64038e-08, 2.543082e-08, 2.530911e-08, 2.473218e-08, 
    2.513731e-08, 2.53471e-08, 2.606725e-08, 2.595107e-08, 2.55315e-08,
  2.027212e-08, 2.169541e-08, 2.324962e-08, 2.445447e-08, 2.631193e-08, 
    2.720805e-08, 2.617941e-08, 2.563137e-08, 2.428059e-08, 2.492456e-08, 
    2.503291e-08, 2.471273e-08, 2.495388e-08, 2.571862e-08, 2.532874e-08,
  2.062967e-08, 2.012607e-08, 2.003219e-08, 2.048031e-08, 2.10604e-08, 
    2.108025e-08, 2.176825e-08, 2.235641e-08, 2.258961e-08, 2.399838e-08, 
    2.600907e-08, 2.416465e-08, 2.330822e-08, 2.197276e-08, 2.103084e-08,
  2.015895e-08, 1.954925e-08, 2.015827e-08, 2.05813e-08, 2.055482e-08, 
    2.105517e-08, 2.20219e-08, 2.248288e-08, 2.298158e-08, 2.330177e-08, 
    2.434246e-08, 2.376873e-08, 2.404108e-08, 2.24588e-08, 2.170506e-08,
  1.873482e-08, 2.024481e-08, 2.06792e-08, 2.030325e-08, 2.112926e-08, 
    2.244771e-08, 2.261691e-08, 2.265595e-08, 2.338345e-08, 2.301635e-08, 
    2.438079e-08, 2.332952e-08, 2.338177e-08, 2.142387e-08, 2.090184e-08,
  2.020949e-08, 2.177976e-08, 2.129911e-08, 2.153115e-08, 2.242501e-08, 
    2.267537e-08, 2.300785e-08, 2.340164e-08, 2.376219e-08, 2.486931e-08, 
    2.78788e-08, 2.669276e-08, 2.473126e-08, 2.145147e-08, 1.985769e-08,
  2.149985e-08, 2.287581e-08, 2.287121e-08, 2.246683e-08, 2.250848e-08, 
    2.377149e-08, 2.477256e-08, 2.453415e-08, 2.507315e-08, 2.513866e-08, 
    2.510843e-08, 2.563902e-08, 2.543217e-08, 2.084101e-08, 2.136808e-08,
  2.249639e-08, 2.269177e-08, 2.212415e-08, 2.189049e-08, 2.217028e-08, 
    2.392314e-08, 2.440587e-08, 2.457419e-08, 2.465308e-08, 2.452507e-08, 
    2.263781e-08, 2.188778e-08, 2.305707e-08, 2.05401e-08, 2.19361e-08,
  2.325909e-08, 2.294718e-08, 2.285185e-08, 2.258485e-08, 2.307826e-08, 
    2.445491e-08, 2.500426e-08, 2.469292e-08, 2.417104e-08, 2.280776e-08, 
    2.245656e-08, 2.187917e-08, 2.17649e-08, 2.163479e-08, 2.166151e-08,
  2.324039e-08, 2.33585e-08, 2.305282e-08, 2.326418e-08, 2.386354e-08, 
    2.487616e-08, 2.493437e-08, 2.433324e-08, 2.378343e-08, 2.349242e-08, 
    2.294216e-08, 2.213591e-08, 2.200194e-08, 2.179948e-08, 1.999123e-08,
  2.287922e-08, 2.258489e-08, 2.319062e-08, 2.454896e-08, 2.514496e-08, 
    2.543634e-08, 2.5084e-08, 2.528133e-08, 2.465397e-08, 2.42871e-08, 
    2.347091e-08, 2.222303e-08, 2.137681e-08, 1.981136e-08, 1.965116e-08,
  2.164269e-08, 2.198922e-08, 2.318349e-08, 2.452726e-08, 2.566711e-08, 
    2.549005e-08, 2.541469e-08, 2.524111e-08, 2.490102e-08, 2.479595e-08, 
    2.403307e-08, 2.230802e-08, 2.064272e-08, 1.938019e-08, 1.89974e-08,
  2.37636e-08, 2.445838e-08, 2.426716e-08, 2.470945e-08, 2.470236e-08, 
    2.50851e-08, 2.553458e-08, 2.557378e-08, 2.485089e-08, 2.472343e-08, 
    2.582181e-08, 2.607269e-08, 2.574184e-08, 2.589345e-08, 2.462101e-08,
  2.408574e-08, 2.459866e-08, 2.444366e-08, 2.445332e-08, 2.43834e-08, 
    2.47777e-08, 2.459072e-08, 2.448675e-08, 2.400465e-08, 2.490251e-08, 
    2.584205e-08, 2.566575e-08, 2.565055e-08, 2.653968e-08, 2.58185e-08,
  2.32226e-08, 2.456777e-08, 2.459413e-08, 2.460711e-08, 2.426785e-08, 
    2.470146e-08, 2.444276e-08, 2.421376e-08, 2.43621e-08, 2.542295e-08, 
    2.597027e-08, 2.520671e-08, 2.607153e-08, 2.688506e-08, 2.610538e-08,
  2.319386e-08, 2.47442e-08, 2.469522e-08, 2.492172e-08, 2.494536e-08, 
    2.455927e-08, 2.444307e-08, 2.39991e-08, 2.378932e-08, 2.558607e-08, 
    2.516875e-08, 2.577978e-08, 2.738982e-08, 2.779056e-08, 2.647873e-08,
  2.34906e-08, 2.418998e-08, 2.506195e-08, 2.474739e-08, 2.458768e-08, 
    2.444708e-08, 2.433832e-08, 2.392296e-08, 2.468032e-08, 2.666225e-08, 
    2.727362e-08, 2.768773e-08, 2.648328e-08, 2.501945e-08, 2.4209e-08,
  2.396414e-08, 2.375399e-08, 2.467585e-08, 2.447291e-08, 2.420557e-08, 
    2.461734e-08, 2.384763e-08, 2.435861e-08, 2.584791e-08, 2.572818e-08, 
    2.90007e-08, 2.708296e-08, 2.457086e-08, 2.065586e-08, 2.258333e-08,
  2.444264e-08, 2.377605e-08, 2.409061e-08, 2.463598e-08, 2.484347e-08, 
    2.496447e-08, 2.484561e-08, 2.442163e-08, 2.713286e-08, 2.648749e-08, 
    2.494152e-08, 2.340886e-08, 2.117222e-08, 1.860794e-08, 2.297049e-08,
  2.383464e-08, 2.395389e-08, 2.377929e-08, 2.398423e-08, 2.425288e-08, 
    2.470898e-08, 2.399424e-08, 2.469674e-08, 2.249516e-08, 2.120535e-08, 
    2.096091e-08, 2.210548e-08, 2.084797e-08, 2.1514e-08, 2.465567e-08,
  2.442133e-08, 2.367912e-08, 2.330407e-08, 2.299599e-08, 2.342977e-08, 
    2.407348e-08, 2.387057e-08, 2.411717e-08, 1.900089e-08, 2.034408e-08, 
    2.071269e-08, 2.252066e-08, 2.071583e-08, 2.316608e-08, 2.290704e-08,
  2.412095e-08, 2.361121e-08, 2.347478e-08, 2.29179e-08, 2.302941e-08, 
    2.300931e-08, 2.223346e-08, 2.163947e-08, 2.069562e-08, 2.143872e-08, 
    2.246692e-08, 2.263749e-08, 2.227319e-08, 1.987169e-08, 2.070164e-08,
  2.69114e-08, 2.538738e-08, 2.406031e-08, 2.326443e-08, 2.394239e-08, 
    2.388683e-08, 2.397995e-08, 2.395506e-08, 2.305432e-08, 2.311952e-08, 
    2.388216e-08, 2.345126e-08, 2.305632e-08, 2.323054e-08, 2.333667e-08,
  2.711951e-08, 2.467653e-08, 2.318622e-08, 2.33185e-08, 2.409196e-08, 
    2.348788e-08, 2.348641e-08, 2.331423e-08, 2.264396e-08, 2.262485e-08, 
    2.318261e-08, 2.307984e-08, 2.315173e-08, 2.363434e-08, 2.405072e-08,
  2.918757e-08, 2.485591e-08, 2.349583e-08, 2.451933e-08, 2.435792e-08, 
    2.387522e-08, 2.368867e-08, 2.314738e-08, 2.281586e-08, 2.241894e-08, 
    2.312565e-08, 2.28502e-08, 2.322159e-08, 2.361425e-08, 2.424255e-08,
  2.485908e-08, 2.393027e-08, 2.392753e-08, 2.423084e-08, 2.397979e-08, 
    2.343535e-08, 2.350982e-08, 2.318007e-08, 2.282649e-08, 2.275962e-08, 
    2.537953e-08, 2.479076e-08, 2.374453e-08, 2.4364e-08, 2.335297e-08,
  2.492517e-08, 2.490725e-08, 2.540821e-08, 2.454832e-08, 2.421098e-08, 
    2.40661e-08, 2.406927e-08, 2.331852e-08, 2.309367e-08, 2.493169e-08, 
    2.431513e-08, 2.297939e-08, 2.339315e-08, 2.417696e-08, 2.191109e-08,
  2.460203e-08, 2.45932e-08, 2.561401e-08, 2.431279e-08, 2.369763e-08, 
    2.335064e-08, 2.299238e-08, 2.247466e-08, 2.338208e-08, 2.338051e-08, 
    2.209288e-08, 2.204026e-08, 2.418752e-08, 2.255223e-08, 2.21333e-08,
  2.437861e-08, 2.57275e-08, 2.58346e-08, 2.436066e-08, 2.358144e-08, 
    2.32458e-08, 2.292949e-08, 2.231745e-08, 2.350749e-08, 2.265741e-08, 
    2.198948e-08, 2.250683e-08, 2.2667e-08, 2.125052e-08, 2.262332e-08,
  2.444697e-08, 2.705314e-08, 2.459712e-08, 2.310549e-08, 2.352754e-08, 
    2.408202e-08, 2.340628e-08, 2.230109e-08, 2.328537e-08, 2.307774e-08, 
    2.229728e-08, 2.252419e-08, 2.240952e-08, 2.148248e-08, 2.402911e-08,
  2.367711e-08, 2.495628e-08, 2.315546e-08, 2.196428e-08, 2.36275e-08, 
    2.474519e-08, 2.343437e-08, 2.327841e-08, 2.157417e-08, 2.241979e-08, 
    2.249776e-08, 2.242316e-08, 2.223456e-08, 2.292234e-08, 2.448073e-08,
  2.1401e-08, 2.07234e-08, 1.979559e-08, 2.094325e-08, 2.458768e-08, 
    2.409874e-08, 2.344745e-08, 2.295442e-08, 2.12364e-08, 2.207148e-08, 
    2.26028e-08, 2.23559e-08, 2.240835e-08, 2.289581e-08, 2.274704e-08,
  2.37496e-08, 2.595292e-08, 2.723833e-08, 2.848186e-08, 2.872265e-08, 
    2.767103e-08, 2.739537e-08, 2.544733e-08, 2.46194e-08, 2.413801e-08, 
    2.427333e-08, 2.442118e-08, 2.298117e-08, 2.282284e-08, 2.243891e-08,
  2.5891e-08, 2.82126e-08, 2.682483e-08, 2.656603e-08, 2.727491e-08, 
    2.808523e-08, 2.606997e-08, 2.477008e-08, 2.453779e-08, 2.456853e-08, 
    2.435685e-08, 2.377525e-08, 2.260661e-08, 2.35786e-08, 2.242043e-08,
  2.249756e-08, 2.643204e-08, 2.496155e-08, 2.378302e-08, 2.49551e-08, 
    2.792012e-08, 2.561981e-08, 2.492944e-08, 2.472755e-08, 2.497352e-08, 
    2.44594e-08, 2.342767e-08, 2.254115e-08, 2.443784e-08, 2.134522e-08,
  1.701279e-08, 1.987389e-08, 2.002625e-08, 2.299972e-08, 2.429946e-08, 
    2.368719e-08, 2.419299e-08, 2.480955e-08, 2.336911e-08, 2.494214e-08, 
    2.348527e-08, 2.331853e-08, 2.26485e-08, 2.441569e-08, 2.14705e-08,
  1.919523e-08, 2.161291e-08, 2.499339e-08, 2.479355e-08, 2.573961e-08, 
    2.515554e-08, 2.589244e-08, 2.461519e-08, 2.51353e-08, 2.553289e-08, 
    2.633049e-08, 2.516958e-08, 2.270519e-08, 2.342057e-08, 2.135136e-08,
  2.128443e-08, 2.108821e-08, 2.582743e-08, 2.402429e-08, 2.366934e-08, 
    2.258026e-08, 2.223245e-08, 2.277133e-08, 2.552595e-08, 2.521352e-08, 
    2.929015e-08, 2.493535e-08, 2.331262e-08, 1.920207e-08, 2.008778e-08,
  1.73186e-08, 2.055839e-08, 2.25229e-08, 2.171006e-08, 2.07926e-08, 
    1.9033e-08, 2.036455e-08, 2.13061e-08, 2.501218e-08, 2.671991e-08, 
    2.613432e-08, 2.363537e-08, 1.964823e-08, 1.731855e-08, 2.332375e-08,
  1.668867e-08, 2.013872e-08, 2.010264e-08, 1.957954e-08, 1.79733e-08, 
    1.758851e-08, 1.910569e-08, 2.033764e-08, 2.194457e-08, 2.117203e-08, 
    2.21189e-08, 2.208853e-08, 1.903286e-08, 2.052849e-08, 2.390389e-08,
  1.653921e-08, 1.770527e-08, 1.837723e-08, 1.698571e-08, 1.653852e-08, 
    1.813913e-08, 1.960784e-08, 1.974252e-08, 1.452962e-08, 1.699503e-08, 
    2.02485e-08, 2.130551e-08, 2.046047e-08, 2.130371e-08, 2.247142e-08,
  1.701323e-08, 1.721942e-08, 1.79107e-08, 1.641494e-08, 1.665935e-08, 
    1.725983e-08, 1.917013e-08, 1.820694e-08, 1.432266e-08, 1.646903e-08, 
    1.966669e-08, 2.047484e-08, 2.020364e-08, 2.038865e-08, 2.106961e-08,
  1.92598e-08, 1.956774e-08, 1.93137e-08, 1.929999e-08, 1.858927e-08, 
    1.853031e-08, 1.866196e-08, 1.896011e-08, 1.903816e-08, 2.065325e-08, 
    2.145734e-08, 2.065449e-08, 1.960251e-08, 2.195809e-08, 2.219293e-08,
  1.967728e-08, 1.975066e-08, 1.941626e-08, 1.904988e-08, 1.772075e-08, 
    1.833045e-08, 1.792263e-08, 1.79619e-08, 1.817673e-08, 1.972335e-08, 
    1.977269e-08, 1.89095e-08, 1.958838e-08, 2.300369e-08, 2.255915e-08,
  2.070921e-08, 1.973222e-08, 1.944209e-08, 1.856077e-08, 1.813391e-08, 
    1.849806e-08, 1.737627e-08, 1.718491e-08, 1.749e-08, 1.945256e-08, 
    1.910562e-08, 1.772356e-08, 1.924096e-08, 2.276847e-08, 2.176292e-08,
  2.112936e-08, 2.019434e-08, 1.933103e-08, 1.885423e-08, 1.89443e-08, 
    1.813273e-08, 1.761533e-08, 1.7507e-08, 1.803796e-08, 2.076491e-08, 
    2.153123e-08, 1.982174e-08, 2.173004e-08, 2.116881e-08, 2.127867e-08,
  2.138971e-08, 2.010229e-08, 1.944685e-08, 1.9432e-08, 1.937226e-08, 
    1.842884e-08, 1.896285e-08, 1.832008e-08, 2.050225e-08, 2.326397e-08, 
    2.318998e-08, 2.331459e-08, 2.114856e-08, 1.933001e-08, 2.018273e-08,
  2.056405e-08, 1.93806e-08, 1.85232e-08, 1.9068e-08, 1.91355e-08, 
    1.883194e-08, 1.916125e-08, 1.922408e-08, 2.143381e-08, 2.217591e-08, 
    2.156383e-08, 2.18457e-08, 2.095801e-08, 1.720233e-08, 1.977942e-08,
  1.980835e-08, 1.916812e-08, 1.864128e-08, 1.904808e-08, 1.907704e-08, 
    1.935026e-08, 1.99169e-08, 2.028481e-08, 2.046286e-08, 2.04242e-08, 
    2.042619e-08, 1.932831e-08, 1.592714e-08, 1.45598e-08, 1.94568e-08,
  1.925067e-08, 1.887384e-08, 1.852514e-08, 1.871185e-08, 1.867378e-08, 
    1.981797e-08, 2.009813e-08, 1.984417e-08, 1.904463e-08, 1.905947e-08, 
    1.831254e-08, 1.797231e-08, 1.580497e-08, 1.69615e-08, 1.951284e-08,
  1.949553e-08, 1.906348e-08, 1.88996e-08, 1.846502e-08, 1.868703e-08, 
    1.964243e-08, 2.027689e-08, 1.977361e-08, 2.017062e-08, 1.945792e-08, 
    1.852774e-08, 1.848657e-08, 1.698092e-08, 1.759711e-08, 1.8697e-08,
  1.939849e-08, 1.87234e-08, 1.821895e-08, 1.795356e-08, 1.860884e-08, 
    1.941248e-08, 1.995507e-08, 2.043356e-08, 2.086792e-08, 2.043262e-08, 
    1.985976e-08, 1.955103e-08, 1.854391e-08, 1.788953e-08, 1.793785e-08,
  1.500515e-08, 1.558278e-08, 1.745266e-08, 1.834069e-08, 1.908401e-08, 
    1.966771e-08, 2.011689e-08, 1.988799e-08, 1.938821e-08, 1.940795e-08, 
    1.982559e-08, 1.906105e-08, 1.827286e-08, 1.816903e-08, 1.866514e-08,
  1.530813e-08, 1.598609e-08, 1.796214e-08, 1.889001e-08, 1.960802e-08, 
    2.023986e-08, 2.010252e-08, 2.000353e-08, 1.936752e-08, 1.970971e-08, 
    1.967153e-08, 1.886138e-08, 1.891692e-08, 1.927381e-08, 2.024145e-08,
  1.616979e-08, 1.660164e-08, 1.846045e-08, 1.906519e-08, 2.047339e-08, 
    2.008103e-08, 1.990239e-08, 1.983804e-08, 1.932033e-08, 1.984044e-08, 
    1.958278e-08, 1.886253e-08, 1.955865e-08, 1.975717e-08, 2.053748e-08,
  1.598399e-08, 1.701071e-08, 1.870252e-08, 1.885621e-08, 1.967359e-08, 
    2.000025e-08, 2.010417e-08, 1.985576e-08, 1.959323e-08, 2.023579e-08, 
    1.997097e-08, 1.974834e-08, 2.088441e-08, 1.992134e-08, 2.017184e-08,
  1.628888e-08, 1.751697e-08, 1.810071e-08, 1.852262e-08, 2.009671e-08, 
    2.036254e-08, 2.031294e-08, 1.98099e-08, 2.019891e-08, 2.003867e-08, 
    2.024108e-08, 2.012951e-08, 1.939208e-08, 1.943495e-08, 1.925961e-08,
  1.647676e-08, 1.767802e-08, 1.794087e-08, 1.8762e-08, 2.036675e-08, 
    2.027103e-08, 2.027462e-08, 2.001074e-08, 2.007708e-08, 1.981423e-08, 
    1.926961e-08, 1.917408e-08, 1.95097e-08, 1.83352e-08, 1.924791e-08,
  1.658131e-08, 1.789071e-08, 1.817265e-08, 1.935924e-08, 2.056791e-08, 
    2.042141e-08, 2.036114e-08, 2.029619e-08, 2.033433e-08, 1.944705e-08, 
    1.91941e-08, 1.977211e-08, 1.854378e-08, 1.792426e-08, 2.006384e-08,
  1.719702e-08, 1.823262e-08, 1.850429e-08, 1.983764e-08, 2.067982e-08, 
    2.085715e-08, 2.098598e-08, 2.063204e-08, 2.041105e-08, 1.986747e-08, 
    2.007774e-08, 1.99931e-08, 1.89631e-08, 2.008056e-08, 2.120969e-08,
  1.740051e-08, 1.843397e-08, 1.895337e-08, 2.021664e-08, 2.08851e-08, 
    2.068525e-08, 2.040023e-08, 2.056501e-08, 2.08082e-08, 2.086665e-08, 
    2.08954e-08, 1.994485e-08, 1.954669e-08, 1.9955e-08, 2.087813e-08,
  1.771955e-08, 1.903855e-08, 1.930351e-08, 1.980422e-08, 2.020841e-08, 
    2.029595e-08, 2.043812e-08, 2.052657e-08, 2.109899e-08, 2.105679e-08, 
    2.088002e-08, 2.013403e-08, 2.031054e-08, 2.026576e-08, 2.076758e-08,
  1.811098e-08, 1.805813e-08, 1.899167e-08, 1.96267e-08, 1.936059e-08, 
    2.018207e-08, 2.07e-08, 2.144698e-08, 2.207439e-08, 2.187051e-08, 
    2.255316e-08, 2.172782e-08, 2.139624e-08, 2.07223e-08, 2.022336e-08,
  1.829129e-08, 1.822455e-08, 1.924964e-08, 2.007712e-08, 2.016394e-08, 
    2.057741e-08, 2.062522e-08, 2.212659e-08, 2.216507e-08, 2.198307e-08, 
    2.278393e-08, 2.21266e-08, 2.160513e-08, 2.109135e-08, 2.096685e-08,
  1.887221e-08, 1.891157e-08, 1.987491e-08, 2.060782e-08, 2.084604e-08, 
    2.055404e-08, 2.057816e-08, 2.222327e-08, 2.233895e-08, 2.229388e-08, 
    2.315063e-08, 2.195801e-08, 2.161895e-08, 2.139169e-08, 2.090296e-08,
  1.877658e-08, 1.932682e-08, 2.002296e-08, 1.977912e-08, 1.990229e-08, 
    2.075527e-08, 2.083441e-08, 2.206819e-08, 2.280658e-08, 2.248303e-08, 
    2.313404e-08, 2.209783e-08, 2.243977e-08, 2.142687e-08, 2.053944e-08,
  1.897751e-08, 1.955418e-08, 1.962405e-08, 1.965794e-08, 2.067548e-08, 
    2.132516e-08, 2.152729e-08, 2.240906e-08, 2.305544e-08, 2.081494e-08, 
    2.144346e-08, 2.328173e-08, 2.341119e-08, 2.074443e-08, 2.078919e-08,
  1.915376e-08, 1.943074e-08, 1.892182e-08, 1.90107e-08, 2.037619e-08, 
    2.118365e-08, 2.10702e-08, 2.121279e-08, 2.092422e-08, 1.985045e-08, 
    2.189743e-08, 2.270012e-08, 2.293863e-08, 2.095447e-08, 2.106935e-08,
  1.903387e-08, 1.913949e-08, 1.858596e-08, 1.894899e-08, 2.055232e-08, 
    2.105017e-08, 2.097949e-08, 2.113269e-08, 2.087548e-08, 2.064821e-08, 
    2.254722e-08, 2.295026e-08, 2.263791e-08, 2.166201e-08, 2.283487e-08,
  1.893461e-08, 1.878262e-08, 1.853994e-08, 1.912485e-08, 2.070029e-08, 
    2.124765e-08, 2.107143e-08, 2.10116e-08, 2.085887e-08, 2.107761e-08, 
    2.242507e-08, 2.292194e-08, 2.279441e-08, 2.322961e-08, 2.228115e-08,
  1.900571e-08, 1.863661e-08, 1.884684e-08, 1.924305e-08, 2.060812e-08, 
    2.061903e-08, 2.004686e-08, 2.04042e-08, 2.087852e-08, 2.177037e-08, 
    2.256428e-08, 2.298044e-08, 2.29674e-08, 2.305914e-08, 2.257731e-08,
  1.926777e-08, 1.876479e-08, 1.892871e-08, 1.877705e-08, 1.980615e-08, 
    2.020632e-08, 2.015874e-08, 2.120816e-08, 2.229294e-08, 2.22821e-08, 
    2.283039e-08, 2.30863e-08, 2.290105e-08, 2.283679e-08, 2.270779e-08,
  2.042537e-08, 2.067023e-08, 2.066447e-08, 2.095845e-08, 2.142732e-08, 
    2.160554e-08, 2.271481e-08, 2.433179e-08, 2.666392e-08, 2.604041e-08, 
    2.67907e-08, 2.365526e-08, 2.441686e-08, 2.204351e-08, 2.166974e-08,
  2.094587e-08, 2.101006e-08, 2.102672e-08, 2.208695e-08, 2.189976e-08, 
    2.198823e-08, 2.282507e-08, 2.50555e-08, 2.633925e-08, 2.508171e-08, 
    2.683853e-08, 2.360428e-08, 2.497122e-08, 2.210973e-08, 2.179722e-08,
  2.279092e-08, 2.132706e-08, 2.179923e-08, 2.291952e-08, 2.253021e-08, 
    2.179974e-08, 2.225568e-08, 2.463817e-08, 2.532595e-08, 2.580381e-08, 
    2.812216e-08, 2.384139e-08, 2.53279e-08, 2.161213e-08, 2.187404e-08,
  2.307343e-08, 2.137302e-08, 2.26573e-08, 2.294599e-08, 2.151243e-08, 
    2.141287e-08, 2.174496e-08, 2.451144e-08, 2.551675e-08, 2.579418e-08, 
    2.671941e-08, 2.396715e-08, 2.555799e-08, 2.116249e-08, 2.23724e-08,
  2.34623e-08, 2.233384e-08, 2.311421e-08, 2.25232e-08, 2.156802e-08, 
    2.131278e-08, 2.202626e-08, 2.458301e-08, 2.289504e-08, 2.220837e-08, 
    2.234264e-08, 2.505314e-08, 2.820403e-08, 2.152834e-08, 2.38333e-08,
  2.363328e-08, 2.349069e-08, 2.246109e-08, 2.155651e-08, 2.144279e-08, 
    2.11866e-08, 2.219901e-08, 2.37298e-08, 2.207736e-08, 2.054222e-08, 
    2.31779e-08, 2.493387e-08, 2.506958e-08, 2.338479e-08, 2.406995e-08,
  2.362385e-08, 2.264901e-08, 2.209256e-08, 2.195162e-08, 2.322834e-08, 
    2.268255e-08, 2.269877e-08, 2.283053e-08, 2.151175e-08, 2.201917e-08, 
    2.42286e-08, 2.50016e-08, 2.531255e-08, 2.471221e-08, 2.287248e-08,
  2.473915e-08, 2.392025e-08, 2.279531e-08, 2.342627e-08, 2.546842e-08, 
    2.30964e-08, 2.233346e-08, 2.209393e-08, 2.108159e-08, 2.280084e-08, 
    2.441628e-08, 2.534779e-08, 2.539227e-08, 2.636638e-08, 2.111804e-08,
  2.479895e-08, 2.465004e-08, 2.35917e-08, 2.551496e-08, 2.453459e-08, 
    2.314446e-08, 2.238729e-08, 1.98105e-08, 2.092227e-08, 2.352554e-08, 
    2.437525e-08, 2.540197e-08, 2.562141e-08, 2.341061e-08, 2.137036e-08,
  2.639053e-08, 2.567667e-08, 2.505942e-08, 2.336713e-08, 2.215081e-08, 
    2.121215e-08, 1.979831e-08, 1.929311e-08, 2.29208e-08, 2.444113e-08, 
    2.51816e-08, 2.583803e-08, 2.525705e-08, 2.313347e-08, 2.110871e-08,
  2.303481e-08, 2.31652e-08, 2.409214e-08, 2.557747e-08, 2.543577e-08, 
    2.526885e-08, 2.648063e-08, 2.815598e-08, 3.182259e-08, 2.852344e-08, 
    2.627816e-08, 2.514648e-08, 2.572232e-08, 2.46301e-08, 2.136323e-08,
  2.372701e-08, 2.386928e-08, 2.432769e-08, 2.593567e-08, 2.625376e-08, 
    2.648211e-08, 2.715382e-08, 2.924075e-08, 3.174186e-08, 2.846634e-08, 
    2.694889e-08, 2.407628e-08, 2.58702e-08, 2.455393e-08, 2.116431e-08,
  2.359483e-08, 2.349553e-08, 2.500928e-08, 2.67949e-08, 2.709096e-08, 
    2.696098e-08, 2.741915e-08, 2.953628e-08, 3.084394e-08, 2.842734e-08, 
    2.84656e-08, 2.429168e-08, 2.655544e-08, 2.418466e-08, 2.220916e-08,
  2.264133e-08, 2.293667e-08, 2.520631e-08, 2.708517e-08, 2.704007e-08, 
    2.676391e-08, 2.751727e-08, 2.929895e-08, 2.968797e-08, 2.674878e-08, 
    2.346768e-08, 2.233756e-08, 2.559516e-08, 2.44537e-08, 2.463892e-08,
  2.289575e-08, 2.37174e-08, 2.583801e-08, 2.665778e-08, 2.64836e-08, 
    2.649297e-08, 2.703311e-08, 2.822328e-08, 2.658236e-08, 2.323549e-08, 
    2.158168e-08, 2.371134e-08, 2.50712e-08, 2.716188e-08, 2.718409e-08,
  2.392103e-08, 2.430024e-08, 2.671388e-08, 2.770412e-08, 2.706312e-08, 
    2.699438e-08, 2.708381e-08, 2.727005e-08, 2.570703e-08, 2.53694e-08, 
    2.609243e-08, 2.439724e-08, 2.255379e-08, 2.920015e-08, 2.74892e-08,
  2.376874e-08, 2.583953e-08, 2.755164e-08, 2.718181e-08, 2.711815e-08, 
    2.77793e-08, 2.753732e-08, 2.767475e-08, 2.774766e-08, 2.956281e-08, 
    2.768833e-08, 2.494657e-08, 2.350528e-08, 3.27963e-08, 2.677274e-08,
  2.383764e-08, 2.630968e-08, 2.726966e-08, 2.732934e-08, 2.783654e-08, 
    2.834206e-08, 2.783468e-08, 2.636905e-08, 2.77871e-08, 2.972644e-08, 
    2.793422e-08, 2.46768e-08, 2.412753e-08, 3.042751e-08, 2.54805e-08,
  2.492568e-08, 2.68912e-08, 2.775182e-08, 2.720731e-08, 2.696952e-08, 
    2.763419e-08, 2.616711e-08, 2.456835e-08, 2.821083e-08, 3.107401e-08, 
    2.90016e-08, 2.530684e-08, 2.468957e-08, 2.741572e-08, 2.567885e-08,
  2.554955e-08, 2.729962e-08, 2.638432e-08, 2.599253e-08, 2.542577e-08, 
    2.350461e-08, 2.207926e-08, 2.329701e-08, 2.912794e-08, 3.01722e-08, 
    2.865783e-08, 2.664118e-08, 2.550652e-08, 2.709722e-08, 2.763887e-08,
  2.394683e-08, 2.474588e-08, 2.422519e-08, 2.536507e-08, 2.42111e-08, 
    2.446387e-08, 2.43719e-08, 2.394887e-08, 2.585335e-08, 2.746288e-08, 
    2.845768e-08, 2.616341e-08, 2.323749e-08, 2.893373e-08, 2.898232e-08,
  2.438214e-08, 2.476721e-08, 2.408161e-08, 2.528808e-08, 2.545796e-08, 
    2.563576e-08, 2.434886e-08, 2.395769e-08, 2.585172e-08, 2.709159e-08, 
    2.828297e-08, 2.519806e-08, 2.283988e-08, 2.764283e-08, 2.700481e-08,
  2.496786e-08, 2.542155e-08, 2.470331e-08, 2.536933e-08, 2.633966e-08, 
    2.609294e-08, 2.398254e-08, 2.36344e-08, 2.499983e-08, 2.738268e-08, 
    2.751022e-08, 2.309581e-08, 2.246525e-08, 2.663317e-08, 2.769782e-08,
  2.476953e-08, 2.482339e-08, 2.448612e-08, 2.538838e-08, 2.538478e-08, 
    2.532253e-08, 2.389225e-08, 2.375499e-08, 2.504492e-08, 2.557792e-08, 
    2.293193e-08, 2.113755e-08, 2.121794e-08, 2.592159e-08, 3.198553e-08,
  2.480442e-08, 2.47151e-08, 2.364293e-08, 2.386936e-08, 2.477074e-08, 
    2.46054e-08, 2.323005e-08, 2.363165e-08, 2.387394e-08, 2.233889e-08, 
    2.19219e-08, 2.281836e-08, 2.22073e-08, 2.85629e-08, 3.177177e-08,
  2.496233e-08, 2.40196e-08, 2.357711e-08, 2.46851e-08, 2.498485e-08, 
    2.458261e-08, 2.36472e-08, 2.394529e-08, 2.294956e-08, 2.45095e-08, 
    2.596717e-08, 2.38816e-08, 2.24328e-08, 3.070917e-08, 2.975096e-08,
  2.457311e-08, 2.404404e-08, 2.41937e-08, 2.473043e-08, 2.475595e-08, 
    2.502998e-08, 2.398025e-08, 2.374078e-08, 2.313465e-08, 2.540266e-08, 
    2.539222e-08, 2.372069e-08, 2.384424e-08, 2.92416e-08, 2.758098e-08,
  2.396147e-08, 2.401383e-08, 2.428774e-08, 2.465595e-08, 2.48687e-08, 
    2.502241e-08, 2.438538e-08, 2.412025e-08, 2.3262e-08, 2.443145e-08, 
    2.493589e-08, 2.324041e-08, 2.378314e-08, 2.636578e-08, 2.693668e-08,
  2.38656e-08, 2.441194e-08, 2.436136e-08, 2.424722e-08, 2.431479e-08, 
    2.427979e-08, 2.350784e-08, 2.265535e-08, 2.218346e-08, 2.418095e-08, 
    2.394929e-08, 2.288443e-08, 2.349846e-08, 2.420087e-08, 2.621177e-08,
  2.408795e-08, 2.376037e-08, 2.391661e-08, 2.333993e-08, 2.320998e-08, 
    2.317307e-08, 2.214493e-08, 2.19001e-08, 2.339106e-08, 2.371845e-08, 
    2.338526e-08, 2.290501e-08, 2.25578e-08, 2.349448e-08, 2.616058e-08,
  2.145947e-08, 2.189978e-08, 2.322327e-08, 2.307199e-08, 2.2411e-08, 
    2.202823e-08, 2.245802e-08, 2.252261e-08, 2.411892e-08, 2.402105e-08, 
    2.377347e-08, 2.436462e-08, 2.436808e-08, 2.387077e-08, 2.309506e-08,
  2.18774e-08, 2.269808e-08, 2.331244e-08, 2.3117e-08, 2.309928e-08, 
    2.26498e-08, 2.259027e-08, 2.278676e-08, 2.414895e-08, 2.373863e-08, 
    2.441671e-08, 2.444249e-08, 2.32361e-08, 2.229296e-08, 2.162631e-08,
  2.232921e-08, 2.304023e-08, 2.39044e-08, 2.375397e-08, 2.303136e-08, 
    2.223261e-08, 2.22283e-08, 2.286126e-08, 2.352667e-08, 2.377909e-08, 
    2.495945e-08, 2.306419e-08, 2.240679e-08, 2.208299e-08, 2.222847e-08,
  2.188242e-08, 2.243642e-08, 2.275725e-08, 2.200683e-08, 2.171851e-08, 
    2.18321e-08, 2.224971e-08, 2.275761e-08, 2.322506e-08, 2.309531e-08, 
    2.19665e-08, 2.012046e-08, 2.142328e-08, 2.169356e-08, 2.379028e-08,
  2.217012e-08, 2.237452e-08, 2.213937e-08, 2.152646e-08, 2.163108e-08, 
    2.162126e-08, 2.210829e-08, 2.262169e-08, 2.22276e-08, 2.118571e-08, 
    2.033332e-08, 2.172217e-08, 2.186376e-08, 2.251164e-08, 2.422749e-08,
  2.217444e-08, 2.206928e-08, 2.16113e-08, 2.107526e-08, 2.106537e-08, 
    2.153762e-08, 2.259924e-08, 2.212716e-08, 2.142522e-08, 2.122009e-08, 
    2.186525e-08, 2.242358e-08, 2.191853e-08, 2.328104e-08, 2.209461e-08,
  2.191053e-08, 2.192934e-08, 2.172019e-08, 2.103339e-08, 2.104053e-08, 
    2.160658e-08, 2.225271e-08, 2.189801e-08, 2.161181e-08, 2.161253e-08, 
    2.173614e-08, 2.241962e-08, 2.24185e-08, 2.256619e-08, 2.08881e-08,
  2.20408e-08, 2.170925e-08, 2.144857e-08, 2.078401e-08, 2.106128e-08, 
    2.192768e-08, 2.236344e-08, 2.176439e-08, 2.128701e-08, 2.150037e-08, 
    2.183792e-08, 2.204292e-08, 2.243222e-08, 2.252431e-08, 2.04214e-08,
  2.183525e-08, 2.155139e-08, 2.169162e-08, 2.073586e-08, 2.100262e-08, 
    2.161187e-08, 2.12474e-08, 2.058452e-08, 2.116354e-08, 2.174179e-08, 
    2.17595e-08, 2.189534e-08, 2.204345e-08, 2.109086e-08, 2.016432e-08,
  2.190325e-08, 2.176249e-08, 2.130682e-08, 2.046959e-08, 2.122997e-08, 
    2.157876e-08, 2.078265e-08, 2.033244e-08, 2.130603e-08, 2.165706e-08, 
    2.160298e-08, 2.15834e-08, 2.142227e-08, 2.107361e-08, 2.102351e-08,
  2.19494e-08, 2.239176e-08, 2.328018e-08, 2.284555e-08, 2.216059e-08, 
    2.215979e-08, 2.297922e-08, 2.280069e-08, 2.173358e-08, 2.117228e-08, 
    2.140418e-08, 2.157896e-08, 2.213123e-08, 2.159764e-08, 2.109628e-08,
  2.239094e-08, 2.351105e-08, 2.31057e-08, 2.275633e-08, 2.282441e-08, 
    2.299649e-08, 2.306626e-08, 2.306752e-08, 2.192836e-08, 2.167647e-08, 
    2.164238e-08, 2.164483e-08, 2.150456e-08, 2.097314e-08, 2.11063e-08,
  2.417087e-08, 2.46596e-08, 2.3758e-08, 2.348467e-08, 2.316401e-08, 
    2.243168e-08, 2.266692e-08, 2.286969e-08, 2.185247e-08, 2.190168e-08, 
    2.197633e-08, 2.138027e-08, 2.13923e-08, 2.097974e-08, 2.191588e-08,
  2.358807e-08, 2.340784e-08, 2.29996e-08, 2.198154e-08, 2.186851e-08, 
    2.208198e-08, 2.262292e-08, 2.239277e-08, 2.201962e-08, 2.197137e-08, 
    2.077107e-08, 1.970953e-08, 2.085274e-08, 2.095193e-08, 2.287697e-08,
  2.343532e-08, 2.314665e-08, 2.180219e-08, 2.128754e-08, 2.17592e-08, 
    2.212168e-08, 2.254408e-08, 2.212356e-08, 2.193403e-08, 2.066454e-08, 
    1.939207e-08, 2.087611e-08, 2.109916e-08, 2.179199e-08, 2.361695e-08,
  2.367447e-08, 2.169885e-08, 2.11276e-08, 2.122666e-08, 2.162574e-08, 
    2.170346e-08, 2.220158e-08, 2.198383e-08, 2.053278e-08, 2.007616e-08, 
    2.16289e-08, 2.166357e-08, 2.246392e-08, 2.264004e-08, 2.289119e-08,
  2.293423e-08, 2.151275e-08, 2.142879e-08, 2.139129e-08, 2.151225e-08, 
    2.14295e-08, 2.215077e-08, 2.215819e-08, 2.106562e-08, 2.116202e-08, 
    2.18594e-08, 2.190326e-08, 2.279011e-08, 2.20483e-08, 2.287223e-08,
  2.249556e-08, 2.107932e-08, 2.115659e-08, 2.127148e-08, 2.137145e-08, 
    2.151664e-08, 2.28017e-08, 2.250984e-08, 2.119324e-08, 2.121471e-08, 
    2.209815e-08, 2.205868e-08, 2.288638e-08, 2.305449e-08, 2.090801e-08,
  2.237408e-08, 2.088768e-08, 2.110666e-08, 2.115047e-08, 2.127077e-08, 
    2.090901e-08, 2.159143e-08, 2.207389e-08, 2.139646e-08, 2.214101e-08, 
    2.228923e-08, 2.211787e-08, 2.225767e-08, 2.181496e-08, 2.135132e-08,
  2.18839e-08, 2.046359e-08, 2.015456e-08, 2.051606e-08, 2.101011e-08, 
    2.098814e-08, 2.255875e-08, 2.281818e-08, 2.228582e-08, 2.275044e-08, 
    2.242532e-08, 2.226559e-08, 2.20815e-08, 2.216983e-08, 2.216635e-08,
  2.091008e-08, 2.15206e-08, 2.125255e-08, 2.159614e-08, 2.161775e-08, 
    2.16161e-08, 2.210735e-08, 2.201275e-08, 2.212002e-08, 2.147816e-08, 
    2.195993e-08, 2.229431e-08, 2.215346e-08, 2.29154e-08, 2.235488e-08,
  2.105841e-08, 2.122171e-08, 2.141234e-08, 2.134643e-08, 2.147582e-08, 
    2.161529e-08, 2.164577e-08, 2.132259e-08, 2.127908e-08, 2.149755e-08, 
    2.131021e-08, 2.034043e-08, 2.056757e-08, 2.114985e-08, 2.022234e-08,
  1.972347e-08, 2.116382e-08, 2.183209e-08, 2.144993e-08, 2.054378e-08, 
    2.073256e-08, 2.066159e-08, 2.063677e-08, 2.152187e-08, 2.097742e-08, 
    2.155616e-08, 2.12053e-08, 2.115857e-08, 2.124941e-08, 2.162774e-08,
  1.97753e-08, 2.078608e-08, 2.105661e-08, 2.036463e-08, 2.009709e-08, 
    1.968594e-08, 2.056062e-08, 2.132886e-08, 2.132576e-08, 2.125471e-08, 
    1.98379e-08, 1.849036e-08, 2.068714e-08, 2.1241e-08, 2.519304e-08,
  2.101437e-08, 2.139615e-08, 2.174736e-08, 2.062682e-08, 2.046034e-08, 
    2.047064e-08, 2.059921e-08, 2.091842e-08, 2.102134e-08, 1.957634e-08, 
    1.92652e-08, 2.155727e-08, 2.161291e-08, 2.259771e-08, 2.747238e-08,
  2.177323e-08, 2.090558e-08, 2.144182e-08, 2.065967e-08, 2.02183e-08, 
    2.039967e-08, 2.056952e-08, 2.125287e-08, 2.061039e-08, 2.018504e-08, 
    2.349689e-08, 2.382816e-08, 2.287568e-08, 2.436778e-08, 2.628497e-08,
  2.2255e-08, 2.087162e-08, 2.208059e-08, 2.08489e-08, 2.069999e-08, 
    2.103404e-08, 2.095523e-08, 2.146202e-08, 2.135346e-08, 2.260242e-08, 
    2.364257e-08, 2.301462e-08, 2.318317e-08, 2.436359e-08, 2.273748e-08,
  2.230852e-08, 2.15126e-08, 2.209129e-08, 2.097965e-08, 2.071291e-08, 
    2.096263e-08, 2.145313e-08, 2.197923e-08, 2.13544e-08, 2.300368e-08, 
    2.276387e-08, 2.277509e-08, 2.418602e-08, 2.389517e-08, 2.142548e-08,
  2.248743e-08, 2.131762e-08, 2.216272e-08, 2.144074e-08, 2.087847e-08, 
    2.091491e-08, 2.178882e-08, 2.216774e-08, 2.192121e-08, 2.427547e-08, 
    2.223571e-08, 2.247853e-08, 2.388482e-08, 2.269176e-08, 2.274985e-08,
  2.248278e-08, 2.141479e-08, 2.256806e-08, 2.212531e-08, 2.213134e-08, 
    2.194786e-08, 2.228117e-08, 2.27145e-08, 2.297814e-08, 2.425446e-08, 
    2.186742e-08, 2.267183e-08, 2.382557e-08, 2.41673e-08, 2.343446e-08,
  2.303138e-08, 2.297308e-08, 2.128728e-08, 1.944245e-08, 1.944898e-08, 
    2.00706e-08, 2.094483e-08, 2.087554e-08, 2.058254e-08, 2.03704e-08, 
    2.047093e-08, 2.094167e-08, 2.066309e-08, 2.270492e-08, 2.41214e-08,
  2.338292e-08, 2.320962e-08, 2.058618e-08, 1.901401e-08, 1.910376e-08, 
    2.00134e-08, 2.082071e-08, 2.090614e-08, 2.069631e-08, 2.081943e-08, 
    2.136596e-08, 2.084688e-08, 2.128759e-08, 2.220541e-08, 2.219207e-08,
  2.579123e-08, 2.325013e-08, 2.058044e-08, 1.926199e-08, 1.929339e-08, 
    2.080677e-08, 2.148835e-08, 2.161436e-08, 2.161251e-08, 2.181653e-08, 
    2.203312e-08, 2.181292e-08, 2.278566e-08, 2.283587e-08, 2.169391e-08,
  2.273868e-08, 2.330819e-08, 2.231345e-08, 2.198314e-08, 2.176695e-08, 
    2.152784e-08, 2.181426e-08, 2.175715e-08, 2.170574e-08, 2.243049e-08, 
    2.172764e-08, 2.03911e-08, 2.178171e-08, 2.255069e-08, 2.276736e-08,
  2.274761e-08, 2.301674e-08, 2.385522e-08, 2.417002e-08, 2.288983e-08, 
    2.205728e-08, 2.224054e-08, 2.189132e-08, 2.245234e-08, 2.205012e-08, 
    2.093394e-08, 2.304856e-08, 2.173568e-08, 2.184061e-08, 2.374708e-08,
  2.211144e-08, 2.251214e-08, 2.263104e-08, 2.321248e-08, 2.31912e-08, 
    2.378911e-08, 2.294598e-08, 2.208835e-08, 2.173449e-08, 2.23083e-08, 
    2.332378e-08, 2.36683e-08, 2.186637e-08, 2.040861e-08, 2.490151e-08,
  2.247211e-08, 2.277003e-08, 2.311072e-08, 2.258176e-08, 2.169743e-08, 
    2.237338e-08, 2.316912e-08, 2.238778e-08, 2.13369e-08, 2.19791e-08, 
    2.197989e-08, 2.13046e-08, 1.992151e-08, 2.056007e-08, 2.304336e-08,
  2.21035e-08, 2.255766e-08, 2.274279e-08, 2.289764e-08, 2.16903e-08, 
    2.220814e-08, 2.291394e-08, 2.305897e-08, 2.200967e-08, 2.16903e-08, 
    2.094309e-08, 2.112069e-08, 2.039892e-08, 2.105931e-08, 2.276642e-08,
  2.267906e-08, 2.261479e-08, 2.276163e-08, 2.288587e-08, 2.1719e-08, 
    2.114453e-08, 2.296258e-08, 2.683773e-08, 2.478659e-08, 2.142498e-08, 
    2.069622e-08, 2.031568e-08, 2.062122e-08, 2.164652e-08, 2.109975e-08,
  2.232244e-08, 2.282271e-08, 2.348075e-08, 2.415175e-08, 2.401596e-08, 
    2.338291e-08, 2.284679e-08, 2.334935e-08, 2.26847e-08, 2.235893e-08, 
    2.137929e-08, 1.990498e-08, 2.056303e-08, 2.142554e-08, 2.160199e-08,
  2.45459e-08, 2.530563e-08, 2.592034e-08, 2.606082e-08, 2.344147e-08, 
    2.188219e-08, 2.102487e-08, 2.139942e-08, 2.087007e-08, 2.142548e-08, 
    2.263938e-08, 2.214688e-08, 2.201079e-08, 2.179524e-08, 2.651104e-08,
  2.372208e-08, 2.486663e-08, 2.670436e-08, 2.619735e-08, 2.32196e-08, 
    2.128844e-08, 2.089207e-08, 2.123392e-08, 2.10873e-08, 2.153731e-08, 
    2.205799e-08, 2.17512e-08, 2.170464e-08, 2.291623e-08, 2.460871e-08,
  2.408774e-08, 2.480792e-08, 2.638954e-08, 2.522598e-08, 2.235556e-08, 
    2.230663e-08, 2.13793e-08, 2.107258e-08, 2.11139e-08, 2.130584e-08, 
    2.21645e-08, 2.19321e-08, 2.153829e-08, 2.356271e-08, 2.2475e-08,
  2.414805e-08, 2.541501e-08, 2.554987e-08, 2.54424e-08, 2.574439e-08, 
    2.291941e-08, 2.158902e-08, 2.191883e-08, 2.165072e-08, 2.347814e-08, 
    2.451663e-08, 2.310508e-08, 2.36973e-08, 2.345774e-08, 2.121548e-08,
  2.48091e-08, 2.482583e-08, 2.66999e-08, 2.718926e-08, 2.529047e-08, 
    2.367407e-08, 2.304207e-08, 2.274551e-08, 2.330211e-08, 2.51758e-08, 
    2.447737e-08, 2.464123e-08, 2.375149e-08, 2.195188e-08, 2.025837e-08,
  2.400114e-08, 2.440587e-08, 2.473809e-08, 2.518608e-08, 2.44635e-08, 
    2.365703e-08, 2.333081e-08, 2.287363e-08, 2.369982e-08, 2.43983e-08, 
    2.249253e-08, 2.211906e-08, 2.212726e-08, 1.932361e-08, 1.937762e-08,
  2.437667e-08, 2.457176e-08, 2.489111e-08, 2.477535e-08, 2.407879e-08, 
    2.342798e-08, 2.294402e-08, 2.299597e-08, 2.397914e-08, 2.324074e-08, 
    2.277503e-08, 2.228948e-08, 2.142151e-08, 1.958614e-08, 2.152967e-08,
  2.434129e-08, 2.447753e-08, 2.444579e-08, 2.42785e-08, 2.39121e-08, 
    2.317454e-08, 2.256483e-08, 2.289393e-08, 2.387164e-08, 2.33659e-08, 
    2.268036e-08, 2.259584e-08, 2.15944e-08, 2.143159e-08, 2.363352e-08,
  2.488232e-08, 2.492866e-08, 2.432469e-08, 2.358601e-08, 2.348602e-08, 
    2.296663e-08, 2.259011e-08, 2.430839e-08, 2.410351e-08, 2.322522e-08, 
    2.272805e-08, 2.261863e-08, 2.254304e-08, 2.259997e-08, 2.235889e-08,
  2.50802e-08, 2.492389e-08, 2.376652e-08, 2.29447e-08, 2.237461e-08, 
    2.243472e-08, 2.290855e-08, 2.321451e-08, 2.315763e-08, 2.317915e-08, 
    2.344266e-08, 2.360084e-08, 2.347562e-08, 2.333222e-08, 2.286764e-08,
  2.085997e-08, 2.109208e-08, 2.187947e-08, 2.18914e-08, 2.25749e-08, 
    2.274186e-08, 2.286312e-08, 2.295628e-08, 2.237424e-08, 2.24525e-08, 
    2.323454e-08, 2.268157e-08, 2.290674e-08, 2.194994e-08, 2.121164e-08,
  2.108101e-08, 2.16213e-08, 2.199424e-08, 2.22031e-08, 2.241835e-08, 
    2.250684e-08, 2.275355e-08, 2.278304e-08, 2.235928e-08, 2.251268e-08, 
    2.232166e-08, 2.211884e-08, 2.239183e-08, 2.139629e-08, 2.126741e-08,
  2.000881e-08, 2.118197e-08, 2.203669e-08, 2.227049e-08, 2.243459e-08, 
    2.269704e-08, 2.265404e-08, 2.251239e-08, 2.258844e-08, 2.207368e-08, 
    2.199264e-08, 2.18408e-08, 2.22929e-08, 2.19113e-08, 2.244791e-08,
  2.060645e-08, 2.185038e-08, 2.201148e-08, 2.2231e-08, 2.233474e-08, 
    2.260129e-08, 2.249138e-08, 2.256565e-08, 2.250811e-08, 2.155916e-08, 
    2.261344e-08, 2.333212e-08, 2.346697e-08, 2.333778e-08, 2.25762e-08,
  2.135231e-08, 2.217503e-08, 2.225195e-08, 2.200167e-08, 2.209504e-08, 
    2.238604e-08, 2.218566e-08, 2.233372e-08, 2.141631e-08, 2.116598e-08, 
    2.199716e-08, 2.266141e-08, 2.228827e-08, 2.228473e-08, 2.200858e-08,
  2.183375e-08, 2.199323e-08, 2.199802e-08, 2.196034e-08, 2.21047e-08, 
    2.210736e-08, 2.237819e-08, 2.189144e-08, 2.093715e-08, 2.148637e-08, 
    2.182101e-08, 2.180514e-08, 2.169338e-08, 2.157189e-08, 2.225851e-08,
  2.199654e-08, 2.184973e-08, 2.191579e-08, 2.187763e-08, 2.215153e-08, 
    2.238978e-08, 2.213383e-08, 2.150363e-08, 2.106749e-08, 2.18692e-08, 
    2.208245e-08, 2.200989e-08, 2.20267e-08, 2.170858e-08, 2.269118e-08,
  2.198448e-08, 2.189181e-08, 2.189756e-08, 2.183948e-08, 2.234378e-08, 
    2.224468e-08, 2.205353e-08, 2.151082e-08, 2.156682e-08, 2.200836e-08, 
    2.197986e-08, 2.198378e-08, 2.203779e-08, 2.153816e-08, 2.199192e-08,
  2.204142e-08, 2.188317e-08, 2.174893e-08, 2.198862e-08, 2.23866e-08, 
    2.225087e-08, 2.187778e-08, 2.144416e-08, 2.185181e-08, 2.219451e-08, 
    2.194882e-08, 2.177453e-08, 2.172468e-08, 2.124129e-08, 2.11564e-08,
  2.23013e-08, 2.204246e-08, 2.242142e-08, 2.234393e-08, 2.226598e-08, 
    2.168736e-08, 2.151861e-08, 2.189591e-08, 2.272022e-08, 2.227965e-08, 
    2.185155e-08, 2.164675e-08, 2.156809e-08, 2.145975e-08, 2.160157e-08,
  2.065065e-08, 2.151396e-08, 2.253404e-08, 2.241235e-08, 2.286337e-08, 
    2.301476e-08, 2.304909e-08, 2.3111e-08, 2.255067e-08, 2.251254e-08, 
    2.241925e-08, 2.254088e-08, 2.259843e-08, 2.254083e-08, 2.192362e-08,
  2.038303e-08, 2.156591e-08, 2.240505e-08, 2.294639e-08, 2.318738e-08, 
    2.316876e-08, 2.307084e-08, 2.316407e-08, 2.311681e-08, 2.238866e-08, 
    2.207197e-08, 2.233479e-08, 2.236396e-08, 2.220434e-08, 2.184819e-08,
  2.063294e-08, 2.119094e-08, 2.221876e-08, 2.305676e-08, 2.334419e-08, 
    2.32575e-08, 2.31179e-08, 2.333481e-08, 2.315409e-08, 2.249274e-08, 
    2.256921e-08, 2.23032e-08, 2.242744e-08, 2.234459e-08, 2.267539e-08,
  2.138386e-08, 2.180812e-08, 2.216961e-08, 2.258031e-08, 2.31718e-08, 
    2.322069e-08, 2.320036e-08, 2.312324e-08, 2.290742e-08, 2.26049e-08, 
    2.211063e-08, 2.15117e-08, 2.195897e-08, 2.214097e-08, 2.36217e-08,
  2.182757e-08, 2.172734e-08, 2.233935e-08, 2.286589e-08, 2.331751e-08, 
    2.356059e-08, 2.316306e-08, 2.287014e-08, 2.239507e-08, 2.145699e-08, 
    2.178903e-08, 2.255904e-08, 2.224838e-08, 2.259e-08, 2.442828e-08,
  2.125799e-08, 2.15709e-08, 2.195569e-08, 2.236821e-08, 2.315256e-08, 
    2.324758e-08, 2.275801e-08, 2.247248e-08, 2.185807e-08, 2.183983e-08, 
    2.313023e-08, 2.306761e-08, 2.289311e-08, 2.337562e-08, 2.378802e-08,
  2.10604e-08, 2.136721e-08, 2.179731e-08, 2.201744e-08, 2.283753e-08, 
    2.301434e-08, 2.270075e-08, 2.239706e-08, 2.221864e-08, 2.25745e-08, 
    2.283085e-08, 2.271807e-08, 2.298908e-08, 2.361758e-08, 2.213046e-08,
  2.046663e-08, 2.124591e-08, 2.159674e-08, 2.162286e-08, 2.252761e-08, 
    2.263269e-08, 2.240366e-08, 2.210481e-08, 2.216328e-08, 2.217382e-08, 
    2.258545e-08, 2.298974e-08, 2.376175e-08, 2.375159e-08, 2.226893e-08,
  2.056043e-08, 2.146292e-08, 2.15e-08, 2.13754e-08, 2.22547e-08, 
    2.257311e-08, 2.212396e-08, 2.193011e-08, 2.192344e-08, 2.23349e-08, 
    2.293922e-08, 2.355704e-08, 2.377723e-08, 2.350227e-08, 2.260493e-08,
  2.013082e-08, 2.109786e-08, 2.145377e-08, 2.115837e-08, 2.21223e-08, 
    2.244763e-08, 2.184836e-08, 2.169426e-08, 2.211259e-08, 2.230751e-08, 
    2.315356e-08, 2.367784e-08, 2.397059e-08, 2.361704e-08, 2.336127e-08,
  1.708222e-08, 1.746225e-08, 1.80063e-08, 1.775199e-08, 1.800036e-08, 
    1.80066e-08, 1.7956e-08, 1.77166e-08, 1.773458e-08, 1.829719e-08, 
    1.890314e-08, 1.874571e-08, 1.864534e-08, 1.869221e-08, 1.921054e-08,
  1.703749e-08, 1.727877e-08, 1.755663e-08, 1.79275e-08, 1.840167e-08, 
    1.803617e-08, 1.752508e-08, 1.750923e-08, 1.787967e-08, 1.813316e-08, 
    1.844703e-08, 1.836587e-08, 1.841845e-08, 1.881081e-08, 1.954961e-08,
  1.817927e-08, 1.712341e-08, 1.763749e-08, 1.82914e-08, 1.852243e-08, 
    1.734794e-08, 1.683559e-08, 1.741069e-08, 1.790038e-08, 1.805694e-08, 
    1.863931e-08, 1.801517e-08, 1.82448e-08, 1.893395e-08, 1.952729e-08,
  1.808269e-08, 1.756726e-08, 1.777095e-08, 1.744622e-08, 1.732379e-08, 
    1.707972e-08, 1.666955e-08, 1.704001e-08, 1.75232e-08, 1.804779e-08, 
    1.866708e-08, 1.823553e-08, 1.877229e-08, 1.940742e-08, 1.937139e-08,
  1.856571e-08, 1.748433e-08, 1.771357e-08, 1.765529e-08, 1.757231e-08, 
    1.704679e-08, 1.672104e-08, 1.706232e-08, 1.729344e-08, 1.657352e-08, 
    1.664486e-08, 1.807424e-08, 1.952396e-08, 2.001851e-08, 1.97791e-08,
  1.734502e-08, 1.740783e-08, 1.753182e-08, 1.730779e-08, 1.716155e-08, 
    1.667669e-08, 1.644165e-08, 1.629544e-08, 1.586632e-08, 1.619077e-08, 
    1.702061e-08, 1.746623e-08, 1.94845e-08, 2.06016e-08, 2.013972e-08,
  1.689315e-08, 1.786682e-08, 1.801129e-08, 1.76409e-08, 1.724005e-08, 
    1.652263e-08, 1.635684e-08, 1.624299e-08, 1.620786e-08, 1.646211e-08, 
    1.72302e-08, 1.759376e-08, 1.975492e-08, 2.067042e-08, 2.006833e-08,
  1.686101e-08, 1.853303e-08, 1.831272e-08, 1.781273e-08, 1.736552e-08, 
    1.672257e-08, 1.638282e-08, 1.582956e-08, 1.570294e-08, 1.619021e-08, 
    1.685661e-08, 1.741016e-08, 1.958643e-08, 1.979826e-08, 1.952235e-08,
  1.738862e-08, 1.915307e-08, 1.863104e-08, 1.818994e-08, 1.737953e-08, 
    1.668815e-08, 1.607099e-08, 1.550704e-08, 1.555912e-08, 1.633753e-08, 
    1.698361e-08, 1.769772e-08, 1.904107e-08, 1.934136e-08, 1.969592e-08,
  1.759797e-08, 1.942687e-08, 1.86442e-08, 1.783639e-08, 1.683669e-08, 
    1.616982e-08, 1.557142e-08, 1.545893e-08, 1.590356e-08, 1.635974e-08, 
    1.710277e-08, 1.809901e-08, 1.91995e-08, 1.971157e-08, 2.074139e-08,
  1.924525e-08, 1.943556e-08, 2.035007e-08, 2.112674e-08, 2.058685e-08, 
    2.13928e-08, 2.191258e-08, 2.235034e-08, 2.166976e-08, 2.107112e-08, 
    1.93512e-08, 1.866596e-08, 1.880945e-08, 1.825122e-08, 1.758679e-08,
  2.056479e-08, 2.032058e-08, 2.110748e-08, 2.201383e-08, 2.185844e-08, 
    2.286967e-08, 2.251399e-08, 2.284409e-08, 2.293128e-08, 2.202801e-08, 
    2.011105e-08, 1.968155e-08, 1.957977e-08, 1.846546e-08, 1.798968e-08,
  2.263623e-08, 2.140511e-08, 2.19489e-08, 2.297605e-08, 2.356016e-08, 
    2.296018e-08, 2.230873e-08, 2.213958e-08, 2.22714e-08, 2.125894e-08, 
    2.117843e-08, 2.051272e-08, 1.946793e-08, 1.798518e-08, 1.854217e-08,
  2.108093e-08, 2.085071e-08, 2.165774e-08, 2.316237e-08, 2.261577e-08, 
    2.21992e-08, 2.220299e-08, 2.182277e-08, 2.150394e-08, 2.022474e-08, 
    1.758841e-08, 1.704443e-08, 1.754039e-08, 1.845789e-08, 1.942209e-08,
  2.082854e-08, 2.051863e-08, 2.102727e-08, 2.177346e-08, 2.207847e-08, 
    2.209967e-08, 2.164264e-08, 2.108086e-08, 2.037584e-08, 1.679478e-08, 
    1.626811e-08, 1.750546e-08, 1.837013e-08, 1.952849e-08, 1.990025e-08,
  1.992596e-08, 2.029783e-08, 2.087634e-08, 2.186572e-08, 2.231887e-08, 
    2.227413e-08, 2.159062e-08, 2.069911e-08, 1.91656e-08, 1.835966e-08, 
    2.002141e-08, 1.952918e-08, 1.877854e-08, 2.044781e-08, 1.973134e-08,
  2.01185e-08, 2.104966e-08, 2.141582e-08, 2.253824e-08, 2.283433e-08, 
    2.270753e-08, 2.16594e-08, 2.081112e-08, 2.015275e-08, 1.961537e-08, 
    1.910829e-08, 1.809367e-08, 1.859843e-08, 2.013968e-08, 1.882255e-08,
  1.969904e-08, 2.172072e-08, 2.258362e-08, 2.355564e-08, 2.374892e-08, 
    2.320863e-08, 2.186154e-08, 2.073137e-08, 1.952613e-08, 1.871549e-08, 
    1.900003e-08, 1.964693e-08, 2.06049e-08, 2.059634e-08, 2.021113e-08,
  2.049311e-08, 2.27134e-08, 2.295631e-08, 2.34591e-08, 2.356474e-08, 
    2.288203e-08, 2.09864e-08, 1.984181e-08, 1.941314e-08, 2.00241e-08, 
    2.062279e-08, 2.072499e-08, 2.069189e-08, 2.08375e-08, 2.101703e-08,
  2.032531e-08, 2.305071e-08, 2.352843e-08, 2.328931e-08, 2.335147e-08, 
    2.216101e-08, 2.038375e-08, 1.982814e-08, 2.028082e-08, 2.024625e-08, 
    2.039815e-08, 2.077962e-08, 2.155051e-08, 2.219164e-08, 2.258241e-08,
  1.885921e-08, 1.914431e-08, 2.029652e-08, 2.221789e-08, 2.273644e-08, 
    2.522744e-08, 2.664591e-08, 2.647383e-08, 2.450954e-08, 2.375847e-08, 
    2.457983e-08, 2.448141e-08, 2.430692e-08, 2.401579e-08, 2.360317e-08,
  1.937314e-08, 1.949908e-08, 2.022166e-08, 2.24569e-08, 2.392543e-08, 
    2.490699e-08, 2.58822e-08, 2.691893e-08, 2.508593e-08, 2.405321e-08, 
    2.468607e-08, 2.435282e-08, 2.434313e-08, 2.441909e-08, 2.437966e-08,
  1.936691e-08, 1.900241e-08, 2.063032e-08, 2.330929e-08, 2.364971e-08, 
    2.422975e-08, 2.539714e-08, 2.647428e-08, 2.487292e-08, 2.429324e-08, 
    2.522888e-08, 2.450418e-08, 2.464874e-08, 2.462581e-08, 2.403969e-08,
  1.804687e-08, 1.879303e-08, 1.955717e-08, 2.111732e-08, 2.191908e-08, 
    2.364884e-08, 2.491945e-08, 2.618495e-08, 2.563391e-08, 2.552377e-08, 
    2.603323e-08, 2.620283e-08, 2.623026e-08, 2.520714e-08, 2.379826e-08,
  1.839908e-08, 1.850901e-08, 1.922236e-08, 2.040198e-08, 2.103793e-08, 
    2.311637e-08, 2.520814e-08, 2.633714e-08, 2.493249e-08, 2.471193e-08, 
    2.574563e-08, 2.69685e-08, 2.72334e-08, 2.432098e-08, 2.352112e-08,
  1.773963e-08, 1.844632e-08, 1.867465e-08, 1.991757e-08, 2.117071e-08, 
    2.270898e-08, 2.446136e-08, 2.538099e-08, 2.373593e-08, 2.479398e-08, 
    2.488276e-08, 2.501773e-08, 2.596674e-08, 2.37192e-08, 2.379729e-08,
  1.777729e-08, 1.831899e-08, 1.903873e-08, 1.998607e-08, 2.114571e-08, 
    2.25942e-08, 2.454797e-08, 2.489176e-08, 2.369504e-08, 2.417285e-08, 
    2.49306e-08, 2.521388e-08, 2.504657e-08, 2.366013e-08, 2.50403e-08,
  1.776018e-08, 1.833221e-08, 1.880638e-08, 1.982445e-08, 2.13266e-08, 
    2.238585e-08, 2.403478e-08, 2.447225e-08, 2.371996e-08, 2.447718e-08, 
    2.512368e-08, 2.537749e-08, 2.526314e-08, 2.568024e-08, 2.569681e-08,
  1.757089e-08, 1.85215e-08, 1.880487e-08, 1.99056e-08, 2.136534e-08, 
    2.235964e-08, 2.381318e-08, 2.441151e-08, 2.431315e-08, 2.489347e-08, 
    2.54107e-08, 2.560252e-08, 2.542466e-08, 2.623575e-08, 2.586662e-08,
  1.730571e-08, 1.854469e-08, 1.824293e-08, 1.930908e-08, 2.086028e-08, 
    2.191848e-08, 2.302438e-08, 2.53325e-08, 2.462611e-08, 2.510934e-08, 
    2.553347e-08, 2.570704e-08, 2.570656e-08, 2.609479e-08, 2.582531e-08,
  1.662215e-08, 1.740653e-08, 1.756645e-08, 1.78719e-08, 1.88286e-08, 
    1.968442e-08, 1.977749e-08, 2.089822e-08, 2.251463e-08, 2.215783e-08, 
    2.237531e-08, 2.122203e-08, 2.213609e-08, 2.185876e-08, 2.272149e-08,
  1.763427e-08, 1.799261e-08, 1.776046e-08, 1.811227e-08, 1.951675e-08, 
    2.009443e-08, 1.971399e-08, 2.134591e-08, 2.276864e-08, 2.17467e-08, 
    2.105148e-08, 2.075565e-08, 2.232756e-08, 2.273439e-08, 2.248778e-08,
  1.745055e-08, 1.843185e-08, 1.903953e-08, 1.976948e-08, 2.007849e-08, 
    1.96357e-08, 1.948977e-08, 2.088042e-08, 2.203565e-08, 2.144618e-08, 
    2.121008e-08, 2.077878e-08, 2.219004e-08, 2.229413e-08, 2.223368e-08,
  1.642316e-08, 1.774406e-08, 1.907076e-08, 1.944619e-08, 1.931705e-08, 
    1.907688e-08, 1.954023e-08, 2.046656e-08, 2.113574e-08, 2.03681e-08, 
    1.977157e-08, 2.144853e-08, 2.353076e-08, 2.285945e-08, 2.228208e-08,
  1.684318e-08, 1.876766e-08, 2.003758e-08, 1.917465e-08, 1.891664e-08, 
    1.84943e-08, 1.884051e-08, 1.960862e-08, 1.909551e-08, 1.722054e-08, 
    1.97154e-08, 2.238398e-08, 2.421562e-08, 2.328361e-08, 2.358565e-08,
  1.890754e-08, 1.950701e-08, 1.949981e-08, 1.891281e-08, 1.878933e-08, 
    1.871907e-08, 1.867968e-08, 1.938693e-08, 1.843058e-08, 1.91624e-08, 
    2.078272e-08, 2.106752e-08, 2.271741e-08, 2.417456e-08, 2.460261e-08,
  1.935143e-08, 1.961027e-08, 2.014703e-08, 1.988281e-08, 1.952448e-08, 
    1.937039e-08, 1.935864e-08, 2.034686e-08, 1.941148e-08, 2.004095e-08, 
    2.090453e-08, 2.102021e-08, 2.310654e-08, 2.440233e-08, 2.506651e-08,
  2.020747e-08, 1.937378e-08, 1.992788e-08, 1.971035e-08, 1.974409e-08, 
    1.968131e-08, 2.025793e-08, 2.061015e-08, 1.967675e-08, 2.038269e-08, 
    2.081739e-08, 2.107309e-08, 2.321584e-08, 2.400705e-08, 2.416626e-08,
  1.909262e-08, 1.899847e-08, 1.965389e-08, 1.999016e-08, 1.977599e-08, 
    1.942051e-08, 2.084286e-08, 2.049958e-08, 2.058689e-08, 2.107919e-08, 
    2.084491e-08, 2.201902e-08, 2.389386e-08, 2.421349e-08, 2.491194e-08,
  1.884653e-08, 1.921954e-08, 2.0046e-08, 2.052792e-08, 1.921986e-08, 
    1.979401e-08, 2.120867e-08, 2.123113e-08, 2.113433e-08, 2.085929e-08, 
    2.114351e-08, 2.295829e-08, 2.407746e-08, 2.41002e-08, 2.477782e-08,
  2.081172e-08, 2.057855e-08, 2.016125e-08, 2.090858e-08, 2.110822e-08, 
    2.129195e-08, 2.1468e-08, 2.185949e-08, 2.166503e-08, 2.123038e-08, 
    2.146816e-08, 2.094716e-08, 2.12824e-08, 2.11387e-08, 2.085479e-08,
  2.131527e-08, 2.089472e-08, 2.048685e-08, 2.055753e-08, 2.126974e-08, 
    2.236942e-08, 2.215683e-08, 2.222028e-08, 2.192283e-08, 2.144108e-08, 
    2.136085e-08, 2.087315e-08, 2.097593e-08, 2.121911e-08, 2.085487e-08,
  2.096389e-08, 2.195555e-08, 2.172904e-08, 2.153374e-08, 2.183147e-08, 
    2.279195e-08, 2.209696e-08, 2.22201e-08, 2.198938e-08, 2.135391e-08, 
    2.113867e-08, 2.025649e-08, 2.066159e-08, 2.107946e-08, 2.14471e-08,
  2.148216e-08, 2.152706e-08, 2.143282e-08, 2.154315e-08, 2.18693e-08, 
    2.160469e-08, 2.238762e-08, 2.234812e-08, 2.149578e-08, 2.168673e-08, 
    2.020923e-08, 1.871249e-08, 2.041581e-08, 2.177664e-08, 2.264712e-08,
  2.231666e-08, 2.201727e-08, 2.225121e-08, 2.226518e-08, 2.190845e-08, 
    2.193515e-08, 2.21733e-08, 2.182722e-08, 2.205045e-08, 2.238336e-08, 
    2.199765e-08, 2.120402e-08, 2.071748e-08, 2.184314e-08, 2.173293e-08,
  2.248502e-08, 2.181994e-08, 2.191199e-08, 2.197252e-08, 2.179856e-08, 
    2.244318e-08, 2.176951e-08, 2.251813e-08, 2.240514e-08, 2.211853e-08, 
    2.273418e-08, 2.258236e-08, 2.17932e-08, 2.097127e-08, 2.277412e-08,
  2.262306e-08, 2.216843e-08, 2.185622e-08, 2.208723e-08, 2.20944e-08, 
    2.241485e-08, 2.207754e-08, 2.278307e-08, 2.214072e-08, 2.232221e-08, 
    2.238628e-08, 2.227151e-08, 2.181394e-08, 2.150689e-08, 2.296928e-08,
  2.257675e-08, 2.224703e-08, 2.178211e-08, 2.20127e-08, 2.185205e-08, 
    2.211719e-08, 2.212036e-08, 2.254965e-08, 2.222892e-08, 2.264032e-08, 
    2.305606e-08, 2.262469e-08, 2.182816e-08, 2.166731e-08, 2.265477e-08,
  2.277139e-08, 2.258105e-08, 2.188733e-08, 2.197209e-08, 2.202249e-08, 
    2.233113e-08, 2.296716e-08, 2.330066e-08, 2.31647e-08, 2.327851e-08, 
    2.274237e-08, 2.194035e-08, 2.172029e-08, 2.199632e-08, 2.262835e-08,
  2.297164e-08, 2.277718e-08, 2.194707e-08, 2.204299e-08, 2.213595e-08, 
    2.304655e-08, 2.314763e-08, 2.333876e-08, 2.283614e-08, 2.226366e-08, 
    2.178871e-08, 2.192101e-08, 2.222875e-08, 2.232276e-08, 2.236488e-08,
  2.361993e-08, 2.442317e-08, 2.472582e-08, 2.447011e-08, 2.412262e-08, 
    2.407224e-08, 2.364455e-08, 2.391664e-08, 2.310348e-08, 2.225938e-08, 
    2.215094e-08, 2.162377e-08, 2.162796e-08, 2.186113e-08, 2.209142e-08,
  2.417237e-08, 2.495761e-08, 2.493818e-08, 2.452045e-08, 2.42504e-08, 
    2.418368e-08, 2.372499e-08, 2.384026e-08, 2.280778e-08, 2.235318e-08, 
    2.156282e-08, 2.13522e-08, 2.138386e-08, 2.189287e-08, 2.189127e-08,
  2.519645e-08, 2.519951e-08, 2.465568e-08, 2.449097e-08, 2.44146e-08, 
    2.399744e-08, 2.342616e-08, 2.327136e-08, 2.252221e-08, 2.168271e-08, 
    2.133535e-08, 2.145818e-08, 2.156222e-08, 2.222251e-08, 2.251372e-08,
  2.516667e-08, 2.493957e-08, 2.449954e-08, 2.425817e-08, 2.416457e-08, 
    2.399879e-08, 2.346112e-08, 2.2921e-08, 2.208681e-08, 2.197292e-08, 
    2.283772e-08, 2.299878e-08, 2.309362e-08, 2.305766e-08, 2.277488e-08,
  2.557023e-08, 2.51822e-08, 2.473455e-08, 2.476616e-08, 2.476304e-08, 
    2.459496e-08, 2.376909e-08, 2.289646e-08, 2.221763e-08, 2.261351e-08, 
    2.301737e-08, 2.329415e-08, 2.266606e-08, 2.217674e-08, 2.186247e-08,
  2.521367e-08, 2.457761e-08, 2.442749e-08, 2.48016e-08, 2.477335e-08, 
    2.434806e-08, 2.311119e-08, 2.243509e-08, 2.221923e-08, 2.263758e-08, 
    2.233298e-08, 2.193934e-08, 2.206637e-08, 2.132126e-08, 2.171019e-08,
  2.455754e-08, 2.462221e-08, 2.501029e-08, 2.523517e-08, 2.505043e-08, 
    2.412128e-08, 2.283636e-08, 2.221396e-08, 2.239918e-08, 2.211026e-08, 
    2.215542e-08, 2.192914e-08, 2.168042e-08, 2.100195e-08, 2.18766e-08,
  2.422249e-08, 2.5179e-08, 2.557068e-08, 2.550942e-08, 2.49747e-08, 
    2.334099e-08, 2.221111e-08, 2.177088e-08, 2.214735e-08, 2.224485e-08, 
    2.219784e-08, 2.176227e-08, 2.160345e-08, 2.135649e-08, 2.165386e-08,
  2.36025e-08, 2.570817e-08, 2.639413e-08, 2.559659e-08, 2.466816e-08, 
    2.261974e-08, 2.170233e-08, 2.222482e-08, 2.238136e-08, 2.212214e-08, 
    2.190092e-08, 2.166442e-08, 2.166823e-08, 2.172786e-08, 2.20547e-08,
  2.389826e-08, 2.574526e-08, 2.655934e-08, 2.516723e-08, 2.335844e-08, 
    2.192077e-08, 2.146763e-08, 2.181301e-08, 2.188426e-08, 2.191841e-08, 
    2.180747e-08, 2.160904e-08, 2.154748e-08, 2.182383e-08, 2.181903e-08,
  2.055949e-08, 2.169707e-08, 2.276465e-08, 2.373187e-08, 2.393993e-08, 
    2.390383e-08, 2.423569e-08, 2.419809e-08, 2.43893e-08, 2.42548e-08, 
    2.529184e-08, 2.546818e-08, 2.600729e-08, 2.554474e-08, 2.474672e-08,
  2.167314e-08, 2.300428e-08, 2.33998e-08, 2.402467e-08, 2.363491e-08, 
    2.397928e-08, 2.393704e-08, 2.433395e-08, 2.477486e-08, 2.563279e-08, 
    2.644726e-08, 2.633438e-08, 2.61125e-08, 2.49798e-08, 2.384101e-08,
  2.302397e-08, 2.390818e-08, 2.41569e-08, 2.434424e-08, 2.342201e-08, 
    2.421998e-08, 2.44776e-08, 2.536115e-08, 2.642971e-08, 2.686856e-08, 
    2.667859e-08, 2.587397e-08, 2.520271e-08, 2.328534e-08, 2.337737e-08,
  2.293951e-08, 2.399198e-08, 2.415037e-08, 2.364258e-08, 2.372679e-08, 
    2.438332e-08, 2.513996e-08, 2.676473e-08, 2.720417e-08, 2.677058e-08, 
    2.543334e-08, 2.412791e-08, 2.333619e-08, 2.251104e-08, 2.304236e-08,
  2.336839e-08, 2.469622e-08, 2.428937e-08, 2.440327e-08, 2.533257e-08, 
    2.628685e-08, 2.761976e-08, 2.8245e-08, 2.766599e-08, 2.548435e-08, 
    2.333324e-08, 2.2947e-08, 2.235341e-08, 2.222884e-08, 2.270192e-08,
  2.440497e-08, 2.443227e-08, 2.414805e-08, 2.536263e-08, 2.618259e-08, 
    2.743434e-08, 2.76247e-08, 2.705118e-08, 2.519109e-08, 2.341002e-08, 
    2.31341e-08, 2.210411e-08, 2.191912e-08, 2.223397e-08, 2.174774e-08,
  2.457737e-08, 2.44844e-08, 2.506568e-08, 2.673321e-08, 2.744104e-08, 
    2.781908e-08, 2.745638e-08, 2.605073e-08, 2.397641e-08, 2.284353e-08, 
    2.234658e-08, 2.181041e-08, 2.19173e-08, 2.200244e-08, 2.169068e-08,
  2.502585e-08, 2.514724e-08, 2.656637e-08, 2.769657e-08, 2.748298e-08, 
    2.740566e-08, 2.597752e-08, 2.420025e-08, 2.296922e-08, 2.246837e-08, 
    2.225752e-08, 2.18762e-08, 2.186736e-08, 2.202208e-08, 2.215802e-08,
  2.459522e-08, 2.629263e-08, 2.758344e-08, 2.765823e-08, 2.716307e-08, 
    2.670052e-08, 2.46143e-08, 2.370722e-08, 2.321861e-08, 2.261574e-08, 
    2.224655e-08, 2.201678e-08, 2.205091e-08, 2.282277e-08, 2.29895e-08,
  2.511112e-08, 2.64218e-08, 2.709558e-08, 2.691555e-08, 2.659015e-08, 
    2.522412e-08, 2.394382e-08, 2.362761e-08, 2.273772e-08, 2.22985e-08, 
    2.23365e-08, 2.253782e-08, 2.270011e-08, 2.325819e-08, 2.367282e-08,
  2.132353e-08, 2.167759e-08, 2.183602e-08, 2.236851e-08, 2.259874e-08, 
    2.304358e-08, 2.38495e-08, 2.42505e-08, 2.448578e-08, 2.428019e-08, 
    2.513226e-08, 2.519329e-08, 2.552924e-08, 2.546625e-08, 2.573509e-08,
  2.254453e-08, 2.273777e-08, 2.258642e-08, 2.309902e-08, 2.316017e-08, 
    2.397706e-08, 2.423385e-08, 2.458127e-08, 2.462758e-08, 2.481094e-08, 
    2.537312e-08, 2.518014e-08, 2.564935e-08, 2.548182e-08, 2.552238e-08,
  2.157101e-08, 2.277425e-08, 2.32737e-08, 2.363558e-08, 2.361549e-08, 
    2.461734e-08, 2.451937e-08, 2.471513e-08, 2.47859e-08, 2.492799e-08, 
    2.53242e-08, 2.510824e-08, 2.548007e-08, 2.520945e-08, 2.522766e-08,
  2.223852e-08, 2.338866e-08, 2.353101e-08, 2.384563e-08, 2.413865e-08, 
    2.461131e-08, 2.441507e-08, 2.476582e-08, 2.46391e-08, 2.554775e-08, 
    2.511904e-08, 2.534007e-08, 2.529447e-08, 2.488119e-08, 2.498632e-08,
  2.338419e-08, 2.422764e-08, 2.450562e-08, 2.462129e-08, 2.475037e-08, 
    2.484389e-08, 2.511705e-08, 2.499077e-08, 2.55057e-08, 2.565952e-08, 
    2.503983e-08, 2.509606e-08, 2.455767e-08, 2.442021e-08, 2.49396e-08,
  2.390398e-08, 2.380562e-08, 2.365662e-08, 2.416935e-08, 2.421827e-08, 
    2.463353e-08, 2.458619e-08, 2.476116e-08, 2.508953e-08, 2.517266e-08, 
    2.472512e-08, 2.441132e-08, 2.448438e-08, 2.413065e-08, 2.469787e-08,
  2.320385e-08, 2.337514e-08, 2.360477e-08, 2.429705e-08, 2.444926e-08, 
    2.456362e-08, 2.455185e-08, 2.477755e-08, 2.520656e-08, 2.452513e-08, 
    2.439383e-08, 2.440397e-08, 2.423326e-08, 2.420176e-08, 2.490962e-08,
  2.378534e-08, 2.356521e-08, 2.381113e-08, 2.427596e-08, 2.3866e-08, 
    2.362285e-08, 2.365014e-08, 2.399486e-08, 2.462202e-08, 2.457925e-08, 
    2.46486e-08, 2.448542e-08, 2.444213e-08, 2.478618e-08, 2.560214e-08,
  2.285501e-08, 2.321534e-08, 2.376298e-08, 2.397194e-08, 2.343765e-08, 
    2.342134e-08, 2.357921e-08, 2.501555e-08, 2.530235e-08, 2.468517e-08, 
    2.44767e-08, 2.433433e-08, 2.454873e-08, 2.521603e-08, 2.520961e-08,
  2.330521e-08, 2.38966e-08, 2.43312e-08, 2.405687e-08, 2.398265e-08, 
    2.426664e-08, 2.440883e-08, 2.490608e-08, 2.417603e-08, 2.401968e-08, 
    2.422974e-08, 2.448541e-08, 2.46922e-08, 2.495451e-08, 2.49206e-08,
  2.205774e-08, 2.148321e-08, 2.103753e-08, 2.066744e-08, 2.086352e-08, 
    2.115173e-08, 2.169496e-08, 2.220533e-08, 2.213272e-08, 2.232483e-08, 
    2.286512e-08, 2.276021e-08, 2.266691e-08, 2.23417e-08, 2.222526e-08,
  2.09074e-08, 2.041489e-08, 2.081296e-08, 2.105174e-08, 2.129063e-08, 
    2.152927e-08, 2.214638e-08, 2.222124e-08, 2.202175e-08, 2.211103e-08, 
    2.233108e-08, 2.207791e-08, 2.193067e-08, 2.214655e-08, 2.25168e-08,
  1.966573e-08, 2.057963e-08, 2.122328e-08, 2.154064e-08, 2.176192e-08, 
    2.231517e-08, 2.239309e-08, 2.199614e-08, 2.196507e-08, 2.200503e-08, 
    2.214197e-08, 2.189161e-08, 2.228813e-08, 2.283057e-08, 2.333991e-08,
  2.07203e-08, 2.205178e-08, 2.182524e-08, 2.197927e-08, 2.242952e-08, 
    2.250281e-08, 2.212579e-08, 2.193983e-08, 2.230991e-08, 2.276448e-08, 
    2.35649e-08, 2.445209e-08, 2.439139e-08, 2.41477e-08, 2.344663e-08,
  2.230444e-08, 2.339347e-08, 2.353261e-08, 2.368167e-08, 2.339693e-08, 
    2.325783e-08, 2.288741e-08, 2.295888e-08, 2.342929e-08, 2.398003e-08, 
    2.449233e-08, 2.452137e-08, 2.41714e-08, 2.353756e-08, 2.301196e-08,
  2.311409e-08, 2.30241e-08, 2.284923e-08, 2.308509e-08, 2.273621e-08, 
    2.280781e-08, 2.300112e-08, 2.342918e-08, 2.362025e-08, 2.398035e-08, 
    2.351146e-08, 2.320793e-08, 2.364878e-08, 2.337752e-08, 2.360376e-08,
  2.317437e-08, 2.346059e-08, 2.346686e-08, 2.320205e-08, 2.30357e-08, 
    2.316948e-08, 2.345304e-08, 2.328674e-08, 2.385917e-08, 2.34114e-08, 
    2.350248e-08, 2.346312e-08, 2.342785e-08, 2.333706e-08, 2.416668e-08,
  2.378585e-08, 2.367079e-08, 2.305769e-08, 2.285876e-08, 2.290047e-08, 
    2.303318e-08, 2.305789e-08, 2.299466e-08, 2.376642e-08, 2.359964e-08, 
    2.375475e-08, 2.336965e-08, 2.331072e-08, 2.339422e-08, 2.38317e-08,
  2.291026e-08, 2.306681e-08, 2.322848e-08, 2.339468e-08, 2.370834e-08, 
    2.359919e-08, 2.354831e-08, 2.43307e-08, 2.444764e-08, 2.367307e-08, 
    2.34106e-08, 2.301833e-08, 2.298475e-08, 2.361051e-08, 2.405166e-08,
  2.278567e-08, 2.310737e-08, 2.361212e-08, 2.348838e-08, 2.39174e-08, 
    2.441738e-08, 2.435677e-08, 2.396528e-08, 2.318587e-08, 2.302185e-08, 
    2.310964e-08, 2.288041e-08, 2.298645e-08, 2.383708e-08, 2.429871e-08,
  2.110937e-08, 2.195915e-08, 2.220436e-08, 2.214769e-08, 2.21468e-08, 
    2.215702e-08, 2.238925e-08, 2.271367e-08, 2.274141e-08, 2.226575e-08, 
    2.28869e-08, 2.261248e-08, 2.283255e-08, 2.26623e-08, 2.237441e-08,
  2.176901e-08, 2.220123e-08, 2.207963e-08, 2.214792e-08, 2.197815e-08, 
    2.209661e-08, 2.243615e-08, 2.270063e-08, 2.264595e-08, 2.234994e-08, 
    2.2612e-08, 2.230087e-08, 2.239969e-08, 2.252584e-08, 2.238031e-08,
  2.247212e-08, 2.259197e-08, 2.22376e-08, 2.215458e-08, 2.184693e-08, 
    2.249528e-08, 2.25186e-08, 2.254862e-08, 2.24891e-08, 2.250693e-08, 
    2.258498e-08, 2.222023e-08, 2.272312e-08, 2.310913e-08, 2.338163e-08,
  2.237616e-08, 2.221443e-08, 2.215925e-08, 2.193557e-08, 2.198771e-08, 
    2.218702e-08, 2.222211e-08, 2.224375e-08, 2.24561e-08, 2.282677e-08, 
    2.256271e-08, 2.312423e-08, 2.361912e-08, 2.400026e-08, 2.448854e-08,
  2.200782e-08, 2.236736e-08, 2.193821e-08, 2.173102e-08, 2.169963e-08, 
    2.176418e-08, 2.211452e-08, 2.275901e-08, 2.338084e-08, 2.315633e-08, 
    2.318085e-08, 2.315504e-08, 2.30847e-08, 2.350329e-08, 2.427033e-08,
  2.279648e-08, 2.191849e-08, 2.112522e-08, 2.129626e-08, 2.120807e-08, 
    2.174358e-08, 2.263926e-08, 2.292924e-08, 2.263377e-08, 2.261623e-08, 
    2.265629e-08, 2.220663e-08, 2.316881e-08, 2.387546e-08, 2.38731e-08,
  2.184558e-08, 2.134101e-08, 2.099643e-08, 2.109407e-08, 2.154537e-08, 
    2.246913e-08, 2.265691e-08, 2.266132e-08, 2.234334e-08, 2.195102e-08, 
    2.224517e-08, 2.239504e-08, 2.394989e-08, 2.485052e-08, 2.373064e-08,
  2.105905e-08, 2.096852e-08, 2.079047e-08, 2.135285e-08, 2.182372e-08, 
    2.223345e-08, 2.203419e-08, 2.198064e-08, 2.148604e-08, 2.213558e-08, 
    2.258743e-08, 2.308078e-08, 2.459876e-08, 2.482402e-08, 2.371559e-08,
  2.104759e-08, 2.097708e-08, 2.118772e-08, 2.167632e-08, 2.163342e-08, 
    2.192332e-08, 2.19122e-08, 2.19037e-08, 2.231657e-08, 2.261215e-08, 
    2.289164e-08, 2.357527e-08, 2.465405e-08, 2.417838e-08, 2.358521e-08,
  2.114888e-08, 2.092414e-08, 2.110823e-08, 2.151451e-08, 2.113501e-08, 
    2.154299e-08, 2.162803e-08, 2.25386e-08, 2.242593e-08, 2.267862e-08, 
    2.355137e-08, 2.42837e-08, 2.443312e-08, 2.416746e-08, 2.429262e-08,
  2.047782e-08, 2.050709e-08, 2.053699e-08, 2.043166e-08, 2.026931e-08, 
    2.043878e-08, 2.046625e-08, 2.073315e-08, 2.085256e-08, 2.03472e-08, 
    2.092282e-08, 2.077136e-08, 2.108205e-08, 2.117096e-08, 2.066545e-08,
  2.029654e-08, 2.035675e-08, 1.996814e-08, 1.99933e-08, 2.03323e-08, 
    2.10229e-08, 2.134251e-08, 2.129969e-08, 2.110409e-08, 2.090261e-08, 
    2.105689e-08, 2.111435e-08, 2.110427e-08, 2.107107e-08, 2.080595e-08,
  1.945131e-08, 1.996387e-08, 2.009041e-08, 2.063521e-08, 2.054577e-08, 
    2.122835e-08, 2.123934e-08, 2.130497e-08, 2.11621e-08, 2.11134e-08, 
    2.115179e-08, 2.107981e-08, 2.105538e-08, 2.106374e-08, 2.12518e-08,
  1.91162e-08, 1.954681e-08, 1.977849e-08, 2.014165e-08, 2.101616e-08, 
    2.148126e-08, 2.152933e-08, 2.163045e-08, 2.110814e-08, 2.179594e-08, 
    2.122652e-08, 2.121661e-08, 2.121459e-08, 2.138032e-08, 2.143623e-08,
  1.929051e-08, 2.029687e-08, 2.10286e-08, 2.21014e-08, 2.259279e-08, 
    2.251265e-08, 2.234261e-08, 2.195759e-08, 2.194417e-08, 2.265851e-08, 
    2.244519e-08, 2.221074e-08, 2.185632e-08, 2.186526e-08, 2.203786e-08,
  1.966121e-08, 2.034533e-08, 2.168514e-08, 2.283332e-08, 2.243411e-08, 
    2.244605e-08, 2.194809e-08, 2.225567e-08, 2.280219e-08, 2.268563e-08, 
    2.249906e-08, 2.210417e-08, 2.215921e-08, 2.194095e-08, 2.286028e-08,
  1.968611e-08, 2.086123e-08, 2.216558e-08, 2.269324e-08, 2.24514e-08, 
    2.246445e-08, 2.247267e-08, 2.300534e-08, 2.288905e-08, 2.245657e-08, 
    2.232765e-08, 2.22584e-08, 2.242332e-08, 2.260322e-08, 2.31106e-08,
  2.015718e-08, 2.16262e-08, 2.257623e-08, 2.31609e-08, 2.251964e-08, 
    2.231788e-08, 2.23968e-08, 2.272788e-08, 2.28469e-08, 2.285507e-08, 
    2.275891e-08, 2.283615e-08, 2.36176e-08, 2.326619e-08, 2.286035e-08,
  2.040277e-08, 2.238628e-08, 2.306578e-08, 2.307853e-08, 2.270422e-08, 
    2.268223e-08, 2.291245e-08, 2.425272e-08, 2.397559e-08, 2.298666e-08, 
    2.325302e-08, 2.357095e-08, 2.406451e-08, 2.355144e-08, 2.307846e-08,
  2.097872e-08, 2.26696e-08, 2.313164e-08, 2.356719e-08, 2.431539e-08, 
    2.423673e-08, 2.444299e-08, 2.440371e-08, 2.320486e-08, 2.353027e-08, 
    2.413672e-08, 2.420989e-08, 2.400344e-08, 2.340754e-08, 2.325812e-08,
  2.114997e-08, 2.029401e-08, 2.019966e-08, 1.978111e-08, 2.004871e-08, 
    2.024771e-08, 2.121247e-08, 2.173456e-08, 2.237708e-08, 2.249923e-08, 
    2.361139e-08, 2.353603e-08, 2.341715e-08, 2.340705e-08, 2.260838e-08,
  2.067105e-08, 2.00024e-08, 2.008659e-08, 1.996163e-08, 2.030079e-08, 
    2.102178e-08, 2.216642e-08, 2.261756e-08, 2.328725e-08, 2.33383e-08, 
    2.386668e-08, 2.361892e-08, 2.330447e-08, 2.356862e-08, 2.298555e-08,
  1.981741e-08, 1.994013e-08, 2.000748e-08, 2.033182e-08, 2.070893e-08, 
    2.238032e-08, 2.308432e-08, 2.319741e-08, 2.391475e-08, 2.379699e-08, 
    2.399273e-08, 2.353127e-08, 2.348697e-08, 2.374773e-08, 2.387567e-08,
  1.984263e-08, 2.006874e-08, 1.989184e-08, 2.031813e-08, 2.182283e-08, 
    2.300987e-08, 2.35309e-08, 2.409634e-08, 2.424184e-08, 2.474272e-08, 
    2.568779e-08, 2.625993e-08, 2.551593e-08, 2.50488e-08, 2.367747e-08,
  2.036971e-08, 2.064998e-08, 2.111361e-08, 2.216738e-08, 2.317826e-08, 
    2.419112e-08, 2.499836e-08, 2.49246e-08, 2.515618e-08, 2.574975e-08, 
    2.609658e-08, 2.606098e-08, 2.507849e-08, 2.452302e-08, 2.389223e-08,
  2.063038e-08, 2.067654e-08, 2.114004e-08, 2.227197e-08, 2.30147e-08, 
    2.416473e-08, 2.429042e-08, 2.415054e-08, 2.432851e-08, 2.523947e-08, 
    2.427169e-08, 2.33274e-08, 2.435474e-08, 2.384769e-08, 2.364338e-08,
  2.078382e-08, 2.113341e-08, 2.150487e-08, 2.225761e-08, 2.328521e-08, 
    2.404632e-08, 2.448636e-08, 2.443708e-08, 2.497094e-08, 2.412868e-08, 
    2.372069e-08, 2.353877e-08, 2.420251e-08, 2.368873e-08, 2.333876e-08,
  2.147401e-08, 2.132206e-08, 2.151286e-08, 2.264487e-08, 2.312606e-08, 
    2.391129e-08, 2.42678e-08, 2.404084e-08, 2.454378e-08, 2.443748e-08, 
    2.408913e-08, 2.376576e-08, 2.419603e-08, 2.309992e-08, 2.322698e-08,
  2.154935e-08, 2.148224e-08, 2.200708e-08, 2.278329e-08, 2.332541e-08, 
    2.400579e-08, 2.436486e-08, 2.582539e-08, 2.571016e-08, 2.428983e-08, 
    2.367969e-08, 2.354588e-08, 2.343043e-08, 2.323949e-08, 2.349008e-08,
  2.180668e-08, 2.193121e-08, 2.225667e-08, 2.342629e-08, 2.4191e-08, 
    2.492334e-08, 2.568408e-08, 2.531037e-08, 2.413809e-08, 2.401876e-08, 
    2.360943e-08, 2.325876e-08, 2.32705e-08, 2.397794e-08, 2.34539e-08,
  2.37377e-08, 2.406801e-08, 2.406992e-08, 2.399907e-08, 2.393014e-08, 
    2.36867e-08, 2.331338e-08, 2.308947e-08, 2.274424e-08, 2.25142e-08, 
    2.293299e-08, 2.254263e-08, 2.289154e-08, 2.307532e-08, 2.272412e-08,
  2.343943e-08, 2.359052e-08, 2.419404e-08, 2.418924e-08, 2.393013e-08, 
    2.369127e-08, 2.333795e-08, 2.318423e-08, 2.298759e-08, 2.267921e-08, 
    2.307097e-08, 2.271969e-08, 2.302305e-08, 2.324587e-08, 2.264325e-08,
  2.394085e-08, 2.378253e-08, 2.39012e-08, 2.370828e-08, 2.36997e-08, 
    2.365485e-08, 2.343553e-08, 2.289693e-08, 2.289833e-08, 2.274608e-08, 
    2.300127e-08, 2.308001e-08, 2.337408e-08, 2.362671e-08, 2.406447e-08,
  2.404933e-08, 2.404986e-08, 2.399636e-08, 2.412291e-08, 2.419058e-08, 
    2.388216e-08, 2.341381e-08, 2.304868e-08, 2.297591e-08, 2.33154e-08, 
    2.350786e-08, 2.414069e-08, 2.408714e-08, 2.420277e-08, 2.415522e-08,
  2.427575e-08, 2.421845e-08, 2.440746e-08, 2.437818e-08, 2.416662e-08, 
    2.386816e-08, 2.369758e-08, 2.335732e-08, 2.346582e-08, 2.390161e-08, 
    2.49286e-08, 2.55231e-08, 2.455163e-08, 2.45458e-08, 2.389695e-08,
  2.359091e-08, 2.406071e-08, 2.416486e-08, 2.435041e-08, 2.416165e-08, 
    2.3809e-08, 2.367003e-08, 2.339891e-08, 2.354821e-08, 2.47685e-08, 
    2.459264e-08, 2.36822e-08, 2.393819e-08, 2.328754e-08, 2.329771e-08,
  2.307164e-08, 2.390857e-08, 2.440339e-08, 2.445839e-08, 2.424856e-08, 
    2.403305e-08, 2.37314e-08, 2.360709e-08, 2.421379e-08, 2.435416e-08, 
    2.409019e-08, 2.366121e-08, 2.404583e-08, 2.318005e-08, 2.330396e-08,
  2.278593e-08, 2.402447e-08, 2.430992e-08, 2.450055e-08, 2.419219e-08, 
    2.383262e-08, 2.339848e-08, 2.351296e-08, 2.409169e-08, 2.470478e-08, 
    2.441369e-08, 2.411411e-08, 2.436239e-08, 2.334978e-08, 2.363318e-08,
  2.264195e-08, 2.374956e-08, 2.432042e-08, 2.441101e-08, 2.416252e-08, 
    2.375075e-08, 2.34987e-08, 2.427281e-08, 2.493485e-08, 2.464549e-08, 
    2.430901e-08, 2.405038e-08, 2.424277e-08, 2.389425e-08, 2.396732e-08,
  2.250644e-08, 2.337818e-08, 2.39851e-08, 2.425499e-08, 2.410187e-08, 
    2.384526e-08, 2.356899e-08, 2.406574e-08, 2.411004e-08, 2.436398e-08, 
    2.464626e-08, 2.439581e-08, 2.437734e-08, 2.459428e-08, 2.451537e-08,
  2.251214e-08, 2.346937e-08, 2.32287e-08, 2.289798e-08, 2.288795e-08, 
    2.311216e-08, 2.348663e-08, 2.360879e-08, 2.437596e-08, 2.427102e-08, 
    2.601802e-08, 2.575235e-08, 2.62114e-08, 2.734388e-08, 2.778794e-08,
  2.265516e-08, 2.288471e-08, 2.294606e-08, 2.275421e-08, 2.2736e-08, 
    2.305599e-08, 2.342672e-08, 2.367915e-08, 2.354949e-08, 2.422397e-08, 
    2.527183e-08, 2.486419e-08, 2.564894e-08, 2.633254e-08, 2.535206e-08,
  2.327228e-08, 2.29212e-08, 2.29318e-08, 2.267783e-08, 2.245073e-08, 
    2.293017e-08, 2.334904e-08, 2.347112e-08, 2.328007e-08, 2.381533e-08, 
    2.358246e-08, 2.374758e-08, 2.462411e-08, 2.51829e-08, 2.439086e-08,
  2.236225e-08, 2.327269e-08, 2.307264e-08, 2.318106e-08, 2.289152e-08, 
    2.264086e-08, 2.317912e-08, 2.349669e-08, 2.347084e-08, 2.423503e-08, 
    2.420076e-08, 2.275976e-08, 2.347107e-08, 2.375135e-08, 2.364125e-08,
  2.246843e-08, 2.315429e-08, 2.389841e-08, 2.423586e-08, 2.297388e-08, 
    2.334066e-08, 2.347281e-08, 2.447833e-08, 2.551389e-08, 2.510555e-08, 
    2.510131e-08, 2.553411e-08, 2.403556e-08, 2.304368e-08, 2.378237e-08,
  2.197459e-08, 2.277369e-08, 2.274703e-08, 2.38104e-08, 2.357581e-08, 
    2.276153e-08, 2.350797e-08, 2.405039e-08, 2.418394e-08, 2.493107e-08, 
    2.375835e-08, 2.339285e-08, 2.325334e-08, 2.316458e-08, 2.619704e-08,
  2.230883e-08, 2.293873e-08, 2.318519e-08, 2.358925e-08, 2.376684e-08, 
    2.241882e-08, 2.294455e-08, 2.374999e-08, 2.367799e-08, 2.360446e-08, 
    2.354764e-08, 2.365234e-08, 2.310535e-08, 2.364368e-08, 2.619954e-08,
  2.207029e-08, 2.281155e-08, 2.300365e-08, 2.371544e-08, 2.430342e-08, 
    2.248861e-08, 2.224465e-08, 2.273492e-08, 2.310349e-08, 2.378213e-08, 
    2.376965e-08, 2.3616e-08, 2.307516e-08, 2.448601e-08, 2.437968e-08,
  2.222982e-08, 2.290889e-08, 2.31591e-08, 2.375927e-08, 2.503645e-08, 
    2.32984e-08, 2.297065e-08, 2.300902e-08, 2.328787e-08, 2.34306e-08, 
    2.366028e-08, 2.365273e-08, 2.344152e-08, 2.374914e-08, 2.360887e-08,
  2.223233e-08, 2.321513e-08, 2.308007e-08, 2.358176e-08, 2.531793e-08, 
    2.327369e-08, 2.225893e-08, 2.313379e-08, 2.271358e-08, 2.341488e-08, 
    2.362815e-08, 2.383426e-08, 2.398623e-08, 2.349004e-08, 2.359705e-08,
  2.503569e-08, 2.518483e-08, 2.504384e-08, 2.409644e-08, 2.403934e-08, 
    2.427e-08, 2.347053e-08, 2.205341e-08, 2.230968e-08, 2.289019e-08, 
    2.24482e-08, 2.194568e-08, 2.371422e-08, 2.582188e-08, 2.581141e-08,
  2.476016e-08, 2.475258e-08, 2.498768e-08, 2.470789e-08, 2.326866e-08, 
    2.295198e-08, 2.354389e-08, 2.259543e-08, 2.221575e-08, 2.240147e-08, 
    2.186762e-08, 2.195016e-08, 2.442935e-08, 2.516593e-08, 2.441792e-08,
  2.371712e-08, 2.506812e-08, 2.53362e-08, 2.489468e-08, 2.380475e-08, 
    2.295731e-08, 2.337387e-08, 2.280731e-08, 2.206989e-08, 2.2213e-08, 
    2.200315e-08, 2.178138e-08, 2.355129e-08, 2.345784e-08, 2.301098e-08,
  2.320749e-08, 2.51189e-08, 2.499896e-08, 2.571286e-08, 2.525821e-08, 
    2.299587e-08, 2.281235e-08, 2.302717e-08, 2.248073e-08, 2.267399e-08, 
    2.395564e-08, 2.230252e-08, 2.330463e-08, 2.240512e-08, 2.522576e-08,
  2.366675e-08, 2.484668e-08, 2.473007e-08, 2.576539e-08, 2.55832e-08, 
    2.321245e-08, 2.236888e-08, 2.250457e-08, 2.361178e-08, 2.401493e-08, 
    2.258694e-08, 2.341241e-08, 2.322326e-08, 2.300653e-08, 2.608782e-08,
  2.419388e-08, 2.520447e-08, 2.477439e-08, 2.577269e-08, 2.603319e-08, 
    2.364138e-08, 2.171309e-08, 2.177067e-08, 2.176557e-08, 2.275328e-08, 
    2.160571e-08, 2.18721e-08, 2.403543e-08, 2.275519e-08, 2.414178e-08,
  2.482022e-08, 2.541991e-08, 2.476635e-08, 2.580853e-08, 2.62168e-08, 
    2.401476e-08, 2.246773e-08, 2.163568e-08, 2.137593e-08, 2.217909e-08, 
    2.248433e-08, 2.189906e-08, 2.097576e-08, 2.095921e-08, 2.248583e-08,
  2.462886e-08, 2.544925e-08, 2.482049e-08, 2.577807e-08, 2.609893e-08, 
    2.384672e-08, 2.219834e-08, 2.066143e-08, 2.019122e-08, 2.274832e-08, 
    2.378214e-08, 2.218539e-08, 2.048193e-08, 2.376502e-08, 2.294889e-08,
  2.501998e-08, 2.5692e-08, 2.488139e-08, 2.561045e-08, 2.606219e-08, 
    2.440607e-08, 2.3345e-08, 2.150547e-08, 2.100156e-08, 2.203281e-08, 
    2.326222e-08, 2.288266e-08, 2.186465e-08, 2.300552e-08, 2.237379e-08,
  2.492495e-08, 2.568799e-08, 2.516644e-08, 2.512038e-08, 2.543661e-08, 
    2.407206e-08, 2.260216e-08, 2.115577e-08, 2.059456e-08, 2.165722e-08, 
    2.286241e-08, 2.317678e-08, 2.201748e-08, 2.213792e-08, 2.212455e-08,
  2.350763e-08, 2.605253e-08, 2.694063e-08, 2.614952e-08, 2.586841e-08, 
    2.545019e-08, 2.560799e-08, 2.434617e-08, 2.284768e-08, 2.294535e-08, 
    2.349582e-08, 2.222736e-08, 2.250628e-08, 2.270673e-08, 2.106128e-08,
  2.288889e-08, 2.533226e-08, 2.662776e-08, 2.677171e-08, 2.633859e-08, 
    2.596471e-08, 2.616912e-08, 2.54477e-08, 2.431867e-08, 2.343827e-08, 
    2.359443e-08, 2.279093e-08, 2.299708e-08, 2.287539e-08, 2.17605e-08,
  2.487907e-08, 2.4809e-08, 2.606876e-08, 2.656019e-08, 2.680204e-08, 
    2.598437e-08, 2.601272e-08, 2.576472e-08, 2.476396e-08, 2.377025e-08, 
    2.345056e-08, 2.268517e-08, 2.306534e-08, 2.276876e-08, 2.20095e-08,
  2.473365e-08, 2.559434e-08, 2.671863e-08, 2.714459e-08, 2.685488e-08, 
    2.594632e-08, 2.610402e-08, 2.593601e-08, 2.534466e-08, 2.415547e-08, 
    2.457278e-08, 2.336169e-08, 2.257018e-08, 2.214619e-08, 2.305051e-08,
  2.530023e-08, 2.527902e-08, 2.666552e-08, 2.732232e-08, 2.689458e-08, 
    2.637436e-08, 2.641494e-08, 2.630984e-08, 2.586461e-08, 2.511329e-08, 
    2.420642e-08, 2.258477e-08, 2.118011e-08, 2.109649e-08, 2.296202e-08,
  2.333211e-08, 2.499255e-08, 2.601513e-08, 2.726198e-08, 2.745461e-08, 
    2.680207e-08, 2.67413e-08, 2.689412e-08, 2.575203e-08, 2.504104e-08, 
    2.444698e-08, 2.26063e-08, 2.181715e-08, 2.08797e-08, 2.238728e-08,
  2.263333e-08, 2.49097e-08, 2.629201e-08, 2.699137e-08, 2.734615e-08, 
    2.706392e-08, 2.685087e-08, 2.652079e-08, 2.543548e-08, 2.489445e-08, 
    2.442956e-08, 2.401229e-08, 2.250643e-08, 2.100562e-08, 2.20363e-08,
  2.219492e-08, 2.548663e-08, 2.650722e-08, 2.698398e-08, 2.766312e-08, 
    2.753666e-08, 2.699784e-08, 2.631472e-08, 2.574735e-08, 2.508707e-08, 
    2.496682e-08, 2.474754e-08, 2.327344e-08, 2.229374e-08, 2.171256e-08,
  2.298312e-08, 2.631969e-08, 2.676901e-08, 2.693046e-08, 2.816589e-08, 
    2.813834e-08, 2.735679e-08, 2.673413e-08, 2.590087e-08, 2.545698e-08, 
    2.526363e-08, 2.472539e-08, 2.380121e-08, 2.298609e-08, 2.149738e-08,
  2.343257e-08, 2.643805e-08, 2.652824e-08, 2.634668e-08, 2.692924e-08, 
    2.699543e-08, 2.680986e-08, 2.630374e-08, 2.624962e-08, 2.584206e-08, 
    2.536712e-08, 2.47531e-08, 2.436284e-08, 2.301575e-08, 2.199753e-08,
  1.722684e-08, 1.932625e-08, 2.11727e-08, 2.285356e-08, 2.33839e-08, 
    2.447405e-08, 2.518791e-08, 2.625668e-08, 2.802604e-08, 2.864617e-08, 
    2.79332e-08, 2.557341e-08, 2.848569e-08, 2.52697e-08, 2.386077e-08,
  1.728091e-08, 1.935739e-08, 2.135098e-08, 2.343067e-08, 2.451996e-08, 
    2.459567e-08, 2.480253e-08, 2.696946e-08, 2.862005e-08, 2.801273e-08, 
    2.732785e-08, 2.575054e-08, 2.957275e-08, 2.488527e-08, 2.268339e-08,
  1.758068e-08, 1.880784e-08, 2.115944e-08, 2.328743e-08, 2.42828e-08, 
    2.361629e-08, 2.416013e-08, 2.639534e-08, 2.824191e-08, 2.882139e-08, 
    2.792473e-08, 2.579128e-08, 2.987858e-08, 2.251497e-08, 2.275587e-08,
  1.74761e-08, 1.881795e-08, 2.048302e-08, 2.22201e-08, 2.298477e-08, 
    2.33961e-08, 2.396921e-08, 2.59532e-08, 2.85746e-08, 2.757915e-08, 
    2.607276e-08, 2.635681e-08, 3.114098e-08, 2.221799e-08, 2.501459e-08,
  1.767102e-08, 1.829605e-08, 1.982465e-08, 2.131556e-08, 2.228919e-08, 
    2.332035e-08, 2.450968e-08, 2.558571e-08, 2.577031e-08, 2.27219e-08, 
    2.233547e-08, 2.846632e-08, 3.156664e-08, 2.487205e-08, 3.068405e-08,
  1.746022e-08, 1.785062e-08, 1.926074e-08, 2.07411e-08, 2.175034e-08, 
    2.266055e-08, 2.377255e-08, 2.405153e-08, 2.289063e-08, 2.301083e-08, 
    2.566868e-08, 2.788119e-08, 2.95119e-08, 3.061195e-08, 3.25123e-08,
  1.713839e-08, 1.817291e-08, 1.959686e-08, 2.072765e-08, 2.180954e-08, 
    2.257935e-08, 2.358057e-08, 2.324816e-08, 2.352644e-08, 2.561275e-08, 
    2.726525e-08, 2.738373e-08, 3.052373e-08, 3.611868e-08, 3.088622e-08,
  1.747353e-08, 1.875722e-08, 1.904347e-08, 2.035009e-08, 2.207182e-08, 
    2.300677e-08, 2.3491e-08, 2.307345e-08, 2.349663e-08, 2.591577e-08, 
    2.767382e-08, 2.789413e-08, 3.106223e-08, 3.547226e-08, 2.727951e-08,
  1.807689e-08, 1.900137e-08, 1.954652e-08, 2.047472e-08, 2.19117e-08, 
    2.237772e-08, 2.177172e-08, 2.097634e-08, 2.345548e-08, 2.764953e-08, 
    2.782824e-08, 2.799527e-08, 3.063023e-08, 3.01297e-08, 2.746181e-08,
  1.83633e-08, 1.920889e-08, 1.953926e-08, 2.022126e-08, 2.087549e-08, 
    2.104367e-08, 2.010409e-08, 2.261418e-08, 2.658502e-08, 2.775467e-08, 
    2.735395e-08, 2.780322e-08, 2.900393e-08, 2.859315e-08, 2.813895e-08,
  1.102756e-08, 1.323064e-08, 1.493489e-08, 1.626658e-08, 1.735635e-08, 
    1.776012e-08, 1.757614e-08, 1.883878e-08, 2.032417e-08, 1.994475e-08, 
    1.993832e-08, 2.144862e-08, 2.257414e-08, 1.976226e-08, 1.921282e-08,
  1.307581e-08, 1.431139e-08, 1.565277e-08, 1.698536e-08, 1.879674e-08, 
    1.896481e-08, 1.889577e-08, 1.987401e-08, 2.108358e-08, 2.099378e-08, 
    2.117051e-08, 2.33296e-08, 2.210284e-08, 2.104485e-08, 2.129584e-08,
  1.585972e-08, 1.662663e-08, 1.691359e-08, 1.907377e-08, 2.005264e-08, 
    1.963625e-08, 1.952477e-08, 2.013875e-08, 2.130421e-08, 2.198722e-08, 
    2.340166e-08, 2.521652e-08, 2.471026e-08, 2.109942e-08, 2.31964e-08,
  1.66391e-08, 1.714232e-08, 1.818559e-08, 1.914929e-08, 1.949391e-08, 
    1.94784e-08, 1.989281e-08, 2.07314e-08, 2.155118e-08, 2.13645e-08, 
    2.270642e-08, 2.46327e-08, 2.524288e-08, 2.473348e-08, 2.330288e-08,
  1.785901e-08, 1.742554e-08, 1.827577e-08, 1.919623e-08, 1.98161e-08, 
    2.030431e-08, 2.057317e-08, 2.174629e-08, 2.221097e-08, 2.118469e-08, 
    2.290941e-08, 2.478591e-08, 2.674229e-08, 2.599255e-08, 2.424698e-08,
  1.943968e-08, 1.91506e-08, 2.018087e-08, 2.071246e-08, 2.169921e-08, 
    2.144615e-08, 2.12129e-08, 2.265637e-08, 2.210724e-08, 2.140437e-08, 
    2.577855e-08, 2.498031e-08, 2.6124e-08, 2.407743e-08, 2.66529e-08,
  1.992234e-08, 2.153502e-08, 2.203968e-08, 2.20895e-08, 2.342969e-08, 
    2.345763e-08, 2.454846e-08, 2.527228e-08, 2.406176e-08, 2.559713e-08, 
    2.500731e-08, 2.309928e-08, 2.582953e-08, 2.475419e-08, 2.533552e-08,
  2.05867e-08, 2.248003e-08, 2.336933e-08, 2.467512e-08, 2.626149e-08, 
    2.68291e-08, 2.690023e-08, 2.496476e-08, 2.307443e-08, 2.36047e-08, 
    2.324636e-08, 2.426357e-08, 2.591407e-08, 2.585923e-08, 2.153614e-08,
  2.247817e-08, 2.386594e-08, 2.547141e-08, 2.731607e-08, 2.828205e-08, 
    2.744164e-08, 2.557456e-08, 2.182551e-08, 2.191921e-08, 2.256203e-08, 
    2.269824e-08, 2.336964e-08, 2.16626e-08, 1.970278e-08, 1.66423e-08,
  2.362799e-08, 2.430045e-08, 2.416087e-08, 2.397272e-08, 2.337029e-08, 
    2.272507e-08, 2.070995e-08, 1.877911e-08, 2.143237e-08, 2.235304e-08, 
    2.259771e-08, 2.325393e-08, 2.233403e-08, 1.83529e-08, 1.807876e-08,
  2.210155e-08, 2.340806e-08, 2.319175e-08, 2.336415e-08, 2.354491e-08, 
    2.38701e-08, 2.348888e-08, 2.420122e-08, 2.377906e-08, 2.492607e-08, 
    2.389839e-08, 2.51468e-08, 2.834172e-08, 2.838525e-08, 2.559545e-08,
  2.402845e-08, 2.423069e-08, 2.370144e-08, 2.443355e-08, 2.499715e-08, 
    2.560427e-08, 2.492336e-08, 2.626094e-08, 2.606669e-08, 2.691518e-08, 
    2.728742e-08, 2.730266e-08, 2.678746e-08, 2.5022e-08, 2.189944e-08,
  2.469636e-08, 2.545525e-08, 2.417985e-08, 2.420461e-08, 2.443278e-08, 
    2.423005e-08, 2.279874e-08, 2.215613e-08, 2.392165e-08, 2.352598e-08, 
    2.426269e-08, 2.355315e-08, 2.325365e-08, 1.991913e-08, 2.037424e-08,
  2.383437e-08, 2.395386e-08, 2.420389e-08, 2.348313e-08, 2.265468e-08, 
    2.251217e-08, 2.198295e-08, 2.150709e-08, 2.101951e-08, 2.077803e-08, 
    1.953577e-08, 1.90205e-08, 2.109803e-08, 2.165824e-08, 2.58789e-08,
  2.32491e-08, 2.400478e-08, 2.429896e-08, 2.267155e-08, 2.245575e-08, 
    2.291104e-08, 2.364192e-08, 2.466284e-08, 2.42208e-08, 2.10898e-08, 
    1.985167e-08, 2.307905e-08, 2.340904e-08, 2.808101e-08, 2.84579e-08,
  2.617388e-08, 2.523317e-08, 2.59668e-08, 2.490443e-08, 2.484423e-08, 
    2.499628e-08, 2.45501e-08, 2.528175e-08, 2.359396e-08, 2.215035e-08, 
    2.603858e-08, 2.757786e-08, 2.66831e-08, 3.077335e-08, 3.081681e-08,
  2.481219e-08, 2.465301e-08, 2.492758e-08, 2.454716e-08, 2.417577e-08, 
    2.438121e-08, 2.390182e-08, 2.517301e-08, 2.392802e-08, 2.488303e-08, 
    2.738736e-08, 2.646477e-08, 2.858113e-08, 3.247082e-08, 2.914697e-08,
  2.428805e-08, 2.463711e-08, 2.463551e-08, 2.465559e-08, 2.42496e-08, 
    2.477857e-08, 2.469081e-08, 2.498993e-08, 2.532663e-08, 2.646432e-08, 
    2.715687e-08, 2.741835e-08, 3.110173e-08, 3.190397e-08, 2.233143e-08,
  2.310149e-08, 2.382202e-08, 2.410538e-08, 2.446614e-08, 2.41179e-08, 
    2.485138e-08, 2.523419e-08, 2.427816e-08, 2.454135e-08, 2.701415e-08, 
    2.850386e-08, 2.926224e-08, 2.79409e-08, 2.637734e-08, 2.159613e-08,
  2.299017e-08, 2.356515e-08, 2.462288e-08, 2.407198e-08, 2.310952e-08, 
    2.312891e-08, 2.346511e-08, 2.463737e-08, 2.682155e-08, 2.822886e-08, 
    2.95159e-08, 2.949253e-08, 2.987283e-08, 2.65555e-08, 2.479538e-08,
  2.419463e-08, 2.416026e-08, 2.374894e-08, 2.39769e-08, 2.407539e-08, 
    2.447766e-08, 2.485736e-08, 2.479847e-08, 2.463955e-08, 2.325251e-08, 
    2.234177e-08, 2.151567e-08, 2.102528e-08, 2.369721e-08, 2.613726e-08,
  2.478051e-08, 2.491616e-08, 2.411376e-08, 2.412961e-08, 2.475935e-08, 
    2.51826e-08, 2.494887e-08, 2.447914e-08, 2.398738e-08, 2.380036e-08, 
    2.370359e-08, 2.279368e-08, 2.000997e-08, 2.32268e-08, 2.255751e-08,
  2.830079e-08, 2.463324e-08, 2.333729e-08, 2.423239e-08, 2.507254e-08, 
    2.526268e-08, 2.45408e-08, 2.382399e-08, 2.363322e-08, 2.3571e-08, 
    2.359636e-08, 2.317018e-08, 2.31473e-08, 2.522659e-08, 2.124661e-08,
  2.733421e-08, 2.412111e-08, 2.35894e-08, 2.420314e-08, 2.44452e-08, 
    2.480007e-08, 2.424514e-08, 2.370125e-08, 2.342805e-08, 2.368369e-08, 
    2.267425e-08, 2.258342e-08, 2.288671e-08, 2.276385e-08, 2.024931e-08,
  2.777903e-08, 2.415127e-08, 2.316485e-08, 2.421384e-08, 2.485418e-08, 
    2.477579e-08, 2.409463e-08, 2.379583e-08, 2.491842e-08, 2.403852e-08, 
    2.286748e-08, 2.214126e-08, 1.995323e-08, 2.030709e-08, 2.247818e-08,
  2.590964e-08, 2.35879e-08, 2.27989e-08, 2.409329e-08, 2.410696e-08, 
    2.395134e-08, 2.35268e-08, 2.405267e-08, 2.481352e-08, 2.311296e-08, 
    2.194136e-08, 2.266927e-08, 1.995251e-08, 1.977281e-08, 2.759253e-08,
  2.483435e-08, 2.308324e-08, 2.280885e-08, 2.372954e-08, 2.372117e-08, 
    2.357259e-08, 2.344962e-08, 2.420163e-08, 2.385725e-08, 2.210156e-08, 
    2.417133e-08, 2.473934e-08, 2.075255e-08, 2.550097e-08, 3.094048e-08,
  2.419129e-08, 2.364717e-08, 2.290085e-08, 2.355816e-08, 2.385821e-08, 
    2.405309e-08, 2.376809e-08, 2.47217e-08, 2.32722e-08, 2.298693e-08, 
    2.394571e-08, 2.365507e-08, 2.332604e-08, 2.261701e-08, 2.183661e-08,
  2.426135e-08, 2.354857e-08, 2.268585e-08, 2.333418e-08, 2.397033e-08, 
    2.424238e-08, 2.361005e-08, 2.404017e-08, 2.364893e-08, 2.371766e-08, 
    2.480733e-08, 2.479729e-08, 2.385029e-08, 2.315749e-08, 2.095618e-08,
  2.450671e-08, 2.351976e-08, 2.305219e-08, 2.359218e-08, 2.442065e-08, 
    2.463001e-08, 2.44965e-08, 2.430248e-08, 2.485674e-08, 2.51581e-08, 
    2.497839e-08, 2.436467e-08, 2.512387e-08, 2.476951e-08, 2.484027e-08,
  2.498241e-08, 2.590573e-08, 2.643331e-08, 2.354556e-08, 2.26202e-08, 
    2.224342e-08, 2.213494e-08, 2.246948e-08, 2.406937e-08, 2.429111e-08, 
    2.258544e-08, 2.103916e-08, 2.007503e-08, 2.160071e-08, 2.256445e-08,
  2.408068e-08, 2.52196e-08, 2.641093e-08, 2.419765e-08, 2.350241e-08, 
    2.284549e-08, 2.227475e-08, 2.280712e-08, 2.380657e-08, 2.300528e-08, 
    2.142942e-08, 2.046105e-08, 2.028688e-08, 2.244932e-08, 2.236993e-08,
  2.565472e-08, 2.440975e-08, 2.592055e-08, 2.391758e-08, 2.387543e-08, 
    2.342779e-08, 2.29039e-08, 2.346644e-08, 2.354635e-08, 2.202625e-08, 
    2.134798e-08, 2.065653e-08, 2.045567e-08, 2.119467e-08, 2.027319e-08,
  2.71103e-08, 2.587049e-08, 2.510047e-08, 2.521528e-08, 2.498506e-08, 
    2.39086e-08, 2.408181e-08, 2.525274e-08, 2.488446e-08, 2.162403e-08, 
    2.299468e-08, 2.407737e-08, 2.005698e-08, 2.156955e-08, 2.435754e-08,
  2.886096e-08, 2.773073e-08, 2.821508e-08, 2.637013e-08, 2.591666e-08, 
    2.609724e-08, 2.558262e-08, 2.60493e-08, 2.671694e-08, 2.138647e-08, 
    2.087658e-08, 2.522926e-08, 2.293227e-08, 2.491048e-08, 3.149144e-08,
  2.605415e-08, 2.609743e-08, 2.60419e-08, 2.689121e-08, 2.593728e-08, 
    2.55996e-08, 2.642992e-08, 2.960514e-08, 2.568531e-08, 1.854307e-08, 
    2.078095e-08, 2.475025e-08, 2.518133e-08, 2.402784e-08, 3.261181e-08,
  2.60276e-08, 2.633486e-08, 2.644208e-08, 2.618043e-08, 2.589953e-08, 
    2.521105e-08, 2.538079e-08, 2.777091e-08, 2.349881e-08, 1.991883e-08, 
    2.374919e-08, 2.449671e-08, 2.482901e-08, 2.334387e-08, 2.672009e-08,
  2.504976e-08, 2.578361e-08, 2.624961e-08, 2.614127e-08, 2.573044e-08, 
    2.565804e-08, 2.585809e-08, 2.698274e-08, 2.550854e-08, 2.369132e-08, 
    2.368774e-08, 2.367518e-08, 2.440741e-08, 2.783474e-08, 2.617179e-08,
  2.523954e-08, 2.631631e-08, 2.645121e-08, 2.695786e-08, 2.801747e-08, 
    2.775279e-08, 2.833138e-08, 2.635633e-08, 2.483969e-08, 2.523974e-08, 
    2.416992e-08, 2.320187e-08, 2.411128e-08, 2.628557e-08, 2.668357e-08,
  2.466722e-08, 2.597312e-08, 2.646408e-08, 2.709814e-08, 2.900181e-08, 
    2.864103e-08, 2.608687e-08, 2.524551e-08, 2.551096e-08, 2.763659e-08, 
    2.487301e-08, 2.250017e-08, 2.328941e-08, 2.532679e-08, 2.544743e-08,
  2.779183e-08, 3.081734e-08, 3.0753e-08, 2.653799e-08, 2.719392e-08, 
    2.441066e-08, 2.171793e-08, 1.72941e-08, 1.811674e-08, 2.258713e-08, 
    2.26494e-08, 2.079057e-08, 1.962176e-08, 1.899204e-08, 2.045627e-08,
  2.670938e-08, 3.159784e-08, 3.257637e-08, 2.790036e-08, 2.753185e-08, 
    2.742168e-08, 2.350333e-08, 1.94603e-08, 1.999219e-08, 2.29162e-08, 
    2.234237e-08, 2.079938e-08, 1.900296e-08, 1.778924e-08, 1.9304e-08,
  2.990067e-08, 3.14169e-08, 3.321841e-08, 2.991491e-08, 2.954792e-08, 
    2.905166e-08, 2.62414e-08, 2.454347e-08, 2.070279e-08, 2.354829e-08, 
    2.395862e-08, 2.28755e-08, 2.031468e-08, 1.655273e-08, 1.551519e-08,
  2.666192e-08, 2.975287e-08, 3.357554e-08, 3.438011e-08, 3.240589e-08, 
    2.938337e-08, 2.831903e-08, 2.659627e-08, 2.313779e-08, 2.568337e-08, 
    2.645517e-08, 2.480776e-08, 2.61846e-08, 2.092781e-08, 1.579192e-08,
  2.596195e-08, 2.766756e-08, 3.303729e-08, 3.64749e-08, 3.287998e-08, 
    3.257935e-08, 2.979239e-08, 2.845055e-08, 3.089128e-08, 2.70906e-08, 
    2.262526e-08, 2.837955e-08, 2.832081e-08, 1.959452e-08, 1.681861e-08,
  2.303615e-08, 2.501607e-08, 2.707842e-08, 3.299142e-08, 3.502439e-08, 
    3.120581e-08, 3.047742e-08, 3.155403e-08, 2.624404e-08, 2.350334e-08, 
    2.276154e-08, 2.667228e-08, 2.55115e-08, 1.897049e-08, 2.214973e-08,
  2.289497e-08, 2.486822e-08, 2.711825e-08, 2.956137e-08, 3.230721e-08, 
    3.14227e-08, 2.917183e-08, 2.653855e-08, 2.43377e-08, 2.404702e-08, 
    2.30319e-08, 2.388948e-08, 2.246873e-08, 2.364981e-08, 2.943865e-08,
  2.183906e-08, 2.368209e-08, 2.531502e-08, 2.77428e-08, 3.085735e-08, 
    3.106773e-08, 3.045875e-08, 2.958851e-08, 2.706174e-08, 2.465018e-08, 
    2.60646e-08, 2.394278e-08, 2.258746e-08, 3.013843e-08, 2.863305e-08,
  2.193215e-08, 2.390985e-08, 2.553233e-08, 2.697208e-08, 3.116568e-08, 
    3.308811e-08, 3.172863e-08, 2.769276e-08, 2.728448e-08, 2.615155e-08, 
    2.770829e-08, 2.587309e-08, 2.422339e-08, 2.344364e-08, 2.685853e-08,
  2.180433e-08, 2.306388e-08, 2.420846e-08, 2.618902e-08, 3.011821e-08, 
    3.500513e-08, 3.077286e-08, 2.73734e-08, 2.686848e-08, 2.787012e-08, 
    2.97272e-08, 2.804476e-08, 2.730895e-08, 2.924725e-08, 2.667472e-08,
  1.930523e-08, 2.053131e-08, 2.428677e-08, 2.518497e-08, 2.84223e-08, 
    3.19771e-08, 2.782143e-08, 2.29051e-08, 2.363302e-08, 2.531714e-08, 
    2.427658e-08, 2.09503e-08, 1.897937e-08, 1.84522e-08, 1.754063e-08,
  1.929316e-08, 2.049833e-08, 2.333264e-08, 2.533935e-08, 2.844272e-08, 
    3.257919e-08, 2.716392e-08, 2.475449e-08, 2.482015e-08, 2.532188e-08, 
    2.236394e-08, 2.050263e-08, 1.918562e-08, 1.783001e-08, 1.874324e-08,
  2.069565e-08, 2.000561e-08, 2.313817e-08, 2.678203e-08, 2.892648e-08, 
    3.191938e-08, 2.703779e-08, 2.556439e-08, 2.174879e-08, 2.445204e-08, 
    2.298393e-08, 2.198297e-08, 2.138639e-08, 1.944641e-08, 1.795632e-08,
  1.96004e-08, 2.064549e-08, 2.237605e-08, 2.651767e-08, 2.960099e-08, 
    3.356749e-08, 2.865766e-08, 2.44406e-08, 2.532373e-08, 2.711258e-08, 
    2.617525e-08, 2.219981e-08, 2.314345e-08, 2.059027e-08, 1.694087e-08,
  1.946155e-08, 2.078774e-08, 2.22333e-08, 2.526018e-08, 3.058458e-08, 
    3.590054e-08, 3.414573e-08, 2.821697e-08, 3.544099e-08, 2.595282e-08, 
    1.898224e-08, 2.754565e-08, 2.757115e-08, 2.016726e-08, 1.984851e-08,
  1.995779e-08, 2.106384e-08, 2.087747e-08, 2.227147e-08, 2.900099e-08, 
    3.73907e-08, 3.669936e-08, 3.179241e-08, 2.635531e-08, 2.391238e-08, 
    2.210783e-08, 2.637878e-08, 2.508862e-08, 2.179959e-08, 2.388028e-08,
  2.090558e-08, 2.114533e-08, 2.115228e-08, 2.149319e-08, 2.541195e-08, 
    3.608488e-08, 3.661519e-08, 2.654648e-08, 2.393726e-08, 2.569496e-08, 
    2.312667e-08, 2.440216e-08, 2.276733e-08, 2.483062e-08, 2.609749e-08,
  2.072134e-08, 2.143055e-08, 2.09777e-08, 2.095152e-08, 2.39388e-08, 
    3.241192e-08, 3.834661e-08, 3.198452e-08, 2.582672e-08, 2.741912e-08, 
    2.76489e-08, 2.450443e-08, 2.533764e-08, 3.074146e-08, 2.561139e-08,
  2.169961e-08, 2.206072e-08, 2.140372e-08, 2.141058e-08, 2.351762e-08, 
    2.884232e-08, 3.565617e-08, 2.866395e-08, 2.623915e-08, 2.648522e-08, 
    2.909787e-08, 2.729816e-08, 2.567032e-08, 2.923987e-08, 2.730911e-08,
  2.201357e-08, 2.162704e-08, 2.092133e-08, 2.119315e-08, 2.337244e-08, 
    2.661951e-08, 3.329181e-08, 2.89057e-08, 2.582724e-08, 2.260595e-08, 
    2.794979e-08, 2.838603e-08, 2.841709e-08, 2.801728e-08, 2.829153e-08,
  2.133868e-08, 2.123536e-08, 2.13406e-08, 2.14003e-08, 2.143262e-08, 
    2.168516e-08, 2.363939e-08, 2.469749e-08, 2.698452e-08, 2.625405e-08, 
    2.533163e-08, 2.359292e-08, 2.298123e-08, 2.133494e-08, 2.121288e-08,
  1.876916e-08, 1.984313e-08, 2.007802e-08, 2.072476e-08, 2.150556e-08, 
    2.192791e-08, 2.396612e-08, 2.574639e-08, 2.813958e-08, 2.733649e-08, 
    2.466824e-08, 2.322034e-08, 2.175672e-08, 2.059373e-08, 2.03387e-08,
  1.791918e-08, 2.071184e-08, 2.196792e-08, 2.166555e-08, 2.163561e-08, 
    2.168721e-08, 2.390644e-08, 2.560778e-08, 2.710152e-08, 2.521428e-08, 
    2.635299e-08, 2.439873e-08, 2.205593e-08, 2.27496e-08, 2.090157e-08,
  1.833914e-08, 2.006639e-08, 2.019427e-08, 2.049051e-08, 2.023962e-08, 
    2.085415e-08, 2.419181e-08, 2.60561e-08, 2.659495e-08, 2.726099e-08, 
    2.969148e-08, 2.042366e-08, 2.309988e-08, 2.520759e-08, 2.053286e-08,
  1.805285e-08, 1.920091e-08, 2.004134e-08, 1.983098e-08, 2.056673e-08, 
    2.121917e-08, 2.583267e-08, 2.795147e-08, 2.731251e-08, 2.591389e-08, 
    1.886385e-08, 2.025189e-08, 3.271064e-08, 2.351446e-08, 2.377249e-08,
  1.975359e-08, 1.987656e-08, 2.003794e-08, 2.035365e-08, 2.074859e-08, 
    2.199558e-08, 2.491e-08, 2.793388e-08, 2.502568e-08, 2.110127e-08, 
    2.047625e-08, 2.331396e-08, 2.743239e-08, 2.287256e-08, 2.871998e-08,
  2.12483e-08, 2.054759e-08, 2.044854e-08, 2.083731e-08, 2.159416e-08, 
    2.227277e-08, 2.316856e-08, 2.62618e-08, 2.55936e-08, 2.495252e-08, 
    2.348828e-08, 2.33489e-08, 2.313739e-08, 2.544157e-08, 2.696657e-08,
  2.135303e-08, 2.130183e-08, 2.153759e-08, 2.231605e-08, 2.189412e-08, 
    2.148843e-08, 2.27392e-08, 2.592385e-08, 2.614769e-08, 2.57915e-08, 
    2.514049e-08, 2.531939e-08, 2.452367e-08, 3.244356e-08, 2.569453e-08,
  2.191461e-08, 2.25487e-08, 2.24647e-08, 2.331685e-08, 2.182691e-08, 
    2.120293e-08, 2.262082e-08, 2.595045e-08, 2.86742e-08, 3.048552e-08, 
    2.708411e-08, 2.633158e-08, 2.543684e-08, 2.777927e-08, 2.403895e-08,
  2.314874e-08, 2.296656e-08, 2.262494e-08, 2.315827e-08, 2.227472e-08, 
    2.327933e-08, 2.544476e-08, 2.737254e-08, 3.125874e-08, 3.178701e-08, 
    2.814656e-08, 2.595655e-08, 2.672612e-08, 2.613536e-08, 2.515011e-08,
  1.922588e-08, 1.95865e-08, 1.933327e-08, 2.00608e-08, 2.030268e-08, 
    2.006703e-08, 2.031772e-08, 2.01262e-08, 2.12804e-08, 2.087683e-08, 
    2.061116e-08, 2.193063e-08, 2.352227e-08, 2.39704e-08, 2.327574e-08,
  1.8086e-08, 1.872128e-08, 1.827519e-08, 1.778928e-08, 1.817541e-08, 
    1.862992e-08, 1.919991e-08, 1.927493e-08, 2.062571e-08, 2.043337e-08, 
    2.101547e-08, 2.334026e-08, 2.429837e-08, 2.355004e-08, 2.303504e-08,
  1.70167e-08, 1.855181e-08, 1.909435e-08, 1.814623e-08, 1.811931e-08, 
    1.906475e-08, 1.935569e-08, 1.945243e-08, 2.045708e-08, 2.050498e-08, 
    2.19243e-08, 2.555431e-08, 2.566888e-08, 2.526041e-08, 2.455559e-08,
  1.909955e-08, 1.99709e-08, 1.911864e-08, 2.012988e-08, 2.033543e-08, 
    2.032187e-08, 2.013601e-08, 1.982466e-08, 2.041286e-08, 2.005657e-08, 
    2.282754e-08, 2.476248e-08, 2.421627e-08, 2.464246e-08, 2.485647e-08,
  2.030977e-08, 2.046109e-08, 2.004523e-08, 1.928853e-08, 1.915693e-08, 
    1.914364e-08, 1.917338e-08, 1.962363e-08, 1.988893e-08, 2.005016e-08, 
    2.105313e-08, 2.166992e-08, 2.428875e-08, 2.745714e-08, 2.68771e-08,
  2.247992e-08, 2.186617e-08, 2.178255e-08, 2.066625e-08, 1.96527e-08, 
    1.951168e-08, 1.977618e-08, 2.006873e-08, 2.036206e-08, 2.123615e-08, 
    2.394811e-08, 2.408487e-08, 2.769766e-08, 2.847264e-08, 2.567976e-08,
  2.393761e-08, 2.267444e-08, 2.172085e-08, 2.029104e-08, 1.965379e-08, 
    1.979943e-08, 2.023926e-08, 2.059821e-08, 2.127005e-08, 2.348212e-08, 
    2.572382e-08, 2.558176e-08, 2.908446e-08, 2.631345e-08, 2.38782e-08,
  2.261764e-08, 2.195299e-08, 2.147345e-08, 2.068136e-08, 1.97547e-08, 
    2.006962e-08, 2.09523e-08, 2.148206e-08, 2.257537e-08, 2.413533e-08, 
    2.596948e-08, 2.725352e-08, 2.800018e-08, 2.655376e-08, 2.750186e-08,
  2.29847e-08, 2.279804e-08, 2.150009e-08, 2.097686e-08, 2.075787e-08, 
    2.170474e-08, 2.18453e-08, 2.257601e-08, 2.282676e-08, 2.584804e-08, 
    2.828282e-08, 2.811938e-08, 2.61686e-08, 2.971574e-08, 2.665222e-08,
  2.221715e-08, 2.221866e-08, 2.207959e-08, 2.332764e-08, 2.419175e-08, 
    2.392032e-08, 2.395952e-08, 2.433876e-08, 2.407044e-08, 2.760162e-08, 
    2.867936e-08, 2.661289e-08, 2.582784e-08, 2.623333e-08, 2.519293e-08,
  2.226687e-08, 2.131609e-08, 2.065535e-08, 2.123975e-08, 2.139547e-08, 
    2.135431e-08, 2.180127e-08, 2.17705e-08, 2.16173e-08, 2.203364e-08, 
    2.135963e-08, 2.098435e-08, 2.054874e-08, 2.085469e-08, 1.971343e-08,
  2.149608e-08, 1.98813e-08, 1.984598e-08, 1.945203e-08, 1.936074e-08, 
    1.969742e-08, 2.020601e-08, 2.063938e-08, 2.060487e-08, 2.051256e-08, 
    2.027375e-08, 1.982563e-08, 1.954714e-08, 1.984981e-08, 1.946879e-08,
  2.160423e-08, 2.015287e-08, 2.0154e-08, 1.966672e-08, 1.915347e-08, 
    1.916407e-08, 1.91612e-08, 1.891249e-08, 1.935019e-08, 1.926811e-08, 
    1.938623e-08, 1.939758e-08, 2.001015e-08, 2.026306e-08, 2.112388e-08,
  2.324549e-08, 2.160164e-08, 1.986401e-08, 2.029839e-08, 2.036982e-08, 
    2.042329e-08, 1.974407e-08, 1.993921e-08, 1.977612e-08, 2.018815e-08, 
    2.006104e-08, 1.982945e-08, 1.979447e-08, 2.001424e-08, 2.321649e-08,
  2.537763e-08, 2.33469e-08, 2.328228e-08, 2.186359e-08, 2.091138e-08, 
    2.064762e-08, 2.000848e-08, 2.011072e-08, 2.080287e-08, 2.223734e-08, 
    2.119913e-08, 2.077618e-08, 1.999348e-08, 2.316941e-08, 2.62493e-08,
  2.821865e-08, 2.457753e-08, 2.325376e-08, 2.312137e-08, 2.205216e-08, 
    2.139295e-08, 2.153443e-08, 2.130751e-08, 2.115076e-08, 2.10361e-08, 
    2.021867e-08, 2.047908e-08, 2.22179e-08, 2.710619e-08, 2.544166e-08,
  2.872154e-08, 2.505111e-08, 2.36021e-08, 2.332641e-08, 2.225556e-08, 
    2.163741e-08, 2.127697e-08, 2.112617e-08, 2.136359e-08, 2.029797e-08, 
    2.086239e-08, 2.10294e-08, 2.462956e-08, 2.476671e-08, 2.29325e-08,
  2.918016e-08, 2.550333e-08, 2.33915e-08, 2.364757e-08, 2.293224e-08, 
    2.17823e-08, 2.094925e-08, 1.967451e-08, 2.015833e-08, 2.102587e-08, 
    2.112615e-08, 2.179333e-08, 2.5783e-08, 2.263072e-08, 2.530431e-08,
  3.14098e-08, 2.756747e-08, 2.477051e-08, 2.395788e-08, 2.35213e-08, 
    2.287043e-08, 2.080055e-08, 2.090339e-08, 2.139123e-08, 2.106551e-08, 
    2.104965e-08, 2.377812e-08, 2.521022e-08, 2.650457e-08, 2.333028e-08,
  3.256988e-08, 2.921838e-08, 2.612924e-08, 2.511461e-08, 2.590512e-08, 
    2.685678e-08, 2.487657e-08, 2.346859e-08, 2.117802e-08, 2.128965e-08, 
    2.294571e-08, 2.589846e-08, 2.548466e-08, 2.516041e-08, 2.268093e-08,
  2.913314e-08, 2.873087e-08, 2.824698e-08, 2.767961e-08, 2.715496e-08, 
    2.654038e-08, 2.644183e-08, 2.48159e-08, 2.28548e-08, 2.186685e-08, 
    2.259683e-08, 2.170619e-08, 2.086434e-08, 2.046547e-08, 1.931756e-08,
  2.917465e-08, 2.911448e-08, 2.875043e-08, 2.846752e-08, 2.837827e-08, 
    2.79003e-08, 2.702312e-08, 2.599467e-08, 2.397549e-08, 2.209921e-08, 
    2.222141e-08, 2.119436e-08, 2.008576e-08, 1.948712e-08, 1.895523e-08,
  3.091589e-08, 2.907117e-08, 2.903416e-08, 2.899023e-08, 2.948323e-08, 
    2.889023e-08, 2.697422e-08, 2.535121e-08, 2.357026e-08, 2.29582e-08, 
    2.360438e-08, 2.051441e-08, 2.00543e-08, 1.925396e-08, 1.98005e-08,
  3.146103e-08, 2.9674e-08, 2.953673e-08, 3.092101e-08, 3.157816e-08, 
    3.042757e-08, 2.774248e-08, 2.598212e-08, 2.532186e-08, 2.535494e-08, 
    2.563716e-08, 2.137411e-08, 2.171862e-08, 1.97252e-08, 2.092446e-08,
  3.146066e-08, 3.070364e-08, 3.147677e-08, 3.304563e-08, 3.249497e-08, 
    3.177859e-08, 2.999796e-08, 2.751615e-08, 2.59615e-08, 2.372023e-08, 
    2.102483e-08, 2.238504e-08, 2.565869e-08, 2.22419e-08, 2.436164e-08,
  2.981577e-08, 3.091741e-08, 3.1664e-08, 3.340697e-08, 3.334578e-08, 
    3.14712e-08, 2.968749e-08, 2.756438e-08, 2.395335e-08, 2.133062e-08, 
    2.217114e-08, 2.324088e-08, 2.631968e-08, 2.485144e-08, 2.622487e-08,
  3.109371e-08, 3.373673e-08, 3.415895e-08, 3.368642e-08, 3.375651e-08, 
    3.204163e-08, 2.957025e-08, 2.736509e-08, 2.400398e-08, 2.28253e-08, 
    2.42688e-08, 2.365679e-08, 2.654239e-08, 2.7111e-08, 2.654353e-08,
  3.171048e-08, 3.376206e-08, 3.272746e-08, 3.231897e-08, 3.385093e-08, 
    3.325645e-08, 3.07529e-08, 2.781061e-08, 2.433733e-08, 2.372642e-08, 
    2.396758e-08, 2.444999e-08, 2.752035e-08, 3.001491e-08, 2.664348e-08,
  2.871162e-08, 3.013005e-08, 3.168888e-08, 3.264318e-08, 3.335805e-08, 
    3.271721e-08, 2.960059e-08, 2.604992e-08, 2.428292e-08, 2.545428e-08, 
    2.481375e-08, 2.531897e-08, 2.759869e-08, 3.075041e-08, 2.775039e-08,
  2.234829e-08, 2.488425e-08, 2.676319e-08, 2.646583e-08, 2.667479e-08, 
    2.582189e-08, 2.405475e-08, 2.323299e-08, 2.462975e-08, 2.527392e-08, 
    2.552202e-08, 2.64369e-08, 2.873896e-08, 3.032915e-08, 2.928075e-08,
  1.865556e-08, 1.873793e-08, 1.909109e-08, 1.97832e-08, 2.163291e-08, 
    2.418689e-08, 2.676448e-08, 2.774136e-08, 2.848848e-08, 2.934067e-08, 
    2.853552e-08, 2.810576e-08, 3.05391e-08, 2.542052e-08, 1.94835e-08,
  1.793635e-08, 1.777121e-08, 1.912378e-08, 1.998987e-08, 2.167132e-08, 
    2.392495e-08, 2.655083e-08, 2.776738e-08, 2.88927e-08, 2.859749e-08, 
    2.872883e-08, 2.834692e-08, 3.054104e-08, 2.300384e-08, 1.992875e-08,
  1.780506e-08, 1.799898e-08, 1.941843e-08, 2.061165e-08, 2.228434e-08, 
    2.502958e-08, 2.723415e-08, 2.840415e-08, 2.914546e-08, 2.789383e-08, 
    2.914821e-08, 2.862736e-08, 2.963146e-08, 2.026264e-08, 2.267788e-08,
  1.83479e-08, 1.872362e-08, 1.989118e-08, 2.140449e-08, 2.351878e-08, 
    2.465062e-08, 2.620218e-08, 2.763401e-08, 2.843148e-08, 2.655963e-08, 
    2.811045e-08, 2.673498e-08, 2.786508e-08, 2.047385e-08, 2.536908e-08,
  1.891303e-08, 1.946591e-08, 2.123201e-08, 2.239969e-08, 2.383e-08, 
    2.440074e-08, 2.476303e-08, 2.511377e-08, 2.63824e-08, 2.601549e-08, 
    2.484156e-08, 2.439943e-08, 2.664668e-08, 2.373823e-08, 2.820914e-08,
  2.001197e-08, 2.0081e-08, 2.121655e-08, 2.214668e-08, 2.195429e-08, 
    2.260875e-08, 2.196846e-08, 2.204293e-08, 2.41656e-08, 2.386978e-08, 
    2.37463e-08, 2.237898e-08, 2.422257e-08, 2.636635e-08, 2.684366e-08,
  2.04258e-08, 2.049101e-08, 2.027553e-08, 2.012093e-08, 1.959019e-08, 
    2.038845e-08, 1.982518e-08, 2.018747e-08, 2.202784e-08, 2.214483e-08, 
    2.233137e-08, 2.133556e-08, 2.383787e-08, 2.618435e-08, 2.334428e-08,
  1.967992e-08, 2.123576e-08, 1.869448e-08, 1.831551e-08, 1.896566e-08, 
    1.827747e-08, 1.756078e-08, 1.733031e-08, 1.833999e-08, 1.991535e-08, 
    2.184658e-08, 2.234647e-08, 2.430547e-08, 2.376578e-08, 2.150416e-08,
  2.104008e-08, 2.15991e-08, 2.043218e-08, 2.019454e-08, 1.976155e-08, 
    1.942369e-08, 1.745939e-08, 1.727418e-08, 1.874592e-08, 2.165776e-08, 
    2.275252e-08, 2.30081e-08, 2.368112e-08, 2.302292e-08, 2.168933e-08,
  2.321361e-08, 2.483514e-08, 2.488315e-08, 2.31962e-08, 2.119299e-08, 
    1.942791e-08, 1.872779e-08, 2.070196e-08, 2.209587e-08, 2.402851e-08, 
    2.387022e-08, 2.406701e-08, 2.450717e-08, 2.278941e-08, 2.305261e-08,
  1.481155e-08, 1.590013e-08, 1.686577e-08, 1.815735e-08, 1.908974e-08, 
    1.963932e-08, 1.886174e-08, 1.938083e-08, 1.938591e-08, 2.152312e-08, 
    2.312113e-08, 2.287026e-08, 2.282926e-08, 2.136577e-08, 1.913123e-08,
  1.536958e-08, 1.644367e-08, 1.742241e-08, 1.831908e-08, 1.928274e-08, 
    1.894061e-08, 1.838173e-08, 1.849259e-08, 1.883752e-08, 2.169739e-08, 
    2.331576e-08, 2.26665e-08, 2.288274e-08, 2.070256e-08, 1.903722e-08,
  1.557454e-08, 1.767361e-08, 1.852312e-08, 1.876215e-08, 1.938914e-08, 
    1.914788e-08, 1.875979e-08, 1.833436e-08, 1.911883e-08, 2.265174e-08, 
    2.37479e-08, 2.262944e-08, 2.257816e-08, 2.000946e-08, 2.066772e-08,
  1.67647e-08, 1.769889e-08, 1.848415e-08, 1.969553e-08, 2.061491e-08, 
    1.944633e-08, 1.87323e-08, 1.863331e-08, 2.039373e-08, 2.402725e-08, 
    2.297651e-08, 2.203884e-08, 2.209829e-08, 1.999405e-08, 2.260235e-08,
  1.647301e-08, 1.742402e-08, 1.951105e-08, 1.84617e-08, 1.920584e-08, 
    1.899445e-08, 1.889265e-08, 1.989597e-08, 2.359283e-08, 2.497754e-08, 
    2.29808e-08, 2.28794e-08, 2.051049e-08, 1.91554e-08, 2.226896e-08,
  1.726515e-08, 1.744743e-08, 1.787179e-08, 1.788841e-08, 1.848912e-08, 
    2.014832e-08, 1.95934e-08, 2.214417e-08, 2.405404e-08, 2.231562e-08, 
    2.456523e-08, 2.230345e-08, 1.913339e-08, 1.904179e-08, 2.280085e-08,
  1.705467e-08, 1.775301e-08, 1.829326e-08, 1.915596e-08, 1.96025e-08, 
    2.119757e-08, 2.168598e-08, 2.357665e-08, 2.414004e-08, 2.250098e-08, 
    2.141572e-08, 1.956838e-08, 2.035889e-08, 2.228182e-08, 2.494096e-08,
  1.747208e-08, 1.921981e-08, 2.035527e-08, 2.080203e-08, 2.169971e-08, 
    2.234573e-08, 2.241222e-08, 2.208093e-08, 2.197926e-08, 2.231623e-08, 
    2.19617e-08, 2.269558e-08, 2.376751e-08, 2.548753e-08, 2.507911e-08,
  1.882918e-08, 2.054569e-08, 2.1373e-08, 2.209122e-08, 2.227538e-08, 
    2.228498e-08, 2.274886e-08, 2.172408e-08, 2.263639e-08, 2.438372e-08, 
    2.495125e-08, 2.603987e-08, 2.547121e-08, 2.709183e-08, 2.502299e-08,
  2.004215e-08, 2.108306e-08, 2.220509e-08, 2.318508e-08, 2.348244e-08, 
    2.27978e-08, 2.379493e-08, 2.479741e-08, 2.731108e-08, 2.810158e-08, 
    2.908957e-08, 2.853588e-08, 2.783945e-08, 2.554908e-08, 2.588644e-08,
  1.808017e-08, 1.928839e-08, 1.860544e-08, 1.817148e-08, 1.800531e-08, 
    1.826174e-08, 1.793418e-08, 1.84058e-08, 1.799256e-08, 1.739242e-08, 
    1.796179e-08, 1.807184e-08, 1.862063e-08, 1.900359e-08, 1.850855e-08,
  1.954296e-08, 1.968466e-08, 1.84731e-08, 1.841616e-08, 1.873013e-08, 
    1.884099e-08, 1.825524e-08, 1.95553e-08, 1.915062e-08, 1.861088e-08, 
    1.831819e-08, 1.777937e-08, 1.822095e-08, 1.887933e-08, 1.883537e-08,
  1.997174e-08, 1.901777e-08, 1.889013e-08, 1.93667e-08, 1.930743e-08, 
    1.932465e-08, 1.919768e-08, 1.958009e-08, 1.985573e-08, 1.95023e-08, 
    1.93409e-08, 1.832257e-08, 1.851912e-08, 1.943682e-08, 1.957518e-08,
  1.889465e-08, 1.847634e-08, 1.933708e-08, 2.010535e-08, 2.002688e-08, 
    1.97616e-08, 2.069772e-08, 1.979975e-08, 1.984167e-08, 1.883905e-08, 
    1.755742e-08, 1.765987e-08, 1.982739e-08, 2.042705e-08, 2.096829e-08,
  1.878412e-08, 1.915121e-08, 1.965764e-08, 1.942803e-08, 1.953228e-08, 
    1.952472e-08, 1.991939e-08, 1.993574e-08, 1.95956e-08, 1.685781e-08, 
    1.780369e-08, 1.893254e-08, 1.904944e-08, 1.941038e-08, 2.076015e-08,
  1.973348e-08, 2.049695e-08, 2.0371e-08, 2.025752e-08, 2.083516e-08, 
    2.056485e-08, 2.059559e-08, 1.978874e-08, 1.802168e-08, 1.823792e-08, 
    2.078973e-08, 2.144535e-08, 2.097042e-08, 1.748046e-08, 2.267157e-08,
  2.024555e-08, 2.146439e-08, 2.096307e-08, 2.089766e-08, 2.163659e-08, 
    2.121227e-08, 2.152839e-08, 2.042592e-08, 2.04289e-08, 2.175958e-08, 
    2.208332e-08, 2.214427e-08, 2.098059e-08, 2.055785e-08, 2.885137e-08,
  2.1372e-08, 2.195589e-08, 2.116366e-08, 2.196859e-08, 2.312262e-08, 
    2.317037e-08, 2.350118e-08, 2.221891e-08, 2.178064e-08, 2.205297e-08, 
    2.171266e-08, 2.192188e-08, 2.198042e-08, 2.689356e-08, 2.69773e-08,
  2.244248e-08, 2.205672e-08, 2.16124e-08, 2.296487e-08, 2.325263e-08, 
    2.257638e-08, 2.201543e-08, 2.0728e-08, 2.095733e-08, 2.230478e-08, 
    2.271418e-08, 2.339649e-08, 2.39002e-08, 2.360928e-08, 1.786786e-08,
  2.236905e-08, 2.209582e-08, 2.155893e-08, 2.198293e-08, 2.151835e-08, 
    2.100778e-08, 2.049101e-08, 2.114329e-08, 2.367871e-08, 2.44435e-08, 
    2.441941e-08, 2.466871e-08, 2.479543e-08, 2.100108e-08, 1.983871e-08,
  2.004293e-08, 2.052018e-08, 2.138925e-08, 2.358079e-08, 2.338348e-08, 
    2.258908e-08, 2.275958e-08, 2.297449e-08, 2.427942e-08, 2.494288e-08, 
    2.432476e-08, 2.526444e-08, 2.393534e-08, 1.938731e-08, 2.005567e-08,
  1.993465e-08, 2.011266e-08, 2.253775e-08, 2.482678e-08, 2.378074e-08, 
    2.30519e-08, 2.376503e-08, 2.464028e-08, 2.656041e-08, 2.620829e-08, 
    2.530713e-08, 2.522135e-08, 2.134381e-08, 2.028799e-08, 2.086021e-08,
  2.227026e-08, 2.273489e-08, 2.501278e-08, 2.602078e-08, 2.522272e-08, 
    2.350394e-08, 2.428096e-08, 2.529529e-08, 2.748214e-08, 2.619375e-08, 
    2.80929e-08, 2.700606e-08, 2.321243e-08, 2.204527e-08, 2.262249e-08,
  2.330559e-08, 2.340647e-08, 2.511941e-08, 2.506629e-08, 2.367515e-08, 
    2.394442e-08, 2.516612e-08, 2.60976e-08, 2.76008e-08, 2.389302e-08, 
    2.186569e-08, 1.943419e-08, 2.083143e-08, 2.195845e-08, 2.417263e-08,
  2.51921e-08, 2.481146e-08, 2.422046e-08, 2.33762e-08, 2.353526e-08, 
    2.520178e-08, 2.556758e-08, 2.683871e-08, 2.471662e-08, 1.871438e-08, 
    1.808473e-08, 2.016824e-08, 2.231286e-08, 2.321705e-08, 2.513818e-08,
  2.539886e-08, 2.48157e-08, 2.327996e-08, 2.326173e-08, 2.544094e-08, 
    2.619417e-08, 2.565938e-08, 2.494277e-08, 2.087198e-08, 2.030285e-08, 
    2.421987e-08, 2.494621e-08, 2.463446e-08, 2.521349e-08, 2.597998e-08,
  2.468602e-08, 2.497453e-08, 2.318172e-08, 2.439898e-08, 2.707567e-08, 
    2.621523e-08, 2.577558e-08, 2.359008e-08, 2.343784e-08, 2.45339e-08, 
    2.538749e-08, 2.473985e-08, 2.491383e-08, 2.519e-08, 2.378051e-08,
  2.508608e-08, 2.503377e-08, 2.432571e-08, 2.617835e-08, 2.834958e-08, 
    2.729967e-08, 2.681164e-08, 2.51269e-08, 2.468797e-08, 2.433403e-08, 
    2.527243e-08, 2.498865e-08, 2.558274e-08, 2.501499e-08, 2.168869e-08,
  2.584682e-08, 2.561401e-08, 2.545462e-08, 2.726383e-08, 2.793927e-08, 
    2.628903e-08, 2.469392e-08, 2.304184e-08, 2.326005e-08, 2.495701e-08, 
    2.532392e-08, 2.445459e-08, 2.449599e-08, 2.192364e-08, 2.102991e-08,
  2.623255e-08, 2.54684e-08, 2.557277e-08, 2.521094e-08, 2.400989e-08, 
    2.320833e-08, 2.294061e-08, 2.426767e-08, 2.5764e-08, 2.545248e-08, 
    2.451379e-08, 2.3712e-08, 2.370983e-08, 2.165786e-08, 2.202098e-08,
  1.804073e-08, 1.875987e-08, 1.911117e-08, 1.989591e-08, 1.991726e-08, 
    2.170896e-08, 2.263352e-08, 2.567854e-08, 2.76341e-08, 2.782514e-08, 
    2.478894e-08, 2.570786e-08, 2.69837e-08, 2.610556e-08, 2.501634e-08,
  1.837436e-08, 1.84096e-08, 1.990556e-08, 2.128403e-08, 2.229594e-08, 
    2.262571e-08, 2.320061e-08, 2.655613e-08, 2.901312e-08, 2.897845e-08, 
    2.799623e-08, 2.764225e-08, 2.702948e-08, 2.440805e-08, 2.393181e-08,
  1.94488e-08, 1.891321e-08, 2.094834e-08, 2.284267e-08, 2.322391e-08, 
    2.203104e-08, 2.32034e-08, 2.638493e-08, 2.946605e-08, 3.005166e-08, 
    3.008332e-08, 2.73533e-08, 2.652882e-08, 2.395366e-08, 2.750008e-08,
  1.915402e-08, 1.878387e-08, 2.045734e-08, 2.121336e-08, 2.105058e-08, 
    2.153102e-08, 2.389263e-08, 2.694328e-08, 2.867058e-08, 2.424099e-08, 
    2.16589e-08, 2.19561e-08, 2.556409e-08, 2.678299e-08, 3.002276e-08,
  1.912657e-08, 1.942278e-08, 1.982215e-08, 2.016632e-08, 2.075682e-08, 
    2.162026e-08, 2.389846e-08, 2.599407e-08, 2.381224e-08, 1.822066e-08, 
    1.950297e-08, 2.526344e-08, 3.081665e-08, 2.958565e-08, 2.867674e-08,
  1.981392e-08, 1.970391e-08, 1.992482e-08, 2.034252e-08, 2.106872e-08, 
    2.273678e-08, 2.513939e-08, 2.471124e-08, 2.175043e-08, 2.120459e-08, 
    2.786184e-08, 2.823793e-08, 3.233777e-08, 3.210854e-08, 2.951863e-08,
  1.939184e-08, 1.993169e-08, 2.016348e-08, 2.100258e-08, 2.249512e-08, 
    2.494101e-08, 2.566629e-08, 2.53278e-08, 2.398254e-08, 2.638312e-08, 
    2.980098e-08, 2.871709e-08, 3.418074e-08, 3.444084e-08, 2.753398e-08,
  1.943051e-08, 2.035164e-08, 2.047962e-08, 2.21407e-08, 2.431699e-08, 
    2.63754e-08, 2.710655e-08, 2.578971e-08, 2.445258e-08, 2.69723e-08, 
    2.863794e-08, 2.91585e-08, 3.313755e-08, 3.201113e-08, 2.229852e-08,
  1.989494e-08, 2.052201e-08, 2.111301e-08, 2.295313e-08, 2.508381e-08, 
    2.61255e-08, 2.483597e-08, 2.284293e-08, 2.43589e-08, 2.867618e-08, 
    2.836332e-08, 2.863101e-08, 2.879375e-08, 2.517749e-08, 2.192853e-08,
  2.055682e-08, 2.108178e-08, 2.154966e-08, 2.235428e-08, 2.325565e-08, 
    2.319714e-08, 2.280016e-08, 2.526938e-08, 2.8353e-08, 2.831632e-08, 
    2.791229e-08, 2.782525e-08, 2.741157e-08, 2.382403e-08, 2.290686e-08,
  1.45982e-08, 1.50531e-08, 1.501822e-08, 1.546078e-08, 1.610898e-08, 
    1.653878e-08, 1.735213e-08, 1.829571e-08, 1.930405e-08, 2.03166e-08, 
    1.959159e-08, 2.084758e-08, 2.341083e-08, 2.428342e-08, 2.289678e-08,
  1.500864e-08, 1.534484e-08, 1.558276e-08, 1.582076e-08, 1.645651e-08, 
    1.736513e-08, 1.802083e-08, 1.885885e-08, 2.051741e-08, 2.165176e-08, 
    2.130362e-08, 2.268503e-08, 2.385356e-08, 2.223027e-08, 2.181134e-08,
  1.546292e-08, 1.601591e-08, 1.610958e-08, 1.648179e-08, 1.712378e-08, 
    1.784344e-08, 1.850757e-08, 1.954263e-08, 2.148325e-08, 2.223997e-08, 
    2.235759e-08, 2.31423e-08, 2.365477e-08, 2.142166e-08, 2.427419e-08,
  1.676401e-08, 1.65877e-08, 1.660206e-08, 1.685685e-08, 1.73738e-08, 
    1.803232e-08, 1.920883e-08, 2.050156e-08, 2.164303e-08, 2.088976e-08, 
    1.947e-08, 2.085331e-08, 2.256354e-08, 2.331084e-08, 2.881722e-08,
  1.707902e-08, 1.682082e-08, 1.70343e-08, 1.716065e-08, 1.772994e-08, 
    1.836144e-08, 1.886717e-08, 2.03505e-08, 2.012162e-08, 1.666484e-08, 
    1.831393e-08, 2.204724e-08, 2.478371e-08, 2.642681e-08, 2.834756e-08,
  1.770506e-08, 1.74545e-08, 1.756228e-08, 1.799145e-08, 1.868879e-08, 
    1.877078e-08, 1.944245e-08, 2.01318e-08, 1.863633e-08, 1.889424e-08, 
    2.357025e-08, 2.372404e-08, 2.60963e-08, 2.854054e-08, 2.68918e-08,
  1.764694e-08, 1.790829e-08, 1.839864e-08, 1.91308e-08, 1.961188e-08, 
    2.031619e-08, 2.104255e-08, 2.117287e-08, 2.054995e-08, 2.258487e-08, 
    2.44618e-08, 2.409307e-08, 2.843038e-08, 3.032145e-08, 2.32593e-08,
  1.780268e-08, 1.9004e-08, 1.980902e-08, 2.025045e-08, 2.077022e-08, 
    2.199248e-08, 2.229746e-08, 2.212755e-08, 2.144804e-08, 2.312216e-08, 
    2.445135e-08, 2.509547e-08, 2.88197e-08, 2.799644e-08, 2.029817e-08,
  1.896168e-08, 2.003999e-08, 2.032947e-08, 2.07625e-08, 2.114219e-08, 
    2.155492e-08, 2.164277e-08, 2.083092e-08, 2.120325e-08, 2.458587e-08, 
    2.489636e-08, 2.519016e-08, 2.620051e-08, 2.384084e-08, 2.253398e-08,
  1.99314e-08, 2.019559e-08, 1.966901e-08, 1.978339e-08, 1.97848e-08, 
    1.893143e-08, 1.939262e-08, 2.056352e-08, 2.394209e-08, 2.504466e-08, 
    2.455701e-08, 2.471942e-08, 2.498422e-08, 2.410631e-08, 2.409066e-08,
  1.622465e-08, 1.66408e-08, 1.700306e-08, 1.736266e-08, 1.775537e-08, 
    1.755777e-08, 1.74262e-08, 1.723131e-08, 1.775372e-08, 1.685488e-08, 
    1.479614e-08, 1.580704e-08, 1.69838e-08, 1.705824e-08, 1.67797e-08,
  1.886482e-08, 1.908502e-08, 1.915869e-08, 1.897394e-08, 1.949807e-08, 
    1.962778e-08, 1.906482e-08, 1.893487e-08, 1.934299e-08, 1.937634e-08, 
    1.764841e-08, 1.764033e-08, 1.768742e-08, 1.812998e-08, 1.80707e-08,
  2.162511e-08, 2.174281e-08, 2.092766e-08, 2.077639e-08, 2.102868e-08, 
    2.120126e-08, 2.094912e-08, 2.13004e-08, 2.15911e-08, 2.108279e-08, 
    2.011568e-08, 2.00006e-08, 2.176365e-08, 2.020858e-08, 2.106585e-08,
  2.244361e-08, 2.189042e-08, 2.151795e-08, 2.207037e-08, 2.151442e-08, 
    2.162946e-08, 2.207897e-08, 2.262204e-08, 2.249869e-08, 2.206025e-08, 
    1.774954e-08, 1.71901e-08, 1.923393e-08, 2.007787e-08, 2.382662e-08,
  2.181103e-08, 2.145345e-08, 2.123844e-08, 2.110185e-08, 2.090283e-08, 
    2.081496e-08, 2.110145e-08, 2.115806e-08, 1.958187e-08, 1.623808e-08, 
    1.638997e-08, 1.893887e-08, 1.7856e-08, 2.160469e-08, 2.403983e-08,
  2.384409e-08, 2.306955e-08, 2.302376e-08, 2.283155e-08, 2.282079e-08, 
    2.234884e-08, 2.107405e-08, 2.046118e-08, 1.776425e-08, 1.717334e-08, 
    2.024221e-08, 2.04212e-08, 1.937033e-08, 2.301998e-08, 2.374957e-08,
  2.343451e-08, 2.342198e-08, 2.372231e-08, 2.343182e-08, 2.335201e-08, 
    2.282788e-08, 2.263468e-08, 2.122611e-08, 2.052411e-08, 2.115326e-08, 
    2.279333e-08, 2.178434e-08, 2.333334e-08, 2.742684e-08, 2.191011e-08,
  2.305559e-08, 2.39878e-08, 2.39903e-08, 2.380924e-08, 2.352293e-08, 
    2.353059e-08, 2.332438e-08, 2.26771e-08, 2.25575e-08, 2.278342e-08, 
    2.281695e-08, 2.275672e-08, 2.42616e-08, 2.298182e-08, 1.576537e-08,
  2.44489e-08, 2.484277e-08, 2.487839e-08, 2.47299e-08, 2.468561e-08, 
    2.397805e-08, 2.399308e-08, 2.267816e-08, 2.247276e-08, 2.272988e-08, 
    2.288311e-08, 2.293624e-08, 2.259004e-08, 2.038823e-08, 1.674396e-08,
  2.519804e-08, 2.521834e-08, 2.469352e-08, 2.462505e-08, 2.423791e-08, 
    2.391902e-08, 2.324201e-08, 2.306445e-08, 2.348911e-08, 2.366284e-08, 
    2.355489e-08, 2.335993e-08, 2.327298e-08, 2.177451e-08, 2.174271e-08,
  2.219221e-08, 2.256144e-08, 2.234753e-08, 2.307743e-08, 2.332183e-08, 
    2.359365e-08, 2.310976e-08, 2.337788e-08, 2.263312e-08, 2.182751e-08, 
    2.067381e-08, 2.098431e-08, 2.281154e-08, 2.188446e-08, 2.256733e-08,
  2.396997e-08, 2.407047e-08, 2.39153e-08, 2.375939e-08, 2.47451e-08, 
    2.551538e-08, 2.481366e-08, 2.477325e-08, 2.454399e-08, 2.421132e-08, 
    2.405295e-08, 2.39926e-08, 2.450372e-08, 2.353927e-08, 2.332913e-08,
  2.417421e-08, 2.527424e-08, 2.544129e-08, 2.560014e-08, 2.6142e-08, 
    2.661815e-08, 2.684136e-08, 2.668719e-08, 2.648101e-08, 2.569611e-08, 
    2.546468e-08, 2.558839e-08, 2.705854e-08, 2.710262e-08, 2.727263e-08,
  2.502558e-08, 2.615115e-08, 2.560709e-08, 2.573648e-08, 2.579264e-08, 
    2.584007e-08, 2.666871e-08, 2.678135e-08, 2.599869e-08, 2.563899e-08, 
    2.28913e-08, 2.229354e-08, 2.469724e-08, 2.767055e-08, 3.115701e-08,
  2.538532e-08, 2.609133e-08, 2.601587e-08, 2.527861e-08, 2.552575e-08, 
    2.583906e-08, 2.655193e-08, 2.598878e-08, 2.617747e-08, 2.260366e-08, 
    2.263041e-08, 2.321546e-08, 2.290688e-08, 2.547317e-08, 2.928561e-08,
  2.725337e-08, 2.77655e-08, 2.791977e-08, 2.757983e-08, 2.753372e-08, 
    2.771626e-08, 2.680863e-08, 2.685016e-08, 2.443415e-08, 2.443711e-08, 
    2.70689e-08, 2.721162e-08, 2.572355e-08, 2.717448e-08, 2.79532e-08,
  2.7373e-08, 2.763917e-08, 2.831407e-08, 2.806132e-08, 2.822998e-08, 
    2.839482e-08, 2.740957e-08, 2.699212e-08, 2.575985e-08, 2.760908e-08, 
    2.808145e-08, 2.724648e-08, 2.794321e-08, 2.807869e-08, 2.599025e-08,
  2.726394e-08, 2.778439e-08, 2.821444e-08, 2.831854e-08, 2.877902e-08, 
    2.925008e-08, 2.866472e-08, 2.766926e-08, 2.672396e-08, 2.740837e-08, 
    2.7163e-08, 2.673656e-08, 2.726936e-08, 2.713223e-08, 2.432908e-08,
  2.571958e-08, 2.701944e-08, 2.744468e-08, 2.730622e-08, 2.811353e-08, 
    2.78463e-08, 2.724929e-08, 2.556477e-08, 2.585598e-08, 2.72059e-08, 
    2.683149e-08, 2.654629e-08, 2.676157e-08, 2.616091e-08, 2.518656e-08,
  2.468245e-08, 2.587812e-08, 2.586451e-08, 2.553598e-08, 2.504114e-08, 
    2.542411e-08, 2.50185e-08, 2.546108e-08, 2.66108e-08, 2.630775e-08, 
    2.604171e-08, 2.59346e-08, 2.639073e-08, 2.619024e-08, 2.62077e-08,
  2.655317e-08, 2.662977e-08, 2.695576e-08, 2.728037e-08, 2.749981e-08, 
    2.724365e-08, 2.715e-08, 2.715417e-08, 2.659889e-08, 2.604223e-08, 
    2.597621e-08, 2.657025e-08, 2.636891e-08, 2.568333e-08, 2.734578e-08,
  2.829683e-08, 2.876076e-08, 2.865141e-08, 2.848849e-08, 2.860076e-08, 
    2.845629e-08, 2.786158e-08, 2.813303e-08, 2.819115e-08, 2.797995e-08, 
    2.829189e-08, 2.75839e-08, 2.707569e-08, 2.647687e-08, 2.638713e-08,
  2.878961e-08, 3.023608e-08, 3.005602e-08, 3.01028e-08, 2.95073e-08, 
    3.06247e-08, 2.969157e-08, 2.928284e-08, 2.905175e-08, 2.933541e-08, 
    2.946243e-08, 2.966415e-08, 2.909604e-08, 2.850998e-08, 2.824222e-08,
  2.935081e-08, 3.010974e-08, 2.903984e-08, 2.886106e-08, 2.816207e-08, 
    2.96612e-08, 2.884052e-08, 3.011012e-08, 3.011184e-08, 3.017244e-08, 
    2.802714e-08, 2.843011e-08, 2.959095e-08, 2.869565e-08, 2.93254e-08,
  2.909446e-08, 2.855452e-08, 2.642902e-08, 2.501603e-08, 2.427765e-08, 
    2.405323e-08, 2.506967e-08, 2.60248e-08, 2.661847e-08, 2.702633e-08, 
    2.779637e-08, 2.685199e-08, 2.643044e-08, 2.714361e-08, 2.898757e-08,
  2.86795e-08, 2.557776e-08, 2.193261e-08, 2.046818e-08, 1.984533e-08, 
    2.012837e-08, 2.084497e-08, 2.237739e-08, 2.347007e-08, 2.257141e-08, 
    2.743556e-08, 2.775278e-08, 2.669997e-08, 2.653709e-08, 2.908893e-08,
  2.591336e-08, 2.095284e-08, 1.770483e-08, 1.689192e-08, 1.754901e-08, 
    1.808179e-08, 1.904827e-08, 2.024953e-08, 2.106701e-08, 2.24559e-08, 
    2.430127e-08, 2.518767e-08, 2.591724e-08, 2.525758e-08, 2.81676e-08,
  2.493489e-08, 2.060583e-08, 1.658645e-08, 1.710864e-08, 1.808556e-08, 
    1.939524e-08, 2.05239e-08, 2.12639e-08, 2.296998e-08, 2.345418e-08, 
    2.35144e-08, 2.431679e-08, 2.431725e-08, 2.436767e-08, 2.447531e-08,
  2.42225e-08, 2.031551e-08, 1.867186e-08, 1.88509e-08, 1.8875e-08, 
    2.038378e-08, 2.200984e-08, 2.354568e-08, 2.311719e-08, 2.346738e-08, 
    2.391712e-08, 2.475977e-08, 2.488572e-08, 2.463232e-08, 2.416328e-08,
  2.593239e-08, 2.273467e-08, 2.15952e-08, 1.94457e-08, 1.967988e-08, 
    2.032818e-08, 2.119627e-08, 2.185095e-08, 2.218117e-08, 2.313168e-08, 
    2.353816e-08, 2.35457e-08, 2.414328e-08, 2.434418e-08, 2.487257e-08,
  2.666932e-08, 2.641989e-08, 2.710345e-08, 2.677039e-08, 2.771727e-08, 
    2.819331e-08, 2.853917e-08, 2.922848e-08, 2.903359e-08, 2.867455e-08, 
    2.856887e-08, 2.796994e-08, 2.841359e-08, 2.71502e-08, 2.739729e-08,
  2.615525e-08, 2.605659e-08, 2.761268e-08, 2.884234e-08, 2.926883e-08, 
    2.93209e-08, 2.953975e-08, 2.984203e-08, 2.937729e-08, 2.964886e-08, 
    2.923656e-08, 2.898709e-08, 2.918681e-08, 2.791247e-08, 2.828126e-08,
  2.568279e-08, 2.796501e-08, 3.023827e-08, 3.073264e-08, 3.001652e-08, 
    2.866208e-08, 2.773669e-08, 2.738353e-08, 2.662737e-08, 2.589908e-08, 
    2.611369e-08, 2.621988e-08, 2.727166e-08, 2.68629e-08, 2.874031e-08,
  2.81733e-08, 3.193398e-08, 3.088839e-08, 2.9833e-08, 2.837047e-08, 
    2.698089e-08, 2.515489e-08, 2.440972e-08, 2.265442e-08, 2.177221e-08, 
    2.305069e-08, 2.509582e-08, 2.644805e-08, 2.702133e-08, 2.901884e-08,
  3.302704e-08, 3.546726e-08, 3.494111e-08, 3.244255e-08, 2.927278e-08, 
    2.719398e-08, 2.469128e-08, 2.276771e-08, 2.045577e-08, 2.071695e-08, 
    2.155387e-08, 2.301609e-08, 2.143467e-08, 2.373078e-08, 2.391659e-08,
  3.538428e-08, 3.608198e-08, 3.241282e-08, 2.96626e-08, 2.73575e-08, 
    2.494919e-08, 2.289718e-08, 2.026767e-08, 1.849862e-08, 1.744293e-08, 
    1.686233e-08, 1.701281e-08, 1.753257e-08, 1.936572e-08, 1.997252e-08,
  3.60636e-08, 3.73178e-08, 3.349271e-08, 3.084254e-08, 2.833913e-08, 
    2.569625e-08, 2.310101e-08, 2.017783e-08, 1.866859e-08, 1.834605e-08, 
    1.850496e-08, 1.70465e-08, 1.797482e-08, 1.760246e-08, 1.606679e-08,
  3.682992e-08, 3.698063e-08, 3.381135e-08, 3.044456e-08, 2.685432e-08, 
    2.48837e-08, 2.252796e-08, 2.039092e-08, 1.971471e-08, 1.999571e-08, 
    2.026923e-08, 1.916155e-08, 1.97629e-08, 1.892106e-08, 1.597203e-08,
  3.60323e-08, 3.610549e-08, 3.411939e-08, 2.88967e-08, 2.506932e-08, 
    2.547402e-08, 2.34444e-08, 2.137255e-08, 2.075561e-08, 2.090421e-08, 
    2.115971e-08, 2.096222e-08, 2.173867e-08, 2.07655e-08, 1.906766e-08,
  3.616494e-08, 3.491337e-08, 3.070369e-08, 2.527596e-08, 2.506045e-08, 
    2.591993e-08, 2.236886e-08, 2.08374e-08, 2.091551e-08, 2.124369e-08, 
    2.161295e-08, 2.212752e-08, 2.259892e-08, 2.205369e-08, 2.142038e-08,
  2.740143e-08, 2.915027e-08, 3.037547e-08, 3.33404e-08, 3.390429e-08, 
    3.484141e-08, 3.570915e-08, 3.743442e-08, 3.966333e-08, 4.060871e-08, 
    3.981865e-08, 3.939777e-08, 4.011228e-08, 3.891809e-08, 3.391548e-08,
  2.868966e-08, 3.127446e-08, 3.281171e-08, 3.481822e-08, 3.444222e-08, 
    3.649508e-08, 3.69299e-08, 3.926259e-08, 3.964056e-08, 3.897375e-08, 
    3.650998e-08, 3.579337e-08, 3.456883e-08, 3.411977e-08, 3.03137e-08,
  2.975557e-08, 3.317163e-08, 3.43402e-08, 3.679408e-08, 3.64523e-08, 
    3.597212e-08, 3.479526e-08, 3.564733e-08, 3.869522e-08, 3.63659e-08, 
    3.424607e-08, 3.300319e-08, 3.169367e-08, 2.881455e-08, 2.817799e-08,
  3.47115e-08, 3.624228e-08, 3.753287e-08, 4.014207e-08, 3.560515e-08, 
    3.412907e-08, 3.32003e-08, 3.044259e-08, 3.002e-08, 3.160556e-08, 
    2.622716e-08, 2.406676e-08, 2.615155e-08, 2.594311e-08, 2.909474e-08,
  3.534241e-08, 3.590882e-08, 3.654275e-08, 3.215548e-08, 3.140581e-08, 
    3.175667e-08, 3.067377e-08, 3.003948e-08, 2.463475e-08, 1.763657e-08, 
    1.747682e-08, 2.114635e-08, 2.165111e-08, 2.890841e-08, 3.142158e-08,
  3.760402e-08, 3.683053e-08, 3.142872e-08, 2.829644e-08, 3.031478e-08, 
    2.940805e-08, 2.808548e-08, 2.788213e-08, 2.277189e-08, 1.890728e-08, 
    2.40002e-08, 2.509497e-08, 2.325573e-08, 2.91451e-08, 2.702066e-08,
  3.769927e-08, 2.931304e-08, 2.564629e-08, 2.874788e-08, 3.09835e-08, 
    2.935554e-08, 2.772684e-08, 2.456364e-08, 2.255147e-08, 2.417108e-08, 
    2.51067e-08, 2.457522e-08, 2.464387e-08, 2.687791e-08, 2.17368e-08,
  3.06843e-08, 2.452355e-08, 2.593047e-08, 3.006561e-08, 3.009428e-08, 
    2.774802e-08, 2.583132e-08, 2.31598e-08, 2.234413e-08, 2.38593e-08, 
    2.438889e-08, 2.510428e-08, 2.567133e-08, 2.276542e-08, 1.851688e-08,
  2.820362e-08, 2.697258e-08, 2.846189e-08, 2.943025e-08, 2.837514e-08, 
    2.735741e-08, 2.649224e-08, 2.360811e-08, 2.290534e-08, 2.58078e-08, 
    2.610329e-08, 2.669309e-08, 2.582453e-08, 2.173363e-08, 1.966323e-08,
  2.885762e-08, 2.892511e-08, 2.859013e-08, 2.884392e-08, 2.725393e-08, 
    2.646776e-08, 2.47465e-08, 2.362705e-08, 2.537715e-08, 2.578574e-08, 
    2.487499e-08, 2.449596e-08, 2.483148e-08, 2.22615e-08, 2.23841e-08,
  2.575862e-08, 2.63144e-08, 2.65343e-08, 2.670467e-08, 2.749847e-08, 
    2.750352e-08, 2.780829e-08, 2.689251e-08, 2.662579e-08, 2.65464e-08, 
    2.798487e-08, 3.157164e-08, 3.501358e-08, 3.70314e-08, 3.953411e-08,
  2.937828e-08, 2.977298e-08, 2.968336e-08, 2.907666e-08, 2.9402e-08, 
    2.978537e-08, 2.933932e-08, 3.016252e-08, 2.93291e-08, 2.874056e-08, 
    2.861194e-08, 2.831796e-08, 2.742322e-08, 2.887556e-08, 2.8364e-08,
  3.187791e-08, 2.896059e-08, 2.749828e-08, 2.767335e-08, 2.673946e-08, 
    2.756484e-08, 2.630897e-08, 2.578273e-08, 2.546841e-08, 2.458707e-08, 
    2.613176e-08, 2.491675e-08, 2.50479e-08, 2.475377e-08, 2.406282e-08,
  2.923456e-08, 2.524488e-08, 2.571687e-08, 2.582498e-08, 2.503006e-08, 
    2.509803e-08, 2.566768e-08, 2.603194e-08, 2.441248e-08, 2.248511e-08, 
    1.984492e-08, 1.905488e-08, 2.125418e-08, 2.07117e-08, 2.241694e-08,
  2.713126e-08, 2.554794e-08, 2.620975e-08, 2.565863e-08, 2.621349e-08, 
    2.57151e-08, 2.690142e-08, 2.62656e-08, 2.597343e-08, 2.169181e-08, 
    2.072665e-08, 2.158767e-08, 2.162474e-08, 2.110589e-08, 2.190392e-08,
  2.870416e-08, 2.738e-08, 2.628127e-08, 2.641218e-08, 2.721668e-08, 
    2.685355e-08, 2.627801e-08, 2.635253e-08, 2.524246e-08, 2.242553e-08, 
    2.794573e-08, 2.782997e-08, 2.60166e-08, 2.205029e-08, 2.341132e-08,
  2.843493e-08, 2.657852e-08, 2.605769e-08, 2.728071e-08, 2.871176e-08, 
    2.774768e-08, 2.747527e-08, 2.759613e-08, 2.711801e-08, 2.979877e-08, 
    3.171484e-08, 3.290415e-08, 3.110641e-08, 2.704314e-08, 2.750854e-08,
  2.801816e-08, 2.976474e-08, 2.846548e-08, 2.976679e-08, 2.97651e-08, 
    2.765495e-08, 2.727164e-08, 2.788298e-08, 2.729746e-08, 2.995126e-08, 
    3.051169e-08, 3.163218e-08, 3.136622e-08, 2.971e-08, 3.031633e-08,
  2.962369e-08, 3.026593e-08, 2.958399e-08, 2.997173e-08, 2.906511e-08, 
    2.619542e-08, 2.579377e-08, 2.406337e-08, 2.161207e-08, 2.341881e-08, 
    2.341659e-08, 2.458168e-08, 2.68169e-08, 2.84271e-08, 2.917423e-08,
  3.063841e-08, 3.219093e-08, 3.035482e-08, 3.092555e-08, 2.811403e-08, 
    2.568387e-08, 2.287372e-08, 1.908809e-08, 1.937314e-08, 1.985369e-08, 
    1.974452e-08, 1.970471e-08, 2.053307e-08, 2.0409e-08, 2.213985e-08,
  2.684482e-08, 2.80121e-08, 2.813446e-08, 2.866611e-08, 2.9109e-08, 
    3.013961e-08, 2.9867e-08, 3.029023e-08, 3.089741e-08, 3.000318e-08, 
    2.842792e-08, 2.89729e-08, 2.798263e-08, 2.411837e-08, 2.53266e-08,
  2.794858e-08, 2.90681e-08, 2.926347e-08, 2.843661e-08, 2.910393e-08, 
    2.942368e-08, 2.929068e-08, 2.894483e-08, 2.939597e-08, 2.894616e-08, 
    2.763276e-08, 2.88428e-08, 2.736035e-08, 2.704052e-08, 2.551375e-08,
  2.956853e-08, 2.783341e-08, 2.628491e-08, 2.813952e-08, 2.794439e-08, 
    2.745881e-08, 2.585763e-08, 2.630135e-08, 2.63388e-08, 2.700306e-08, 
    2.617909e-08, 2.69982e-08, 2.585491e-08, 2.643536e-08, 2.570937e-08,
  2.723845e-08, 2.66494e-08, 2.851591e-08, 2.871503e-08, 2.741919e-08, 
    2.603836e-08, 2.525822e-08, 2.661086e-08, 2.613068e-08, 2.628857e-08, 
    2.335686e-08, 2.559052e-08, 2.423103e-08, 2.59499e-08, 2.331227e-08,
  2.753478e-08, 2.752389e-08, 2.805032e-08, 2.708215e-08, 2.637267e-08, 
    2.628174e-08, 2.638655e-08, 2.640258e-08, 2.475545e-08, 2.406592e-08, 
    2.162812e-08, 2.485808e-08, 2.499782e-08, 2.518962e-08, 2.252361e-08,
  2.753756e-08, 2.718426e-08, 2.685235e-08, 2.624484e-08, 2.6861e-08, 
    2.662264e-08, 2.730364e-08, 2.658392e-08, 2.573933e-08, 2.306593e-08, 
    2.290618e-08, 2.247005e-08, 2.255632e-08, 2.155161e-08, 2.449068e-08,
  2.650465e-08, 2.63629e-08, 2.676908e-08, 2.6295e-08, 2.666291e-08, 
    2.600874e-08, 2.630122e-08, 2.577388e-08, 2.532187e-08, 2.255626e-08, 
    2.216597e-08, 2.185712e-08, 2.232778e-08, 2.205165e-08, 2.395339e-08,
  2.635624e-08, 2.662543e-08, 2.661806e-08, 2.644914e-08, 2.694721e-08, 
    2.684024e-08, 2.798712e-08, 2.749383e-08, 2.462691e-08, 2.301132e-08, 
    2.346202e-08, 2.284904e-08, 2.308644e-08, 2.226523e-08, 2.291684e-08,
  2.60372e-08, 2.621312e-08, 2.616856e-08, 2.691961e-08, 2.792439e-08, 
    2.755068e-08, 2.772501e-08, 2.755421e-08, 2.576806e-08, 2.577942e-08, 
    2.699803e-08, 2.576733e-08, 2.485348e-08, 2.263241e-08, 2.142518e-08,
  2.6332e-08, 2.645482e-08, 2.576823e-08, 2.684891e-08, 2.822338e-08, 
    2.804783e-08, 2.806826e-08, 2.659559e-08, 2.580569e-08, 2.771991e-08, 
    2.884759e-08, 2.697574e-08, 2.572483e-08, 2.466074e-08, 2.283503e-08,
  2.582187e-08, 2.591642e-08, 2.606861e-08, 2.644149e-08, 2.6728e-08, 
    2.673397e-08, 2.688824e-08, 2.710444e-08, 2.780967e-08, 2.664843e-08, 
    2.658244e-08, 2.599587e-08, 2.689797e-08, 2.638181e-08, 2.643355e-08,
  2.531715e-08, 2.533433e-08, 2.579401e-08, 2.590043e-08, 2.624437e-08, 
    2.592777e-08, 2.585249e-08, 2.615395e-08, 2.59298e-08, 2.526403e-08, 
    2.524369e-08, 2.496165e-08, 2.551365e-08, 2.459079e-08, 2.444976e-08,
  2.594764e-08, 2.503213e-08, 2.487422e-08, 2.454367e-08, 2.520651e-08, 
    2.533845e-08, 2.517702e-08, 2.49552e-08, 2.487582e-08, 2.480452e-08, 
    2.500886e-08, 2.517051e-08, 2.591623e-08, 2.560703e-08, 2.658962e-08,
  2.695591e-08, 2.50985e-08, 2.488588e-08, 2.544104e-08, 2.60366e-08, 
    2.527037e-08, 2.478476e-08, 2.479151e-08, 2.541719e-08, 2.493293e-08, 
    2.716422e-08, 2.74099e-08, 2.824946e-08, 2.907685e-08, 3.080903e-08,
  2.684045e-08, 2.719953e-08, 2.713853e-08, 2.561931e-08, 2.565532e-08, 
    2.578623e-08, 2.527217e-08, 2.529405e-08, 2.653294e-08, 2.77172e-08, 
    2.723266e-08, 2.810064e-08, 2.93145e-08, 2.947352e-08, 2.780642e-08,
  2.653452e-08, 2.595823e-08, 2.568353e-08, 2.585347e-08, 2.63417e-08, 
    2.616757e-08, 2.600014e-08, 2.725245e-08, 2.849557e-08, 2.756456e-08, 
    2.712981e-08, 2.737898e-08, 3.052337e-08, 2.825196e-08, 2.423423e-08,
  2.625924e-08, 2.601235e-08, 2.542109e-08, 2.527882e-08, 2.548213e-08, 
    2.595123e-08, 2.603836e-08, 2.683941e-08, 2.706302e-08, 2.627401e-08, 
    2.729465e-08, 2.793421e-08, 2.96265e-08, 2.661561e-08, 2.603421e-08,
  2.666967e-08, 2.554693e-08, 2.543831e-08, 2.512447e-08, 2.496139e-08, 
    2.512734e-08, 2.502702e-08, 2.580129e-08, 2.647379e-08, 2.632438e-08, 
    2.719958e-08, 2.757696e-08, 2.817158e-08, 2.952275e-08, 2.858513e-08,
  2.652686e-08, 2.60161e-08, 2.536954e-08, 2.530301e-08, 2.525152e-08, 
    2.591725e-08, 2.628124e-08, 2.64175e-08, 2.547519e-08, 2.550218e-08, 
    2.611416e-08, 2.638258e-08, 2.720884e-08, 2.968521e-08, 2.662892e-08,
  2.624182e-08, 2.626755e-08, 2.582165e-08, 2.579416e-08, 2.580833e-08, 
    2.591816e-08, 2.561829e-08, 2.525407e-08, 2.439927e-08, 2.495065e-08, 
    2.539167e-08, 2.543198e-08, 2.641164e-08, 2.668867e-08, 2.636093e-08,
  2.511051e-08, 2.446562e-08, 2.574789e-08, 2.553486e-08, 2.534248e-08, 
    2.481188e-08, 2.465672e-08, 2.578924e-08, 2.486465e-08, 2.442822e-08, 
    2.510504e-08, 2.506685e-08, 2.514574e-08, 2.499822e-08, 2.566281e-08,
  2.327097e-08, 2.307085e-08, 2.506559e-08, 2.469149e-08, 2.408215e-08, 
    2.429382e-08, 2.518732e-08, 2.560401e-08, 2.437754e-08, 2.437164e-08, 
    2.459892e-08, 2.420699e-08, 2.44256e-08, 2.446215e-08, 2.50505e-08,
  2.302887e-08, 2.299807e-08, 2.415958e-08, 2.374193e-08, 2.414237e-08, 
    2.474948e-08, 2.423186e-08, 2.427559e-08, 2.454264e-08, 2.426553e-08, 
    2.32543e-08, 2.310904e-08, 2.302409e-08, 2.372123e-08, 2.364589e-08,
  2.409068e-08, 2.413439e-08, 2.434257e-08, 2.464266e-08, 2.626751e-08, 
    2.441264e-08, 2.365593e-08, 2.40425e-08, 2.391429e-08, 2.345168e-08, 
    2.835485e-08, 2.945355e-08, 2.677908e-08, 2.727478e-08, 2.471771e-08,
  2.46187e-08, 2.444016e-08, 2.536393e-08, 2.555415e-08, 2.478845e-08, 
    2.546472e-08, 2.451929e-08, 2.331286e-08, 2.354013e-08, 2.748238e-08, 
    2.670673e-08, 2.597409e-08, 2.642571e-08, 2.58095e-08, 2.276007e-08,
  2.474402e-08, 2.393525e-08, 2.325563e-08, 2.347041e-08, 2.393595e-08, 
    2.384729e-08, 2.304209e-08, 2.141356e-08, 2.223957e-08, 2.229975e-08, 
    2.142195e-08, 2.160558e-08, 2.427766e-08, 2.303997e-08, 2.219243e-08,
  2.486162e-08, 2.414139e-08, 2.352242e-08, 2.37109e-08, 2.369993e-08, 
    2.342478e-08, 2.208735e-08, 2.000959e-08, 2.025715e-08, 2.044477e-08, 
    2.10901e-08, 2.115603e-08, 2.186362e-08, 2.157646e-08, 2.193484e-08,
  2.5415e-08, 2.445869e-08, 2.344419e-08, 2.340051e-08, 2.369022e-08, 
    2.305728e-08, 2.116e-08, 1.918156e-08, 1.969433e-08, 2.026249e-08, 
    2.087356e-08, 2.079033e-08, 2.147601e-08, 2.245428e-08, 2.179644e-08,
  2.51688e-08, 2.512304e-08, 2.402584e-08, 2.414818e-08, 2.454507e-08, 
    2.339416e-08, 2.043034e-08, 1.948659e-08, 2.024061e-08, 2.040691e-08, 
    2.080195e-08, 2.081322e-08, 2.064906e-08, 1.970199e-08, 1.819499e-08,
  2.46649e-08, 2.482724e-08, 2.39275e-08, 2.428335e-08, 2.471887e-08, 
    2.204952e-08, 1.874852e-08, 1.914807e-08, 2.058079e-08, 2.065714e-08, 
    2.104348e-08, 2.029811e-08, 1.957388e-08, 1.705539e-08, 1.584131e-08,
  2.43558e-08, 2.35797e-08, 2.285881e-08, 2.251191e-08, 2.227264e-08, 
    2.238124e-08, 2.293287e-08, 2.312157e-08, 2.221318e-08, 2.231694e-08, 
    2.086525e-08, 2.258067e-08, 2.217576e-08, 2.156651e-08, 2.234522e-08,
  2.346689e-08, 2.235963e-08, 2.261172e-08, 2.245879e-08, 2.2008e-08, 
    2.253104e-08, 2.304817e-08, 2.277364e-08, 2.275816e-08, 2.229963e-08, 
    2.112759e-08, 2.258489e-08, 2.164469e-08, 2.159236e-08, 2.207942e-08,
  2.275388e-08, 2.27677e-08, 2.272334e-08, 2.242347e-08, 2.309051e-08, 
    2.379449e-08, 2.36349e-08, 2.323414e-08, 2.290754e-08, 2.150288e-08, 
    2.223477e-08, 2.323548e-08, 2.13046e-08, 2.341685e-08, 2.241603e-08,
  2.385597e-08, 2.441275e-08, 2.416509e-08, 2.382221e-08, 2.550662e-08, 
    2.562131e-08, 2.487655e-08, 2.436826e-08, 2.332662e-08, 2.21394e-08, 
    2.520512e-08, 2.430302e-08, 2.201316e-08, 2.399014e-08, 2.077006e-08,
  2.529333e-08, 2.596274e-08, 2.639589e-08, 2.685702e-08, 2.691691e-08, 
    2.766331e-08, 2.724767e-08, 2.558312e-08, 2.378987e-08, 2.17669e-08, 
    2.156877e-08, 2.205001e-08, 2.451197e-08, 2.365137e-08, 1.98769e-08,
  2.51132e-08, 2.575511e-08, 2.586662e-08, 2.687913e-08, 2.826154e-08, 
    2.852985e-08, 2.718242e-08, 2.489864e-08, 2.301644e-08, 2.213244e-08, 
    2.241825e-08, 2.170504e-08, 2.50641e-08, 2.395243e-08, 2.095773e-08,
  2.561581e-08, 2.646195e-08, 2.689131e-08, 2.7859e-08, 2.936902e-08, 
    2.79661e-08, 2.554655e-08, 2.352327e-08, 2.301687e-08, 2.288242e-08, 
    2.360211e-08, 2.272198e-08, 2.537694e-08, 2.413676e-08, 2.265512e-08,
  2.632419e-08, 2.730853e-08, 2.747161e-08, 2.740109e-08, 2.785505e-08, 
    2.520179e-08, 2.300688e-08, 2.173128e-08, 2.245348e-08, 2.325394e-08, 
    2.355859e-08, 2.32632e-08, 2.553813e-08, 2.42387e-08, 2.349909e-08,
  2.637631e-08, 2.771754e-08, 2.69493e-08, 2.563129e-08, 2.454473e-08, 
    2.149161e-08, 2.04121e-08, 2.032975e-08, 2.263365e-08, 2.398116e-08, 
    2.393055e-08, 2.343087e-08, 2.436641e-08, 2.424871e-08, 2.293653e-08,
  2.620436e-08, 2.473198e-08, 2.26977e-08, 2.146197e-08, 2.07179e-08, 
    2.029294e-08, 1.983318e-08, 2.11516e-08, 2.476852e-08, 2.486306e-08, 
    2.449267e-08, 2.35049e-08, 2.335645e-08, 2.290913e-08, 2.353043e-08,
  1.932511e-08, 2.01399e-08, 2.055869e-08, 2.115975e-08, 2.204722e-08, 
    2.338029e-08, 2.401382e-08, 2.491336e-08, 2.519013e-08, 2.554669e-08, 
    2.664543e-08, 2.637801e-08, 2.549523e-08, 2.372748e-08, 2.161878e-08,
  1.974371e-08, 2.064876e-08, 2.106375e-08, 2.167939e-08, 2.238395e-08, 
    2.370637e-08, 2.453493e-08, 2.522242e-08, 2.533401e-08, 2.597028e-08, 
    2.667442e-08, 2.538307e-08, 2.452852e-08, 2.252395e-08, 2.184118e-08,
  1.971944e-08, 2.07757e-08, 2.182074e-08, 2.238111e-08, 2.319049e-08, 
    2.455685e-08, 2.537535e-08, 2.570481e-08, 2.600099e-08, 2.628762e-08, 
    2.572039e-08, 2.401787e-08, 2.31145e-08, 2.223458e-08, 2.4027e-08,
  2.024325e-08, 2.127824e-08, 2.199063e-08, 2.250792e-08, 2.32648e-08, 
    2.423914e-08, 2.500454e-08, 2.521806e-08, 2.566453e-08, 2.534258e-08, 
    2.333463e-08, 2.289549e-08, 2.284138e-08, 2.372737e-08, 2.601695e-08,
  2.055293e-08, 2.149602e-08, 2.212873e-08, 2.235874e-08, 2.309425e-08, 
    2.409165e-08, 2.420803e-08, 2.413535e-08, 2.428524e-08, 2.180207e-08, 
    2.23274e-08, 2.269112e-08, 2.292618e-08, 2.400854e-08, 2.530303e-08,
  2.120104e-08, 2.182828e-08, 2.190952e-08, 2.212027e-08, 2.251407e-08, 
    2.333806e-08, 2.311089e-08, 2.367761e-08, 2.167269e-08, 2.098483e-08, 
    2.213666e-08, 2.185547e-08, 2.456087e-08, 2.586427e-08, 2.682988e-08,
  2.150815e-08, 2.155198e-08, 2.173593e-08, 2.169569e-08, 2.243062e-08, 
    2.288636e-08, 2.271926e-08, 2.241013e-08, 2.10994e-08, 2.117954e-08, 
    2.249108e-08, 2.389422e-08, 2.834481e-08, 2.679945e-08, 2.754963e-08,
  2.104492e-08, 2.131963e-08, 2.139448e-08, 2.175779e-08, 2.266304e-08, 
    2.221265e-08, 2.207804e-08, 2.117345e-08, 2.053523e-08, 2.236138e-08, 
    2.465683e-08, 2.739545e-08, 2.855893e-08, 2.738399e-08, 2.3016e-08,
  2.061577e-08, 2.130984e-08, 2.115569e-08, 2.22258e-08, 2.259948e-08, 
    2.26459e-08, 2.309843e-08, 2.196477e-08, 2.293736e-08, 2.587324e-08, 
    2.695485e-08, 2.786214e-08, 2.506328e-08, 2.212191e-08, 1.917585e-08,
  2.040078e-08, 2.062265e-08, 2.120545e-08, 2.172093e-08, 2.234316e-08, 
    2.296691e-08, 2.360859e-08, 2.398848e-08, 2.585656e-08, 2.657353e-08, 
    2.635942e-08, 2.398798e-08, 2.012279e-08, 1.747338e-08, 1.765162e-08,
  2.024307e-08, 2.036981e-08, 2.053314e-08, 2.027458e-08, 2.067678e-08, 
    2.101547e-08, 2.137622e-08, 2.19633e-08, 2.19453e-08, 2.192737e-08, 
    2.175007e-08, 2.177196e-08, 2.227604e-08, 2.262438e-08, 2.25904e-08,
  2.005428e-08, 2.061152e-08, 2.026366e-08, 2.046578e-08, 2.106798e-08, 
    2.153665e-08, 2.173264e-08, 2.242078e-08, 2.238625e-08, 2.254511e-08, 
    2.215715e-08, 2.259157e-08, 2.305848e-08, 2.321229e-08, 2.293556e-08,
  2.005386e-08, 2.03384e-08, 2.037548e-08, 2.116422e-08, 2.178714e-08, 
    2.228206e-08, 2.224282e-08, 2.277723e-08, 2.292909e-08, 2.304661e-08, 
    2.25941e-08, 2.324479e-08, 2.354807e-08, 2.339405e-08, 2.331698e-08,
  2.058914e-08, 2.04596e-08, 2.067898e-08, 2.140297e-08, 2.198059e-08, 
    2.24585e-08, 2.262111e-08, 2.304259e-08, 2.324401e-08, 2.268396e-08, 
    2.283706e-08, 2.351883e-08, 2.442256e-08, 2.484243e-08, 2.387643e-08,
  2.090418e-08, 2.099453e-08, 2.16559e-08, 2.240544e-08, 2.299225e-08, 
    2.328626e-08, 2.316895e-08, 2.338352e-08, 2.249923e-08, 2.159989e-08, 
    2.213017e-08, 2.337404e-08, 2.46083e-08, 2.418183e-08, 2.282972e-08,
  2.124664e-08, 2.196669e-08, 2.229394e-08, 2.277673e-08, 2.307001e-08, 
    2.303198e-08, 2.3074e-08, 2.256212e-08, 2.203851e-08, 2.180449e-08, 
    2.319585e-08, 2.316889e-08, 2.509993e-08, 2.415585e-08, 2.596888e-08,
  2.156562e-08, 2.266038e-08, 2.321749e-08, 2.324071e-08, 2.356615e-08, 
    2.33823e-08, 2.310026e-08, 2.268504e-08, 2.287416e-08, 2.283592e-08, 
    2.367982e-08, 2.367392e-08, 2.572747e-08, 2.656618e-08, 2.696765e-08,
  2.292288e-08, 2.384372e-08, 2.363601e-08, 2.34055e-08, 2.34986e-08, 
    2.273757e-08, 2.277792e-08, 2.271793e-08, 2.30495e-08, 2.313145e-08, 
    2.397377e-08, 2.428461e-08, 2.627658e-08, 2.64039e-08, 2.491368e-08,
  2.396113e-08, 2.37054e-08, 2.311513e-08, 2.23142e-08, 2.173917e-08, 
    2.168544e-08, 2.241124e-08, 2.297454e-08, 2.323537e-08, 2.359582e-08, 
    2.421609e-08, 2.466104e-08, 2.464257e-08, 2.425018e-08, 2.297416e-08,
  2.38223e-08, 2.259451e-08, 2.200762e-08, 2.094711e-08, 2.082462e-08, 
    2.163543e-08, 2.249382e-08, 2.337655e-08, 2.372655e-08, 2.364115e-08, 
    2.436412e-08, 2.408955e-08, 2.379188e-08, 2.311144e-08, 2.307131e-08,
  2.373506e-08, 2.343318e-08, 2.284792e-08, 2.256234e-08, 2.256567e-08, 
    2.270576e-08, 2.229008e-08, 2.280591e-08, 2.271987e-08, 2.328061e-08, 
    2.411859e-08, 2.415394e-08, 2.392451e-08, 2.273889e-08, 2.200943e-08,
  2.266157e-08, 2.269501e-08, 2.272665e-08, 2.226925e-08, 2.238451e-08, 
    2.265167e-08, 2.225006e-08, 2.267457e-08, 2.343192e-08, 2.427758e-08, 
    2.471291e-08, 2.399832e-08, 2.270486e-08, 2.170115e-08, 2.17963e-08,
  2.291057e-08, 2.34217e-08, 2.337723e-08, 2.274455e-08, 2.270898e-08, 
    2.247647e-08, 2.220015e-08, 2.277117e-08, 2.447375e-08, 2.509738e-08, 
    2.42602e-08, 2.184677e-08, 2.165435e-08, 2.194565e-08, 2.274748e-08,
  2.295284e-08, 2.35407e-08, 2.33014e-08, 2.283266e-08, 2.218102e-08, 
    2.194341e-08, 2.219658e-08, 2.327751e-08, 2.454298e-08, 2.341024e-08, 
    2.196915e-08, 2.125079e-08, 2.216899e-08, 2.239472e-08, 2.467894e-08,
  2.244833e-08, 2.320349e-08, 2.309613e-08, 2.258322e-08, 2.214311e-08, 
    2.199116e-08, 2.25276e-08, 2.326549e-08, 2.26403e-08, 2.086887e-08, 
    2.062538e-08, 2.141467e-08, 2.235073e-08, 2.318511e-08, 2.494956e-08,
  2.308888e-08, 2.374219e-08, 2.325472e-08, 2.294005e-08, 2.263019e-08, 
    2.271047e-08, 2.306641e-08, 2.268424e-08, 2.126299e-08, 2.074165e-08, 
    2.091705e-08, 2.161477e-08, 2.309321e-08, 2.375646e-08, 2.387726e-08,
  2.391717e-08, 2.363412e-08, 2.390477e-08, 2.397944e-08, 2.361167e-08, 
    2.354266e-08, 2.298867e-08, 2.187596e-08, 2.10317e-08, 2.086063e-08, 
    2.174945e-08, 2.234502e-08, 2.334761e-08, 2.325033e-08, 2.357471e-08,
  2.393298e-08, 2.372986e-08, 2.429316e-08, 2.425067e-08, 2.386525e-08, 
    2.316646e-08, 2.201314e-08, 2.145398e-08, 2.093172e-08, 2.162079e-08, 
    2.247383e-08, 2.266972e-08, 2.340624e-08, 2.279886e-08, 2.274179e-08,
  2.364899e-08, 2.366243e-08, 2.398152e-08, 2.378751e-08, 2.303721e-08, 
    2.209231e-08, 2.126994e-08, 2.070381e-08, 2.149213e-08, 2.253039e-08, 
    2.282082e-08, 2.301759e-08, 2.364676e-08, 2.360625e-08, 2.328926e-08,
  2.33459e-08, 2.309252e-08, 2.32445e-08, 2.243514e-08, 2.2018e-08, 
    2.107491e-08, 2.055401e-08, 2.108125e-08, 2.222074e-08, 2.282136e-08, 
    2.335607e-08, 2.360126e-08, 2.420325e-08, 2.4027e-08, 2.390404e-08,
  2.452264e-08, 2.453941e-08, 2.416255e-08, 2.411375e-08, 2.437777e-08, 
    2.477002e-08, 2.540473e-08, 2.505083e-08, 2.495662e-08, 2.483664e-08, 
    2.466271e-08, 2.36365e-08, 2.2974e-08, 2.256045e-08, 2.177639e-08,
  2.437365e-08, 2.405644e-08, 2.416513e-08, 2.401957e-08, 2.405814e-08, 
    2.432603e-08, 2.506126e-08, 2.480985e-08, 2.510109e-08, 2.448487e-08, 
    2.418124e-08, 2.356004e-08, 2.300992e-08, 2.260908e-08, 2.207846e-08,
  2.317554e-08, 2.368822e-08, 2.397906e-08, 2.423706e-08, 2.458843e-08, 
    2.511947e-08, 2.557024e-08, 2.51274e-08, 2.526594e-08, 2.459013e-08, 
    2.460947e-08, 2.381927e-08, 2.341457e-08, 2.297877e-08, 2.231887e-08,
  2.404616e-08, 2.405395e-08, 2.430261e-08, 2.461781e-08, 2.488034e-08, 
    2.489859e-08, 2.545446e-08, 2.526529e-08, 2.523547e-08, 2.491153e-08, 
    2.461443e-08, 2.406311e-08, 2.307242e-08, 2.228095e-08, 2.271031e-08,
  2.394468e-08, 2.422216e-08, 2.493659e-08, 2.508681e-08, 2.476556e-08, 
    2.49325e-08, 2.546319e-08, 2.543348e-08, 2.541841e-08, 2.449017e-08, 
    2.449483e-08, 2.353416e-08, 2.204922e-08, 2.226282e-08, 2.338119e-08,
  2.428795e-08, 2.502556e-08, 2.49709e-08, 2.448478e-08, 2.422342e-08, 
    2.448418e-08, 2.466138e-08, 2.489115e-08, 2.428152e-08, 2.457617e-08, 
    2.362722e-08, 2.236811e-08, 2.179931e-08, 2.268489e-08, 2.329044e-08,
  2.432923e-08, 2.485361e-08, 2.44441e-08, 2.416119e-08, 2.413851e-08, 
    2.424128e-08, 2.451471e-08, 2.45454e-08, 2.416256e-08, 2.360857e-08, 
    2.293922e-08, 2.238455e-08, 2.223882e-08, 2.288177e-08, 2.348973e-08,
  2.404839e-08, 2.458002e-08, 2.43796e-08, 2.416462e-08, 2.410019e-08, 
    2.432298e-08, 2.450279e-08, 2.445491e-08, 2.335526e-08, 2.305871e-08, 
    2.289786e-08, 2.241559e-08, 2.268489e-08, 2.303078e-08, 2.345902e-08,
  2.355855e-08, 2.407801e-08, 2.405178e-08, 2.392252e-08, 2.406684e-08, 
    2.440393e-08, 2.433754e-08, 2.391078e-08, 2.349793e-08, 2.359146e-08, 
    2.299611e-08, 2.266748e-08, 2.322289e-08, 2.405044e-08, 2.475043e-08,
  2.324341e-08, 2.351314e-08, 2.377137e-08, 2.328543e-08, 2.346049e-08, 
    2.400088e-08, 2.3933e-08, 2.421734e-08, 2.431563e-08, 2.374597e-08, 
    2.297288e-08, 2.320349e-08, 2.399244e-08, 2.485018e-08, 2.534099e-08,
  2.496168e-08, 2.56034e-08, 2.575963e-08, 2.474922e-08, 2.392894e-08, 
    2.224612e-08, 2.179438e-08, 2.140258e-08, 2.211968e-08, 2.293768e-08, 
    2.298479e-08, 2.320152e-08, 2.412011e-08, 2.370654e-08, 2.315264e-08,
  2.47548e-08, 2.509094e-08, 2.520188e-08, 2.469089e-08, 2.344157e-08, 
    2.208226e-08, 2.171446e-08, 2.143622e-08, 2.207501e-08, 2.248253e-08, 
    2.245287e-08, 2.310156e-08, 2.387716e-08, 2.342974e-08, 2.321773e-08,
  2.374363e-08, 2.305233e-08, 2.377669e-08, 2.383998e-08, 2.34122e-08, 
    2.210974e-08, 2.142383e-08, 2.134844e-08, 2.21186e-08, 2.174077e-08, 
    2.236592e-08, 2.32898e-08, 2.376393e-08, 2.322687e-08, 2.351649e-08,
  2.309328e-08, 2.302817e-08, 2.32483e-08, 2.340068e-08, 2.269507e-08, 
    2.170837e-08, 2.147014e-08, 2.132826e-08, 2.172649e-08, 2.10687e-08, 
    2.275635e-08, 2.33694e-08, 2.367765e-08, 2.378381e-08, 2.444414e-08,
  2.317953e-08, 2.284244e-08, 2.30428e-08, 2.253549e-08, 2.203594e-08, 
    2.152337e-08, 2.137367e-08, 2.123024e-08, 2.095171e-08, 2.054044e-08, 
    2.186756e-08, 2.322459e-08, 2.359702e-08, 2.365121e-08, 2.511928e-08,
  2.262646e-08, 2.293079e-08, 2.256085e-08, 2.221147e-08, 2.165108e-08, 
    2.109673e-08, 2.109536e-08, 2.087549e-08, 2.03791e-08, 2.10282e-08, 
    2.266149e-08, 2.279296e-08, 2.345362e-08, 2.484584e-08, 2.593441e-08,
  2.197824e-08, 2.196177e-08, 2.191442e-08, 2.20289e-08, 2.153647e-08, 
    2.09982e-08, 2.092679e-08, 2.050132e-08, 2.068784e-08, 2.194658e-08, 
    2.280955e-08, 2.284395e-08, 2.384487e-08, 2.524062e-08, 2.514331e-08,
  2.1456e-08, 2.146399e-08, 2.152957e-08, 2.154276e-08, 2.115556e-08, 
    2.101951e-08, 2.10156e-08, 2.061819e-08, 2.094938e-08, 2.195412e-08, 
    2.262079e-08, 2.284051e-08, 2.403276e-08, 2.451534e-08, 2.417567e-08,
  2.127968e-08, 2.140046e-08, 2.132771e-08, 2.131456e-08, 2.084328e-08, 
    2.118237e-08, 2.113845e-08, 2.064616e-08, 2.117148e-08, 2.221718e-08, 
    2.267032e-08, 2.294435e-08, 2.37456e-08, 2.388588e-08, 2.436293e-08,
  2.170517e-08, 2.124686e-08, 2.088845e-08, 2.056332e-08, 2.032998e-08, 
    2.039425e-08, 2.022611e-08, 2.064775e-08, 2.173638e-08, 2.227091e-08, 
    2.259536e-08, 2.309323e-08, 2.332815e-08, 2.362812e-08, 2.586638e-08,
  2.301074e-08, 2.41806e-08, 2.453791e-08, 2.494807e-08, 2.600332e-08, 
    2.772728e-08, 2.722055e-08, 2.813791e-08, 2.903546e-08, 2.524742e-08, 
    2.145486e-08, 2.046709e-08, 2.208071e-08, 2.251739e-08, 2.12744e-08,
  2.497942e-08, 2.5666e-08, 2.592272e-08, 2.695482e-08, 2.886042e-08, 
    2.876499e-08, 2.760223e-08, 2.889417e-08, 2.881855e-08, 2.43898e-08, 
    2.219729e-08, 2.145356e-08, 2.253494e-08, 2.196611e-08, 2.075426e-08,
  2.786587e-08, 2.925515e-08, 2.830139e-08, 3.056076e-08, 3.048902e-08, 
    2.877754e-08, 2.715861e-08, 2.817742e-08, 2.667372e-08, 2.371785e-08, 
    2.289598e-08, 2.164244e-08, 2.276424e-08, 2.193076e-08, 2.290886e-08,
  3.037656e-08, 3.15993e-08, 3.025612e-08, 3.047569e-08, 2.839509e-08, 
    2.641074e-08, 2.615458e-08, 2.561304e-08, 2.472177e-08, 2.219571e-08, 
    2.002712e-08, 1.989327e-08, 2.207661e-08, 2.177049e-08, 2.577748e-08,
  2.927051e-08, 2.816413e-08, 2.910158e-08, 2.699344e-08, 2.598188e-08, 
    2.508667e-08, 2.404127e-08, 2.344328e-08, 2.269757e-08, 1.960305e-08, 
    1.934892e-08, 2.078771e-08, 2.226228e-08, 2.364683e-08, 2.70384e-08,
  2.923865e-08, 2.684886e-08, 2.881399e-08, 2.732948e-08, 2.560692e-08, 
    2.401555e-08, 2.274151e-08, 2.319694e-08, 2.27456e-08, 2.053787e-08, 
    2.10244e-08, 2.157022e-08, 2.394559e-08, 2.539928e-08, 2.488903e-08,
  2.901391e-08, 2.93977e-08, 2.933018e-08, 2.815015e-08, 2.579596e-08, 
    2.386754e-08, 2.434889e-08, 2.52153e-08, 2.447012e-08, 2.150521e-08, 
    2.146453e-08, 2.183576e-08, 2.49216e-08, 2.624412e-08, 2.355335e-08,
  2.944042e-08, 3.098296e-08, 2.882848e-08, 2.598735e-08, 2.373745e-08, 
    2.368554e-08, 2.447329e-08, 2.496614e-08, 2.232496e-08, 2.007511e-08, 
    2.091248e-08, 2.202692e-08, 2.452638e-08, 2.421117e-08, 2.269885e-08,
  2.372598e-08, 2.58331e-08, 2.370449e-08, 2.186886e-08, 2.173384e-08, 
    2.187142e-08, 2.266961e-08, 2.141979e-08, 1.98793e-08, 2.028558e-08, 
    2.120224e-08, 2.296304e-08, 2.37545e-08, 2.25284e-08, 2.36085e-08,
  1.76429e-08, 1.778308e-08, 1.662812e-08, 1.57122e-08, 1.684323e-08, 
    1.781426e-08, 1.86317e-08, 1.891453e-08, 2.041475e-08, 2.079286e-08, 
    2.126658e-08, 2.306973e-08, 2.337069e-08, 2.259353e-08, 2.505976e-08,
  1.74031e-08, 1.943451e-08, 2.057628e-08, 2.259958e-08, 2.562475e-08, 
    2.689793e-08, 2.625677e-08, 2.718329e-08, 2.556478e-08, 2.420971e-08, 
    2.129678e-08, 1.866007e-08, 1.933365e-08, 1.879079e-08, 1.773742e-08,
  1.857986e-08, 1.9573e-08, 2.120323e-08, 2.341735e-08, 2.536351e-08, 
    2.601104e-08, 2.625647e-08, 2.695604e-08, 2.593714e-08, 2.524269e-08, 
    2.107869e-08, 1.922774e-08, 1.85894e-08, 1.725274e-08, 1.724483e-08,
  1.857598e-08, 2.063471e-08, 2.222501e-08, 2.467363e-08, 2.578509e-08, 
    2.641728e-08, 2.714977e-08, 2.695996e-08, 2.671023e-08, 2.47452e-08, 
    1.986059e-08, 1.822485e-08, 1.811849e-08, 1.769503e-08, 2.127525e-08,
  1.965234e-08, 2.134424e-08, 2.276969e-08, 2.428178e-08, 2.556702e-08, 
    2.650445e-08, 2.761756e-08, 2.670928e-08, 2.508013e-08, 2.05513e-08, 
    1.616933e-08, 1.594457e-08, 1.721351e-08, 1.732641e-08, 2.408556e-08,
  1.955851e-08, 2.132717e-08, 2.274553e-08, 2.41112e-08, 2.531857e-08, 
    2.57977e-08, 2.574865e-08, 2.439818e-08, 2.134318e-08, 1.538347e-08, 
    1.522876e-08, 1.657338e-08, 1.653598e-08, 1.842904e-08, 2.575762e-08,
  2.131366e-08, 2.292147e-08, 2.37683e-08, 2.583953e-08, 2.638893e-08, 
    2.597451e-08, 2.47555e-08, 2.243956e-08, 1.707176e-08, 1.586728e-08, 
    1.727545e-08, 1.727404e-08, 1.796347e-08, 2.128131e-08, 2.427476e-08,
  2.17622e-08, 2.364139e-08, 2.550753e-08, 2.663242e-08, 2.68174e-08, 
    2.6095e-08, 2.427054e-08, 2.024944e-08, 1.765814e-08, 1.740464e-08, 
    1.666037e-08, 1.729442e-08, 1.930526e-08, 2.25845e-08, 2.2792e-08,
  2.265428e-08, 2.54809e-08, 2.626497e-08, 2.640369e-08, 2.71185e-08, 
    2.638549e-08, 2.350126e-08, 2.036548e-08, 1.742051e-08, 1.617627e-08, 
    1.619409e-08, 1.842211e-08, 2.064e-08, 2.278768e-08, 2.225594e-08,
  2.31702e-08, 2.51867e-08, 2.455924e-08, 2.380802e-08, 2.348805e-08, 
    2.205037e-08, 1.848407e-08, 1.650867e-08, 1.52436e-08, 1.59267e-08, 
    1.751916e-08, 1.996803e-08, 2.136937e-08, 2.164621e-08, 2.27461e-08,
  2.338225e-08, 2.22486e-08, 2.04711e-08, 1.869487e-08, 1.811098e-08, 
    1.619219e-08, 1.534191e-08, 1.479959e-08, 1.653259e-08, 1.812094e-08, 
    2.01202e-08, 2.11992e-08, 2.213044e-08, 2.239122e-08, 2.358541e-08,
  2.257166e-08, 2.304049e-08, 2.272212e-08, 2.291571e-08, 2.268662e-08, 
    2.235821e-08, 2.171474e-08, 2.128971e-08, 2.083519e-08, 2.031588e-08, 
    2.073222e-08, 2.119896e-08, 2.118968e-08, 2.062477e-08, 1.897816e-08,
  2.376938e-08, 2.405408e-08, 2.365322e-08, 2.375071e-08, 2.266914e-08, 
    2.22618e-08, 2.111231e-08, 2.114641e-08, 2.035314e-08, 2.090983e-08, 
    2.135024e-08, 2.170063e-08, 2.143372e-08, 2.020109e-08, 1.859014e-08,
  2.538182e-08, 2.476797e-08, 2.365973e-08, 2.318273e-08, 2.214495e-08, 
    2.192697e-08, 2.112419e-08, 2.140637e-08, 2.083144e-08, 2.152786e-08, 
    2.176625e-08, 2.150938e-08, 2.104642e-08, 1.987445e-08, 1.871154e-08,
  2.620832e-08, 2.458276e-08, 2.377572e-08, 2.291544e-08, 2.205448e-08, 
    2.184548e-08, 2.18469e-08, 2.181025e-08, 2.135039e-08, 2.168623e-08, 
    2.057712e-08, 1.943359e-08, 2.009873e-08, 1.935952e-08, 1.910576e-08,
  2.534726e-08, 2.379053e-08, 2.304283e-08, 2.209624e-08, 2.200332e-08, 
    2.146304e-08, 2.176943e-08, 2.17148e-08, 2.206943e-08, 2.042717e-08, 
    1.997513e-08, 1.914506e-08, 1.806339e-08, 1.753285e-08, 1.885573e-08,
  2.460923e-08, 2.378911e-08, 2.350487e-08, 2.254669e-08, 2.17697e-08, 
    2.095873e-08, 2.087516e-08, 2.123743e-08, 2.010386e-08, 1.904e-08, 
    2.077705e-08, 2.007133e-08, 1.773613e-08, 1.620553e-08, 1.844623e-08,
  2.401764e-08, 2.384903e-08, 2.304404e-08, 2.128871e-08, 2.08636e-08, 
    2.070536e-08, 2.110998e-08, 2.035445e-08, 2.025578e-08, 1.976276e-08, 
    1.936386e-08, 1.833146e-08, 1.69707e-08, 1.673398e-08, 1.771676e-08,
  2.327623e-08, 2.267106e-08, 2.106598e-08, 2.082113e-08, 2.113891e-08, 
    2.206208e-08, 2.220679e-08, 2.118593e-08, 2.136517e-08, 1.979292e-08, 
    1.837384e-08, 1.781484e-08, 1.613548e-08, 1.650349e-08, 1.757731e-08,
  2.264257e-08, 2.113121e-08, 2.073851e-08, 2.112059e-08, 2.173313e-08, 
    2.251868e-08, 2.242501e-08, 2.160809e-08, 2.029814e-08, 1.97284e-08, 
    1.942303e-08, 1.839221e-08, 1.751197e-08, 1.741624e-08, 1.783258e-08,
  2.158534e-08, 2.125705e-08, 2.135348e-08, 2.177139e-08, 2.226647e-08, 
    2.228781e-08, 2.208055e-08, 2.169617e-08, 2.135557e-08, 2.048343e-08, 
    2.051515e-08, 1.963071e-08, 1.97105e-08, 1.931311e-08, 2.005211e-08,
  2.616238e-08, 2.529702e-08, 2.440806e-08, 2.414176e-08, 2.456049e-08, 
    2.486978e-08, 2.459833e-08, 2.474653e-08, 2.48678e-08, 2.445291e-08, 
    2.485063e-08, 2.509031e-08, 2.5177e-08, 2.568101e-08, 2.485327e-08,
  2.643954e-08, 2.43892e-08, 2.392212e-08, 2.406294e-08, 2.507314e-08, 
    2.519321e-08, 2.499265e-08, 2.537024e-08, 2.50445e-08, 2.493604e-08, 
    2.449743e-08, 2.459231e-08, 2.491282e-08, 2.565676e-08, 2.406827e-08,
  2.597143e-08, 2.423743e-08, 2.42618e-08, 2.484405e-08, 2.557783e-08, 
    2.505032e-08, 2.453119e-08, 2.474251e-08, 2.454592e-08, 2.470243e-08, 
    2.450946e-08, 2.460397e-08, 2.461799e-08, 2.496554e-08, 2.382616e-08,
  2.534197e-08, 2.411812e-08, 2.512415e-08, 2.562117e-08, 2.528894e-08, 
    2.474875e-08, 2.491835e-08, 2.507296e-08, 2.447739e-08, 2.43575e-08, 
    2.483861e-08, 2.459221e-08, 2.590076e-08, 2.559046e-08, 2.38089e-08,
  2.458119e-08, 2.504684e-08, 2.52059e-08, 2.486435e-08, 2.475461e-08, 
    2.474375e-08, 2.526478e-08, 2.457781e-08, 2.464043e-08, 2.612447e-08, 
    2.390742e-08, 2.427184e-08, 2.437354e-08, 2.331662e-08, 2.2704e-08,
  2.52596e-08, 2.517134e-08, 2.483537e-08, 2.500546e-08, 2.554235e-08, 
    2.584269e-08, 2.516309e-08, 2.448079e-08, 2.517596e-08, 2.367272e-08, 
    2.281873e-08, 2.322287e-08, 2.318889e-08, 1.896833e-08, 2.213697e-08,
  2.446011e-08, 2.516351e-08, 2.524456e-08, 2.577043e-08, 2.625861e-08, 
    2.595915e-08, 2.484738e-08, 2.426877e-08, 2.402304e-08, 2.301399e-08, 
    2.263156e-08, 2.210871e-08, 2.179327e-08, 1.873907e-08, 2.469067e-08,
  2.485751e-08, 2.543757e-08, 2.603705e-08, 2.665813e-08, 2.692993e-08, 
    2.626408e-08, 2.531776e-08, 2.498709e-08, 2.42494e-08, 2.396466e-08, 
    2.338502e-08, 2.268832e-08, 2.10256e-08, 2.073535e-08, 2.415151e-08,
  2.492616e-08, 2.552583e-08, 2.710644e-08, 2.743624e-08, 2.730463e-08, 
    2.627909e-08, 2.497704e-08, 2.466175e-08, 2.396841e-08, 2.369956e-08, 
    2.40546e-08, 2.375504e-08, 2.298344e-08, 2.313091e-08, 2.281329e-08,
  2.52273e-08, 2.677941e-08, 2.816547e-08, 2.775229e-08, 2.683559e-08, 
    2.511527e-08, 2.383758e-08, 2.372888e-08, 2.438208e-08, 2.444749e-08, 
    2.471561e-08, 2.385804e-08, 2.412568e-08, 2.414397e-08, 2.179561e-08,
  2.560115e-08, 2.563015e-08, 2.488241e-08, 2.516383e-08, 2.549032e-08, 
    2.555909e-08, 2.505627e-08, 2.57076e-08, 2.595354e-08, 2.532897e-08, 
    2.506751e-08, 2.53701e-08, 2.54648e-08, 2.543807e-08, 2.514569e-08,
  2.701674e-08, 2.558543e-08, 2.443077e-08, 2.483113e-08, 2.609703e-08, 
    2.584226e-08, 2.550544e-08, 2.620119e-08, 2.640381e-08, 2.633332e-08, 
    2.583649e-08, 2.605108e-08, 2.578252e-08, 2.568224e-08, 2.478047e-08,
  2.904093e-08, 2.479647e-08, 2.454017e-08, 2.572529e-08, 2.642758e-08, 
    2.625471e-08, 2.604058e-08, 2.63754e-08, 2.699419e-08, 2.67583e-08, 
    2.688607e-08, 2.667561e-08, 2.602601e-08, 2.594807e-08, 2.52354e-08,
  2.472703e-08, 2.272635e-08, 2.403524e-08, 2.538195e-08, 2.532951e-08, 
    2.569825e-08, 2.637474e-08, 2.672387e-08, 2.687511e-08, 2.734574e-08, 
    2.717843e-08, 2.644143e-08, 2.613818e-08, 2.605293e-08, 2.541105e-08,
  2.417889e-08, 2.328816e-08, 2.415911e-08, 2.44863e-08, 2.493605e-08, 
    2.543149e-08, 2.612554e-08, 2.642337e-08, 2.652999e-08, 2.613879e-08, 
    2.548978e-08, 2.601509e-08, 2.620258e-08, 2.582167e-08, 2.487637e-08,
  2.424803e-08, 2.401815e-08, 2.450361e-08, 2.530134e-08, 2.612662e-08, 
    2.62072e-08, 2.633764e-08, 2.657536e-08, 2.600328e-08, 2.60327e-08, 
    2.716074e-08, 2.695594e-08, 2.686162e-08, 2.512451e-08, 2.610625e-08,
  2.362554e-08, 2.421832e-08, 2.525343e-08, 2.589181e-08, 2.60952e-08, 
    2.618457e-08, 2.594046e-08, 2.630073e-08, 2.596692e-08, 2.6534e-08, 
    2.650542e-08, 2.615562e-08, 2.608278e-08, 2.389425e-08, 2.665656e-08,
  2.405967e-08, 2.521993e-08, 2.558949e-08, 2.605722e-08, 2.586378e-08, 
    2.590749e-08, 2.563478e-08, 2.606525e-08, 2.56083e-08, 2.539133e-08, 
    2.524512e-08, 2.517415e-08, 2.503493e-08, 2.502606e-08, 2.707767e-08,
  2.480715e-08, 2.548537e-08, 2.604854e-08, 2.605042e-08, 2.558065e-08, 
    2.570457e-08, 2.559211e-08, 2.570466e-08, 2.460518e-08, 2.531435e-08, 
    2.507217e-08, 2.491393e-08, 2.502459e-08, 2.512287e-08, 2.56962e-08,
  2.525752e-08, 2.577902e-08, 2.632019e-08, 2.546762e-08, 2.510699e-08, 
    2.449992e-08, 2.465663e-08, 2.514252e-08, 2.587878e-08, 2.590276e-08, 
    2.572514e-08, 2.505728e-08, 2.507813e-08, 2.516342e-08, 2.480974e-08,
  2.46161e-08, 2.477801e-08, 2.51704e-08, 2.565564e-08, 2.568067e-08, 
    2.570429e-08, 2.552696e-08, 2.52711e-08, 2.471294e-08, 2.201516e-08, 
    2.070948e-08, 2.152411e-08, 2.269082e-08, 2.191813e-08, 2.166087e-08,
  2.528196e-08, 2.491378e-08, 2.503383e-08, 2.582842e-08, 2.608386e-08, 
    2.585958e-08, 2.479115e-08, 2.465001e-08, 2.429124e-08, 2.286353e-08, 
    2.16208e-08, 2.053059e-08, 2.114602e-08, 1.996606e-08, 1.98107e-08,
  2.852749e-08, 2.556247e-08, 2.558053e-08, 2.600187e-08, 2.61345e-08, 
    2.520241e-08, 2.425538e-08, 2.444545e-08, 2.477881e-08, 2.373687e-08, 
    2.366242e-08, 2.276544e-08, 2.257474e-08, 2.116816e-08, 2.179915e-08,
  2.63574e-08, 2.478524e-08, 2.565789e-08, 2.567192e-08, 2.518049e-08, 
    2.457957e-08, 2.454198e-08, 2.505405e-08, 2.473996e-08, 2.501892e-08, 
    2.382804e-08, 2.324661e-08, 2.425902e-08, 2.371457e-08, 2.4865e-08,
  2.613699e-08, 2.542831e-08, 2.554044e-08, 2.529231e-08, 2.463515e-08, 
    2.439001e-08, 2.473252e-08, 2.515639e-08, 2.538756e-08, 2.4437e-08, 
    2.300393e-08, 2.392983e-08, 2.382962e-08, 2.442722e-08, 2.520373e-08,
  2.499938e-08, 2.524251e-08, 2.504891e-08, 2.549368e-08, 2.540873e-08, 
    2.535148e-08, 2.570168e-08, 2.527276e-08, 2.462691e-08, 2.298238e-08, 
    2.532134e-08, 2.515389e-08, 2.45178e-08, 2.373134e-08, 2.628762e-08,
  2.43277e-08, 2.526891e-08, 2.517614e-08, 2.529776e-08, 2.540756e-08, 
    2.567679e-08, 2.539934e-08, 2.451397e-08, 2.421987e-08, 2.409158e-08, 
    2.413391e-08, 2.342494e-08, 2.365763e-08, 2.345865e-08, 2.600289e-08,
  2.378219e-08, 2.531979e-08, 2.512948e-08, 2.541318e-08, 2.558028e-08, 
    2.562969e-08, 2.501509e-08, 2.444597e-08, 2.445035e-08, 2.356414e-08, 
    2.327883e-08, 2.282299e-08, 2.297123e-08, 2.31898e-08, 2.456941e-08,
  2.413743e-08, 2.553521e-08, 2.530528e-08, 2.50411e-08, 2.548616e-08, 
    2.53384e-08, 2.429075e-08, 2.478586e-08, 2.401219e-08, 2.428494e-08, 
    2.425644e-08, 2.369765e-08, 2.433611e-08, 2.471137e-08, 2.388453e-08,
  2.42812e-08, 2.53969e-08, 2.446442e-08, 2.398188e-08, 2.504787e-08, 
    2.534633e-08, 2.502387e-08, 2.443152e-08, 2.436083e-08, 2.443177e-08, 
    2.470608e-08, 2.403369e-08, 2.538668e-08, 2.591587e-08, 2.592049e-08,
  2.108769e-08, 2.081222e-08, 2.074545e-08, 2.281582e-08, 2.311148e-08, 
    2.44367e-08, 2.617279e-08, 2.831884e-08, 2.691908e-08, 2.494419e-08, 
    2.353688e-08, 2.428732e-08, 2.429884e-08, 2.383502e-08, 2.404082e-08,
  2.2414e-08, 2.180807e-08, 2.183531e-08, 2.382031e-08, 2.451834e-08, 
    2.563768e-08, 2.66039e-08, 2.816971e-08, 2.655959e-08, 2.460585e-08, 
    2.493731e-08, 2.477739e-08, 2.447556e-08, 2.401731e-08, 2.381883e-08,
  2.385067e-08, 2.197614e-08, 2.268615e-08, 2.501955e-08, 2.54293e-08, 
    2.487406e-08, 2.631798e-08, 2.778977e-08, 2.534417e-08, 2.56746e-08, 
    2.605678e-08, 2.487915e-08, 2.441113e-08, 2.419912e-08, 2.410239e-08,
  2.21725e-08, 2.086007e-08, 2.232971e-08, 2.345783e-08, 2.374223e-08, 
    2.453369e-08, 2.634217e-08, 2.671685e-08, 2.560181e-08, 2.619391e-08, 
    2.415476e-08, 2.275732e-08, 2.442526e-08, 2.436112e-08, 2.405118e-08,
  2.178633e-08, 2.079058e-08, 2.134605e-08, 2.233515e-08, 2.343055e-08, 
    2.398985e-08, 2.52472e-08, 2.535063e-08, 2.488603e-08, 2.407143e-08, 
    2.310605e-08, 2.412162e-08, 2.603776e-08, 2.441429e-08, 2.52192e-08,
  2.127316e-08, 2.062058e-08, 2.082623e-08, 2.150355e-08, 2.330003e-08, 
    2.39837e-08, 2.518253e-08, 2.537396e-08, 2.435486e-08, 2.37989e-08, 
    2.428635e-08, 2.38743e-08, 2.539917e-08, 2.193018e-08, 2.568467e-08,
  2.064273e-08, 2.076893e-08, 2.100408e-08, 2.131054e-08, 2.314307e-08, 
    2.360242e-08, 2.438422e-08, 2.493049e-08, 2.42926e-08, 2.45515e-08, 
    2.403015e-08, 2.370381e-08, 2.387593e-08, 2.219863e-08, 2.649002e-08,
  2.100136e-08, 2.100534e-08, 2.073307e-08, 2.091085e-08, 2.311903e-08, 
    2.377534e-08, 2.5054e-08, 2.483144e-08, 2.437036e-08, 2.479344e-08, 
    2.426135e-08, 2.369341e-08, 2.373731e-08, 2.64916e-08, 2.624303e-08,
  2.129871e-08, 2.108921e-08, 2.062312e-08, 2.091544e-08, 2.27991e-08, 
    2.303872e-08, 2.361522e-08, 2.407643e-08, 2.413228e-08, 2.508023e-08, 
    2.431553e-08, 2.354917e-08, 2.413407e-08, 2.5051e-08, 2.658978e-08,
  2.165109e-08, 2.11055e-08, 2.030074e-08, 2.029292e-08, 2.149526e-08, 
    2.196637e-08, 2.334338e-08, 2.382119e-08, 2.453808e-08, 2.545918e-08, 
    2.478054e-08, 2.361004e-08, 2.409857e-08, 2.523167e-08, 2.633922e-08,
  2.261413e-08, 2.34425e-08, 2.426108e-08, 2.532067e-08, 2.948491e-08, 
    3.204188e-08, 2.864358e-08, 2.624732e-08, 2.66255e-08, 2.518009e-08, 
    2.578886e-08, 2.676088e-08, 2.580114e-08, 2.386309e-08, 2.409263e-08,
  2.406261e-08, 2.532904e-08, 2.497141e-08, 2.837403e-08, 3.26787e-08, 
    3.170924e-08, 2.562297e-08, 2.586168e-08, 2.69999e-08, 2.641551e-08, 
    2.708725e-08, 2.690596e-08, 2.4385e-08, 2.339817e-08, 2.478737e-08,
  2.592989e-08, 2.640722e-08, 2.638328e-08, 3.235458e-08, 3.182356e-08, 
    2.752575e-08, 2.362933e-08, 2.509134e-08, 2.710425e-08, 2.643645e-08, 
    2.831709e-08, 2.596087e-08, 2.394406e-08, 2.426711e-08, 2.521891e-08,
  2.176957e-08, 2.246858e-08, 2.492634e-08, 2.755479e-08, 2.639961e-08, 
    2.490904e-08, 2.299585e-08, 2.412861e-08, 2.675492e-08, 2.637069e-08, 
    2.618455e-08, 2.458733e-08, 2.464776e-08, 2.596892e-08, 2.494633e-08,
  2.020316e-08, 2.158673e-08, 2.299184e-08, 2.456659e-08, 2.573362e-08, 
    2.417855e-08, 2.270675e-08, 2.402665e-08, 2.42045e-08, 2.22819e-08, 
    2.277121e-08, 2.507852e-08, 2.700765e-08, 2.436031e-08, 2.410116e-08,
  2.087949e-08, 2.169439e-08, 2.24835e-08, 2.387057e-08, 2.572849e-08, 
    2.333548e-08, 2.215856e-08, 2.359816e-08, 2.228274e-08, 2.234328e-08, 
    2.4907e-08, 2.47313e-08, 2.604908e-08, 2.307394e-08, 2.459496e-08,
  2.142256e-08, 2.16008e-08, 2.312643e-08, 2.506069e-08, 2.651048e-08, 
    2.379027e-08, 2.192514e-08, 2.311694e-08, 2.315096e-08, 2.385728e-08, 
    2.542176e-08, 2.496592e-08, 2.402306e-08, 2.288162e-08, 2.387703e-08,
  2.14574e-08, 2.208049e-08, 2.360146e-08, 2.554059e-08, 2.785677e-08, 
    2.44287e-08, 2.215423e-08, 2.316599e-08, 2.296562e-08, 2.377396e-08, 
    2.522889e-08, 2.503935e-08, 2.361108e-08, 2.500407e-08, 2.426201e-08,
  2.236652e-08, 2.274769e-08, 2.424356e-08, 2.582106e-08, 2.813429e-08, 
    2.471381e-08, 2.148299e-08, 2.15551e-08, 2.252228e-08, 2.410271e-08, 
    2.525878e-08, 2.538213e-08, 2.406772e-08, 2.346859e-08, 2.349021e-08,
  2.305775e-08, 2.331394e-08, 2.434156e-08, 2.484909e-08, 2.620937e-08, 
    2.423916e-08, 2.185671e-08, 2.154579e-08, 2.322713e-08, 2.423941e-08, 
    2.468206e-08, 2.52723e-08, 2.464907e-08, 2.347717e-08, 2.21041e-08,
  2.189427e-08, 2.238341e-08, 2.23969e-08, 2.232848e-08, 2.119851e-08, 
    2.069821e-08, 2.044285e-08, 2.055494e-08, 2.08815e-08, 2.173619e-08, 
    2.238069e-08, 2.476708e-08, 2.650918e-08, 2.461829e-08, 2.300308e-08,
  2.212285e-08, 2.177304e-08, 2.179958e-08, 2.182809e-08, 2.058578e-08, 
    2.02333e-08, 2.029487e-08, 2.006127e-08, 2.083589e-08, 2.357529e-08, 
    2.515659e-08, 2.613819e-08, 2.578343e-08, 2.294072e-08, 2.14562e-08,
  2.213346e-08, 2.211434e-08, 2.224555e-08, 2.123655e-08, 2.026202e-08, 
    2.04485e-08, 1.999545e-08, 2.023102e-08, 2.260418e-08, 2.446017e-08, 
    2.568993e-08, 2.545196e-08, 2.408705e-08, 2.240918e-08, 2.196715e-08,
  2.235465e-08, 2.306972e-08, 2.301848e-08, 2.31414e-08, 2.295231e-08, 
    2.170355e-08, 2.117365e-08, 2.126454e-08, 2.313929e-08, 2.334872e-08, 
    2.067402e-08, 1.998831e-08, 2.102928e-08, 2.202998e-08, 2.494576e-08,
  2.220646e-08, 2.291218e-08, 2.291903e-08, 2.283362e-08, 2.232386e-08, 
    2.145315e-08, 2.07774e-08, 2.131823e-08, 2.14309e-08, 1.972428e-08, 
    1.920927e-08, 2.08644e-08, 2.227956e-08, 2.428054e-08, 2.627786e-08,
  2.343411e-08, 2.40964e-08, 2.380161e-08, 2.297968e-08, 2.149065e-08, 
    2.063464e-08, 2.046442e-08, 2.049826e-08, 2.039841e-08, 2.17947e-08, 
    2.415791e-08, 2.367771e-08, 2.453938e-08, 2.611715e-08, 2.472988e-08,
  2.389553e-08, 2.369589e-08, 2.348911e-08, 2.205319e-08, 2.063886e-08, 
    2.029301e-08, 2.053153e-08, 2.091849e-08, 2.246687e-08, 2.540488e-08, 
    2.516877e-08, 2.39406e-08, 2.525847e-08, 2.464853e-08, 2.147525e-08,
  2.326831e-08, 2.301399e-08, 2.343948e-08, 2.189089e-08, 2.024631e-08, 
    2.034321e-08, 2.05773e-08, 2.212013e-08, 2.412606e-08, 2.490015e-08, 
    2.373337e-08, 2.310542e-08, 2.383375e-08, 2.280725e-08, 2.146799e-08,
  2.284722e-08, 2.296573e-08, 2.376558e-08, 2.194219e-08, 2.108615e-08, 
    2.110246e-08, 2.110734e-08, 2.239135e-08, 2.252554e-08, 2.414346e-08, 
    2.269926e-08, 2.302788e-08, 2.301201e-08, 2.252708e-08, 2.150232e-08,
  2.336587e-08, 2.296625e-08, 2.396674e-08, 2.260454e-08, 2.229117e-08, 
    2.160209e-08, 2.216337e-08, 2.215511e-08, 2.340255e-08, 2.486781e-08, 
    2.376713e-08, 2.362444e-08, 2.351282e-08, 2.282267e-08, 2.157002e-08,
  2.430168e-08, 2.426312e-08, 2.339025e-08, 2.39136e-08, 2.402728e-08, 
    2.349236e-08, 2.318461e-08, 2.294937e-08, 2.248347e-08, 2.014518e-08, 
    1.940594e-08, 2.00131e-08, 2.169936e-08, 2.600758e-08, 2.762472e-08,
  2.4234e-08, 2.289732e-08, 2.236823e-08, 2.206043e-08, 2.249318e-08, 
    2.307326e-08, 2.370656e-08, 2.323695e-08, 2.356185e-08, 2.205365e-08, 
    2.05681e-08, 1.902617e-08, 1.938909e-08, 2.118473e-08, 2.22595e-08,
  2.373217e-08, 2.216323e-08, 2.298828e-08, 2.157558e-08, 2.075165e-08, 
    2.123638e-08, 2.245078e-08, 2.232207e-08, 2.303963e-08, 2.288376e-08, 
    2.247139e-08, 2.107082e-08, 1.98304e-08, 1.928781e-08, 1.935547e-08,
  2.230207e-08, 2.29724e-08, 2.137849e-08, 2.188209e-08, 2.225917e-08, 
    2.219578e-08, 2.209905e-08, 2.206222e-08, 2.298408e-08, 2.317971e-08, 
    2.359216e-08, 2.322563e-08, 2.232114e-08, 2.125952e-08, 1.990488e-08,
  2.31201e-08, 2.394419e-08, 2.367078e-08, 2.316585e-08, 2.305315e-08, 
    2.264995e-08, 2.193111e-08, 2.195394e-08, 2.257591e-08, 2.461142e-08, 
    2.385602e-08, 2.258961e-08, 2.215751e-08, 2.15688e-08, 1.992137e-08,
  2.363118e-08, 2.398454e-08, 2.416415e-08, 2.447996e-08, 2.402762e-08, 
    2.346095e-08, 2.314827e-08, 2.248774e-08, 2.240598e-08, 2.198442e-08, 
    2.19224e-08, 2.215911e-08, 2.154099e-08, 2.133306e-08, 2.292624e-08,
  2.493287e-08, 2.449129e-08, 2.514265e-08, 2.47697e-08, 2.417736e-08, 
    2.373175e-08, 2.332593e-08, 2.272068e-08, 2.23571e-08, 2.14325e-08, 
    2.140886e-08, 2.161958e-08, 2.179486e-08, 2.252517e-08, 2.332513e-08,
  2.47361e-08, 2.397891e-08, 2.493595e-08, 2.587979e-08, 2.446032e-08, 
    2.30462e-08, 2.253278e-08, 2.15648e-08, 2.140874e-08, 2.092328e-08, 
    2.137196e-08, 2.114057e-08, 2.192847e-08, 2.181017e-08, 2.183083e-08,
  2.457056e-08, 2.376229e-08, 2.470187e-08, 2.596261e-08, 2.451118e-08, 
    2.346603e-08, 2.170019e-08, 2.085669e-08, 2.033155e-08, 2.039002e-08, 
    2.04391e-08, 2.107711e-08, 2.212304e-08, 2.185497e-08, 2.134266e-08,
  2.457413e-08, 2.4191e-08, 2.480118e-08, 2.464476e-08, 2.466028e-08, 
    2.226074e-08, 2.047801e-08, 2.13434e-08, 2.163194e-08, 2.181715e-08, 
    2.256106e-08, 2.359397e-08, 2.34289e-08, 2.282191e-08, 2.274072e-08,
  2.563579e-08, 2.472103e-08, 2.371064e-08, 2.397503e-08, 2.449824e-08, 
    2.399524e-08, 2.278746e-08, 2.253666e-08, 2.101818e-08, 2.23609e-08, 
    2.708775e-08, 2.560272e-08, 2.812366e-08, 3.305411e-08, 3.604428e-08,
  2.481212e-08, 2.332453e-08, 2.363463e-08, 2.339491e-08, 2.319718e-08, 
    2.323964e-08, 2.36388e-08, 2.369715e-08, 2.252634e-08, 2.066453e-08, 
    2.206475e-08, 2.232718e-08, 2.194157e-08, 2.781352e-08, 2.852576e-08,
  2.387759e-08, 2.306452e-08, 2.366092e-08, 2.262433e-08, 2.213328e-08, 
    2.28741e-08, 2.344275e-08, 2.338147e-08, 2.346384e-08, 2.291238e-08, 
    2.142907e-08, 2.063441e-08, 1.796103e-08, 1.974582e-08, 2.225754e-08,
  2.330527e-08, 2.388749e-08, 2.248572e-08, 2.241072e-08, 2.34506e-08, 
    2.270544e-08, 2.323339e-08, 2.388576e-08, 2.408237e-08, 2.314445e-08, 
    2.365188e-08, 2.32885e-08, 2.040914e-08, 1.933482e-08, 1.901609e-08,
  2.376142e-08, 2.43248e-08, 2.458756e-08, 2.421434e-08, 2.39809e-08, 
    2.360795e-08, 2.33149e-08, 2.275319e-08, 2.251336e-08, 2.653203e-08, 
    2.880749e-08, 2.675462e-08, 2.370537e-08, 2.14107e-08, 1.963202e-08,
  2.417279e-08, 2.383791e-08, 2.461879e-08, 2.452856e-08, 2.413261e-08, 
    2.393125e-08, 2.370601e-08, 2.300891e-08, 2.414649e-08, 2.394529e-08, 
    2.293781e-08, 2.466653e-08, 2.458645e-08, 2.355357e-08, 2.253442e-08,
  2.461497e-08, 2.38975e-08, 2.454138e-08, 2.474815e-08, 2.5009e-08, 
    2.514514e-08, 2.469614e-08, 2.373068e-08, 2.326313e-08, 2.185902e-08, 
    2.205287e-08, 2.192859e-08, 2.368748e-08, 2.317999e-08, 2.322139e-08,
  2.469392e-08, 2.365582e-08, 2.450298e-08, 2.465452e-08, 2.471705e-08, 
    2.413815e-08, 2.374215e-08, 2.272508e-08, 2.225004e-08, 2.177891e-08, 
    2.205594e-08, 2.179693e-08, 2.336347e-08, 2.322841e-08, 2.389707e-08,
  2.504882e-08, 2.398473e-08, 2.440816e-08, 2.432222e-08, 2.442973e-08, 
    2.324213e-08, 2.343756e-08, 2.212819e-08, 2.226415e-08, 2.188486e-08, 
    2.179139e-08, 2.127859e-08, 2.156406e-08, 2.198088e-08, 2.239197e-08,
  2.512654e-08, 2.409779e-08, 2.484754e-08, 2.412086e-08, 2.419387e-08, 
    2.407063e-08, 2.289729e-08, 2.329821e-08, 2.34518e-08, 2.327536e-08, 
    2.302142e-08, 2.250924e-08, 2.185043e-08, 2.152532e-08, 2.133736e-08,
  2.462691e-08, 2.486357e-08, 2.63014e-08, 2.579027e-08, 2.550489e-08, 
    2.494884e-08, 2.467455e-08, 2.452636e-08, 2.368139e-08, 2.355815e-08, 
    2.462301e-08, 2.485359e-08, 2.350769e-08, 2.547112e-08, 2.922667e-08,
  2.492038e-08, 2.504906e-08, 2.614831e-08, 2.633711e-08, 2.56705e-08, 
    2.509592e-08, 2.460425e-08, 2.426056e-08, 2.405648e-08, 2.373394e-08, 
    2.413333e-08, 2.502622e-08, 2.458953e-08, 2.427369e-08, 2.571013e-08,
  2.716455e-08, 2.559915e-08, 2.590259e-08, 2.592995e-08, 2.582365e-08, 
    2.503754e-08, 2.446232e-08, 2.412992e-08, 2.372669e-08, 2.292321e-08, 
    2.204259e-08, 2.345729e-08, 2.46606e-08, 2.308149e-08, 2.385933e-08,
  2.664818e-08, 2.60797e-08, 2.641344e-08, 2.628702e-08, 2.579637e-08, 
    2.519431e-08, 2.471285e-08, 2.434173e-08, 2.306057e-08, 2.138433e-08, 
    2.327965e-08, 2.503541e-08, 2.540644e-08, 2.419926e-08, 2.385592e-08,
  2.675497e-08, 2.590579e-08, 2.604768e-08, 2.613278e-08, 2.571463e-08, 
    2.537977e-08, 2.505881e-08, 2.423005e-08, 2.288725e-08, 2.490399e-08, 
    2.777278e-08, 2.735166e-08, 2.260848e-08, 2.244284e-08, 2.227367e-08,
  2.558094e-08, 2.559408e-08, 2.557246e-08, 2.622311e-08, 2.638467e-08, 
    2.585409e-08, 2.52436e-08, 2.421569e-08, 2.497232e-08, 2.422832e-08, 
    2.213932e-08, 2.323735e-08, 2.366931e-08, 2.239089e-08, 2.23171e-08,
  2.517059e-08, 2.547948e-08, 2.561796e-08, 2.588634e-08, 2.614484e-08, 
    2.604828e-08, 2.568552e-08, 2.529017e-08, 2.420502e-08, 2.209209e-08, 
    2.266258e-08, 2.220452e-08, 2.478949e-08, 2.29286e-08, 2.079159e-08,
  2.461044e-08, 2.557727e-08, 2.561413e-08, 2.596385e-08, 2.630607e-08, 
    2.609249e-08, 2.549463e-08, 2.481094e-08, 2.304596e-08, 2.280698e-08, 
    2.331863e-08, 2.28001e-08, 2.500865e-08, 2.378091e-08, 2.275982e-08,
  2.438765e-08, 2.571767e-08, 2.572982e-08, 2.57844e-08, 2.640401e-08, 
    2.624329e-08, 2.553842e-08, 2.50055e-08, 2.451313e-08, 2.436452e-08, 
    2.419921e-08, 2.323233e-08, 2.388049e-08, 2.341314e-08, 2.373682e-08,
  2.43328e-08, 2.557038e-08, 2.547807e-08, 2.557467e-08, 2.585261e-08, 
    2.592147e-08, 2.568282e-08, 2.536604e-08, 2.538425e-08, 2.457078e-08, 
    2.419596e-08, 2.323292e-08, 2.33652e-08, 2.325917e-08, 2.315678e-08,
  2.166719e-08, 2.290009e-08, 2.386045e-08, 2.407161e-08, 2.416974e-08, 
    2.534299e-08, 2.622713e-08, 2.660724e-08, 2.559601e-08, 2.56975e-08, 
    2.54166e-08, 2.565075e-08, 2.579022e-08, 2.657241e-08, 2.751913e-08,
  2.1373e-08, 2.257891e-08, 2.380388e-08, 2.457527e-08, 2.452316e-08, 
    2.528034e-08, 2.586287e-08, 2.660896e-08, 2.637772e-08, 2.590614e-08, 
    2.562988e-08, 2.528556e-08, 2.505318e-08, 2.55643e-08, 2.550863e-08,
  2.337674e-08, 2.270128e-08, 2.391589e-08, 2.537616e-08, 2.559645e-08, 
    2.513376e-08, 2.549711e-08, 2.625647e-08, 2.620013e-08, 2.621523e-08, 
    2.550607e-08, 2.531654e-08, 2.473797e-08, 2.477411e-08, 2.456061e-08,
  2.252503e-08, 2.281762e-08, 2.396461e-08, 2.4289e-08, 2.473474e-08, 
    2.51018e-08, 2.560716e-08, 2.611728e-08, 2.674226e-08, 2.654184e-08, 
    2.747869e-08, 2.730083e-08, 2.530907e-08, 2.531006e-08, 2.497043e-08,
  2.300717e-08, 2.308244e-08, 2.317648e-08, 2.394292e-08, 2.47798e-08, 
    2.525045e-08, 2.631886e-08, 2.608371e-08, 2.708887e-08, 2.704435e-08, 
    2.535856e-08, 2.559504e-08, 2.502426e-08, 2.505421e-08, 2.439729e-08,
  2.251471e-08, 2.289153e-08, 2.248248e-08, 2.300523e-08, 2.418402e-08, 
    2.443376e-08, 2.52035e-08, 2.553119e-08, 2.498573e-08, 2.470038e-08, 
    2.474022e-08, 2.424738e-08, 2.578558e-08, 2.552026e-08, 2.421739e-08,
  2.23042e-08, 2.311121e-08, 2.267713e-08, 2.337171e-08, 2.408389e-08, 
    2.423013e-08, 2.477453e-08, 2.457487e-08, 2.465093e-08, 2.445382e-08, 
    2.549281e-08, 2.490366e-08, 2.626343e-08, 2.571744e-08, 2.392395e-08,
  2.239484e-08, 2.305395e-08, 2.27847e-08, 2.356846e-08, 2.41953e-08, 
    2.472511e-08, 2.472619e-08, 2.421806e-08, 2.369739e-08, 2.439933e-08, 
    2.540851e-08, 2.534301e-08, 2.63268e-08, 2.59005e-08, 2.526337e-08,
  2.258246e-08, 2.330564e-08, 2.322367e-08, 2.382443e-08, 2.433396e-08, 
    2.474806e-08, 2.39868e-08, 2.317116e-08, 2.364126e-08, 2.518457e-08, 
    2.550917e-08, 2.555793e-08, 2.582996e-08, 2.577681e-08, 2.498987e-08,
  2.305384e-08, 2.33505e-08, 2.313571e-08, 2.306021e-08, 2.345017e-08, 
    2.34946e-08, 2.276967e-08, 2.313419e-08, 2.46302e-08, 2.541941e-08, 
    2.541253e-08, 2.539593e-08, 2.556203e-08, 2.500999e-08, 2.446353e-08,
  1.534016e-08, 1.704235e-08, 1.838143e-08, 2.025849e-08, 2.099316e-08, 
    2.244315e-08, 2.285998e-08, 2.316554e-08, 2.400514e-08, 2.478505e-08, 
    2.508003e-08, 2.525727e-08, 2.568603e-08, 2.637823e-08, 2.898289e-08,
  1.715538e-08, 1.846249e-08, 1.98776e-08, 2.194909e-08, 2.289912e-08, 
    2.305159e-08, 2.270172e-08, 2.332253e-08, 2.451617e-08, 2.506028e-08, 
    2.493658e-08, 2.550795e-08, 2.536939e-08, 2.628614e-08, 2.667937e-08,
  2.000376e-08, 2.07291e-08, 2.216293e-08, 2.482687e-08, 2.455014e-08, 
    2.35434e-08, 2.294243e-08, 2.358789e-08, 2.475102e-08, 2.495883e-08, 
    2.575164e-08, 2.643242e-08, 2.565067e-08, 2.603818e-08, 2.50373e-08,
  2.178344e-08, 2.147497e-08, 2.293102e-08, 2.354586e-08, 2.323718e-08, 
    2.352044e-08, 2.333659e-08, 2.388587e-08, 2.490652e-08, 2.513245e-08, 
    2.839434e-08, 2.790823e-08, 2.527729e-08, 2.644547e-08, 2.605505e-08,
  2.253712e-08, 2.216319e-08, 2.296563e-08, 2.33321e-08, 2.401193e-08, 
    2.414872e-08, 2.406588e-08, 2.467164e-08, 2.501044e-08, 2.584256e-08, 
    2.708374e-08, 2.623177e-08, 2.585942e-08, 2.603875e-08, 2.400081e-08,
  2.318981e-08, 2.281857e-08, 2.32274e-08, 2.313717e-08, 2.38153e-08, 
    2.379838e-08, 2.437653e-08, 2.47892e-08, 2.452021e-08, 2.600939e-08, 
    2.609118e-08, 2.552203e-08, 2.789018e-08, 2.688448e-08, 2.424204e-08,
  2.225488e-08, 2.297319e-08, 2.341093e-08, 2.341516e-08, 2.431943e-08, 
    2.443454e-08, 2.427821e-08, 2.363156e-08, 2.31598e-08, 2.396586e-08, 
    2.561546e-08, 2.640541e-08, 2.870375e-08, 2.798316e-08, 2.592211e-08,
  2.228512e-08, 2.330177e-08, 2.301403e-08, 2.359259e-08, 2.480815e-08, 
    2.51497e-08, 2.435767e-08, 2.28568e-08, 2.184623e-08, 2.359607e-08, 
    2.480933e-08, 2.55289e-08, 2.779972e-08, 2.75495e-08, 2.43842e-08,
  2.228746e-08, 2.300428e-08, 2.300395e-08, 2.497995e-08, 2.528987e-08, 
    2.47387e-08, 2.268679e-08, 2.088686e-08, 2.166307e-08, 2.381801e-08, 
    2.411223e-08, 2.489869e-08, 2.624989e-08, 2.552305e-08, 2.430921e-08,
  2.258076e-08, 2.274123e-08, 2.328633e-08, 2.225475e-08, 2.155907e-08, 
    2.076388e-08, 2.00479e-08, 2.086992e-08, 2.307601e-08, 2.362305e-08, 
    2.372764e-08, 2.446397e-08, 2.491947e-08, 2.490676e-08, 2.548101e-08,
  1.824685e-08, 1.846612e-08, 1.898686e-08, 1.911928e-08, 1.912677e-08, 
    1.904222e-08, 1.894528e-08, 1.979192e-08, 2.087406e-08, 2.066518e-08, 
    2.103443e-08, 2.228253e-08, 2.315229e-08, 2.098916e-08, 2.045442e-08,
  2.094229e-08, 2.069725e-08, 1.994121e-08, 1.972054e-08, 1.98319e-08, 
    2.008208e-08, 2.006097e-08, 2.040736e-08, 2.147117e-08, 2.098343e-08, 
    2.152071e-08, 2.23041e-08, 2.275274e-08, 2.048828e-08, 1.943012e-08,
  2.275829e-08, 2.168822e-08, 2.018078e-08, 2.036161e-08, 2.052894e-08, 
    2.034496e-08, 2.050919e-08, 2.023113e-08, 2.107059e-08, 2.058298e-08, 
    2.100997e-08, 2.104761e-08, 2.234079e-08, 2.076596e-08, 2.051616e-08,
  2.492225e-08, 2.292881e-08, 2.167862e-08, 2.147888e-08, 2.097368e-08, 
    2.022469e-08, 1.981982e-08, 1.97654e-08, 1.964595e-08, 2.006649e-08, 
    1.996459e-08, 2.009996e-08, 2.173783e-08, 2.178713e-08, 2.379774e-08,
  2.41753e-08, 2.201265e-08, 2.101462e-08, 2.142471e-08, 2.141425e-08, 
    2.101582e-08, 2.015921e-08, 2.006262e-08, 1.960459e-08, 1.855518e-08, 
    1.92486e-08, 2.072792e-08, 2.132187e-08, 2.335366e-08, 2.403186e-08,
  2.332741e-08, 2.213763e-08, 2.088659e-08, 2.119061e-08, 2.092568e-08, 
    2.11277e-08, 2.077015e-08, 2.102228e-08, 2.134365e-08, 2.03772e-08, 
    2.227914e-08, 2.128102e-08, 2.026993e-08, 2.594932e-08, 2.226001e-08,
  2.192233e-08, 2.278302e-08, 2.292145e-08, 2.210078e-08, 2.137586e-08, 
    2.136907e-08, 2.098741e-08, 2.176617e-08, 2.206675e-08, 2.156095e-08, 
    2.172398e-08, 2.060476e-08, 2.078696e-08, 2.255983e-08, 1.990894e-08,
  2.200498e-08, 2.359139e-08, 2.419556e-08, 2.269849e-08, 2.244529e-08, 
    2.128283e-08, 2.072917e-08, 2.081821e-08, 2.141065e-08, 2.109563e-08, 
    2.038226e-08, 1.974322e-08, 2.01198e-08, 1.804347e-08, 1.685534e-08,
  2.292324e-08, 2.371668e-08, 2.365436e-08, 2.291115e-08, 2.304878e-08, 
    2.288031e-08, 2.218325e-08, 2.038189e-08, 2.049898e-08, 2.068896e-08, 
    2.038646e-08, 1.985223e-08, 1.956204e-08, 1.852289e-08, 1.891903e-08,
  2.374874e-08, 2.331385e-08, 2.220121e-08, 2.108178e-08, 2.087316e-08, 
    2.093858e-08, 2.082365e-08, 2.090635e-08, 2.199639e-08, 2.165434e-08, 
    2.117075e-08, 2.04291e-08, 2.041412e-08, 2.033859e-08, 2.207278e-08,
  2.404847e-08, 2.405293e-08, 2.330817e-08, 2.371596e-08, 2.241886e-08, 
    2.170383e-08, 2.045376e-08, 2.027164e-08, 1.92334e-08, 1.906698e-08, 
    2.046977e-08, 2.205275e-08, 2.238973e-08, 2.12455e-08, 2.108091e-08,
  2.589778e-08, 2.67617e-08, 2.692849e-08, 2.718859e-08, 2.631627e-08, 
    2.446083e-08, 2.227685e-08, 2.110113e-08, 1.971923e-08, 2.018189e-08, 
    2.065951e-08, 2.130149e-08, 2.179762e-08, 2.105241e-08, 2.037699e-08,
  2.688307e-08, 2.798662e-08, 2.735999e-08, 2.721418e-08, 2.669239e-08, 
    2.577604e-08, 2.467534e-08, 2.251905e-08, 2.116544e-08, 2.113338e-08, 
    2.185331e-08, 2.113959e-08, 2.147277e-08, 2.160362e-08, 2.12057e-08,
  2.746495e-08, 2.73083e-08, 2.741497e-08, 2.67917e-08, 2.528577e-08, 
    2.535506e-08, 2.366634e-08, 2.166923e-08, 2.31723e-08, 2.344517e-08, 
    2.278746e-08, 2.357789e-08, 2.327837e-08, 2.636992e-08, 2.500694e-08,
  2.43483e-08, 2.416341e-08, 2.371063e-08, 2.306336e-08, 2.311956e-08, 
    2.509834e-08, 2.589356e-08, 2.410789e-08, 2.342084e-08, 2.608369e-08, 
    2.605932e-08, 2.544209e-08, 2.41113e-08, 2.819945e-08, 2.765584e-08,
  2.250073e-08, 2.267121e-08, 2.341897e-08, 2.224303e-08, 2.173148e-08, 
    2.241145e-08, 2.583731e-08, 2.914666e-08, 3.016843e-08, 2.535234e-08, 
    2.594336e-08, 2.582396e-08, 2.418153e-08, 2.598823e-08, 2.769529e-08,
  2.21859e-08, 2.188879e-08, 2.261165e-08, 2.288537e-08, 2.203613e-08, 
    2.256018e-08, 2.631156e-08, 3.168091e-08, 3.106116e-08, 2.495606e-08, 
    2.475508e-08, 2.439007e-08, 2.358011e-08, 2.530678e-08, 2.423663e-08,
  2.39226e-08, 2.306706e-08, 2.24863e-08, 2.251841e-08, 2.162537e-08, 
    1.877194e-08, 2.478612e-08, 3.455338e-08, 3.541636e-08, 2.891243e-08, 
    2.602131e-08, 2.391051e-08, 2.347756e-08, 2.304027e-08, 2.344083e-08,
  2.367374e-08, 2.408395e-08, 2.290109e-08, 2.213131e-08, 2.207492e-08, 
    1.842851e-08, 2.038959e-08, 2.955276e-08, 3.268523e-08, 2.965069e-08, 
    2.576509e-08, 2.439886e-08, 2.329724e-08, 2.314951e-08, 2.18363e-08,
  2.372557e-08, 2.431288e-08, 2.413293e-08, 2.309122e-08, 1.947324e-08, 
    1.704859e-08, 2.055778e-08, 2.686593e-08, 2.59617e-08, 2.998592e-08, 
    2.723139e-08, 2.537765e-08, 2.467589e-08, 2.369871e-08, 2.284442e-08,
  2.615186e-08, 2.77978e-08, 2.808432e-08, 2.911616e-08, 2.983051e-08, 
    2.928357e-08, 2.88122e-08, 2.845183e-08, 2.675914e-08, 2.574857e-08, 
    2.615972e-08, 2.607909e-08, 2.495434e-08, 2.463482e-08, 2.468037e-08,
  2.615477e-08, 2.767266e-08, 2.795566e-08, 2.822368e-08, 2.957592e-08, 
    2.97878e-08, 2.967302e-08, 2.74162e-08, 2.665327e-08, 2.787061e-08, 
    2.74028e-08, 2.705934e-08, 2.591908e-08, 2.620515e-08, 2.446449e-08,
  2.495793e-08, 2.703159e-08, 2.914653e-08, 2.937768e-08, 3.02024e-08, 
    3.152587e-08, 3.187483e-08, 2.836192e-08, 2.750382e-08, 2.693323e-08, 
    2.741096e-08, 2.783494e-08, 2.72672e-08, 2.727e-08, 2.51449e-08,
  2.395251e-08, 2.51478e-08, 2.578182e-08, 2.87526e-08, 3.01493e-08, 
    3.20427e-08, 3.049834e-08, 2.865572e-08, 2.867147e-08, 2.855051e-08, 
    2.523466e-08, 2.670605e-08, 2.971898e-08, 2.99165e-08, 2.687294e-08,
  2.31426e-08, 2.297612e-08, 2.338352e-08, 2.439342e-08, 2.700612e-08, 
    2.968302e-08, 3.148686e-08, 3.011376e-08, 2.871639e-08, 3.196087e-08, 
    2.732988e-08, 2.282419e-08, 2.55817e-08, 2.893809e-08, 2.77801e-08,
  2.2443e-08, 2.206042e-08, 2.254206e-08, 2.231216e-08, 2.389556e-08, 
    2.627225e-08, 2.938843e-08, 3.154807e-08, 3.384564e-08, 3.21418e-08, 
    2.89458e-08, 2.587029e-08, 2.494654e-08, 2.608729e-08, 2.933214e-08,
  2.328877e-08, 2.27656e-08, 2.273032e-08, 2.136421e-08, 2.030577e-08, 
    2.094107e-08, 2.515968e-08, 2.799907e-08, 3.212725e-08, 3.121418e-08, 
    3.393702e-08, 3.103609e-08, 2.560679e-08, 2.511324e-08, 3.141695e-08,
  2.389394e-08, 2.391144e-08, 2.276799e-08, 2.19603e-08, 2.180489e-08, 
    1.981891e-08, 2.136007e-08, 2.416605e-08, 3.072299e-08, 2.954221e-08, 
    3.190226e-08, 3.019816e-08, 2.601172e-08, 2.394148e-08, 2.892626e-08,
  2.555455e-08, 2.426904e-08, 2.268522e-08, 2.219901e-08, 2.196748e-08, 
    2.019851e-08, 1.964341e-08, 1.913161e-08, 2.039179e-08, 2.546208e-08, 
    2.942256e-08, 3.053093e-08, 2.872279e-08, 2.470693e-08, 2.542091e-08,
  2.617545e-08, 2.494857e-08, 2.282918e-08, 2.204435e-08, 2.188907e-08, 
    2.098708e-08, 1.971624e-08, 1.836868e-08, 1.852247e-08, 2.121425e-08, 
    2.433844e-08, 2.794616e-08, 2.908019e-08, 2.655861e-08, 2.411022e-08,
  2.329895e-08, 2.323032e-08, 2.325911e-08, 2.262672e-08, 2.228471e-08, 
    2.393396e-08, 2.473665e-08, 2.436865e-08, 2.355303e-08, 2.41666e-08, 
    2.337639e-08, 2.32014e-08, 2.385209e-08, 2.747948e-08, 2.806365e-08,
  2.32842e-08, 2.285093e-08, 2.298794e-08, 2.24056e-08, 2.187448e-08, 
    2.35191e-08, 2.550292e-08, 2.561436e-08, 2.445559e-08, 2.557012e-08, 
    2.487775e-08, 2.342754e-08, 2.236808e-08, 2.521173e-08, 2.625728e-08,
  2.418926e-08, 2.371372e-08, 2.366589e-08, 2.308808e-08, 2.223438e-08, 
    2.378267e-08, 2.569053e-08, 2.600884e-08, 2.532591e-08, 2.66795e-08, 
    2.724563e-08, 2.488449e-08, 2.269312e-08, 2.404927e-08, 2.440247e-08,
  2.497436e-08, 2.426077e-08, 2.359386e-08, 2.272865e-08, 2.222952e-08, 
    2.260616e-08, 2.411707e-08, 2.701067e-08, 2.772973e-08, 2.859021e-08, 
    2.758336e-08, 2.559284e-08, 2.20191e-08, 2.255404e-08, 2.270343e-08,
  2.558305e-08, 2.474903e-08, 2.484652e-08, 2.384312e-08, 2.272386e-08, 
    2.241912e-08, 2.329405e-08, 2.63064e-08, 2.890953e-08, 3.183577e-08, 
    2.693265e-08, 2.461016e-08, 2.069403e-08, 1.995291e-08, 2.028185e-08,
  2.503871e-08, 2.4879e-08, 2.399209e-08, 2.395337e-08, 2.311095e-08, 
    2.221206e-08, 2.262419e-08, 2.495837e-08, 3.05614e-08, 2.951976e-08, 
    2.782897e-08, 2.752055e-08, 2.399649e-08, 2.015689e-08, 2.229247e-08,
  2.484179e-08, 2.59461e-08, 2.517019e-08, 2.504318e-08, 2.361691e-08, 
    2.288195e-08, 2.191562e-08, 2.295566e-08, 2.796826e-08, 2.811991e-08, 
    2.967152e-08, 3.112506e-08, 2.64877e-08, 2.20333e-08, 2.589655e-08,
  2.628673e-08, 2.732543e-08, 2.645847e-08, 2.560475e-08, 2.359929e-08, 
    2.264558e-08, 2.175648e-08, 2.123141e-08, 2.580793e-08, 2.81879e-08, 
    2.956572e-08, 3.001404e-08, 2.863066e-08, 2.462742e-08, 2.508039e-08,
  2.605048e-08, 2.730164e-08, 2.71063e-08, 2.578789e-08, 2.326178e-08, 
    2.164421e-08, 2.116663e-08, 2.020836e-08, 2.014762e-08, 2.534008e-08, 
    2.924082e-08, 2.986278e-08, 3.023264e-08, 2.967853e-08, 2.847729e-08,
  2.64195e-08, 2.695035e-08, 2.645399e-08, 2.525228e-08, 2.348848e-08, 
    2.232659e-08, 2.128708e-08, 2.081447e-08, 1.914223e-08, 2.089959e-08, 
    2.63469e-08, 2.888506e-08, 3.001107e-08, 3.174526e-08, 3.032687e-08,
  2.557134e-08, 2.604765e-08, 2.561813e-08, 2.605206e-08, 2.524019e-08, 
    2.557268e-08, 2.409704e-08, 2.508423e-08, 2.383301e-08, 2.367893e-08, 
    2.467118e-08, 2.394219e-08, 2.199522e-08, 2.26282e-08, 2.327503e-08,
  2.550208e-08, 2.584906e-08, 2.543361e-08, 2.553447e-08, 2.505307e-08, 
    2.502459e-08, 2.38534e-08, 2.464326e-08, 2.375455e-08, 2.370463e-08, 
    2.399839e-08, 2.359797e-08, 2.201929e-08, 2.200262e-08, 2.293053e-08,
  2.575016e-08, 2.675911e-08, 2.669103e-08, 2.582293e-08, 2.479519e-08, 
    2.454442e-08, 2.40283e-08, 2.400778e-08, 2.288082e-08, 2.374594e-08, 
    2.428334e-08, 2.463824e-08, 2.312395e-08, 2.310395e-08, 2.205408e-08,
  2.658637e-08, 2.763628e-08, 2.758994e-08, 2.678869e-08, 2.587757e-08, 
    2.539641e-08, 2.465065e-08, 2.486152e-08, 2.370516e-08, 2.367473e-08, 
    2.555786e-08, 2.691318e-08, 2.543862e-08, 2.326818e-08, 2.030922e-08,
  2.715751e-08, 2.817231e-08, 2.833572e-08, 2.782015e-08, 2.640715e-08, 
    2.569022e-08, 2.487911e-08, 2.533708e-08, 2.433393e-08, 2.821782e-08, 
    2.451783e-08, 2.183634e-08, 2.644377e-08, 2.104364e-08, 1.707286e-08,
  2.889917e-08, 2.923641e-08, 2.93317e-08, 2.84984e-08, 2.718977e-08, 
    2.615334e-08, 2.477852e-08, 2.526313e-08, 2.4804e-08, 2.504457e-08, 
    2.250178e-08, 2.116529e-08, 2.079339e-08, 1.738871e-08, 1.769335e-08,
  3.025837e-08, 3.017225e-08, 2.96135e-08, 2.863935e-08, 2.725155e-08, 
    2.646059e-08, 2.529134e-08, 2.520618e-08, 2.47479e-08, 2.283291e-08, 
    2.200595e-08, 2.160399e-08, 1.925127e-08, 1.589922e-08, 2.112767e-08,
  3.106273e-08, 3.242867e-08, 3.133656e-08, 2.962197e-08, 2.756118e-08, 
    2.66532e-08, 2.570727e-08, 2.521515e-08, 2.519342e-08, 2.32935e-08, 
    2.20073e-08, 2.145171e-08, 1.903254e-08, 1.763264e-08, 2.160858e-08,
  2.899544e-08, 3.1544e-08, 3.257902e-08, 3.125876e-08, 2.86164e-08, 
    2.724753e-08, 2.646933e-08, 2.593657e-08, 2.479585e-08, 2.35053e-08, 
    2.185007e-08, 2.144509e-08, 2.017071e-08, 1.987395e-08, 1.998354e-08,
  2.580106e-08, 2.78265e-08, 3.168307e-08, 3.293307e-08, 3.017689e-08, 
    2.793879e-08, 2.725601e-08, 2.50867e-08, 2.404202e-08, 2.369228e-08, 
    2.22488e-08, 2.179955e-08, 2.13668e-08, 2.131703e-08, 2.061791e-08,
  2.379916e-08, 2.378378e-08, 2.322701e-08, 2.360951e-08, 2.390592e-08, 
    2.410808e-08, 2.470308e-08, 2.446413e-08, 2.419271e-08, 2.433023e-08, 
    2.530477e-08, 2.527373e-08, 2.405522e-08, 2.371326e-08, 2.538922e-08,
  2.351387e-08, 2.312861e-08, 2.262511e-08, 2.359969e-08, 2.410475e-08, 
    2.46486e-08, 2.476922e-08, 2.500386e-08, 2.462491e-08, 2.480689e-08, 
    2.525161e-08, 2.521014e-08, 2.38766e-08, 2.337256e-08, 2.571938e-08,
  2.233811e-08, 2.367456e-08, 2.342777e-08, 2.407301e-08, 2.434396e-08, 
    2.527876e-08, 2.434243e-08, 2.390136e-08, 2.423777e-08, 2.515944e-08, 
    2.554843e-08, 2.53392e-08, 2.356599e-08, 2.381574e-08, 2.437129e-08,
  2.260428e-08, 2.389186e-08, 2.443673e-08, 2.443846e-08, 2.531142e-08, 
    2.596596e-08, 2.600745e-08, 2.478376e-08, 2.485616e-08, 2.556519e-08, 
    2.674893e-08, 2.580854e-08, 2.37115e-08, 2.424334e-08, 2.295731e-08,
  2.30859e-08, 2.500135e-08, 2.73635e-08, 2.818679e-08, 2.766456e-08, 
    2.685575e-08, 2.619803e-08, 2.571085e-08, 2.536729e-08, 2.815819e-08, 
    2.80396e-08, 2.519196e-08, 2.477996e-08, 2.261096e-08, 2.213279e-08,
  2.501716e-08, 2.636352e-08, 2.835746e-08, 2.866543e-08, 2.957374e-08, 
    2.84247e-08, 2.686333e-08, 2.645348e-08, 2.655845e-08, 2.757905e-08, 
    2.647544e-08, 2.438805e-08, 2.215897e-08, 2.060826e-08, 2.269621e-08,
  2.515503e-08, 2.649915e-08, 2.920881e-08, 2.979262e-08, 3.068076e-08, 
    2.992475e-08, 2.796949e-08, 2.758946e-08, 2.687383e-08, 2.619577e-08, 
    2.600427e-08, 2.369105e-08, 2.051513e-08, 2.068264e-08, 2.562096e-08,
  2.559523e-08, 2.7064e-08, 3.041274e-08, 3.057379e-08, 3.104596e-08, 
    3.018704e-08, 2.832923e-08, 2.770719e-08, 2.680276e-08, 2.613703e-08, 
    2.548578e-08, 2.274756e-08, 1.983831e-08, 2.22635e-08, 2.518379e-08,
  2.505153e-08, 2.713086e-08, 3.003299e-08, 3.105065e-08, 3.169992e-08, 
    3.226716e-08, 2.93497e-08, 2.863053e-08, 2.70612e-08, 2.520082e-08, 
    2.468376e-08, 2.185467e-08, 2.035168e-08, 2.284817e-08, 2.175312e-08,
  2.545e-08, 2.769471e-08, 2.875922e-08, 3.222515e-08, 3.339957e-08, 
    3.364724e-08, 3.132309e-08, 2.800387e-08, 2.587407e-08, 2.499807e-08, 
    2.424672e-08, 2.171563e-08, 2.063696e-08, 2.104415e-08, 2.022655e-08,
  2.816774e-08, 2.749226e-08, 2.692431e-08, 2.645709e-08, 2.617455e-08, 
    2.596934e-08, 2.609067e-08, 2.621348e-08, 2.557363e-08, 2.615982e-08, 
    2.813349e-08, 2.820585e-08, 2.730549e-08, 2.754484e-08, 2.970698e-08,
  2.771199e-08, 2.582703e-08, 2.516459e-08, 2.525271e-08, 2.486505e-08, 
    2.460289e-08, 2.428047e-08, 2.466213e-08, 2.42144e-08, 2.602038e-08, 
    2.724204e-08, 2.825817e-08, 2.714889e-08, 2.725614e-08, 2.979875e-08,
  2.707671e-08, 2.45965e-08, 2.398538e-08, 2.410391e-08, 2.327586e-08, 
    2.360112e-08, 2.272221e-08, 2.286266e-08, 2.379465e-08, 2.499003e-08, 
    2.671216e-08, 2.772865e-08, 2.704277e-08, 2.797776e-08, 2.809907e-08,
  2.557457e-08, 2.360792e-08, 2.419902e-08, 2.484447e-08, 2.455024e-08, 
    2.414998e-08, 2.347289e-08, 2.244447e-08, 2.264154e-08, 2.389859e-08, 
    2.641195e-08, 3.001239e-08, 3.024654e-08, 2.8847e-08, 2.553947e-08,
  2.558165e-08, 2.48466e-08, 2.585948e-08, 2.618462e-08, 2.621837e-08, 
    2.568946e-08, 2.427972e-08, 2.333829e-08, 2.270367e-08, 2.690481e-08, 
    2.440826e-08, 2.451964e-08, 2.908589e-08, 2.544261e-08, 2.495404e-08,
  2.604284e-08, 2.599441e-08, 2.648159e-08, 2.619943e-08, 2.55856e-08, 
    2.586746e-08, 2.570754e-08, 2.478072e-08, 2.393095e-08, 2.393577e-08, 
    2.46852e-08, 2.577561e-08, 2.636114e-08, 2.214344e-08, 2.651887e-08,
  2.588483e-08, 2.57383e-08, 2.584467e-08, 2.498188e-08, 2.545461e-08, 
    2.521888e-08, 2.445938e-08, 2.403901e-08, 2.383063e-08, 2.207185e-08, 
    2.50404e-08, 2.676707e-08, 2.485128e-08, 2.165462e-08, 3.015754e-08,
  2.540411e-08, 2.548403e-08, 2.566169e-08, 2.497766e-08, 2.492504e-08, 
    2.550669e-08, 2.513327e-08, 2.471834e-08, 2.405636e-08, 2.273509e-08, 
    2.541334e-08, 2.651518e-08, 2.358821e-08, 2.524419e-08, 3.082533e-08,
  2.565452e-08, 2.635949e-08, 2.529621e-08, 2.460034e-08, 2.530965e-08, 
    2.683319e-08, 2.607125e-08, 2.498154e-08, 2.467035e-08, 2.33058e-08, 
    2.543282e-08, 2.636172e-08, 2.474312e-08, 2.72926e-08, 2.625987e-08,
  2.607215e-08, 2.584342e-08, 2.508411e-08, 2.61246e-08, 2.680257e-08, 
    2.822723e-08, 2.830367e-08, 2.536466e-08, 2.439033e-08, 2.402897e-08, 
    2.559499e-08, 2.62554e-08, 2.533728e-08, 2.577514e-08, 2.399771e-08,
  2.779323e-08, 2.753496e-08, 2.744921e-08, 2.691137e-08, 2.700864e-08, 
    2.680381e-08, 2.59406e-08, 2.605464e-08, 2.586078e-08, 2.618942e-08, 
    2.712621e-08, 2.814362e-08, 2.823315e-08, 2.993264e-08, 3.264031e-08,
  2.874961e-08, 2.811269e-08, 2.708627e-08, 2.684324e-08, 2.769688e-08, 
    2.707349e-08, 2.611247e-08, 2.621713e-08, 2.507867e-08, 2.566285e-08, 
    2.663596e-08, 2.734282e-08, 2.780064e-08, 3.091891e-08, 3.242331e-08,
  3.09376e-08, 2.867145e-08, 2.710202e-08, 2.699659e-08, 2.833478e-08, 
    2.706295e-08, 2.584772e-08, 2.552849e-08, 2.576619e-08, 2.570809e-08, 
    2.640992e-08, 2.751021e-08, 2.855511e-08, 3.204863e-08, 3.118515e-08,
  2.973786e-08, 2.758053e-08, 2.765661e-08, 2.796864e-08, 2.770171e-08, 
    2.697278e-08, 2.644862e-08, 2.522108e-08, 2.447049e-08, 2.47038e-08, 
    2.619695e-08, 2.84944e-08, 3.14303e-08, 3.329168e-08, 3.032748e-08,
  2.898374e-08, 2.797001e-08, 2.786831e-08, 2.674926e-08, 2.621519e-08, 
    2.632045e-08, 2.569514e-08, 2.462393e-08, 2.366194e-08, 2.585565e-08, 
    2.570906e-08, 2.506778e-08, 2.923143e-08, 2.921759e-08, 2.87544e-08,
  2.965897e-08, 2.875967e-08, 2.799321e-08, 2.619729e-08, 2.592825e-08, 
    2.537293e-08, 2.4824e-08, 2.394692e-08, 2.306078e-08, 2.329091e-08, 
    2.532293e-08, 2.647783e-08, 2.810305e-08, 2.451165e-08, 3.183322e-08,
  2.890242e-08, 2.847978e-08, 2.765818e-08, 2.639351e-08, 2.618173e-08, 
    2.56147e-08, 2.417432e-08, 2.380164e-08, 2.244667e-08, 2.128614e-08, 
    2.488028e-08, 2.737866e-08, 2.634854e-08, 2.542977e-08, 3.507932e-08,
  2.860961e-08, 2.865693e-08, 2.732819e-08, 2.633356e-08, 2.641104e-08, 
    2.490328e-08, 2.358097e-08, 2.372962e-08, 2.25121e-08, 2.100613e-08, 
    2.48988e-08, 2.725293e-08, 2.56085e-08, 2.92738e-08, 3.724049e-08,
  2.789732e-08, 2.793534e-08, 2.736727e-08, 2.635446e-08, 2.601156e-08, 
    2.467183e-08, 2.265002e-08, 2.209308e-08, 2.204795e-08, 2.104635e-08, 
    2.478979e-08, 2.808654e-08, 2.758546e-08, 3.260224e-08, 3.093529e-08,
  2.632589e-08, 2.706133e-08, 2.776482e-08, 2.688993e-08, 2.615017e-08, 
    2.67549e-08, 2.589586e-08, 2.323172e-08, 2.205647e-08, 2.102946e-08, 
    2.500297e-08, 2.868645e-08, 2.888548e-08, 3.014848e-08, 2.84811e-08,
  2.72768e-08, 2.813272e-08, 2.814079e-08, 2.904278e-08, 2.898373e-08, 
    2.984986e-08, 2.925681e-08, 2.915666e-08, 2.87969e-08, 2.802333e-08, 
    2.748303e-08, 2.664877e-08, 2.597043e-08, 2.517997e-08, 2.619744e-08,
  2.82656e-08, 2.853446e-08, 2.863064e-08, 2.920051e-08, 3.017719e-08, 
    3.118471e-08, 3.036358e-08, 3.005147e-08, 2.972414e-08, 2.837714e-08, 
    2.751045e-08, 2.622938e-08, 2.498978e-08, 2.509676e-08, 2.610033e-08,
  2.819714e-08, 2.960163e-08, 2.963599e-08, 3.073105e-08, 3.153248e-08, 
    3.189344e-08, 3.059818e-08, 3.012726e-08, 2.958728e-08, 2.829576e-08, 
    2.697616e-08, 2.604872e-08, 2.499049e-08, 2.498375e-08, 2.625405e-08,
  2.84926e-08, 2.849739e-08, 2.960082e-08, 3.060581e-08, 3.090129e-08, 
    2.994525e-08, 2.962634e-08, 2.920097e-08, 2.735364e-08, 2.747067e-08, 
    2.764603e-08, 2.694489e-08, 2.699444e-08, 2.731077e-08, 2.720784e-08,
  2.934947e-08, 2.931823e-08, 3.049903e-08, 3.068511e-08, 3.049475e-08, 
    2.952958e-08, 2.904436e-08, 2.876514e-08, 2.789941e-08, 2.874889e-08, 
    2.64198e-08, 2.432887e-08, 2.447674e-08, 2.431946e-08, 2.846351e-08,
  2.79977e-08, 2.835213e-08, 2.863479e-08, 2.990269e-08, 2.991786e-08, 
    2.953714e-08, 2.846291e-08, 2.795229e-08, 2.788548e-08, 2.537667e-08, 
    2.573439e-08, 2.45008e-08, 2.404528e-08, 2.173071e-08, 2.770236e-08,
  2.778602e-08, 2.831226e-08, 2.825718e-08, 2.879903e-08, 2.826187e-08, 
    2.817423e-08, 2.685436e-08, 2.731341e-08, 2.642931e-08, 2.456822e-08, 
    2.515536e-08, 2.516262e-08, 2.390031e-08, 2.412221e-08, 3.051276e-08,
  2.685143e-08, 2.790759e-08, 2.805258e-08, 2.740821e-08, 2.738747e-08, 
    2.769978e-08, 2.682051e-08, 2.715086e-08, 2.65666e-08, 2.42195e-08, 
    2.466554e-08, 2.536124e-08, 2.437392e-08, 2.618293e-08, 2.808191e-08,
  2.746015e-08, 2.831838e-08, 2.780728e-08, 2.731647e-08, 2.688655e-08, 
    2.721428e-08, 2.570189e-08, 2.574998e-08, 2.504754e-08, 2.361713e-08, 
    2.442378e-08, 2.605046e-08, 2.458777e-08, 2.505266e-08, 2.604286e-08,
  2.738773e-08, 2.826104e-08, 2.784315e-08, 2.6943e-08, 2.648434e-08, 
    2.698179e-08, 2.585418e-08, 2.35462e-08, 2.394642e-08, 2.277404e-08, 
    2.444653e-08, 2.688837e-08, 2.53412e-08, 2.539117e-08, 2.671955e-08,
  2.971779e-08, 2.741551e-08, 2.664519e-08, 2.781601e-08, 2.941058e-08, 
    2.990575e-08, 3.032048e-08, 2.828267e-08, 2.732687e-08, 2.670624e-08, 
    2.733747e-08, 2.704318e-08, 2.732319e-08, 2.662172e-08, 2.415594e-08,
  2.832684e-08, 2.787239e-08, 2.574552e-08, 2.582208e-08, 2.812092e-08, 
    3.010426e-08, 3.163271e-08, 3.12245e-08, 2.916203e-08, 2.902066e-08, 
    2.80532e-08, 2.728244e-08, 2.670278e-08, 2.564493e-08, 2.388916e-08,
  3.042765e-08, 2.861302e-08, 2.661548e-08, 2.482428e-08, 2.731012e-08, 
    3.03651e-08, 3.146404e-08, 3.366153e-08, 3.204179e-08, 3.208492e-08, 
    3.031775e-08, 2.835968e-08, 2.729102e-08, 2.532705e-08, 2.557187e-08,
  3.184816e-08, 3.0653e-08, 2.881592e-08, 2.553606e-08, 2.681619e-08, 
    2.826296e-08, 3.07436e-08, 3.245003e-08, 3.238522e-08, 3.400959e-08, 
    3.311855e-08, 2.954599e-08, 2.86568e-08, 2.410797e-08, 2.605385e-08,
  3.122519e-08, 3.10494e-08, 3.199318e-08, 3.023703e-08, 2.712227e-08, 
    2.792087e-08, 2.850615e-08, 2.989927e-08, 3.052686e-08, 3.106508e-08, 
    3.031457e-08, 2.515223e-08, 2.286266e-08, 2.325221e-08, 2.480195e-08,
  2.778253e-08, 2.860262e-08, 2.783133e-08, 2.971849e-08, 2.799075e-08, 
    2.613718e-08, 2.679004e-08, 2.732556e-08, 2.737812e-08, 2.764669e-08, 
    2.68108e-08, 2.307051e-08, 2.309838e-08, 2.292855e-08, 2.502715e-08,
  2.68778e-08, 2.842865e-08, 2.92821e-08, 2.738354e-08, 2.795181e-08, 
    2.588525e-08, 2.517682e-08, 2.579863e-08, 2.631675e-08, 2.675945e-08, 
    2.494824e-08, 2.306642e-08, 2.243219e-08, 2.205658e-08, 2.61649e-08,
  2.563405e-08, 2.699076e-08, 2.773711e-08, 2.72603e-08, 2.685574e-08, 
    2.68177e-08, 2.500764e-08, 2.443001e-08, 2.553529e-08, 2.66883e-08, 
    2.490109e-08, 2.428365e-08, 2.230024e-08, 2.368371e-08, 2.691221e-08,
  2.375821e-08, 2.675909e-08, 2.712319e-08, 2.756338e-08, 2.80759e-08, 
    2.721715e-08, 2.562109e-08, 2.357725e-08, 2.481989e-08, 2.518591e-08, 
    2.469552e-08, 2.44554e-08, 2.256273e-08, 2.396087e-08, 2.695665e-08,
  2.16452e-08, 2.462031e-08, 2.617603e-08, 2.711387e-08, 2.818044e-08, 
    2.768105e-08, 2.520716e-08, 2.345745e-08, 2.321564e-08, 2.380543e-08, 
    2.415993e-08, 2.295086e-08, 2.295729e-08, 2.46558e-08, 2.63493e-08,
  2.266607e-08, 2.38353e-08, 2.560083e-08, 2.611693e-08, 2.76372e-08, 
    2.838349e-08, 2.926128e-08, 2.850567e-08, 2.802393e-08, 2.82058e-08, 
    2.777877e-08, 2.852462e-08, 2.868287e-08, 2.76118e-08, 2.877416e-08,
  2.190036e-08, 2.242655e-08, 2.443485e-08, 2.453984e-08, 2.608189e-08, 
    2.757571e-08, 2.854512e-08, 2.788916e-08, 2.785104e-08, 2.731138e-08, 
    2.80926e-08, 2.765587e-08, 2.824102e-08, 2.855743e-08, 2.834869e-08,
  2.188983e-08, 2.13274e-08, 2.329099e-08, 2.408144e-08, 2.565325e-08, 
    2.678815e-08, 2.744175e-08, 2.781313e-08, 2.779921e-08, 2.70568e-08, 
    2.743655e-08, 2.615105e-08, 2.771301e-08, 2.896383e-08, 2.642958e-08,
  1.917128e-08, 2.095163e-08, 2.30728e-08, 2.483559e-08, 2.495265e-08, 
    2.554005e-08, 2.665123e-08, 2.820192e-08, 2.927323e-08, 2.886996e-08, 
    2.92875e-08, 3.175944e-08, 3.233352e-08, 2.894284e-08, 2.581021e-08,
  1.922076e-08, 2.011485e-08, 2.273481e-08, 2.495536e-08, 2.462679e-08, 
    2.554579e-08, 2.610112e-08, 2.681811e-08, 2.782537e-08, 2.813295e-08, 
    2.637957e-08, 2.441387e-08, 2.408095e-08, 2.539138e-08, 2.776639e-08,
  1.939817e-08, 2.011299e-08, 2.089082e-08, 2.306437e-08, 2.509904e-08, 
    2.393906e-08, 2.484887e-08, 2.549449e-08, 2.579591e-08, 2.385765e-08, 
    2.266085e-08, 2.424445e-08, 2.649857e-08, 2.526554e-08, 2.65815e-08,
  2.068278e-08, 2.026077e-08, 2.118897e-08, 2.180273e-08, 2.375996e-08, 
    2.430222e-08, 2.430107e-08, 2.430336e-08, 2.38235e-08, 2.324938e-08, 
    2.312574e-08, 2.450337e-08, 2.523848e-08, 2.490849e-08, 2.625855e-08,
  2.092849e-08, 2.031217e-08, 2.042427e-08, 2.158924e-08, 2.395673e-08, 
    2.407951e-08, 2.48823e-08, 2.466456e-08, 2.343989e-08, 2.309177e-08, 
    2.334817e-08, 2.465071e-08, 2.49163e-08, 2.513913e-08, 2.469302e-08,
  2.139102e-08, 2.102968e-08, 2.112613e-08, 2.087293e-08, 2.316502e-08, 
    2.453073e-08, 2.466231e-08, 2.510658e-08, 2.340408e-08, 2.26706e-08, 
    2.30362e-08, 2.452384e-08, 2.443291e-08, 2.363298e-08, 2.44878e-08,
  2.158974e-08, 2.14787e-08, 2.139949e-08, 2.052533e-08, 2.162959e-08, 
    2.39487e-08, 2.545222e-08, 2.554083e-08, 2.340641e-08, 2.295734e-08, 
    2.341165e-08, 2.534231e-08, 2.51026e-08, 2.37963e-08, 2.4194e-08,
  2.049769e-08, 2.084234e-08, 2.055443e-08, 1.995084e-08, 1.997293e-08, 
    2.085849e-08, 2.178875e-08, 2.342797e-08, 2.387298e-08, 2.442228e-08, 
    2.590225e-08, 2.630858e-08, 2.722269e-08, 2.783228e-08, 2.973284e-08,
  2.044077e-08, 2.037761e-08, 2.027159e-08, 1.983202e-08, 2.008566e-08, 
    2.060911e-08, 2.167379e-08, 2.285082e-08, 2.428825e-08, 2.573693e-08, 
    2.53205e-08, 2.5309e-08, 2.633276e-08, 2.703707e-08, 2.736918e-08,
  2.001357e-08, 2.115235e-08, 2.113742e-08, 2.053193e-08, 2.086391e-08, 
    2.119411e-08, 2.151927e-08, 2.284427e-08, 2.441339e-08, 2.419691e-08, 
    2.362204e-08, 2.490133e-08, 2.550688e-08, 2.571295e-08, 2.48592e-08,
  2.065703e-08, 2.160143e-08, 2.125925e-08, 2.169247e-08, 2.176371e-08, 
    2.134194e-08, 2.106247e-08, 2.240819e-08, 2.428524e-08, 2.275507e-08, 
    2.725971e-08, 2.946369e-08, 2.713216e-08, 2.749985e-08, 2.628582e-08,
  2.198335e-08, 2.289076e-08, 2.268918e-08, 2.231886e-08, 2.196238e-08, 
    2.1562e-08, 2.13984e-08, 2.270201e-08, 2.290727e-08, 2.592391e-08, 
    2.415109e-08, 2.470252e-08, 2.496098e-08, 2.673941e-08, 2.698481e-08,
  2.481586e-08, 2.449259e-08, 2.330829e-08, 2.3208e-08, 2.207694e-08, 
    2.169341e-08, 2.181729e-08, 2.181642e-08, 2.317394e-08, 2.328892e-08, 
    2.274353e-08, 2.271515e-08, 2.662023e-08, 2.555255e-08, 2.486733e-08,
  2.536324e-08, 2.462483e-08, 2.401267e-08, 2.344302e-08, 2.283001e-08, 
    2.259181e-08, 2.253292e-08, 2.237259e-08, 2.297823e-08, 2.297677e-08, 
    2.306464e-08, 2.29294e-08, 2.597833e-08, 2.344842e-08, 2.377543e-08,
  2.558158e-08, 2.531115e-08, 2.506087e-08, 2.374951e-08, 2.330093e-08, 
    2.302949e-08, 2.316248e-08, 2.25223e-08, 2.233015e-08, 2.311023e-08, 
    2.317599e-08, 2.331071e-08, 2.552679e-08, 2.434131e-08, 2.561787e-08,
  2.540729e-08, 2.565188e-08, 2.55676e-08, 2.490739e-08, 2.377492e-08, 
    2.366938e-08, 2.373941e-08, 2.32806e-08, 2.276754e-08, 2.315127e-08, 
    2.34794e-08, 2.385884e-08, 2.511807e-08, 2.413726e-08, 2.414002e-08,
  2.503482e-08, 2.564266e-08, 2.575714e-08, 2.514539e-08, 2.485094e-08, 
    2.380332e-08, 2.301188e-08, 2.31084e-08, 2.230463e-08, 2.259981e-08, 
    2.280432e-08, 2.376608e-08, 2.437788e-08, 2.405939e-08, 2.410108e-08,
  2.404712e-08, 2.485562e-08, 2.428088e-08, 2.42691e-08, 2.353266e-08, 
    2.291928e-08, 2.266886e-08, 2.237133e-08, 2.24029e-08, 2.235738e-08, 
    2.257405e-08, 2.172757e-08, 2.208609e-08, 2.092268e-08, 2.134263e-08,
  2.44275e-08, 2.419911e-08, 2.386371e-08, 2.34923e-08, 2.316308e-08, 
    2.27826e-08, 2.317551e-08, 2.258026e-08, 2.274609e-08, 2.260917e-08, 
    2.286351e-08, 2.197561e-08, 2.247079e-08, 2.115769e-08, 2.14197e-08,
  2.468192e-08, 2.706908e-08, 2.727481e-08, 2.458841e-08, 2.325289e-08, 
    2.349402e-08, 2.308078e-08, 2.254467e-08, 2.283385e-08, 2.325324e-08, 
    2.320497e-08, 2.23883e-08, 2.293401e-08, 2.243099e-08, 2.272924e-08,
  2.662261e-08, 2.775072e-08, 2.725373e-08, 2.765528e-08, 2.728579e-08, 
    2.599102e-08, 2.471838e-08, 2.394194e-08, 2.36821e-08, 2.351779e-08, 
    2.282093e-08, 2.336736e-08, 2.367176e-08, 2.396202e-08, 2.457665e-08,
  2.751588e-08, 2.911102e-08, 2.933926e-08, 2.798092e-08, 2.647831e-08, 
    2.504036e-08, 2.416528e-08, 2.352794e-08, 2.329642e-08, 2.24853e-08, 
    2.264399e-08, 2.366897e-08, 2.344279e-08, 2.498358e-08, 2.580786e-08,
  2.891715e-08, 3.053054e-08, 3.133497e-08, 2.906502e-08, 2.76468e-08, 
    2.628092e-08, 2.405832e-08, 2.299523e-08, 2.226761e-08, 2.272735e-08, 
    2.21107e-08, 2.19819e-08, 2.359145e-08, 2.49305e-08, 2.272355e-08,
  2.86419e-08, 3.030598e-08, 3.047833e-08, 2.958259e-08, 2.852799e-08, 
    2.701265e-08, 2.52319e-08, 2.374603e-08, 2.324433e-08, 2.236921e-08, 
    2.281472e-08, 2.20426e-08, 2.407561e-08, 2.446393e-08, 2.296938e-08,
  2.86331e-08, 3.096107e-08, 3.145421e-08, 2.990327e-08, 2.820047e-08, 
    2.707414e-08, 2.623251e-08, 2.453384e-08, 2.396854e-08, 2.257301e-08, 
    2.293319e-08, 2.238165e-08, 2.384727e-08, 2.194028e-08, 2.397225e-08,
  2.853657e-08, 3.082553e-08, 3.165788e-08, 2.97637e-08, 2.845604e-08, 
    2.749973e-08, 2.749801e-08, 2.577602e-08, 2.568478e-08, 2.415936e-08, 
    2.383063e-08, 2.284508e-08, 2.350637e-08, 2.408366e-08, 2.383407e-08,
  2.855579e-08, 3.03117e-08, 3.119985e-08, 2.984695e-08, 2.915128e-08, 
    2.67929e-08, 2.664368e-08, 2.512806e-08, 2.470077e-08, 2.453669e-08, 
    2.448729e-08, 2.40042e-08, 2.318582e-08, 2.330684e-08, 2.36855e-08,
  2.407941e-08, 2.413156e-08, 2.362896e-08, 2.383389e-08, 2.362271e-08, 
    2.350775e-08, 2.333293e-08, 2.318895e-08, 2.301804e-08, 2.272589e-08, 
    2.325392e-08, 2.276261e-08, 2.316629e-08, 2.280625e-08, 2.270717e-08,
  2.457883e-08, 2.495389e-08, 2.465831e-08, 2.421556e-08, 2.365936e-08, 
    2.356836e-08, 2.359773e-08, 2.398165e-08, 2.393781e-08, 2.400089e-08, 
    2.38684e-08, 2.39264e-08, 2.362093e-08, 2.354937e-08, 2.250166e-08,
  2.681297e-08, 2.753249e-08, 2.81686e-08, 2.682102e-08, 2.60966e-08, 
    2.614364e-08, 2.47785e-08, 2.343906e-08, 2.392476e-08, 2.472558e-08, 
    2.490882e-08, 2.505526e-08, 2.469672e-08, 2.460404e-08, 2.296769e-08,
  2.813619e-08, 2.844042e-08, 2.784676e-08, 2.829783e-08, 2.887614e-08, 
    2.946923e-08, 2.807379e-08, 2.647005e-08, 2.558386e-08, 2.567353e-08, 
    2.605954e-08, 2.580407e-08, 2.517332e-08, 2.471239e-08, 2.318671e-08,
  2.978517e-08, 2.9572e-08, 3.148646e-08, 3.119811e-08, 2.984462e-08, 
    2.941649e-08, 2.876247e-08, 2.880554e-08, 2.828613e-08, 2.852824e-08, 
    2.626452e-08, 2.560923e-08, 2.446689e-08, 2.459457e-08, 2.423815e-08,
  2.766822e-08, 2.834912e-08, 3.026466e-08, 3.161069e-08, 3.141574e-08, 
    2.990205e-08, 2.930675e-08, 2.828498e-08, 2.903976e-08, 2.735133e-08, 
    2.494442e-08, 2.480283e-08, 2.47856e-08, 2.478928e-08, 2.418412e-08,
  2.738679e-08, 2.852936e-08, 2.990239e-08, 3.09472e-08, 3.118321e-08, 
    3.165745e-08, 3.093926e-08, 3.002939e-08, 2.842468e-08, 2.631002e-08, 
    2.503403e-08, 2.410431e-08, 2.527196e-08, 2.507421e-08, 2.309636e-08,
  2.591673e-08, 2.714778e-08, 2.873059e-08, 3.108113e-08, 3.011417e-08, 
    3.15777e-08, 3.092609e-08, 3.017179e-08, 2.875605e-08, 2.60064e-08, 
    2.507381e-08, 2.33493e-08, 2.495755e-08, 2.361966e-08, 2.326204e-08,
  2.599113e-08, 2.71882e-08, 2.778234e-08, 3.020694e-08, 2.965782e-08, 
    3.022559e-08, 3.210694e-08, 3.001124e-08, 2.860096e-08, 2.584175e-08, 
    2.509866e-08, 2.326282e-08, 2.420079e-08, 2.38043e-08, 2.371169e-08,
  2.508099e-08, 2.653769e-08, 2.742621e-08, 2.916508e-08, 2.856703e-08, 
    2.679211e-08, 2.822742e-08, 2.650974e-08, 2.753472e-08, 2.684818e-08, 
    2.606531e-08, 2.457089e-08, 2.468673e-08, 2.460925e-08, 2.468337e-08,
  2.589752e-08, 2.645116e-08, 2.745394e-08, 2.738756e-08, 2.691148e-08, 
    2.681696e-08, 2.598101e-08, 2.538947e-08, 2.384584e-08, 2.359084e-08, 
    2.379188e-08, 2.357308e-08, 2.336616e-08, 2.317799e-08, 2.198056e-08,
  2.529251e-08, 2.588754e-08, 2.707723e-08, 2.691626e-08, 2.635033e-08, 
    2.661297e-08, 2.615104e-08, 2.577311e-08, 2.452623e-08, 2.505115e-08, 
    2.510365e-08, 2.451114e-08, 2.367429e-08, 2.290859e-08, 2.151839e-08,
  2.714261e-08, 2.526219e-08, 2.684959e-08, 2.719464e-08, 2.705562e-08, 
    2.735242e-08, 2.625682e-08, 2.511936e-08, 2.44989e-08, 2.514244e-08, 
    2.520271e-08, 2.477121e-08, 2.420653e-08, 2.296344e-08, 2.188997e-08,
  2.658901e-08, 2.562795e-08, 2.659179e-08, 2.784099e-08, 2.833154e-08, 
    2.800038e-08, 2.726709e-08, 2.700226e-08, 2.60574e-08, 2.54862e-08, 
    2.526912e-08, 2.502177e-08, 2.484831e-08, 2.425869e-08, 2.280083e-08,
  2.673266e-08, 2.590863e-08, 2.802767e-08, 2.857445e-08, 2.849258e-08, 
    2.799275e-08, 2.764835e-08, 2.802206e-08, 2.839571e-08, 2.926181e-08, 
    2.632942e-08, 2.458135e-08, 2.352096e-08, 2.337807e-08, 2.330922e-08,
  2.442594e-08, 2.469463e-08, 2.468317e-08, 2.616869e-08, 2.703985e-08, 
    2.739659e-08, 2.784317e-08, 2.80537e-08, 2.936425e-08, 2.811257e-08, 
    2.589352e-08, 2.584277e-08, 2.500801e-08, 2.327408e-08, 2.405569e-08,
  2.37419e-08, 2.474632e-08, 2.538445e-08, 2.600408e-08, 2.670557e-08, 
    2.686218e-08, 2.760368e-08, 2.897329e-08, 2.828478e-08, 2.62455e-08, 
    2.619234e-08, 2.647547e-08, 2.574906e-08, 2.48859e-08, 2.622813e-08,
  2.337492e-08, 2.488246e-08, 2.49959e-08, 2.506297e-08, 2.553283e-08, 
    2.600734e-08, 2.558573e-08, 2.598301e-08, 2.546917e-08, 2.648056e-08, 
    2.694982e-08, 2.645147e-08, 2.618436e-08, 2.649553e-08, 2.640491e-08,
  2.356531e-08, 2.50582e-08, 2.562641e-08, 2.52053e-08, 2.552831e-08, 
    2.542112e-08, 2.510733e-08, 2.433357e-08, 2.573839e-08, 2.600688e-08, 
    2.664464e-08, 2.64681e-08, 2.645373e-08, 2.648646e-08, 2.587773e-08,
  2.438559e-08, 2.5297e-08, 2.528889e-08, 2.483417e-08, 2.436523e-08, 
    2.463332e-08, 2.369646e-08, 2.34952e-08, 2.421036e-08, 2.434476e-08, 
    2.548427e-08, 2.537647e-08, 2.585092e-08, 2.592739e-08, 2.553745e-08,
  1.970406e-08, 2.066523e-08, 2.135742e-08, 2.172315e-08, 2.196611e-08, 
    2.272135e-08, 2.363033e-08, 2.539891e-08, 2.535033e-08, 2.606674e-08, 
    2.714362e-08, 2.623382e-08, 2.544181e-08, 2.529269e-08, 2.47985e-08,
  2.039397e-08, 2.062649e-08, 2.17408e-08, 2.178193e-08, 2.18917e-08, 
    2.244393e-08, 2.367601e-08, 2.469698e-08, 2.485376e-08, 2.587331e-08, 
    2.704649e-08, 2.774775e-08, 2.677113e-08, 2.570563e-08, 2.322507e-08,
  2.262397e-08, 2.215227e-08, 2.205609e-08, 2.164106e-08, 2.272659e-08, 
    2.295113e-08, 2.309483e-08, 2.388989e-08, 2.444083e-08, 2.490622e-08, 
    2.579132e-08, 2.708796e-08, 2.78838e-08, 2.658584e-08, 2.467705e-08,
  2.360216e-08, 2.335055e-08, 2.279583e-08, 2.225645e-08, 2.34314e-08, 
    2.35083e-08, 2.291013e-08, 2.360304e-08, 2.412325e-08, 2.476366e-08, 
    2.622842e-08, 2.692647e-08, 2.732783e-08, 2.62339e-08, 2.479135e-08,
  2.349529e-08, 2.332391e-08, 2.286807e-08, 2.39356e-08, 2.352361e-08, 
    2.412176e-08, 2.380654e-08, 2.40145e-08, 2.381394e-08, 2.53136e-08, 
    2.592806e-08, 2.667388e-08, 2.606067e-08, 2.525802e-08, 2.436573e-08,
  2.421804e-08, 2.482849e-08, 2.462852e-08, 2.484389e-08, 2.43942e-08, 
    2.413099e-08, 2.367599e-08, 2.337134e-08, 2.35385e-08, 2.390416e-08, 
    2.427305e-08, 2.546138e-08, 2.537198e-08, 2.453686e-08, 2.696452e-08,
  2.583838e-08, 2.709287e-08, 2.794996e-08, 2.684786e-08, 2.606055e-08, 
    2.504317e-08, 2.42973e-08, 2.3437e-08, 2.340871e-08, 2.318134e-08, 
    2.352964e-08, 2.359417e-08, 2.478641e-08, 2.590102e-08, 2.826202e-08,
  2.891898e-08, 3.088138e-08, 3.122293e-08, 2.986322e-08, 2.834311e-08, 
    2.652823e-08, 2.541608e-08, 2.437897e-08, 2.395077e-08, 2.360874e-08, 
    2.364804e-08, 2.297161e-08, 2.425426e-08, 2.446038e-08, 2.490404e-08,
  2.511518e-08, 2.839498e-08, 3.08827e-08, 3.244799e-08, 3.138809e-08, 
    2.935188e-08, 2.739136e-08, 2.620449e-08, 2.549243e-08, 2.44358e-08, 
    2.368649e-08, 2.306811e-08, 2.403027e-08, 2.387762e-08, 2.385017e-08,
  2.537634e-08, 2.281597e-08, 2.496495e-08, 2.684308e-08, 2.759059e-08, 
    2.900004e-08, 2.923649e-08, 2.940664e-08, 2.97997e-08, 2.698471e-08, 
    2.474323e-08, 2.276708e-08, 2.326693e-08, 2.310152e-08, 2.310692e-08,
  2.30149e-08, 2.226203e-08, 2.188695e-08, 2.270883e-08, 2.220836e-08, 
    2.217015e-08, 2.181429e-08, 2.236281e-08, 2.244421e-08, 2.263283e-08, 
    2.283309e-08, 2.22158e-08, 2.260329e-08, 2.206414e-08, 2.360903e-08,
  2.714326e-08, 2.740688e-08, 2.565472e-08, 2.597575e-08, 2.344111e-08, 
    2.290903e-08, 2.217422e-08, 2.28433e-08, 2.335481e-08, 2.306086e-08, 
    2.330975e-08, 2.308909e-08, 2.322104e-08, 2.322656e-08, 2.321053e-08,
  2.961209e-08, 3.000001e-08, 2.761043e-08, 2.650489e-08, 2.608916e-08, 
    2.45761e-08, 2.270936e-08, 2.24704e-08, 2.333137e-08, 2.384594e-08, 
    2.403485e-08, 2.371847e-08, 2.340684e-08, 2.390859e-08, 2.300446e-08,
  2.975331e-08, 3.10879e-08, 2.965466e-08, 2.770348e-08, 2.630913e-08, 
    2.549083e-08, 2.400097e-08, 2.293224e-08, 2.327551e-08, 2.392001e-08, 
    2.399866e-08, 2.398144e-08, 2.354068e-08, 2.382254e-08, 2.258995e-08,
  2.574792e-08, 2.78059e-08, 2.683994e-08, 2.547238e-08, 2.432442e-08, 
    2.5362e-08, 2.582776e-08, 2.576503e-08, 2.466793e-08, 2.53664e-08, 
    2.464642e-08, 2.477392e-08, 2.399919e-08, 2.362761e-08, 2.267517e-08,
  2.473574e-08, 2.568138e-08, 2.745473e-08, 2.730517e-08, 2.537111e-08, 
    2.46805e-08, 2.491339e-08, 2.670397e-08, 2.752729e-08, 2.712795e-08, 
    2.599241e-08, 2.503297e-08, 2.477956e-08, 2.364865e-08, 2.324272e-08,
  2.321955e-08, 2.4744e-08, 2.70472e-08, 2.800187e-08, 2.831914e-08, 
    2.715346e-08, 2.551907e-08, 2.631106e-08, 2.713277e-08, 2.759182e-08, 
    2.768037e-08, 2.617645e-08, 2.556347e-08, 2.345119e-08, 2.379241e-08,
  2.093253e-08, 2.437069e-08, 2.720732e-08, 2.807104e-08, 2.852796e-08, 
    2.800765e-08, 2.757207e-08, 2.793404e-08, 2.823543e-08, 2.838958e-08, 
    2.926277e-08, 2.840764e-08, 2.738598e-08, 2.515179e-08, 2.438148e-08,
  2.025909e-08, 2.334224e-08, 2.731726e-08, 3.016586e-08, 3.055707e-08, 
    3.121871e-08, 3.052895e-08, 2.976702e-08, 2.843069e-08, 2.821244e-08, 
    2.939989e-08, 2.904988e-08, 2.851284e-08, 2.683412e-08, 2.557167e-08,
  1.939739e-08, 2.202993e-08, 2.554139e-08, 3.000327e-08, 3.16845e-08, 
    3.231655e-08, 3.495013e-08, 3.197814e-08, 2.925746e-08, 2.91701e-08, 
    2.961949e-08, 2.880143e-08, 2.811786e-08, 2.690461e-08, 2.605494e-08,
  2.283376e-08, 2.263366e-08, 2.280994e-08, 2.346127e-08, 2.321966e-08, 
    2.312203e-08, 2.326258e-08, 2.302816e-08, 2.279497e-08, 2.077315e-08, 
    2.047165e-08, 2.151318e-08, 2.469003e-08, 2.40108e-08, 2.29853e-08,
  2.471596e-08, 2.669799e-08, 2.605749e-08, 2.718976e-08, 2.800782e-08, 
    2.694892e-08, 2.471279e-08, 2.403467e-08, 2.294845e-08, 2.118253e-08, 
    1.881918e-08, 1.788411e-08, 1.862912e-08, 2.150688e-08, 2.188028e-08,
  2.83791e-08, 2.924933e-08, 3.005359e-08, 3.057559e-08, 3.040376e-08, 
    3.050026e-08, 2.984025e-08, 2.795576e-08, 2.687917e-08, 2.321594e-08, 
    2.078143e-08, 1.875606e-08, 1.733481e-08, 1.89401e-08, 2.005147e-08,
  3.079137e-08, 2.907193e-08, 2.979609e-08, 3.136186e-08, 3.025958e-08, 
    2.858507e-08, 2.891434e-08, 2.728064e-08, 2.569128e-08, 2.368843e-08, 
    2.031203e-08, 2.020001e-08, 1.989589e-08, 1.870556e-08, 1.924778e-08,
  2.828066e-08, 2.684183e-08, 2.72241e-08, 2.661744e-08, 2.801621e-08, 
    2.86272e-08, 3.047813e-08, 2.942165e-08, 2.665099e-08, 2.442086e-08, 
    2.350808e-08, 2.213785e-08, 2.106295e-08, 2.150647e-08, 2.169831e-08,
  2.418525e-08, 2.123935e-08, 2.33415e-08, 2.174807e-08, 2.260793e-08, 
    2.406879e-08, 2.42031e-08, 2.655988e-08, 2.610671e-08, 2.325462e-08, 
    2.577525e-08, 2.40972e-08, 2.304955e-08, 2.301887e-08, 2.446579e-08,
  2.236775e-08, 1.940905e-08, 1.997042e-08, 2.021455e-08, 1.885844e-08, 
    1.978004e-08, 2.108682e-08, 2.177501e-08, 2.236438e-08, 2.269782e-08, 
    2.573411e-08, 2.625876e-08, 2.563511e-08, 2.423948e-08, 2.62819e-08,
  2.3403e-08, 2.111912e-08, 1.660409e-08, 1.712477e-08, 1.782228e-08, 
    1.698563e-08, 1.857468e-08, 1.965569e-08, 1.967164e-08, 1.988458e-08, 
    2.15926e-08, 2.403175e-08, 2.442506e-08, 2.491417e-08, 2.730348e-08,
  2.254186e-08, 2.102986e-08, 1.707879e-08, 1.373312e-08, 1.481189e-08, 
    1.495612e-08, 1.501091e-08, 1.759568e-08, 1.586765e-08, 1.691411e-08, 
    1.806449e-08, 1.95386e-08, 2.096016e-08, 2.33861e-08, 2.433103e-08,
  1.840674e-08, 1.76381e-08, 1.658995e-08, 1.377808e-08, 1.264639e-08, 
    1.2239e-08, 1.368432e-08, 1.583635e-08, 1.645275e-08, 1.787086e-08, 
    1.824539e-08, 1.839617e-08, 1.993377e-08, 1.965301e-08, 2.15028e-08,
  2.552235e-08, 2.620712e-08, 2.610934e-08, 2.607311e-08, 2.627919e-08, 
    2.627513e-08, 2.64217e-08, 2.644418e-08, 2.659742e-08, 2.722005e-08, 
    2.660754e-08, 2.760465e-08, 2.771333e-08, 2.710032e-08, 2.596893e-08,
  2.625948e-08, 2.721458e-08, 2.717131e-08, 2.740095e-08, 2.712368e-08, 
    2.651552e-08, 2.661276e-08, 2.658428e-08, 2.673436e-08, 2.774647e-08, 
    2.81158e-08, 2.770966e-08, 2.978738e-08, 2.98729e-08, 2.893271e-08,
  2.7869e-08, 2.92828e-08, 2.910948e-08, 2.906664e-08, 2.886517e-08, 
    2.833973e-08, 2.728971e-08, 2.684427e-08, 2.813589e-08, 2.784848e-08, 
    2.880539e-08, 2.828029e-08, 2.907432e-08, 2.874034e-08, 2.923334e-08,
  2.857443e-08, 2.87567e-08, 2.887061e-08, 2.85149e-08, 2.754512e-08, 
    2.729005e-08, 2.628136e-08, 2.465069e-08, 2.327171e-08, 2.407593e-08, 
    2.470825e-08, 2.557473e-08, 2.753519e-08, 2.706617e-08, 2.941931e-08,
  2.76587e-08, 2.790993e-08, 2.73294e-08, 2.693448e-08, 2.660033e-08, 
    2.643105e-08, 2.663981e-08, 2.558759e-08, 2.273882e-08, 2.326113e-08, 
    2.211195e-08, 2.172706e-08, 2.239525e-08, 2.392827e-08, 2.598211e-08,
  2.582467e-08, 2.618461e-08, 2.522884e-08, 2.469811e-08, 2.49656e-08, 
    2.544794e-08, 2.68039e-08, 2.64557e-08, 2.529333e-08, 2.173327e-08, 
    2.361691e-08, 2.347489e-08, 2.215763e-08, 2.367327e-08, 2.377484e-08,
  2.45377e-08, 2.481678e-08, 2.35437e-08, 2.30155e-08, 2.281386e-08, 
    2.359565e-08, 2.606016e-08, 2.580292e-08, 2.629421e-08, 2.530438e-08, 
    2.4634e-08, 2.365464e-08, 2.254129e-08, 2.352662e-08, 2.419694e-08,
  2.390695e-08, 2.465916e-08, 2.456048e-08, 2.359849e-08, 2.321408e-08, 
    2.450199e-08, 2.481188e-08, 2.502456e-08, 2.543578e-08, 2.486887e-08, 
    2.443191e-08, 2.417258e-08, 2.447136e-08, 2.059255e-08, 2.208183e-08,
  2.323669e-08, 2.537205e-08, 2.616371e-08, 2.442858e-08, 2.318068e-08, 
    2.26583e-08, 2.278673e-08, 2.206308e-08, 2.018977e-08, 2.305258e-08, 
    2.321762e-08, 2.297239e-08, 2.333004e-08, 2.017885e-08, 1.99244e-08,
  2.484465e-08, 2.546871e-08, 2.579748e-08, 2.47332e-08, 2.262938e-08, 
    2.139644e-08, 2.063725e-08, 1.948096e-08, 1.851397e-08, 1.844889e-08, 
    1.793678e-08, 1.838308e-08, 1.892063e-08, 1.777096e-08, 1.750425e-08,
  2.306514e-08, 2.46259e-08, 2.627662e-08, 2.406985e-08, 2.365027e-08, 
    2.321405e-08, 2.262735e-08, 2.280351e-08, 2.319167e-08, 2.233813e-08, 
    2.198617e-08, 2.183606e-08, 2.207993e-08, 2.198088e-08, 2.077235e-08,
  2.211627e-08, 2.387835e-08, 2.45715e-08, 2.541722e-08, 2.341771e-08, 
    2.212243e-08, 2.191746e-08, 2.243744e-08, 2.221426e-08, 2.268801e-08, 
    2.287016e-08, 2.28955e-08, 2.303956e-08, 2.246977e-08, 2.128976e-08,
  2.925092e-08, 2.576087e-08, 2.71421e-08, 2.569311e-08, 2.377923e-08, 
    2.411844e-08, 2.437628e-08, 2.452521e-08, 2.380186e-08, 2.371906e-08, 
    2.41968e-08, 2.43096e-08, 2.518846e-08, 2.445977e-08, 2.493723e-08,
  3.439091e-08, 2.993712e-08, 2.850208e-08, 2.737777e-08, 2.739561e-08, 
    2.650031e-08, 2.555348e-08, 2.622259e-08, 2.571594e-08, 2.514659e-08, 
    2.623546e-08, 2.671989e-08, 2.72149e-08, 2.629768e-08, 2.71564e-08,
  3.423979e-08, 3.149934e-08, 3.335199e-08, 3.294483e-08, 2.933936e-08, 
    2.731316e-08, 2.727041e-08, 2.782271e-08, 2.707902e-08, 2.809859e-08, 
    2.637685e-08, 2.611523e-08, 2.602655e-08, 2.649973e-08, 2.783529e-08,
  3.116523e-08, 3.059985e-08, 3.031257e-08, 3.080308e-08, 2.972202e-08, 
    2.836121e-08, 2.766156e-08, 2.700959e-08, 2.770764e-08, 2.57279e-08, 
    2.435821e-08, 2.458403e-08, 2.493941e-08, 2.55123e-08, 2.822684e-08,
  2.875917e-08, 2.866793e-08, 3.028871e-08, 3.193108e-08, 2.997357e-08, 
    2.710007e-08, 2.702819e-08, 2.653073e-08, 2.713579e-08, 2.510703e-08, 
    2.469264e-08, 2.435318e-08, 2.442848e-08, 2.542378e-08, 2.655196e-08,
  2.62645e-08, 2.766603e-08, 2.91195e-08, 3.111061e-08, 2.980817e-08, 
    2.850982e-08, 2.709407e-08, 2.56062e-08, 2.633321e-08, 2.605888e-08, 
    2.59354e-08, 2.469884e-08, 2.49822e-08, 2.583047e-08, 2.514028e-08,
  2.527589e-08, 2.557828e-08, 2.731412e-08, 2.909368e-08, 2.929719e-08, 
    3.017115e-08, 2.872229e-08, 2.588378e-08, 2.417235e-08, 2.651785e-08, 
    2.766188e-08, 2.628539e-08, 2.63765e-08, 2.543781e-08, 2.307238e-08,
  2.491599e-08, 2.464968e-08, 2.479649e-08, 2.653773e-08, 2.798288e-08, 
    3.113979e-08, 3.018413e-08, 2.538455e-08, 2.393049e-08, 2.772423e-08, 
    3.026552e-08, 2.823679e-08, 2.695126e-08, 2.325876e-08, 2.088771e-08,
  2.530296e-08, 2.543125e-08, 2.540174e-08, 2.545025e-08, 2.657083e-08, 
    2.678647e-08, 2.703698e-08, 2.751251e-08, 2.619644e-08, 2.515751e-08, 
    2.460546e-08, 2.568487e-08, 2.717895e-08, 2.590621e-08, 2.530098e-08,
  2.474022e-08, 2.582449e-08, 2.639416e-08, 2.818908e-08, 2.938793e-08, 
    2.877722e-08, 2.90157e-08, 2.82255e-08, 2.836517e-08, 2.804576e-08, 
    2.659967e-08, 2.561884e-08, 2.415754e-08, 2.206347e-08, 2.112517e-08,
  2.81137e-08, 2.954522e-08, 3.027712e-08, 3.111528e-08, 3.193417e-08, 
    3.003525e-08, 2.972476e-08, 2.975559e-08, 3.056681e-08, 3.031539e-08, 
    3.086904e-08, 3.006217e-08, 2.6923e-08, 2.390625e-08, 2.156087e-08,
  2.863653e-08, 2.949219e-08, 3.218143e-08, 3.359519e-08, 3.179106e-08, 
    2.960422e-08, 2.876412e-08, 3.022209e-08, 3.320712e-08, 3.521713e-08, 
    3.947656e-08, 3.777971e-08, 3.461837e-08, 2.959698e-08, 2.504019e-08,
  2.773727e-08, 2.796411e-08, 3.155603e-08, 3.15619e-08, 2.92424e-08, 
    2.856999e-08, 2.871204e-08, 3.049551e-08, 3.358772e-08, 3.469713e-08, 
    3.352217e-08, 3.50607e-08, 3.532179e-08, 2.813604e-08, 2.362072e-08,
  2.766442e-08, 2.78071e-08, 2.763072e-08, 2.899573e-08, 2.953555e-08, 
    2.865267e-08, 2.802354e-08, 2.784694e-08, 2.813017e-08, 3.168047e-08, 
    2.852767e-08, 2.834962e-08, 3.356907e-08, 2.679949e-08, 2.489756e-08,
  2.782946e-08, 2.683292e-08, 2.550519e-08, 2.590161e-08, 3.007954e-08, 
    2.941872e-08, 2.833408e-08, 2.749223e-08, 2.7491e-08, 2.893653e-08, 
    2.892511e-08, 2.964757e-08, 3.258776e-08, 2.867389e-08, 3.067596e-08,
  2.72027e-08, 2.626178e-08, 2.548949e-08, 2.607725e-08, 2.919651e-08, 
    2.886647e-08, 2.970975e-08, 2.776097e-08, 2.578087e-08, 2.66158e-08, 
    2.714642e-08, 2.870439e-08, 3.066004e-08, 3.250497e-08, 3.142705e-08,
  2.807097e-08, 2.665744e-08, 2.620838e-08, 2.676176e-08, 2.775013e-08, 
    2.853464e-08, 3.078942e-08, 2.848724e-08, 2.729658e-08, 2.700462e-08, 
    2.704717e-08, 2.728604e-08, 2.799314e-08, 2.987164e-08, 2.784993e-08,
  2.857171e-08, 2.603798e-08, 2.537095e-08, 2.595575e-08, 2.602674e-08, 
    2.768407e-08, 3.072861e-08, 2.882171e-08, 2.853282e-08, 2.577183e-08, 
    2.501609e-08, 2.585096e-08, 2.721748e-08, 2.801491e-08, 2.792689e-08,
  2.274956e-08, 2.523672e-08, 2.436366e-08, 2.36598e-08, 2.349142e-08, 
    2.450886e-08, 2.559599e-08, 2.627322e-08, 2.603043e-08, 2.659257e-08, 
    2.700787e-08, 2.70083e-08, 2.884615e-08, 2.819841e-08, 2.766163e-08,
  2.286716e-08, 2.434677e-08, 2.431636e-08, 2.335873e-08, 2.370656e-08, 
    2.462545e-08, 2.504712e-08, 2.584312e-08, 2.612119e-08, 2.661358e-08, 
    2.65881e-08, 2.672441e-08, 2.730976e-08, 2.657191e-08, 2.593687e-08,
  2.562185e-08, 2.576727e-08, 2.463847e-08, 2.406913e-08, 2.291948e-08, 
    2.296342e-08, 2.316363e-08, 2.32765e-08, 2.405612e-08, 2.472101e-08, 
    2.421014e-08, 2.527423e-08, 2.583378e-08, 2.593098e-08, 2.595737e-08,
  2.784269e-08, 2.640285e-08, 2.432046e-08, 2.221407e-08, 2.103203e-08, 
    2.248498e-08, 2.257907e-08, 2.143472e-08, 2.112398e-08, 2.128948e-08, 
    1.96923e-08, 2.05112e-08, 2.303219e-08, 2.541034e-08, 2.840192e-08,
  2.838968e-08, 2.539585e-08, 2.225464e-08, 2.032841e-08, 2.06538e-08, 
    2.279384e-08, 2.215063e-08, 2.031028e-08, 2.052452e-08, 1.88487e-08, 
    1.814906e-08, 2.142664e-08, 2.325319e-08, 2.519643e-08, 2.885166e-08,
  2.662731e-08, 2.288239e-08, 2.039218e-08, 2.076576e-08, 2.249477e-08, 
    2.350007e-08, 2.198697e-08, 2.157988e-08, 2.06289e-08, 1.975009e-08, 
    2.269419e-08, 2.468206e-08, 2.523213e-08, 2.568783e-08, 2.784482e-08,
  2.487438e-08, 2.159654e-08, 2.037898e-08, 2.167629e-08, 2.24277e-08, 
    2.149768e-08, 2.122996e-08, 2.072792e-08, 1.95714e-08, 2.08399e-08, 
    2.262513e-08, 2.404547e-08, 2.501717e-08, 2.672395e-08, 2.669652e-08,
  2.389205e-08, 2.20972e-08, 2.121796e-08, 2.19848e-08, 2.210408e-08, 
    2.216405e-08, 2.307101e-08, 2.081425e-08, 2.041397e-08, 2.190895e-08, 
    2.345043e-08, 2.463991e-08, 2.511434e-08, 2.517317e-08, 2.421164e-08,
  2.415123e-08, 2.338754e-08, 2.226257e-08, 2.18985e-08, 2.113942e-08, 
    2.230156e-08, 2.163793e-08, 2.016142e-08, 2.195056e-08, 2.379537e-08, 
    2.475376e-08, 2.513046e-08, 2.60411e-08, 2.572718e-08, 2.45082e-08,
  2.453105e-08, 2.472407e-08, 2.244905e-08, 2.010895e-08, 1.966671e-08, 
    2.054445e-08, 2.030335e-08, 2.153823e-08, 2.449782e-08, 2.529422e-08, 
    2.592273e-08, 2.593227e-08, 2.651115e-08, 2.632999e-08, 2.598322e-08,
  1.605045e-08, 1.661041e-08, 1.721056e-08, 1.719374e-08, 1.679131e-08, 
    1.716275e-08, 1.823236e-08, 1.949248e-08, 2.002556e-08, 1.951746e-08, 
    1.807194e-08, 1.719421e-08, 1.767588e-08, 1.777807e-08, 1.810415e-08,
  1.722556e-08, 1.750353e-08, 1.754655e-08, 1.766663e-08, 1.762975e-08, 
    1.818331e-08, 1.893066e-08, 2.050194e-08, 2.058694e-08, 2.013509e-08, 
    1.917662e-08, 1.887243e-08, 1.873708e-08, 1.814457e-08, 1.884105e-08,
  1.899908e-08, 1.803206e-08, 1.785678e-08, 1.863797e-08, 1.868852e-08, 
    1.898724e-08, 1.938102e-08, 2.071124e-08, 2.038931e-08, 1.98209e-08, 
    1.942767e-08, 1.945337e-08, 1.910376e-08, 1.903888e-08, 2.195875e-08,
  1.917585e-08, 1.813593e-08, 1.829935e-08, 1.857917e-08, 1.807115e-08, 
    1.804094e-08, 1.907316e-08, 2.011813e-08, 2.005192e-08, 1.884621e-08, 
    1.88178e-08, 1.901341e-08, 1.910666e-08, 2.126135e-08, 2.414202e-08,
  1.92802e-08, 1.847171e-08, 1.906596e-08, 1.84757e-08, 1.830175e-08, 
    1.800174e-08, 1.863293e-08, 1.933929e-08, 1.829483e-08, 1.818276e-08, 
    1.858431e-08, 2.011839e-08, 2.133444e-08, 2.403434e-08, 2.296315e-08,
  1.926883e-08, 1.958475e-08, 1.975653e-08, 1.902394e-08, 1.908795e-08, 
    1.824414e-08, 1.899586e-08, 1.86253e-08, 1.870985e-08, 1.956161e-08, 
    2.12437e-08, 2.132481e-08, 2.30938e-08, 2.448565e-08, 2.26669e-08,
  1.964336e-08, 2.014216e-08, 2.011544e-08, 2.0156e-08, 1.967013e-08, 
    1.921016e-08, 1.952217e-08, 1.908846e-08, 1.911106e-08, 2.061315e-08, 
    2.165241e-08, 2.160019e-08, 2.421828e-08, 2.443847e-08, 2.239427e-08,
  1.980862e-08, 2.072918e-08, 2.116346e-08, 2.146683e-08, 2.075733e-08, 
    2.052617e-08, 2.043143e-08, 1.969619e-08, 1.970791e-08, 2.071537e-08, 
    2.172689e-08, 2.2266e-08, 2.458181e-08, 2.282077e-08, 2.22162e-08,
  2.122801e-08, 2.204103e-08, 2.212427e-08, 2.232481e-08, 2.174726e-08, 
    2.145365e-08, 2.036071e-08, 1.963915e-08, 1.961557e-08, 2.083901e-08, 
    2.168146e-08, 2.207396e-08, 2.300813e-08, 2.347758e-08, 2.277062e-08,
  2.187901e-08, 2.162471e-08, 2.18232e-08, 2.214813e-08, 2.220854e-08, 
    2.175924e-08, 2.024654e-08, 1.980384e-08, 2.048603e-08, 2.065861e-08, 
    2.107867e-08, 2.18214e-08, 2.295011e-08, 2.314469e-08, 2.352934e-08,
  1.876797e-08, 2.007125e-08, 2.088989e-08, 2.255072e-08, 2.395311e-08, 
    2.451508e-08, 2.310217e-08, 2.288079e-08, 2.141539e-08, 2.056962e-08, 
    1.976857e-08, 1.956065e-08, 1.954804e-08, 1.969353e-08, 1.956771e-08,
  2.013729e-08, 2.149601e-08, 2.151789e-08, 2.371082e-08, 2.506756e-08, 
    2.405089e-08, 2.214206e-08, 2.229442e-08, 2.113462e-08, 2.053262e-08, 
    2.009568e-08, 2.014148e-08, 2.024263e-08, 2.031788e-08, 2.021673e-08,
  2.187352e-08, 2.102421e-08, 2.132497e-08, 2.349788e-08, 2.224411e-08, 
    2.073507e-08, 2.016291e-08, 2.193486e-08, 2.211899e-08, 2.129565e-08, 
    2.111654e-08, 2.109466e-08, 2.108902e-08, 2.080155e-08, 2.104893e-08,
  2.038833e-08, 2.052363e-08, 2.138663e-08, 2.242522e-08, 2.117748e-08, 
    2.065672e-08, 2.100517e-08, 2.206101e-08, 2.175579e-08, 2.138218e-08, 
    2.135875e-08, 2.172687e-08, 2.160741e-08, 2.136076e-08, 2.165748e-08,
  2.030054e-08, 2.085005e-08, 2.257546e-08, 2.234714e-08, 2.125013e-08, 
    2.08342e-08, 2.11582e-08, 2.206361e-08, 2.153051e-08, 2.088193e-08, 
    2.116624e-08, 2.1553e-08, 2.083449e-08, 2.118399e-08, 2.164617e-08,
  2.16136e-08, 2.271459e-08, 2.339123e-08, 2.281252e-08, 2.232722e-08, 
    2.213397e-08, 2.231367e-08, 2.270567e-08, 2.130518e-08, 2.060139e-08, 
    2.187781e-08, 2.172884e-08, 2.102926e-08, 2.098012e-08, 2.156378e-08,
  2.278191e-08, 2.292982e-08, 2.241044e-08, 2.27785e-08, 2.38858e-08, 
    2.335405e-08, 2.368606e-08, 2.218257e-08, 2.133131e-08, 2.100724e-08, 
    2.155619e-08, 2.185669e-08, 2.159496e-08, 2.140938e-08, 2.074217e-08,
  2.32113e-08, 2.239008e-08, 2.213838e-08, 2.363608e-08, 2.543727e-08, 
    2.418933e-08, 2.426977e-08, 2.244102e-08, 2.221609e-08, 2.186239e-08, 
    2.231075e-08, 2.267022e-08, 2.250379e-08, 2.200974e-08, 2.081703e-08,
  2.226874e-08, 2.179913e-08, 2.212288e-08, 2.466468e-08, 2.542669e-08, 
    2.445202e-08, 2.416739e-08, 2.284691e-08, 2.249145e-08, 2.29872e-08, 
    2.31853e-08, 2.337655e-08, 2.344386e-08, 2.28594e-08, 2.185383e-08,
  2.201467e-08, 2.195081e-08, 2.267768e-08, 2.333047e-08, 2.329264e-08, 
    2.324564e-08, 2.3059e-08, 2.343501e-08, 2.443335e-08, 2.430048e-08, 
    2.396809e-08, 2.385104e-08, 2.385142e-08, 2.333771e-08, 2.253419e-08,
  2.034815e-08, 2.092576e-08, 2.160182e-08, 2.200337e-08, 2.22816e-08, 
    2.184134e-08, 2.156969e-08, 2.148654e-08, 2.167114e-08, 2.106405e-08, 
    2.110397e-08, 2.076978e-08, 2.164901e-08, 2.112666e-08, 2.067702e-08,
  2.168151e-08, 2.267165e-08, 2.269205e-08, 2.290829e-08, 2.301441e-08, 
    2.225903e-08, 2.142081e-08, 2.149544e-08, 2.157017e-08, 2.11994e-08, 
    2.064393e-08, 2.052746e-08, 2.079971e-08, 2.05271e-08, 2.048071e-08,
  2.372723e-08, 2.31187e-08, 2.261692e-08, 2.302171e-08, 2.296438e-08, 
    2.234781e-08, 2.203127e-08, 2.142756e-08, 2.185711e-08, 2.074422e-08, 
    2.033867e-08, 2.040823e-08, 2.033245e-08, 2.010717e-08, 2.115965e-08,
  2.324066e-08, 2.266238e-08, 2.273986e-08, 2.320238e-08, 2.289695e-08, 
    2.301001e-08, 2.355389e-08, 2.335727e-08, 2.239931e-08, 2.118253e-08, 
    1.93548e-08, 1.834164e-08, 1.877798e-08, 1.883043e-08, 2.120894e-08,
  2.362336e-08, 2.3089e-08, 2.299966e-08, 2.290051e-08, 2.313539e-08, 
    2.304595e-08, 2.338146e-08, 2.301381e-08, 2.134307e-08, 1.865471e-08, 
    1.826009e-08, 1.835802e-08, 1.847168e-08, 2.022272e-08, 2.247164e-08,
  2.402121e-08, 2.323138e-08, 2.326414e-08, 2.362878e-08, 2.386558e-08, 
    2.411375e-08, 2.379345e-08, 2.314648e-08, 2.103726e-08, 1.988183e-08, 
    2.190195e-08, 2.157014e-08, 2.01489e-08, 2.209188e-08, 2.259961e-08,
  2.38307e-08, 2.32927e-08, 2.401579e-08, 2.415387e-08, 2.428609e-08, 
    2.511482e-08, 2.481024e-08, 2.440582e-08, 2.296477e-08, 2.380539e-08, 
    2.396976e-08, 2.299444e-08, 2.210463e-08, 2.267679e-08, 2.107658e-08,
  2.391234e-08, 2.441752e-08, 2.489917e-08, 2.43641e-08, 2.494786e-08, 
    2.600758e-08, 2.576513e-08, 2.533203e-08, 2.420273e-08, 2.47661e-08, 
    2.439481e-08, 2.364009e-08, 2.29884e-08, 2.195931e-08, 1.932128e-08,
  2.467555e-08, 2.5519e-08, 2.556464e-08, 2.48181e-08, 2.509977e-08, 
    2.499416e-08, 2.465798e-08, 2.406401e-08, 2.392079e-08, 2.583919e-08, 
    2.578925e-08, 2.484125e-08, 2.423896e-08, 2.311512e-08, 2.124599e-08,
  2.525e-08, 2.590662e-08, 2.592133e-08, 2.486537e-08, 2.458513e-08, 
    2.388354e-08, 2.414331e-08, 2.453611e-08, 2.599723e-08, 2.719696e-08, 
    2.710549e-08, 2.623686e-08, 2.564633e-08, 2.462804e-08, 2.381681e-08,
  2.204298e-08, 2.233367e-08, 2.256969e-08, 2.317621e-08, 2.354126e-08, 
    2.376536e-08, 2.402124e-08, 2.365212e-08, 2.399882e-08, 2.278686e-08, 
    2.273542e-08, 2.266545e-08, 2.389406e-08, 2.398619e-08, 2.457497e-08,
  2.258506e-08, 2.322429e-08, 2.340591e-08, 2.334508e-08, 2.394482e-08, 
    2.383427e-08, 2.400029e-08, 2.424762e-08, 2.311064e-08, 2.287599e-08, 
    2.153568e-08, 2.076934e-08, 1.909189e-08, 1.917739e-08, 2.009673e-08,
  2.299985e-08, 2.413015e-08, 2.395169e-08, 2.399113e-08, 2.432027e-08, 
    2.445239e-08, 2.434281e-08, 2.441046e-08, 2.484603e-08, 2.343942e-08, 
    2.298916e-08, 2.176423e-08, 2.051861e-08, 1.917027e-08, 1.966214e-08,
  2.28402e-08, 2.368448e-08, 2.432154e-08, 2.489127e-08, 2.46671e-08, 
    2.450042e-08, 2.452415e-08, 2.487126e-08, 2.535112e-08, 2.516037e-08, 
    2.39301e-08, 2.36381e-08, 2.317423e-08, 2.209188e-08, 2.188735e-08,
  2.33714e-08, 2.43307e-08, 2.452812e-08, 2.4004e-08, 2.373228e-08, 
    2.387605e-08, 2.4155e-08, 2.462008e-08, 2.467198e-08, 2.304457e-08, 
    2.202197e-08, 2.335691e-08, 2.34294e-08, 2.335623e-08, 2.406177e-08,
  2.414988e-08, 2.437607e-08, 2.427e-08, 2.433689e-08, 2.424703e-08, 
    2.44314e-08, 2.444534e-08, 2.508156e-08, 2.390319e-08, 2.329429e-08, 
    2.569389e-08, 2.541742e-08, 2.471167e-08, 2.458091e-08, 2.606031e-08,
  2.44854e-08, 2.444496e-08, 2.459211e-08, 2.490617e-08, 2.489571e-08, 
    2.516448e-08, 2.527404e-08, 2.494115e-08, 2.461061e-08, 2.534814e-08, 
    2.624084e-08, 2.600334e-08, 2.607239e-08, 2.618607e-08, 2.627145e-08,
  2.47036e-08, 2.413314e-08, 2.474903e-08, 2.55391e-08, 2.572876e-08, 
    2.624723e-08, 2.589221e-08, 2.516935e-08, 2.513677e-08, 2.551609e-08, 
    2.614462e-08, 2.648554e-08, 2.662802e-08, 2.614966e-08, 2.525189e-08,
  2.480474e-08, 2.473329e-08, 2.572795e-08, 2.629611e-08, 2.596403e-08, 
    2.63937e-08, 2.584832e-08, 2.450266e-08, 2.489688e-08, 2.609164e-08, 
    2.704453e-08, 2.740694e-08, 2.735895e-08, 2.575847e-08, 2.542952e-08,
  2.479655e-08, 2.582428e-08, 2.600357e-08, 2.585271e-08, 2.55379e-08, 
    2.577189e-08, 2.433753e-08, 2.443602e-08, 2.643008e-08, 2.695665e-08, 
    2.769384e-08, 2.798587e-08, 2.828153e-08, 2.697012e-08, 2.655956e-08,
  2.435529e-08, 2.463619e-08, 2.517423e-08, 2.592071e-08, 2.590795e-08, 
    2.566291e-08, 2.515338e-08, 2.474543e-08, 2.414333e-08, 2.244588e-08, 
    2.293694e-08, 2.526373e-08, 2.77944e-08, 2.697891e-08, 2.683447e-08,
  2.426933e-08, 2.518429e-08, 2.591859e-08, 2.639669e-08, 2.617599e-08, 
    2.629327e-08, 2.571829e-08, 2.564313e-08, 2.575711e-08, 2.49741e-08, 
    2.343747e-08, 2.259902e-08, 2.426645e-08, 2.570391e-08, 2.617486e-08,
  2.719767e-08, 2.65894e-08, 2.701321e-08, 2.778409e-08, 2.803471e-08, 
    2.811682e-08, 2.659473e-08, 2.402954e-08, 2.545916e-08, 2.770988e-08, 
    2.691553e-08, 2.487429e-08, 2.138123e-08, 2.083133e-08, 2.307707e-08,
  2.748039e-08, 2.680187e-08, 2.746116e-08, 2.806118e-08, 2.829585e-08, 
    2.826309e-08, 2.807244e-08, 2.588355e-08, 2.439093e-08, 2.573355e-08, 
    2.540938e-08, 2.568073e-08, 2.452388e-08, 2.205891e-08, 2.073216e-08,
  2.761706e-08, 2.726768e-08, 2.767371e-08, 2.806948e-08, 2.82709e-08, 
    2.796513e-08, 2.776618e-08, 2.799406e-08, 2.523142e-08, 2.612941e-08, 
    2.4386e-08, 2.449196e-08, 2.431372e-08, 2.316694e-08, 2.042247e-08,
  2.766089e-08, 2.721653e-08, 2.70228e-08, 2.769751e-08, 2.796302e-08, 
    2.817103e-08, 2.796379e-08, 2.810077e-08, 2.799982e-08, 2.436278e-08, 
    2.448363e-08, 2.498492e-08, 2.479104e-08, 2.341282e-08, 2.471178e-08,
  2.784003e-08, 2.705888e-08, 2.769962e-08, 2.891278e-08, 2.942528e-08, 
    2.996468e-08, 2.959556e-08, 2.886782e-08, 2.847404e-08, 2.624131e-08, 
    2.484501e-08, 2.44223e-08, 2.364097e-08, 2.302629e-08, 2.501033e-08,
  2.761188e-08, 2.779483e-08, 2.886552e-08, 2.976741e-08, 3.029943e-08, 
    3.059876e-08, 3.081018e-08, 3.073537e-08, 2.99857e-08, 2.782238e-08, 
    2.554157e-08, 2.449871e-08, 2.354622e-08, 2.320579e-08, 2.352819e-08,
  2.797206e-08, 2.865708e-08, 3.024784e-08, 3.068029e-08, 3.070307e-08, 
    3.049217e-08, 3.04811e-08, 3.135501e-08, 2.991013e-08, 2.8709e-08, 
    2.679709e-08, 2.510163e-08, 2.388721e-08, 2.262016e-08, 2.190174e-08,
  2.911754e-08, 2.942602e-08, 3.032831e-08, 2.933734e-08, 2.874385e-08, 
    2.835201e-08, 2.882891e-08, 2.848363e-08, 2.894649e-08, 2.920991e-08, 
    2.795194e-08, 2.591624e-08, 2.474895e-08, 2.351619e-08, 2.278426e-08,
  2.305304e-08, 2.403826e-08, 2.37969e-08, 2.44091e-08, 2.480153e-08, 
    2.46128e-08, 2.460236e-08, 2.507269e-08, 2.560118e-08, 2.538092e-08, 
    2.464735e-08, 2.460666e-08, 2.546836e-08, 2.500347e-08, 2.56365e-08,
  2.534895e-08, 2.617318e-08, 2.546221e-08, 2.593058e-08, 2.646119e-08, 
    2.677863e-08, 2.55146e-08, 2.612579e-08, 2.677124e-08, 2.643315e-08, 
    2.436013e-08, 2.331009e-08, 2.311254e-08, 2.439345e-08, 2.517192e-08,
  2.533102e-08, 2.672099e-08, 2.557952e-08, 2.459942e-08, 2.496371e-08, 
    2.575999e-08, 2.502201e-08, 2.484071e-08, 2.589854e-08, 2.604108e-08, 
    2.632758e-08, 2.458795e-08, 2.254703e-08, 2.330453e-08, 2.296815e-08,
  2.451602e-08, 2.445009e-08, 2.546997e-08, 2.45954e-08, 2.279262e-08, 
    2.206869e-08, 2.213108e-08, 2.14852e-08, 2.163159e-08, 2.337166e-08, 
    2.466928e-08, 2.51141e-08, 2.445087e-08, 2.442279e-08, 2.275212e-08,
  2.514465e-08, 2.753594e-08, 2.805431e-08, 2.753453e-08, 2.594771e-08, 
    2.394962e-08, 2.309172e-08, 2.189163e-08, 1.986074e-08, 2.144716e-08, 
    2.341865e-08, 2.388312e-08, 2.382873e-08, 2.376923e-08, 2.193496e-08,
  2.934999e-08, 3.00379e-08, 3.002106e-08, 2.961843e-08, 2.89942e-08, 
    2.763119e-08, 2.516263e-08, 2.380756e-08, 2.261705e-08, 2.057038e-08, 
    2.158598e-08, 2.415615e-08, 2.446262e-08, 2.365212e-08, 2.454074e-08,
  2.938022e-08, 3.036287e-08, 3.074458e-08, 2.998671e-08, 2.992924e-08, 
    2.958735e-08, 2.797011e-08, 2.584376e-08, 2.543349e-08, 2.253385e-08, 
    2.172171e-08, 2.326966e-08, 2.421295e-08, 2.340486e-08, 2.59919e-08,
  3.026185e-08, 3.178185e-08, 3.087193e-08, 2.944639e-08, 2.975404e-08, 
    3.017952e-08, 3.0567e-08, 2.901082e-08, 2.911471e-08, 2.613215e-08, 
    2.350524e-08, 2.286835e-08, 2.372894e-08, 2.408882e-08, 2.582722e-08,
  3.006005e-08, 3.085563e-08, 3.064134e-08, 3.000819e-08, 2.944256e-08, 
    3.117746e-08, 3.343742e-08, 3.119657e-08, 3.014301e-08, 2.853928e-08, 
    2.643603e-08, 2.377166e-08, 2.43934e-08, 2.516896e-08, 2.441594e-08,
  2.878799e-08, 2.997346e-08, 3.140926e-08, 3.091131e-08, 3.12404e-08, 
    3.056101e-08, 3.192461e-08, 2.89936e-08, 2.921545e-08, 2.866035e-08, 
    2.759204e-08, 2.503383e-08, 2.524077e-08, 2.582738e-08, 2.476545e-08,
  2.658453e-08, 2.873176e-08, 2.853722e-08, 2.97263e-08, 2.908419e-08, 
    2.870387e-08, 2.792279e-08, 2.836721e-08, 2.607282e-08, 2.415924e-08, 
    2.328767e-08, 2.38092e-08, 2.192892e-08, 2.181777e-08, 2.01512e-08,
  2.738118e-08, 2.858037e-08, 2.804877e-08, 2.775013e-08, 2.850407e-08, 
    2.784448e-08, 2.720786e-08, 2.793203e-08, 2.637602e-08, 2.461404e-08, 
    2.286943e-08, 2.25766e-08, 2.134839e-08, 2.085818e-08, 2.074438e-08,
  2.931844e-08, 2.899387e-08, 2.920564e-08, 2.741684e-08, 2.64524e-08, 
    2.853929e-08, 2.799049e-08, 2.754913e-08, 2.633927e-08, 2.486559e-08, 
    2.3713e-08, 2.212486e-08, 2.275484e-08, 2.182079e-08, 2.197183e-08,
  3.015178e-08, 2.951953e-08, 2.936117e-08, 2.857173e-08, 2.710609e-08, 
    2.734255e-08, 2.776836e-08, 2.873952e-08, 2.899981e-08, 2.710366e-08, 
    2.563885e-08, 2.463141e-08, 2.382449e-08, 2.348982e-08, 2.2454e-08,
  3.156418e-08, 3.026103e-08, 2.989937e-08, 2.949558e-08, 2.818534e-08, 
    2.682238e-08, 2.558835e-08, 2.764474e-08, 2.932722e-08, 3.290264e-08, 
    2.989368e-08, 2.300569e-08, 2.368446e-08, 2.363276e-08, 2.201043e-08,
  2.974547e-08, 2.947216e-08, 2.89001e-08, 2.953481e-08, 2.815436e-08, 
    2.831673e-08, 2.687038e-08, 2.713564e-08, 2.743105e-08, 2.644777e-08, 
    2.653267e-08, 2.456417e-08, 2.25372e-08, 2.254501e-08, 2.421514e-08,
  3.012202e-08, 2.903121e-08, 2.902363e-08, 2.972122e-08, 2.738816e-08, 
    2.834336e-08, 2.851957e-08, 2.807547e-08, 2.649507e-08, 2.352396e-08, 
    2.433093e-08, 2.578424e-08, 2.22951e-08, 2.232145e-08, 2.631585e-08,
  2.830715e-08, 2.983148e-08, 2.945087e-08, 2.98549e-08, 2.741463e-08, 
    2.692527e-08, 2.819928e-08, 2.889005e-08, 2.749439e-08, 2.456637e-08, 
    2.296622e-08, 2.316961e-08, 2.121034e-08, 2.20268e-08, 2.584408e-08,
  2.850473e-08, 3.148455e-08, 2.999831e-08, 2.980222e-08, 2.804837e-08, 
    2.707056e-08, 2.948924e-08, 3.146326e-08, 2.738144e-08, 2.495108e-08, 
    2.345579e-08, 2.162902e-08, 2.007889e-08, 2.095125e-08, 2.416857e-08,
  2.861364e-08, 3.139771e-08, 3.028961e-08, 2.894759e-08, 2.804386e-08, 
    2.721648e-08, 2.870515e-08, 2.753334e-08, 2.738593e-08, 2.632662e-08, 
    2.428949e-08, 2.237949e-08, 2.001798e-08, 2.003631e-08, 2.254621e-08,
  2.303227e-08, 2.57936e-08, 2.830753e-08, 2.826393e-08, 2.613629e-08, 
    2.51351e-08, 2.55131e-08, 2.712205e-08, 2.745546e-08, 2.991472e-08, 
    2.747595e-08, 2.661831e-08, 2.459818e-08, 2.414961e-08, 1.945644e-08,
  2.442803e-08, 2.681328e-08, 2.727855e-08, 2.865918e-08, 2.597884e-08, 
    2.480354e-08, 2.525405e-08, 2.555651e-08, 2.716234e-08, 2.69361e-08, 
    2.845364e-08, 2.837771e-08, 2.766014e-08, 2.69406e-08, 2.618594e-08,
  2.932778e-08, 2.716821e-08, 2.885035e-08, 2.800608e-08, 2.74633e-08, 
    2.594336e-08, 2.527253e-08, 2.523688e-08, 2.569855e-08, 2.554278e-08, 
    2.615464e-08, 2.736261e-08, 2.827439e-08, 2.832961e-08, 2.828951e-08,
  2.999393e-08, 2.807986e-08, 2.917237e-08, 2.942411e-08, 2.884989e-08, 
    2.742165e-08, 2.552269e-08, 2.56515e-08, 2.526653e-08, 2.614551e-08, 
    2.911133e-08, 2.829671e-08, 2.83946e-08, 2.881841e-08, 2.922049e-08,
  3.138535e-08, 2.9425e-08, 3.003954e-08, 3.055318e-08, 2.977363e-08, 
    2.742341e-08, 2.545174e-08, 2.59074e-08, 2.614839e-08, 3.069943e-08, 
    2.758677e-08, 2.714781e-08, 2.761409e-08, 2.919653e-08, 2.967384e-08,
  2.963811e-08, 2.859274e-08, 2.718775e-08, 2.784534e-08, 2.740092e-08, 
    2.719222e-08, 2.741353e-08, 2.730424e-08, 2.777963e-08, 2.712074e-08, 
    2.756441e-08, 2.828287e-08, 2.773079e-08, 2.972899e-08, 2.991985e-08,
  2.726195e-08, 2.828293e-08, 2.802527e-08, 2.851124e-08, 2.948981e-08, 
    2.829177e-08, 2.759051e-08, 2.604651e-08, 2.772457e-08, 2.716306e-08, 
    2.737719e-08, 2.811243e-08, 2.724528e-08, 2.720243e-08, 2.902452e-08,
  2.571575e-08, 2.77591e-08, 2.794163e-08, 2.764881e-08, 2.760252e-08, 
    2.748473e-08, 2.596504e-08, 2.440214e-08, 2.476266e-08, 2.57679e-08, 
    2.664127e-08, 2.722988e-08, 2.548306e-08, 2.824476e-08, 2.9038e-08,
  2.422667e-08, 2.721628e-08, 2.745799e-08, 2.837354e-08, 2.80994e-08, 
    2.854005e-08, 2.600689e-08, 2.531846e-08, 2.433556e-08, 2.690357e-08, 
    2.682014e-08, 2.772378e-08, 2.639319e-08, 2.76601e-08, 2.778616e-08,
  2.413958e-08, 2.612962e-08, 2.657338e-08, 2.672225e-08, 2.618273e-08, 
    2.590514e-08, 2.510295e-08, 2.259118e-08, 2.36336e-08, 2.66068e-08, 
    2.679858e-08, 2.806812e-08, 2.76027e-08, 2.627258e-08, 2.701005e-08,
  2.155426e-08, 2.234245e-08, 2.30452e-08, 2.333724e-08, 2.494643e-08, 
    2.584722e-08, 2.787688e-08, 2.999672e-08, 3.031656e-08, 2.812415e-08, 
    2.559656e-08, 2.452041e-08, 2.279752e-08, 2.331691e-08, 2.494897e-08,
  2.152266e-08, 2.212576e-08, 2.34082e-08, 2.427093e-08, 2.577849e-08, 
    2.657891e-08, 2.773139e-08, 3.07179e-08, 3.162291e-08, 2.941886e-08, 
    2.645734e-08, 2.593217e-08, 2.413974e-08, 2.375412e-08, 2.493957e-08,
  2.443443e-08, 2.205722e-08, 2.379839e-08, 2.628668e-08, 2.766593e-08, 
    2.767623e-08, 2.771496e-08, 2.957544e-08, 3.061107e-08, 2.897767e-08, 
    2.875542e-08, 2.760104e-08, 2.480517e-08, 2.449111e-08, 2.537176e-08,
  2.388714e-08, 2.29268e-08, 2.417157e-08, 2.580198e-08, 2.697626e-08, 
    2.815669e-08, 2.784238e-08, 2.925241e-08, 3.043645e-08, 2.859076e-08, 
    2.907553e-08, 2.716678e-08, 2.719078e-08, 2.466389e-08, 2.552858e-08,
  2.36167e-08, 2.306128e-08, 2.424084e-08, 2.582203e-08, 2.696966e-08, 
    2.850035e-08, 2.914077e-08, 2.889889e-08, 2.687242e-08, 2.761587e-08, 
    2.676998e-08, 2.749945e-08, 2.960525e-08, 2.471756e-08, 2.52235e-08,
  2.276592e-08, 2.345945e-08, 2.477705e-08, 2.55027e-08, 2.731659e-08, 
    2.767339e-08, 2.825962e-08, 2.661398e-08, 2.682713e-08, 2.77264e-08, 
    3.183422e-08, 3.146781e-08, 3.125034e-08, 2.66371e-08, 2.849195e-08,
  2.414757e-08, 2.533951e-08, 2.531614e-08, 2.55625e-08, 2.765102e-08, 
    2.765852e-08, 2.77301e-08, 2.596419e-08, 2.505239e-08, 2.644577e-08, 
    2.991203e-08, 2.989777e-08, 3.09225e-08, 2.85237e-08, 3.115405e-08,
  2.51465e-08, 2.641941e-08, 2.509903e-08, 2.490469e-08, 2.734877e-08, 
    2.795237e-08, 2.738159e-08, 2.593259e-08, 2.467554e-08, 2.594732e-08, 
    2.849903e-08, 3.069149e-08, 3.058654e-08, 3.109796e-08, 2.853434e-08,
  2.144369e-08, 2.653576e-08, 2.414363e-08, 2.589583e-08, 2.628814e-08, 
    2.649513e-08, 2.482332e-08, 2.396436e-08, 2.471019e-08, 2.680291e-08, 
    2.827237e-08, 2.948162e-08, 2.966838e-08, 3.017406e-08, 2.639007e-08,
  1.865293e-08, 2.018406e-08, 2.050413e-08, 2.214636e-08, 2.309038e-08, 
    2.262073e-08, 2.210575e-08, 2.323329e-08, 2.435415e-08, 2.431865e-08, 
    2.556851e-08, 2.719946e-08, 2.812574e-08, 2.831312e-08, 2.70609e-08,
  1.604155e-08, 1.76448e-08, 2.0047e-08, 2.079096e-08, 1.922651e-08, 
    1.743727e-08, 1.663177e-08, 1.971719e-08, 2.383986e-08, 2.709864e-08, 
    3.05339e-08, 3.021561e-08, 3.153481e-08, 2.727517e-08, 2.209031e-08,
  1.869103e-08, 2.090146e-08, 2.221041e-08, 2.364061e-08, 2.188878e-08, 
    1.940757e-08, 1.739345e-08, 1.850462e-08, 2.173982e-08, 2.434567e-08, 
    2.906767e-08, 2.96172e-08, 3.112907e-08, 2.680428e-08, 2.14944e-08,
  2.450873e-08, 2.394712e-08, 2.418916e-08, 2.653424e-08, 2.512677e-08, 
    2.122178e-08, 1.823872e-08, 1.795031e-08, 2.062189e-08, 2.310333e-08, 
    2.854851e-08, 2.816617e-08, 2.87163e-08, 2.391043e-08, 2.340139e-08,
  2.454113e-08, 2.119167e-08, 2.264867e-08, 2.533725e-08, 2.403805e-08, 
    2.22835e-08, 1.996735e-08, 1.912573e-08, 2.008425e-08, 2.042576e-08, 
    2.228766e-08, 2.55755e-08, 2.793514e-08, 2.468009e-08, 2.915221e-08,
  2.19843e-08, 1.977982e-08, 2.069964e-08, 2.070592e-08, 2.171057e-08, 
    2.217077e-08, 2.112002e-08, 2.047116e-08, 1.930265e-08, 1.722161e-08, 
    1.94425e-08, 2.450632e-08, 2.759528e-08, 2.879633e-08, 3.349359e-08,
  2.237843e-08, 2.074452e-08, 2.062836e-08, 2.014659e-08, 2.030032e-08, 
    2.049755e-08, 2.038184e-08, 1.972209e-08, 1.961061e-08, 1.8808e-08, 
    2.126141e-08, 2.280962e-08, 2.576993e-08, 3.26434e-08, 3.136612e-08,
  2.314046e-08, 2.328564e-08, 2.311313e-08, 2.198551e-08, 2.097097e-08, 
    2.019131e-08, 2.062398e-08, 1.981161e-08, 2.100519e-08, 2.101844e-08, 
    2.280934e-08, 2.157856e-08, 2.625917e-08, 3.346939e-08, 2.480473e-08,
  2.464153e-08, 2.542527e-08, 2.500104e-08, 2.384936e-08, 2.336159e-08, 
    2.154621e-08, 2.089833e-08, 1.949447e-08, 1.980301e-08, 2.010444e-08, 
    2.114214e-08, 2.161199e-08, 2.626176e-08, 2.59109e-08, 2.13324e-08,
  2.364989e-08, 2.579515e-08, 2.524434e-08, 2.543161e-08, 2.69974e-08, 
    2.467316e-08, 2.176454e-08, 1.982037e-08, 1.940084e-08, 2.083326e-08, 
    2.057554e-08, 2.089833e-08, 2.266688e-08, 2.271172e-08, 2.209123e-08,
  2.765889e-08, 2.651688e-08, 2.41232e-08, 2.121204e-08, 2.149837e-08, 
    2.253412e-08, 2.129844e-08, 2.335934e-08, 2.463753e-08, 2.313427e-08, 
    2.073352e-08, 2.039978e-08, 2.073112e-08, 2.075768e-08, 2.218255e-08,
  1.626092e-08, 1.512029e-08, 1.4667e-08, 1.508516e-08, 1.508388e-08, 
    1.633209e-08, 1.623138e-08, 1.599743e-08, 1.69357e-08, 1.659475e-08, 
    1.793378e-08, 2.180505e-08, 2.627624e-08, 2.370351e-08, 2.4483e-08,
  1.686549e-08, 1.612585e-08, 1.541981e-08, 1.54769e-08, 1.626205e-08, 
    1.711107e-08, 1.675089e-08, 1.680338e-08, 1.678591e-08, 1.698202e-08, 
    1.713237e-08, 2.202034e-08, 2.658838e-08, 2.115542e-08, 2.326052e-08,
  1.733985e-08, 1.755515e-08, 1.713634e-08, 1.682998e-08, 1.75991e-08, 
    1.709047e-08, 1.711151e-08, 1.771871e-08, 1.7358e-08, 1.729219e-08, 
    1.746763e-08, 2.191595e-08, 2.539633e-08, 1.859079e-08, 2.314609e-08,
  1.777734e-08, 1.771232e-08, 1.731997e-08, 1.825913e-08, 1.863294e-08, 
    1.884541e-08, 1.884699e-08, 1.889097e-08, 1.92671e-08, 1.733586e-08, 
    1.850686e-08, 2.245877e-08, 2.595363e-08, 2.054721e-08, 2.655301e-08,
  1.939188e-08, 1.823273e-08, 1.667068e-08, 1.528888e-08, 1.695574e-08, 
    2.009048e-08, 2.06791e-08, 2.08965e-08, 2.085047e-08, 1.876503e-08, 
    2.043396e-08, 2.335881e-08, 2.440308e-08, 2.495929e-08, 2.961127e-08,
  2.246407e-08, 2.088365e-08, 1.960489e-08, 1.686915e-08, 1.653586e-08, 
    1.747546e-08, 1.861922e-08, 1.99777e-08, 1.903894e-08, 1.994068e-08, 
    2.141973e-08, 2.06066e-08, 2.193075e-08, 2.650032e-08, 2.57116e-08,
  2.307846e-08, 2.293391e-08, 2.176963e-08, 2.029246e-08, 1.826556e-08, 
    1.846438e-08, 1.903377e-08, 1.972106e-08, 1.917095e-08, 2.088081e-08, 
    2.223113e-08, 2.016343e-08, 2.108323e-08, 2.550331e-08, 2.217434e-08,
  2.32961e-08, 2.456522e-08, 2.312848e-08, 2.194537e-08, 1.983985e-08, 
    1.992221e-08, 1.978365e-08, 2.058051e-08, 1.961955e-08, 1.974626e-08, 
    2.083097e-08, 1.979841e-08, 2.096048e-08, 2.15069e-08, 1.984133e-08,
  2.653668e-08, 2.711473e-08, 2.708915e-08, 2.503566e-08, 2.220726e-08, 
    2.086805e-08, 1.999715e-08, 1.915656e-08, 1.900715e-08, 2.039808e-08, 
    1.998199e-08, 1.868775e-08, 1.880034e-08, 1.892531e-08, 1.858362e-08,
  3.038422e-08, 2.928295e-08, 2.874448e-08, 2.702193e-08, 2.34172e-08, 
    1.974309e-08, 2.000586e-08, 2.259231e-08, 2.317392e-08, 2.211029e-08, 
    2.013148e-08, 1.896061e-08, 1.793872e-08, 1.737296e-08, 1.804618e-08,
  1.720154e-08, 1.705842e-08, 1.659581e-08, 1.612804e-08, 1.566779e-08, 
    1.569847e-08, 1.563179e-08, 1.604917e-08, 1.745479e-08, 1.800347e-08, 
    2.202038e-08, 2.458501e-08, 2.403089e-08, 2.380707e-08, 2.476858e-08,
  1.808898e-08, 1.802391e-08, 1.7264e-08, 1.668994e-08, 1.623702e-08, 
    1.589375e-08, 1.596907e-08, 1.638072e-08, 1.781757e-08, 1.841914e-08, 
    2.083927e-08, 2.410704e-08, 2.549891e-08, 2.355604e-08, 2.302438e-08,
  1.990989e-08, 1.962605e-08, 1.835476e-08, 1.751037e-08, 1.723959e-08, 
    1.684865e-08, 1.64029e-08, 1.67513e-08, 1.722968e-08, 1.91382e-08, 
    2.058125e-08, 2.39445e-08, 2.528542e-08, 2.267102e-08, 2.251531e-08,
  2.197358e-08, 1.995602e-08, 1.886172e-08, 1.830568e-08, 1.852234e-08, 
    1.819448e-08, 1.76052e-08, 1.714688e-08, 1.739419e-08, 1.780281e-08, 
    1.858139e-08, 2.364697e-08, 2.66328e-08, 2.393691e-08, 2.364028e-08,
  2.27607e-08, 2.105502e-08, 1.968294e-08, 1.813901e-08, 1.773248e-08, 
    1.863805e-08, 1.844306e-08, 1.758752e-08, 1.704837e-08, 1.559614e-08, 
    1.71121e-08, 2.329791e-08, 2.384096e-08, 2.178418e-08, 2.693262e-08,
  2.271798e-08, 2.234124e-08, 2.1407e-08, 1.982535e-08, 1.837307e-08, 
    1.76685e-08, 1.789776e-08, 1.781084e-08, 1.778591e-08, 1.745126e-08, 
    1.827273e-08, 1.801941e-08, 2.163474e-08, 2.122333e-08, 2.563559e-08,
  2.243014e-08, 2.238415e-08, 2.268624e-08, 2.186874e-08, 2.073378e-08, 
    1.925352e-08, 1.792617e-08, 1.772497e-08, 1.757368e-08, 1.780439e-08, 
    1.785406e-08, 1.765851e-08, 1.961166e-08, 2.148076e-08, 2.24566e-08,
  2.304077e-08, 2.342665e-08, 2.331933e-08, 2.298116e-08, 2.208651e-08, 
    2.170864e-08, 2.043268e-08, 1.953174e-08, 1.941723e-08, 1.862523e-08, 
    1.829357e-08, 1.755008e-08, 1.747298e-08, 2.037937e-08, 1.797969e-08,
  2.618149e-08, 2.551187e-08, 2.535551e-08, 2.422904e-08, 2.29792e-08, 
    2.165461e-08, 2.184112e-08, 1.98993e-08, 1.906087e-08, 1.90925e-08, 
    1.899754e-08, 1.855701e-08, 1.707492e-08, 1.79832e-08, 1.788471e-08,
  2.978239e-08, 2.861957e-08, 2.7668e-08, 2.66154e-08, 2.492177e-08, 
    2.302978e-08, 2.271039e-08, 2.1517e-08, 1.970311e-08, 1.886466e-08, 
    1.859515e-08, 1.890891e-08, 1.798573e-08, 1.729614e-08, 1.767704e-08,
  1.697241e-08, 1.641626e-08, 1.568889e-08, 1.572656e-08, 1.542982e-08, 
    1.593497e-08, 1.64332e-08, 1.768433e-08, 1.794497e-08, 1.952365e-08, 
    2.037319e-08, 1.912593e-08, 2.20978e-08, 2.159586e-08, 2.241581e-08,
  2.137482e-08, 2.082039e-08, 1.909097e-08, 1.846387e-08, 1.755727e-08, 
    1.745112e-08, 1.765272e-08, 1.838394e-08, 1.899815e-08, 2.117338e-08, 
    2.141291e-08, 1.946803e-08, 2.19994e-08, 2.096292e-08, 2.179939e-08,
  2.530284e-08, 2.40241e-08, 2.218909e-08, 2.051457e-08, 2.001553e-08, 
    1.948772e-08, 1.928299e-08, 1.939872e-08, 2.019414e-08, 2.115093e-08, 
    2.416462e-08, 2.165626e-08, 2.223038e-08, 2.067011e-08, 2.177205e-08,
  2.853816e-08, 2.668816e-08, 2.487091e-08, 2.248465e-08, 2.178697e-08, 
    2.105248e-08, 2.077938e-08, 2.069535e-08, 2.102219e-08, 2.109063e-08, 
    1.938653e-08, 2.286121e-08, 2.45973e-08, 2.077201e-08, 2.249076e-08,
  2.816113e-08, 2.771471e-08, 2.611751e-08, 2.42141e-08, 2.193245e-08, 
    2.100526e-08, 2.025675e-08, 2.080031e-08, 2.027733e-08, 1.961504e-08, 
    1.785096e-08, 2.053572e-08, 2.489682e-08, 2.1596e-08, 2.242382e-08,
  2.817526e-08, 2.821715e-08, 2.811626e-08, 2.694601e-08, 2.37874e-08, 
    2.152076e-08, 2.090907e-08, 2.119914e-08, 2.141494e-08, 2.021438e-08, 
    2.064971e-08, 2.010859e-08, 2.086195e-08, 2.205009e-08, 2.364831e-08,
  2.774999e-08, 2.756947e-08, 2.768957e-08, 2.775214e-08, 2.671521e-08, 
    2.452622e-08, 2.286293e-08, 2.267093e-08, 2.184537e-08, 2.02615e-08, 
    2.007912e-08, 1.962692e-08, 1.987658e-08, 2.195278e-08, 2.074853e-08,
  2.784003e-08, 2.867321e-08, 2.887219e-08, 2.830645e-08, 2.720125e-08, 
    2.663798e-08, 2.624988e-08, 2.681375e-08, 2.647542e-08, 2.334114e-08, 
    2.1891e-08, 2.056118e-08, 2.061107e-08, 2.069828e-08, 2.042118e-08,
  2.689955e-08, 2.897126e-08, 3.004225e-08, 2.976061e-08, 2.86702e-08, 
    2.762324e-08, 2.682726e-08, 2.581787e-08, 2.45453e-08, 2.396665e-08, 
    2.39485e-08, 2.296592e-08, 2.170304e-08, 2.062481e-08, 1.970062e-08,
  2.645642e-08, 2.878981e-08, 3.035262e-08, 3.024897e-08, 2.956908e-08, 
    2.906919e-08, 2.904843e-08, 2.722983e-08, 2.546635e-08, 2.529389e-08, 
    2.442555e-08, 2.434746e-08, 2.335827e-08, 2.170031e-08, 2.024139e-08,
  1.88044e-08, 1.796753e-08, 1.643573e-08, 1.604008e-08, 1.494161e-08, 
    1.397897e-08, 1.313508e-08, 1.268997e-08, 1.228429e-08, 1.259575e-08, 
    1.2438e-08, 1.4812e-08, 1.588343e-08, 1.880908e-08, 1.947574e-08,
  2.575715e-08, 2.59412e-08, 2.313437e-08, 2.049976e-08, 1.880415e-08, 
    1.684741e-08, 1.519723e-08, 1.434286e-08, 1.337218e-08, 1.362092e-08, 
    1.348777e-08, 1.508453e-08, 1.591053e-08, 1.882431e-08, 1.893206e-08,
  3.317778e-08, 3.171949e-08, 2.834599e-08, 2.617988e-08, 2.357779e-08, 
    2.147737e-08, 1.90007e-08, 1.715481e-08, 1.540889e-08, 1.521225e-08, 
    1.444776e-08, 1.561049e-08, 1.66662e-08, 2.007594e-08, 1.884811e-08,
  3.898875e-08, 3.589464e-08, 3.417999e-08, 3.229977e-08, 2.890063e-08, 
    2.643325e-08, 2.410423e-08, 2.234473e-08, 1.935993e-08, 1.812151e-08, 
    1.552545e-08, 1.495426e-08, 1.734734e-08, 2.160584e-08, 2.023969e-08,
  3.209418e-08, 3.241136e-08, 3.214222e-08, 3.132577e-08, 3.034381e-08, 
    2.905658e-08, 2.761017e-08, 2.559442e-08, 2.34686e-08, 2.094941e-08, 
    1.905906e-08, 1.84689e-08, 1.929648e-08, 2.193264e-08, 2.246541e-08,
  2.78621e-08, 2.748025e-08, 2.800411e-08, 2.795974e-08, 2.929802e-08, 
    2.981449e-08, 2.947144e-08, 2.809422e-08, 2.768525e-08, 2.528657e-08, 
    2.369443e-08, 2.15143e-08, 2.125037e-08, 2.282002e-08, 2.281838e-08,
  1.955167e-08, 1.940161e-08, 2.11254e-08, 2.257537e-08, 2.526519e-08, 
    2.72945e-08, 2.909923e-08, 2.940487e-08, 2.938655e-08, 2.680906e-08, 
    2.578255e-08, 2.39978e-08, 2.412299e-08, 2.377585e-08, 2.201859e-08,
  1.709962e-08, 1.805858e-08, 1.908189e-08, 1.972853e-08, 2.088095e-08, 
    2.281199e-08, 2.572002e-08, 2.762709e-08, 2.960747e-08, 2.907646e-08, 
    2.760356e-08, 2.681396e-08, 2.777344e-08, 2.674438e-08, 2.441146e-08,
  1.919486e-08, 1.880412e-08, 2.207877e-08, 2.346181e-08, 2.35162e-08, 
    2.327805e-08, 2.344583e-08, 2.447928e-08, 2.511431e-08, 2.681984e-08, 
    2.727448e-08, 2.769135e-08, 2.847723e-08, 2.847249e-08, 2.577844e-08,
  2.163951e-08, 1.811241e-08, 2.246266e-08, 2.740003e-08, 2.851337e-08, 
    2.757645e-08, 2.503674e-08, 2.371315e-08, 2.333202e-08, 2.436234e-08, 
    2.512889e-08, 2.59059e-08, 2.705471e-08, 2.727096e-08, 2.674338e-08,
  2.10099e-08, 2.147351e-08, 2.121311e-08, 2.12133e-08, 2.075153e-08, 
    1.989194e-08, 1.909508e-08, 1.851551e-08, 1.818522e-08, 1.755658e-08, 
    1.735986e-08, 1.649306e-08, 1.640013e-08, 1.615327e-08, 1.526338e-08,
  2.458565e-08, 2.488838e-08, 2.401636e-08, 2.32522e-08, 2.215318e-08, 
    2.173503e-08, 2.072311e-08, 2.040507e-08, 1.999889e-08, 2.012994e-08, 
    2.017521e-08, 1.946322e-08, 1.860875e-08, 1.771958e-08, 1.628362e-08,
  2.661024e-08, 2.838065e-08, 2.748934e-08, 2.672284e-08, 2.572936e-08, 
    2.471238e-08, 2.381042e-08, 2.21015e-08, 2.139172e-08, 2.107587e-08, 
    2.137653e-08, 2.137629e-08, 2.089168e-08, 1.892594e-08, 1.752835e-08,
  2.762359e-08, 2.862014e-08, 2.853161e-08, 2.996363e-08, 2.934089e-08, 
    2.916691e-08, 2.735808e-08, 2.658351e-08, 2.470139e-08, 2.401078e-08, 
    2.139986e-08, 2.157975e-08, 2.301979e-08, 2.195355e-08, 2.112863e-08,
  2.090726e-08, 2.209237e-08, 2.318166e-08, 2.549293e-08, 2.72578e-08, 
    2.889215e-08, 2.959101e-08, 2.929371e-08, 2.810974e-08, 2.5524e-08, 
    2.420003e-08, 2.445596e-08, 2.425562e-08, 2.482079e-08, 2.354123e-08,
  1.590602e-08, 1.722322e-08, 1.855696e-08, 1.978803e-08, 2.231646e-08, 
    2.498041e-08, 2.708149e-08, 2.788351e-08, 2.777963e-08, 2.587596e-08, 
    3.004276e-08, 2.85936e-08, 2.590352e-08, 2.363225e-08, 2.4181e-08,
  1.439695e-08, 1.575559e-08, 1.639965e-08, 1.736111e-08, 1.869594e-08, 
    1.97285e-08, 2.167212e-08, 2.267671e-08, 2.345123e-08, 2.488378e-08, 
    2.766398e-08, 2.758024e-08, 2.772796e-08, 2.47198e-08, 2.428611e-08,
  1.599503e-08, 1.671372e-08, 1.754424e-08, 1.835259e-08, 1.854783e-08, 
    1.910632e-08, 2.022082e-08, 2.085973e-08, 2.244208e-08, 2.336135e-08, 
    2.371895e-08, 2.45409e-08, 2.55846e-08, 2.438594e-08, 2.25511e-08,
  1.424831e-08, 1.680303e-08, 1.854917e-08, 2.153278e-08, 2.351071e-08, 
    2.389376e-08, 2.322115e-08, 2.221795e-08, 2.051367e-08, 2.188353e-08, 
    2.243176e-08, 2.331775e-08, 2.393427e-08, 2.416402e-08, 2.327011e-08,
  1.473136e-08, 1.914586e-08, 2.096295e-08, 2.262501e-08, 2.642425e-08, 
    2.994923e-08, 2.998451e-08, 2.6807e-08, 2.498153e-08, 2.433908e-08, 
    2.381198e-08, 2.380174e-08, 2.422544e-08, 2.437495e-08, 2.483987e-08,
  2.38869e-08, 2.406364e-08, 2.352575e-08, 2.352588e-08, 2.30795e-08, 
    2.254019e-08, 2.156149e-08, 2.091467e-08, 2.008079e-08, 1.96062e-08, 
    2.057752e-08, 1.976681e-08, 1.996747e-08, 2.05404e-08, 2.061393e-08,
  2.437441e-08, 2.442662e-08, 2.3824e-08, 2.355587e-08, 2.298045e-08, 
    2.279611e-08, 2.270574e-08, 2.188275e-08, 2.072474e-08, 2.079821e-08, 
    2.149564e-08, 2.147002e-08, 2.210937e-08, 2.223015e-08, 2.062671e-08,
  2.49192e-08, 2.471295e-08, 2.515752e-08, 2.364817e-08, 2.287267e-08, 
    2.316276e-08, 2.292198e-08, 2.216337e-08, 2.134218e-08, 2.193469e-08, 
    2.275277e-08, 2.281361e-08, 2.392155e-08, 2.456967e-08, 2.283617e-08,
  2.641708e-08, 2.608721e-08, 2.579053e-08, 2.643853e-08, 2.589475e-08, 
    2.584366e-08, 2.384525e-08, 2.421887e-08, 2.369213e-08, 2.344751e-08, 
    2.380957e-08, 2.355986e-08, 2.429144e-08, 2.275901e-08, 2.381625e-08,
  2.718308e-08, 2.824976e-08, 2.713825e-08, 2.719752e-08, 2.596943e-08, 
    2.586185e-08, 2.536482e-08, 2.534628e-08, 2.580037e-08, 2.662643e-08, 
    2.396634e-08, 2.392219e-08, 2.325817e-08, 2.170391e-08, 2.313698e-08,
  2.272619e-08, 2.505813e-08, 2.577964e-08, 2.555365e-08, 2.494879e-08, 
    2.47692e-08, 2.462738e-08, 2.419423e-08, 2.396763e-08, 2.222379e-08, 
    2.394015e-08, 2.448057e-08, 2.425302e-08, 2.257434e-08, 2.46373e-08,
  1.50323e-08, 1.730143e-08, 1.855366e-08, 1.991603e-08, 2.11466e-08, 
    2.194888e-08, 2.237422e-08, 2.186725e-08, 2.168773e-08, 2.256832e-08, 
    2.317351e-08, 2.443998e-08, 2.492501e-08, 2.507153e-08, 2.549813e-08,
  1.312973e-08, 1.497641e-08, 1.573068e-08, 1.618212e-08, 1.659266e-08, 
    1.787076e-08, 1.840074e-08, 1.961399e-08, 2.003285e-08, 2.102802e-08, 
    2.128792e-08, 2.166381e-08, 2.186784e-08, 2.12125e-08, 2.005256e-08,
  1.186256e-08, 1.495019e-08, 1.630261e-08, 1.879279e-08, 1.994122e-08, 
    1.886119e-08, 1.826612e-08, 1.957527e-08, 1.837168e-08, 1.951649e-08, 
    2.010178e-08, 2.04282e-08, 2.085423e-08, 2.073471e-08, 2.013895e-08,
  1.910883e-08, 1.822212e-08, 1.970452e-08, 2.224771e-08, 2.723214e-08, 
    3.030046e-08, 3.073168e-08, 2.706167e-08, 2.553895e-08, 2.635369e-08, 
    2.616878e-08, 2.603409e-08, 2.635617e-08, 2.632905e-08, 2.612583e-08,
  2.324222e-08, 2.406778e-08, 2.387112e-08, 2.358225e-08, 2.292487e-08, 
    2.261029e-08, 2.188266e-08, 2.173063e-08, 2.133002e-08, 2.014875e-08, 
    2.0549e-08, 2.021728e-08, 2.133078e-08, 2.132079e-08, 2.338749e-08,
  2.526684e-08, 2.525189e-08, 2.535607e-08, 2.496126e-08, 2.443168e-08, 
    2.399575e-08, 2.360327e-08, 2.317805e-08, 2.272244e-08, 2.146141e-08, 
    2.110685e-08, 1.95619e-08, 1.960344e-08, 2.0413e-08, 2.080187e-08,
  2.611392e-08, 2.622047e-08, 2.79492e-08, 2.676655e-08, 2.442754e-08, 
    2.433352e-08, 2.451051e-08, 2.373385e-08, 2.407966e-08, 2.334741e-08, 
    2.28572e-08, 2.165822e-08, 2.024349e-08, 2.041795e-08, 1.806613e-08,
  2.511184e-08, 2.57472e-08, 2.614754e-08, 2.80985e-08, 2.846053e-08, 
    2.615413e-08, 2.540098e-08, 2.50898e-08, 2.484935e-08, 2.446394e-08, 
    2.3694e-08, 2.3852e-08, 2.25718e-08, 2.114088e-08, 1.954942e-08,
  2.243672e-08, 2.529275e-08, 2.5686e-08, 2.579074e-08, 2.653646e-08, 
    2.640657e-08, 2.573851e-08, 2.601917e-08, 2.555659e-08, 2.619627e-08, 
    2.583974e-08, 2.443178e-08, 2.369892e-08, 2.207443e-08, 1.958813e-08,
  1.983786e-08, 2.288702e-08, 2.54334e-08, 2.679242e-08, 2.764134e-08, 
    2.625099e-08, 2.547212e-08, 2.68788e-08, 2.723152e-08, 2.59642e-08, 
    2.520027e-08, 2.488108e-08, 2.395603e-08, 2.162668e-08, 2.297919e-08,
  1.758236e-08, 1.948733e-08, 2.189081e-08, 2.479722e-08, 2.595798e-08, 
    2.613392e-08, 2.662595e-08, 2.64693e-08, 2.640606e-08, 2.468708e-08, 
    2.464232e-08, 2.476474e-08, 2.359144e-08, 2.247997e-08, 2.432771e-08,
  1.747265e-08, 1.867018e-08, 1.955259e-08, 2.144498e-08, 2.301533e-08, 
    2.361927e-08, 2.417263e-08, 2.504661e-08, 2.689195e-08, 2.569502e-08, 
    2.556738e-08, 2.497618e-08, 2.442586e-08, 2.3805e-08, 2.32936e-08,
  1.960178e-08, 1.899734e-08, 1.845666e-08, 2.000365e-08, 2.169641e-08, 
    2.201281e-08, 2.169732e-08, 2.263118e-08, 2.298149e-08, 2.349387e-08, 
    2.349607e-08, 2.295154e-08, 2.359138e-08, 2.300449e-08, 2.256776e-08,
  2.084559e-08, 2.373137e-08, 2.288358e-08, 1.957511e-08, 2.115653e-08, 
    2.453717e-08, 2.448899e-08, 2.380072e-08, 2.344265e-08, 2.390907e-08, 
    2.344453e-08, 2.321217e-08, 2.348429e-08, 2.377602e-08, 2.375381e-08,
  1.912293e-08, 1.971321e-08, 2.026486e-08, 2.032895e-08, 2.063022e-08, 
    2.078458e-08, 2.087381e-08, 2.116698e-08, 2.103297e-08, 2.045698e-08, 
    2.015002e-08, 1.996117e-08, 1.993783e-08, 1.951665e-08, 1.925847e-08,
  1.664234e-08, 1.716981e-08, 1.920582e-08, 2.15069e-08, 2.206929e-08, 
    2.278796e-08, 2.263439e-08, 2.347164e-08, 2.363735e-08, 2.314368e-08, 
    2.264834e-08, 2.212453e-08, 2.179291e-08, 2.098481e-08, 2.071546e-08,
  1.733908e-08, 1.916931e-08, 2.176313e-08, 2.334782e-08, 2.489966e-08, 
    2.525832e-08, 2.583269e-08, 2.623556e-08, 2.58021e-08, 2.54443e-08, 
    2.510666e-08, 2.450178e-08, 2.406865e-08, 2.362584e-08, 2.26764e-08,
  1.820523e-08, 1.829138e-08, 1.912056e-08, 2.171961e-08, 2.691997e-08, 
    2.846384e-08, 2.708817e-08, 2.701215e-08, 2.642463e-08, 2.612486e-08, 
    2.638387e-08, 2.658119e-08, 2.605544e-08, 2.557157e-08, 2.408654e-08,
  1.498502e-08, 1.550812e-08, 1.819815e-08, 2.161982e-08, 2.397105e-08, 
    2.408027e-08, 2.489604e-08, 2.641059e-08, 2.599586e-08, 2.745696e-08, 
    2.988601e-08, 2.977634e-08, 2.658709e-08, 2.659607e-08, 2.462372e-08,
  1.404484e-08, 1.48776e-08, 1.673053e-08, 1.963973e-08, 2.182768e-08, 
    2.290652e-08, 2.442784e-08, 2.610134e-08, 2.845777e-08, 2.790406e-08, 
    2.482916e-08, 2.740924e-08, 2.860232e-08, 2.451986e-08, 2.286507e-08,
  1.50188e-08, 1.500362e-08, 1.625621e-08, 1.935602e-08, 2.179672e-08, 
    2.226263e-08, 2.41203e-08, 2.672148e-08, 2.783528e-08, 2.475277e-08, 
    2.43166e-08, 2.525213e-08, 2.643986e-08, 2.243864e-08, 2.38854e-08,
  1.987191e-08, 1.797896e-08, 1.826968e-08, 2.077438e-08, 2.196374e-08, 
    2.261194e-08, 2.359372e-08, 2.47148e-08, 2.817054e-08, 2.609018e-08, 
    2.403394e-08, 2.349632e-08, 2.448057e-08, 2.270952e-08, 2.621696e-08,
  2.479483e-08, 2.301033e-08, 2.301818e-08, 2.436397e-08, 2.349865e-08, 
    2.36398e-08, 2.372173e-08, 2.486125e-08, 2.366862e-08, 2.421729e-08, 
    2.478624e-08, 2.337374e-08, 2.322489e-08, 2.393008e-08, 2.430612e-08,
  2.771471e-08, 2.762189e-08, 2.870514e-08, 2.811434e-08, 2.642052e-08, 
    2.569566e-08, 2.469227e-08, 2.22232e-08, 2.080003e-08, 2.114399e-08, 
    2.280386e-08, 2.344867e-08, 2.413371e-08, 2.470839e-08, 2.292564e-08,
  1.71211e-08, 1.612551e-08, 1.537129e-08, 1.498051e-08, 1.504626e-08, 
    1.691595e-08, 1.88144e-08, 2.065139e-08, 2.135381e-08, 2.17368e-08, 
    2.202732e-08, 2.221407e-08, 2.234048e-08, 2.180306e-08, 2.274151e-08,
  1.624088e-08, 1.480621e-08, 1.430862e-08, 1.427578e-08, 1.479951e-08, 
    1.718296e-08, 1.933215e-08, 2.08871e-08, 2.247661e-08, 2.305759e-08, 
    2.251689e-08, 2.227587e-08, 2.193574e-08, 2.092127e-08, 2.199672e-08,
  1.616067e-08, 1.451184e-08, 1.341697e-08, 1.395986e-08, 1.565914e-08, 
    1.77462e-08, 1.899563e-08, 2.058411e-08, 2.37782e-08, 2.396339e-08, 
    2.375077e-08, 2.347084e-08, 2.334525e-08, 2.320138e-08, 2.260724e-08,
  1.724048e-08, 1.509301e-08, 1.367604e-08, 1.41706e-08, 1.524347e-08, 
    1.662174e-08, 1.836448e-08, 2.060399e-08, 2.505541e-08, 2.501381e-08, 
    2.98828e-08, 2.784212e-08, 2.747162e-08, 3.000751e-08, 2.581334e-08,
  1.885311e-08, 1.670168e-08, 1.544007e-08, 1.51404e-08, 1.588113e-08, 
    1.754606e-08, 1.858592e-08, 2.158029e-08, 2.505356e-08, 3.266733e-08, 
    2.874404e-08, 2.7745e-08, 3.033406e-08, 2.742737e-08, 2.369881e-08,
  2.158129e-08, 1.945035e-08, 1.856628e-08, 1.774673e-08, 1.808191e-08, 
    1.84776e-08, 1.85528e-08, 2.089677e-08, 2.734172e-08, 2.884861e-08, 
    2.500663e-08, 2.609943e-08, 2.816333e-08, 2.072616e-08, 2.300981e-08,
  2.317196e-08, 2.244506e-08, 2.186492e-08, 2.064402e-08, 2.016571e-08, 
    1.93668e-08, 1.94223e-08, 2.232633e-08, 2.567286e-08, 2.576197e-08, 
    2.603275e-08, 2.458926e-08, 2.580398e-08, 1.891791e-08, 2.630577e-08,
  2.596284e-08, 2.737247e-08, 2.673207e-08, 2.553721e-08, 2.372546e-08, 
    2.173904e-08, 2.162179e-08, 2.227038e-08, 2.410764e-08, 2.546034e-08, 
    2.46798e-08, 2.437544e-08, 2.596438e-08, 2.309102e-08, 2.675331e-08,
  2.4959e-08, 2.768836e-08, 2.90019e-08, 2.842135e-08, 2.711215e-08, 
    2.513367e-08, 2.396591e-08, 2.599065e-08, 2.676202e-08, 2.548214e-08, 
    2.447033e-08, 2.370798e-08, 2.471264e-08, 2.395278e-08, 2.367947e-08,
  2.32907e-08, 2.639074e-08, 2.892196e-08, 2.977921e-08, 3.047428e-08, 
    2.980858e-08, 2.739311e-08, 2.592405e-08, 2.454397e-08, 2.382414e-08, 
    2.295877e-08, 2.190841e-08, 2.234494e-08, 2.377053e-08, 2.348745e-08,
  2.099796e-08, 2.088027e-08, 2.098286e-08, 2.13553e-08, 2.123215e-08, 
    1.972148e-08, 1.703598e-08, 1.601103e-08, 1.534963e-08, 1.66783e-08, 
    2.066568e-08, 2.304147e-08, 2.446118e-08, 2.331238e-08, 2.376597e-08,
  2.052853e-08, 2.054487e-08, 2.070121e-08, 2.119915e-08, 2.086522e-08, 
    1.871357e-08, 1.732432e-08, 1.677404e-08, 1.645918e-08, 1.904047e-08, 
    2.283374e-08, 2.465208e-08, 2.423916e-08, 2.443629e-08, 2.575547e-08,
  1.989698e-08, 1.998831e-08, 2.139645e-08, 2.157473e-08, 2.08528e-08, 
    1.857704e-08, 1.774154e-08, 1.706762e-08, 1.689745e-08, 2.048084e-08, 
    2.478607e-08, 2.672727e-08, 2.724694e-08, 3.176818e-08, 2.458542e-08,
  2.017569e-08, 1.974227e-08, 2.069736e-08, 2.077817e-08, 2.027514e-08, 
    1.904158e-08, 1.855177e-08, 1.83981e-08, 1.826185e-08, 2.308041e-08, 
    2.806664e-08, 2.846288e-08, 2.954895e-08, 3.024804e-08, 2.35694e-08,
  2.068656e-08, 2.098636e-08, 2.159631e-08, 2.159108e-08, 2.099043e-08, 
    2.14548e-08, 2.10565e-08, 2.099964e-08, 1.914539e-08, 2.772533e-08, 
    2.897721e-08, 2.481707e-08, 2.406677e-08, 2.27402e-08, 2.103985e-08,
  2.183728e-08, 2.177359e-08, 2.163507e-08, 2.148774e-08, 2.171285e-08, 
    2.206964e-08, 2.217013e-08, 2.119095e-08, 2.176477e-08, 2.2045e-08, 
    2.312493e-08, 2.83679e-08, 2.861291e-08, 2.056127e-08, 2.014415e-08,
  2.1783e-08, 2.12093e-08, 2.099749e-08, 2.176973e-08, 2.246832e-08, 
    2.370814e-08, 2.361756e-08, 2.326403e-08, 2.142334e-08, 2.067257e-08, 
    2.290058e-08, 2.50477e-08, 2.812362e-08, 1.899827e-08, 2.048145e-08,
  2.189271e-08, 2.130469e-08, 2.121279e-08, 2.232753e-08, 2.352002e-08, 
    2.492754e-08, 2.562829e-08, 2.500845e-08, 2.214709e-08, 2.142902e-08, 
    2.254233e-08, 2.354107e-08, 2.507166e-08, 2.162979e-08, 2.349341e-08,
  2.19206e-08, 2.127466e-08, 2.107971e-08, 2.217505e-08, 2.366252e-08, 
    2.474133e-08, 2.549612e-08, 2.58896e-08, 2.552435e-08, 2.468423e-08, 
    2.48218e-08, 2.459959e-08, 2.461706e-08, 2.465331e-08, 2.463469e-08,
  2.240923e-08, 2.137466e-08, 2.137055e-08, 2.184087e-08, 2.326333e-08, 
    2.480094e-08, 2.704422e-08, 2.809071e-08, 2.691219e-08, 2.638953e-08, 
    2.524723e-08, 2.363219e-08, 2.330461e-08, 2.40391e-08, 2.4331e-08,
  2.452505e-08, 2.433929e-08, 2.332224e-08, 2.275822e-08, 2.25109e-08, 
    2.276153e-08, 2.224572e-08, 2.215725e-08, 2.171914e-08, 2.042738e-08, 
    1.814439e-08, 1.846238e-08, 2.002422e-08, 2.195801e-08, 2.110715e-08,
  2.409226e-08, 2.348789e-08, 2.217607e-08, 2.161399e-08, 2.193371e-08, 
    2.28644e-08, 2.196169e-08, 2.233348e-08, 2.1578e-08, 2.009171e-08, 
    1.894579e-08, 2.072115e-08, 2.229835e-08, 2.517349e-08, 2.314683e-08,
  2.288494e-08, 2.299484e-08, 2.173913e-08, 2.170044e-08, 2.247679e-08, 
    2.299767e-08, 2.138114e-08, 2.092022e-08, 1.9878e-08, 2.023298e-08, 
    2.022706e-08, 2.375618e-08, 2.797245e-08, 3.097825e-08, 2.437202e-08,
  2.366965e-08, 2.272153e-08, 2.202133e-08, 2.232911e-08, 2.25038e-08, 
    2.220527e-08, 2.118437e-08, 2.091736e-08, 2.178822e-08, 2.442709e-08, 
    2.307377e-08, 2.50103e-08, 2.731965e-08, 2.817935e-08, 2.260385e-08,
  2.235424e-08, 2.256093e-08, 2.235058e-08, 2.269807e-08, 2.26412e-08, 
    2.254597e-08, 2.201174e-08, 2.164889e-08, 2.238973e-08, 2.605424e-08, 
    2.697038e-08, 2.677774e-08, 2.323634e-08, 2.251855e-08, 2.220772e-08,
  2.348244e-08, 2.317746e-08, 2.318629e-08, 2.293033e-08, 2.309216e-08, 
    2.276262e-08, 2.256448e-08, 2.175515e-08, 2.323244e-08, 2.373492e-08, 
    2.356058e-08, 2.345842e-08, 2.379997e-08, 2.33193e-08, 2.192652e-08,
  2.26944e-08, 2.274044e-08, 2.28723e-08, 2.323056e-08, 2.351212e-08, 
    2.287901e-08, 2.255021e-08, 2.196444e-08, 2.277969e-08, 2.324724e-08, 
    2.2558e-08, 2.149431e-08, 2.284747e-08, 2.42222e-08, 2.085897e-08,
  2.252463e-08, 2.376046e-08, 2.36057e-08, 2.395184e-08, 2.41267e-08, 
    2.399092e-08, 2.312876e-08, 2.20639e-08, 2.262535e-08, 2.344449e-08, 
    2.298796e-08, 2.155254e-08, 2.221969e-08, 2.195313e-08, 2.042925e-08,
  2.22228e-08, 2.421187e-08, 2.43959e-08, 2.411229e-08, 2.43878e-08, 
    2.454908e-08, 2.361165e-08, 2.260541e-08, 2.229051e-08, 2.310221e-08, 
    2.343978e-08, 2.210458e-08, 2.228652e-08, 2.200682e-08, 2.136767e-08,
  2.37327e-08, 2.461085e-08, 2.461394e-08, 2.417449e-08, 2.365639e-08, 
    2.308851e-08, 2.207712e-08, 2.110552e-08, 2.143238e-08, 2.211932e-08, 
    2.376303e-08, 2.343599e-08, 2.334928e-08, 2.344781e-08, 2.300635e-08,
  2.398554e-08, 2.504809e-08, 2.565042e-08, 2.540765e-08, 2.536542e-08, 
    2.470428e-08, 2.451983e-08, 2.471432e-08, 2.459935e-08, 2.590197e-08, 
    2.571232e-08, 2.400616e-08, 2.351553e-08, 2.240169e-08, 2.238638e-08,
  2.368779e-08, 2.471395e-08, 2.508131e-08, 2.477548e-08, 2.510178e-08, 
    2.498306e-08, 2.527488e-08, 2.366158e-08, 2.338878e-08, 2.456739e-08, 
    2.376086e-08, 2.341463e-08, 2.2767e-08, 2.337269e-08, 2.123118e-08,
  2.27368e-08, 2.167643e-08, 2.280733e-08, 2.312231e-08, 2.385747e-08, 
    2.481295e-08, 2.554059e-08, 2.464947e-08, 2.333369e-08, 2.3901e-08, 
    2.299022e-08, 2.448664e-08, 2.382222e-08, 2.400789e-08, 2.265353e-08,
  2.07697e-08, 2.01507e-08, 2.248158e-08, 2.329726e-08, 2.374635e-08, 
    2.425856e-08, 2.448685e-08, 2.537141e-08, 2.359817e-08, 2.434524e-08, 
    2.63497e-08, 2.663056e-08, 2.77902e-08, 2.617174e-08, 2.255565e-08,
  2.063609e-08, 2.094264e-08, 2.276163e-08, 2.341362e-08, 2.2892e-08, 
    2.291851e-08, 2.25637e-08, 2.395208e-08, 2.430584e-08, 2.715114e-08, 
    2.525365e-08, 2.513876e-08, 2.473637e-08, 2.256216e-08, 2.078538e-08,
  2.129266e-08, 2.086344e-08, 2.179942e-08, 2.322233e-08, 2.346513e-08, 
    2.303457e-08, 2.302891e-08, 2.281117e-08, 2.366875e-08, 2.153321e-08, 
    2.073277e-08, 2.290269e-08, 2.475406e-08, 2.2237e-08, 2.355303e-08,
  2.185491e-08, 2.059036e-08, 2.040977e-08, 2.078788e-08, 2.221525e-08, 
    2.265751e-08, 2.33652e-08, 2.341017e-08, 2.34276e-08, 2.257641e-08, 
    2.052148e-08, 2.094617e-08, 2.07514e-08, 2.143477e-08, 2.236909e-08,
  2.052857e-08, 2.10389e-08, 2.114452e-08, 2.069475e-08, 2.135644e-08, 
    2.301387e-08, 2.400049e-08, 2.445629e-08, 2.492448e-08, 2.420033e-08, 
    2.283204e-08, 2.177999e-08, 1.936533e-08, 1.992164e-08, 2.055739e-08,
  2.123617e-08, 2.129475e-08, 2.248971e-08, 2.177702e-08, 2.217562e-08, 
    2.430627e-08, 2.557329e-08, 2.678969e-08, 2.519083e-08, 2.502851e-08, 
    2.479229e-08, 2.4259e-08, 2.219484e-08, 2.120318e-08, 2.071827e-08,
  2.232306e-08, 2.190964e-08, 2.293755e-08, 2.209907e-08, 2.299966e-08, 
    2.386289e-08, 2.425194e-08, 2.463342e-08, 2.451665e-08, 2.485792e-08, 
    2.490448e-08, 2.451935e-08, 2.395628e-08, 2.344641e-08, 2.203211e-08,
  2.022722e-08, 2.002827e-08, 2.12319e-08, 2.190438e-08, 2.304509e-08, 
    2.441227e-08, 2.517771e-08, 2.571473e-08, 2.532664e-08, 2.48395e-08, 
    2.666062e-08, 2.588347e-08, 3.112788e-08, 3.002497e-08, 3.062323e-08,
  1.948802e-08, 1.836622e-08, 1.933229e-08, 2.022807e-08, 2.132722e-08, 
    2.339621e-08, 2.567119e-08, 2.66162e-08, 2.649967e-08, 2.658888e-08, 
    2.665874e-08, 2.67513e-08, 3.077622e-08, 2.885786e-08, 3.060786e-08,
  1.95912e-08, 1.879796e-08, 1.948728e-08, 1.945009e-08, 2.081912e-08, 
    2.212945e-08, 2.531381e-08, 2.547576e-08, 2.559066e-08, 2.624923e-08, 
    2.690867e-08, 2.797586e-08, 2.991391e-08, 2.801716e-08, 3.039575e-08,
  1.966212e-08, 1.866445e-08, 1.920338e-08, 2.063904e-08, 2.215161e-08, 
    2.227214e-08, 2.244598e-08, 2.434513e-08, 2.623563e-08, 2.726692e-08, 
    2.795518e-08, 2.812182e-08, 2.812146e-08, 2.802104e-08, 2.647484e-08,
  2.104758e-08, 2.006312e-08, 2.087493e-08, 2.140831e-08, 2.158594e-08, 
    2.216465e-08, 2.094377e-08, 2.207783e-08, 2.489031e-08, 2.954509e-08, 
    2.679863e-08, 2.353366e-08, 2.103545e-08, 1.906817e-08, 1.961093e-08,
  2.105523e-08, 2.114684e-08, 2.096288e-08, 2.084041e-08, 2.102848e-08, 
    2.170757e-08, 2.18948e-08, 2.203299e-08, 2.38677e-08, 2.382334e-08, 
    2.462892e-08, 2.459577e-08, 2.157261e-08, 1.824269e-08, 2.015099e-08,
  2.131734e-08, 2.141429e-08, 2.181646e-08, 2.163477e-08, 2.137747e-08, 
    2.073878e-08, 2.069896e-08, 2.10107e-08, 2.208022e-08, 2.122239e-08, 
    2.159324e-08, 2.343843e-08, 2.13007e-08, 1.922828e-08, 2.206966e-08,
  2.250736e-08, 2.17253e-08, 2.110386e-08, 2.146325e-08, 2.151012e-08, 
    2.028965e-08, 2.005447e-08, 1.994683e-08, 2.178243e-08, 2.208623e-08, 
    2.144482e-08, 2.223193e-08, 2.130443e-08, 2.013552e-08, 2.142274e-08,
  2.181824e-08, 2.126433e-08, 2.052924e-08, 2.147594e-08, 2.199871e-08, 
    2.121215e-08, 2.070082e-08, 2.057932e-08, 2.029989e-08, 2.132992e-08, 
    2.221467e-08, 2.213998e-08, 2.211973e-08, 2.137959e-08, 2.169942e-08,
  2.144995e-08, 2.10888e-08, 2.038734e-08, 2.105268e-08, 2.17548e-08, 
    2.213911e-08, 2.192013e-08, 2.167556e-08, 2.143411e-08, 2.096293e-08, 
    2.185948e-08, 2.230226e-08, 2.312905e-08, 2.318643e-08, 2.315034e-08,
  2.066437e-08, 2.053366e-08, 2.012759e-08, 1.904551e-08, 1.909392e-08, 
    1.913139e-08, 1.930546e-08, 2.063343e-08, 2.102985e-08, 2.089875e-08, 
    2.202666e-08, 2.278254e-08, 2.283903e-08, 2.695153e-08, 2.735042e-08,
  2.085352e-08, 1.996648e-08, 1.92151e-08, 1.894304e-08, 1.821257e-08, 
    1.855424e-08, 1.949957e-08, 2.074897e-08, 2.123316e-08, 2.177102e-08, 
    2.448326e-08, 2.457169e-08, 2.178985e-08, 3.113855e-08, 2.784211e-08,
  2.05376e-08, 1.951363e-08, 1.960309e-08, 1.940829e-08, 1.839459e-08, 
    1.847914e-08, 1.927672e-08, 2.07856e-08, 2.057211e-08, 2.227894e-08, 
    2.577305e-08, 2.62198e-08, 2.326708e-08, 3.260953e-08, 2.687205e-08,
  2.00398e-08, 1.950352e-08, 1.914334e-08, 1.86764e-08, 1.869641e-08, 
    1.919051e-08, 1.936413e-08, 2.02811e-08, 2.08138e-08, 2.291019e-08, 
    2.451011e-08, 2.69692e-08, 2.523476e-08, 2.918396e-08, 2.68291e-08,
  1.982302e-08, 1.880573e-08, 1.882518e-08, 1.963966e-08, 2.020257e-08, 
    2.072694e-08, 2.080961e-08, 2.133153e-08, 2.107454e-08, 2.403372e-08, 
    2.441959e-08, 2.35747e-08, 2.299413e-08, 2.001424e-08, 2.185598e-08,
  1.954854e-08, 1.90244e-08, 1.874854e-08, 1.956026e-08, 2.045101e-08, 
    2.065131e-08, 2.083206e-08, 2.068971e-08, 2.060015e-08, 2.143594e-08, 
    2.267664e-08, 2.476816e-08, 2.423653e-08, 1.964766e-08, 2.076366e-08,
  1.973973e-08, 1.906119e-08, 1.949958e-08, 1.992033e-08, 2.130363e-08, 
    2.200973e-08, 2.157781e-08, 2.056565e-08, 2.04554e-08, 2.002444e-08, 
    2.043889e-08, 2.238447e-08, 2.354874e-08, 2.033345e-08, 2.144432e-08,
  2.031849e-08, 2.053989e-08, 2.076855e-08, 2.09539e-08, 2.254348e-08, 
    2.384322e-08, 2.275114e-08, 2.109461e-08, 2.06566e-08, 2.060333e-08, 
    1.999593e-08, 1.96696e-08, 2.072309e-08, 2.072687e-08, 2.163325e-08,
  2.286009e-08, 2.137233e-08, 2.091313e-08, 2.078747e-08, 2.105855e-08, 
    2.168467e-08, 2.140965e-08, 2.089312e-08, 2.194581e-08, 2.166591e-08, 
    2.074006e-08, 1.978498e-08, 1.951939e-08, 1.984639e-08, 2.126198e-08,
  2.408725e-08, 2.285893e-08, 2.101607e-08, 2.051663e-08, 1.985391e-08, 
    2.044132e-08, 2.098117e-08, 2.292585e-08, 2.388412e-08, 2.31103e-08, 
    2.179335e-08, 2.08141e-08, 2.047895e-08, 2.006602e-08, 2.095829e-08,
  1.619957e-08, 1.7656e-08, 1.842282e-08, 1.764061e-08, 1.732892e-08, 
    1.751693e-08, 1.750667e-08, 1.819952e-08, 1.843415e-08, 1.906381e-08, 
    1.936291e-08, 2.031264e-08, 1.975805e-08, 1.986536e-08, 2.080194e-08,
  1.783523e-08, 1.81676e-08, 1.808614e-08, 1.845893e-08, 1.757286e-08, 
    1.701999e-08, 1.712942e-08, 1.792876e-08, 1.828798e-08, 1.911437e-08, 
    1.897244e-08, 1.956855e-08, 1.967365e-08, 2.044946e-08, 2.090333e-08,
  1.995087e-08, 1.931814e-08, 1.863842e-08, 1.816707e-08, 1.824302e-08, 
    1.726449e-08, 1.723325e-08, 1.812328e-08, 1.856019e-08, 1.905864e-08, 
    1.936303e-08, 1.947192e-08, 1.949211e-08, 2.047279e-08, 2.077166e-08,
  2.054909e-08, 1.938974e-08, 1.871835e-08, 1.794853e-08, 1.707284e-08, 
    1.688567e-08, 1.717803e-08, 1.773873e-08, 1.831266e-08, 1.902298e-08, 
    2.093017e-08, 2.307998e-08, 2.208402e-08, 2.215417e-08, 2.155129e-08,
  2.199378e-08, 2.129979e-08, 2.012182e-08, 1.859173e-08, 1.789456e-08, 
    1.737394e-08, 1.717987e-08, 1.79035e-08, 1.819494e-08, 1.853316e-08, 
    1.989472e-08, 2.203031e-08, 2.201136e-08, 2.112674e-08, 2.127632e-08,
  2.39772e-08, 2.337168e-08, 2.207871e-08, 2.091908e-08, 1.950546e-08, 
    1.836786e-08, 1.745906e-08, 1.76715e-08, 1.728707e-08, 1.752776e-08, 
    1.874252e-08, 1.882474e-08, 2.013943e-08, 1.981268e-08, 2.232289e-08,
  2.543867e-08, 2.598173e-08, 2.52645e-08, 2.433941e-08, 2.287503e-08, 
    2.11499e-08, 1.95598e-08, 1.86053e-08, 1.767227e-08, 1.79865e-08, 
    1.945819e-08, 1.953786e-08, 2.104952e-08, 2.000196e-08, 2.206066e-08,
  2.837344e-08, 2.971477e-08, 2.779025e-08, 2.645461e-08, 2.572254e-08, 
    2.394251e-08, 2.267372e-08, 2.193003e-08, 2.08879e-08, 2.081443e-08, 
    2.093228e-08, 2.07594e-08, 2.25239e-08, 2.042004e-08, 2.084753e-08,
  2.720228e-08, 2.833093e-08, 2.819937e-08, 2.783267e-08, 2.747011e-08, 
    2.584328e-08, 2.334733e-08, 2.231244e-08, 2.276429e-08, 2.282525e-08, 
    2.216613e-08, 2.158966e-08, 2.287073e-08, 2.165379e-08, 2.176939e-08,
  2.59835e-08, 2.292552e-08, 2.346554e-08, 2.329632e-08, 2.477032e-08, 
    2.577038e-08, 2.482925e-08, 2.388454e-08, 2.455501e-08, 2.428436e-08, 
    2.407117e-08, 2.389112e-08, 2.421464e-08, 2.37196e-08, 2.398826e-08,
  1.909739e-08, 1.881338e-08, 1.854702e-08, 1.866055e-08, 1.844637e-08, 
    1.826375e-08, 1.783101e-08, 1.758029e-08, 1.727195e-08, 1.672911e-08, 
    1.636989e-08, 1.616324e-08, 1.646891e-08, 1.672781e-08, 1.706164e-08,
  2.030477e-08, 2.101038e-08, 2.02881e-08, 1.985019e-08, 1.980591e-08, 
    1.943642e-08, 1.876196e-08, 1.86015e-08, 1.799101e-08, 1.747319e-08, 
    1.704677e-08, 1.666043e-08, 1.645722e-08, 1.622527e-08, 1.69206e-08,
  2.26221e-08, 2.179108e-08, 2.131834e-08, 2.115675e-08, 2.064668e-08, 
    2.037919e-08, 1.991501e-08, 1.944874e-08, 1.894583e-08, 1.838622e-08, 
    1.782582e-08, 1.696096e-08, 1.64527e-08, 1.604514e-08, 1.708822e-08,
  2.325405e-08, 2.287438e-08, 2.219327e-08, 2.186402e-08, 2.060384e-08, 
    2.002549e-08, 1.948901e-08, 1.947008e-08, 1.867359e-08, 1.814841e-08, 
    1.735765e-08, 1.63858e-08, 1.627773e-08, 1.60508e-08, 1.722058e-08,
  2.432694e-08, 2.476515e-08, 2.471289e-08, 2.388444e-08, 2.319252e-08, 
    2.208491e-08, 2.11515e-08, 2.018927e-08, 1.956438e-08, 1.872881e-08, 
    1.763598e-08, 1.749024e-08, 1.679352e-08, 1.721861e-08, 1.843839e-08,
  2.398821e-08, 2.475177e-08, 2.495191e-08, 2.445948e-08, 2.422294e-08, 
    2.344633e-08, 2.260323e-08, 2.16948e-08, 2.053544e-08, 2.002349e-08, 
    2.04707e-08, 1.99888e-08, 1.836164e-08, 1.825781e-08, 1.881875e-08,
  2.488687e-08, 2.597238e-08, 2.615954e-08, 2.557709e-08, 2.521727e-08, 
    2.472089e-08, 2.389775e-08, 2.318385e-08, 2.208689e-08, 2.177609e-08, 
    2.070455e-08, 2.057342e-08, 1.916294e-08, 1.858135e-08, 1.807491e-08,
  2.643633e-08, 2.626684e-08, 2.544316e-08, 2.579905e-08, 2.577775e-08, 
    2.59314e-08, 2.55661e-08, 2.490554e-08, 2.462355e-08, 2.482478e-08, 
    2.385205e-08, 2.249621e-08, 2.175154e-08, 1.979092e-08, 1.78763e-08,
  2.649793e-08, 2.511569e-08, 2.51741e-08, 2.605086e-08, 2.615588e-08, 
    2.595834e-08, 2.551529e-08, 2.459045e-08, 2.404621e-08, 2.44599e-08, 
    2.452286e-08, 2.393391e-08, 2.329067e-08, 2.178056e-08, 1.932731e-08,
  2.594411e-08, 2.628928e-08, 2.708918e-08, 2.736922e-08, 2.721638e-08, 
    2.708254e-08, 2.72185e-08, 2.702286e-08, 2.630669e-08, 2.540958e-08, 
    2.452779e-08, 2.381258e-08, 2.347213e-08, 2.232242e-08, 2.129016e-08,
  1.875055e-08, 1.890515e-08, 1.840656e-08, 1.817651e-08, 1.811246e-08, 
    1.864841e-08, 1.841299e-08, 1.88696e-08, 1.941313e-08, 1.859953e-08, 
    1.918037e-08, 1.863499e-08, 1.837597e-08, 1.793403e-08, 1.8116e-08,
  1.863088e-08, 1.876515e-08, 1.859576e-08, 1.857742e-08, 1.861938e-08, 
    1.912018e-08, 1.871981e-08, 1.95994e-08, 1.943116e-08, 1.895114e-08, 
    1.879185e-08, 1.814412e-08, 1.804986e-08, 1.812962e-08, 1.792001e-08,
  1.882469e-08, 1.801766e-08, 1.796809e-08, 1.820015e-08, 1.839279e-08, 
    1.831803e-08, 1.837647e-08, 1.897752e-08, 1.968466e-08, 1.910425e-08, 
    1.892078e-08, 1.799016e-08, 1.823768e-08, 1.792802e-08, 1.753728e-08,
  1.826931e-08, 1.711578e-08, 1.712031e-08, 1.742678e-08, 1.76064e-08, 
    1.810498e-08, 1.865766e-08, 1.974468e-08, 1.978496e-08, 1.927907e-08, 
    1.877849e-08, 1.849659e-08, 1.810873e-08, 1.784136e-08, 1.662134e-08,
  1.67028e-08, 1.561847e-08, 1.601114e-08, 1.672717e-08, 1.76912e-08, 
    1.857489e-08, 1.923527e-08, 2.016872e-08, 1.997965e-08, 1.941316e-08, 
    1.90581e-08, 2.034353e-08, 1.958734e-08, 1.834381e-08, 1.720193e-08,
  1.505786e-08, 1.498594e-08, 1.593906e-08, 1.699789e-08, 1.794842e-08, 
    1.86783e-08, 1.938698e-08, 2.00934e-08, 2.036528e-08, 2.047301e-08, 
    2.193449e-08, 2.196117e-08, 2.1556e-08, 1.913381e-08, 2.095293e-08,
  1.574656e-08, 1.616456e-08, 1.661656e-08, 1.728582e-08, 1.800207e-08, 
    1.905951e-08, 1.927645e-08, 2.013359e-08, 2.077856e-08, 2.226574e-08, 
    2.29469e-08, 2.255052e-08, 2.241649e-08, 1.987953e-08, 2.435264e-08,
  1.76937e-08, 1.836148e-08, 1.794997e-08, 1.851647e-08, 1.980222e-08, 
    2.022923e-08, 2.020546e-08, 2.065878e-08, 2.140751e-08, 2.21893e-08, 
    2.379336e-08, 2.331815e-08, 2.370591e-08, 2.267699e-08, 2.504533e-08,
  1.961656e-08, 1.961409e-08, 1.906744e-08, 1.985712e-08, 2.083653e-08, 
    2.098931e-08, 2.06523e-08, 2.077619e-08, 2.070688e-08, 2.168147e-08, 
    2.28793e-08, 2.359415e-08, 2.401715e-08, 2.488427e-08, 2.438217e-08,
  2.048945e-08, 2.04225e-08, 2.012963e-08, 1.980291e-08, 2.09401e-08, 
    2.172906e-08, 2.20021e-08, 2.144733e-08, 2.166205e-08, 2.172848e-08, 
    2.229841e-08, 2.284351e-08, 2.353073e-08, 2.418662e-08, 2.491406e-08,
  1.859687e-08, 1.882449e-08, 1.867903e-08, 1.867773e-08, 1.866355e-08, 
    1.849611e-08, 1.851529e-08, 1.858742e-08, 1.866971e-08, 1.917112e-08, 
    1.958658e-08, 1.906521e-08, 1.896755e-08, 1.79901e-08, 1.85355e-08,
  1.872058e-08, 1.857421e-08, 1.863063e-08, 1.846113e-08, 1.853165e-08, 
    1.864245e-08, 1.8774e-08, 1.897643e-08, 1.927944e-08, 1.938148e-08, 
    1.934774e-08, 1.888714e-08, 1.869942e-08, 1.854237e-08, 1.863268e-08,
  1.729969e-08, 1.762725e-08, 1.808326e-08, 1.817761e-08, 1.822231e-08, 
    1.886315e-08, 1.900213e-08, 1.904105e-08, 1.965826e-08, 1.973042e-08, 
    1.969315e-08, 1.916537e-08, 1.863975e-08, 1.927051e-08, 1.907889e-08,
  1.716789e-08, 1.753702e-08, 1.778131e-08, 1.835257e-08, 1.845667e-08, 
    1.85721e-08, 1.843128e-08, 1.852392e-08, 1.861088e-08, 1.888054e-08, 
    1.858611e-08, 1.894095e-08, 1.925853e-08, 1.955949e-08, 1.927418e-08,
  1.809578e-08, 1.80838e-08, 1.890664e-08, 1.937561e-08, 1.941849e-08, 
    1.869317e-08, 1.851448e-08, 1.777445e-08, 1.765413e-08, 1.714081e-08, 
    1.638898e-08, 1.653854e-08, 1.636564e-08, 1.692629e-08, 1.805357e-08,
  1.859009e-08, 1.885659e-08, 1.948228e-08, 2.027394e-08, 2.057473e-08, 
    2.016725e-08, 2.020052e-08, 1.957017e-08, 1.908574e-08, 1.746241e-08, 
    1.75513e-08, 1.722012e-08, 1.643016e-08, 1.565873e-08, 1.754924e-08,
  1.888573e-08, 1.93416e-08, 1.947642e-08, 2.034877e-08, 2.071583e-08, 
    2.064415e-08, 2.061129e-08, 1.978553e-08, 2.011266e-08, 1.966871e-08, 
    2.018732e-08, 1.95214e-08, 1.878103e-08, 1.702664e-08, 1.747109e-08,
  1.983063e-08, 1.941948e-08, 1.943747e-08, 2.057488e-08, 2.052962e-08, 
    2.015307e-08, 2.038883e-08, 2.021573e-08, 2.098295e-08, 2.033114e-08, 
    2.107893e-08, 2.093481e-08, 2.096988e-08, 2.038724e-08, 1.871457e-08,
  1.998934e-08, 2.025719e-08, 2.06156e-08, 2.112515e-08, 2.040015e-08, 
    2.020879e-08, 2.043244e-08, 2.220271e-08, 2.131483e-08, 2.095459e-08, 
    2.030987e-08, 2.077788e-08, 2.149554e-08, 2.109653e-08, 2.0195e-08,
  1.827552e-08, 1.976593e-08, 2.189579e-08, 2.27035e-08, 2.358279e-08, 
    2.328666e-08, 2.219838e-08, 2.08551e-08, 2.094821e-08, 2.180787e-08, 
    2.182924e-08, 2.084121e-08, 2.110451e-08, 2.178448e-08, 2.132002e-08,
  1.8773e-08, 1.855582e-08, 1.867627e-08, 1.80895e-08, 1.827409e-08, 
    1.87327e-08, 1.890192e-08, 1.90921e-08, 1.941124e-08, 1.933474e-08, 
    1.95806e-08, 1.926806e-08, 1.952558e-08, 1.923603e-08, 1.999488e-08,
  1.767106e-08, 1.790719e-08, 1.913222e-08, 1.873579e-08, 1.886794e-08, 
    1.961109e-08, 1.951415e-08, 1.931329e-08, 1.92799e-08, 1.897706e-08, 
    1.892454e-08, 2.057568e-08, 2.094962e-08, 2.090528e-08, 1.990379e-08,
  1.963905e-08, 1.902316e-08, 1.992696e-08, 1.973411e-08, 2.00341e-08, 
    2.136408e-08, 2.059242e-08, 1.96969e-08, 1.904484e-08, 1.881582e-08, 
    1.99112e-08, 2.300286e-08, 2.177151e-08, 2.200287e-08, 2.006598e-08,
  2.186409e-08, 1.971578e-08, 1.966544e-08, 2.183323e-08, 2.318549e-08, 
    2.181936e-08, 2.127429e-08, 2.086035e-08, 2.003516e-08, 2.022601e-08, 
    2.033996e-08, 1.934348e-08, 2.011183e-08, 2.085154e-08, 2.051031e-08,
  2.135947e-08, 2.177214e-08, 2.2116e-08, 2.374433e-08, 2.29788e-08, 
    2.249604e-08, 2.302857e-08, 2.113939e-08, 2.115683e-08, 2.217362e-08, 
    2.031427e-08, 1.904101e-08, 1.783866e-08, 1.765369e-08, 1.986826e-08,
  2.004554e-08, 2.061265e-08, 2.163612e-08, 2.165922e-08, 2.364608e-08, 
    2.337253e-08, 2.308123e-08, 2.314359e-08, 2.271899e-08, 2.21816e-08, 
    1.991756e-08, 1.941871e-08, 1.932786e-08, 1.809191e-08, 1.952704e-08,
  2.167192e-08, 2.207639e-08, 2.369802e-08, 2.204534e-08, 2.202848e-08, 
    2.263964e-08, 2.358167e-08, 2.374107e-08, 2.273532e-08, 2.243002e-08, 
    2.09963e-08, 1.995473e-08, 2.063749e-08, 2.177602e-08, 2.094957e-08,
  2.252337e-08, 2.298507e-08, 2.306965e-08, 2.24827e-08, 2.190654e-08, 
    2.330553e-08, 2.394283e-08, 2.341463e-08, 2.306517e-08, 2.435232e-08, 
    2.419693e-08, 2.282586e-08, 2.234453e-08, 2.162773e-08, 2.058283e-08,
  2.343443e-08, 2.588397e-08, 2.635804e-08, 2.525061e-08, 2.386121e-08, 
    2.43501e-08, 2.605756e-08, 2.397723e-08, 2.30105e-08, 2.313482e-08, 
    2.462968e-08, 2.463598e-08, 2.256025e-08, 2.205315e-08, 2.115311e-08,
  2.418287e-08, 2.316936e-08, 2.292559e-08, 2.46333e-08, 2.533356e-08, 
    2.480432e-08, 2.417333e-08, 2.247167e-08, 2.227718e-08, 2.369367e-08, 
    2.415309e-08, 2.473111e-08, 2.478052e-08, 2.331311e-08, 2.210484e-08,
  2.186477e-08, 2.427698e-08, 2.216568e-08, 1.968411e-08, 2.194403e-08, 
    2.163928e-08, 1.687895e-08, 1.430786e-08, 1.834747e-08, 2.205467e-08, 
    2.362704e-08, 2.669044e-08, 2.848274e-08, 2.439494e-08, 2.332462e-08,
  2.079756e-08, 2.322069e-08, 2.298422e-08, 1.970614e-08, 2.243824e-08, 
    2.442407e-08, 1.901446e-08, 1.366317e-08, 1.740097e-08, 2.190225e-08, 
    2.166163e-08, 2.37245e-08, 2.779021e-08, 2.142561e-08, 2.252093e-08,
  2.497944e-08, 2.323991e-08, 2.301019e-08, 2.206796e-08, 2.048662e-08, 
    2.474806e-08, 2.355986e-08, 1.883853e-08, 1.774496e-08, 2.160304e-08, 
    2.188128e-08, 2.199344e-08, 2.312527e-08, 1.705641e-08, 2.067897e-08,
  2.508414e-08, 2.30725e-08, 2.192435e-08, 2.465688e-08, 2.326513e-08, 
    2.185879e-08, 2.243193e-08, 2.097185e-08, 1.974862e-08, 2.19916e-08, 
    2.241973e-08, 2.287544e-08, 2.181948e-08, 1.748055e-08, 2.202433e-08,
  2.193882e-08, 2.205692e-08, 2.249906e-08, 2.308633e-08, 2.256878e-08, 
    2.24404e-08, 2.16966e-08, 1.919341e-08, 2.146798e-08, 2.378654e-08, 
    2.28427e-08, 2.227298e-08, 2.094051e-08, 2.033606e-08, 2.239228e-08,
  2.133763e-08, 2.090785e-08, 2.120501e-08, 2.108406e-08, 2.251072e-08, 
    2.193645e-08, 2.227168e-08, 2.041216e-08, 1.790446e-08, 1.969216e-08, 
    2.067382e-08, 2.264888e-08, 2.309674e-08, 2.121376e-08, 2.154518e-08,
  2.10193e-08, 2.108389e-08, 2.16985e-08, 1.885345e-08, 2.005352e-08, 
    2.137643e-08, 2.100704e-08, 1.999712e-08, 1.835506e-08, 1.836341e-08, 
    2.017265e-08, 2.266228e-08, 2.255291e-08, 2.080472e-08, 2.215461e-08,
  2.092495e-08, 2.027432e-08, 1.939732e-08, 1.890481e-08, 1.934155e-08, 
    2.072904e-08, 2.053121e-08, 1.927416e-08, 1.807839e-08, 1.864196e-08, 
    1.948684e-08, 2.150821e-08, 2.282335e-08, 2.452457e-08, 2.351855e-08,
  2.004686e-08, 2.030832e-08, 1.889501e-08, 1.902984e-08, 1.882269e-08, 
    1.839594e-08, 1.841144e-08, 1.714794e-08, 1.799736e-08, 1.99381e-08, 
    1.973332e-08, 2.07573e-08, 2.302348e-08, 2.378525e-08, 2.293211e-08,
  1.760189e-08, 1.85215e-08, 1.751429e-08, 1.879091e-08, 1.836662e-08, 
    1.778862e-08, 1.774681e-08, 1.710027e-08, 1.803059e-08, 2.065769e-08, 
    2.01525e-08, 2.052181e-08, 2.23352e-08, 2.338747e-08, 2.447208e-08,
  1.657527e-08, 1.757483e-08, 1.996971e-08, 1.952206e-08, 1.861014e-08, 
    1.869854e-08, 1.754083e-08, 1.442878e-08, 1.422236e-08, 1.663306e-08, 
    1.752725e-08, 1.868068e-08, 2.014561e-08, 2.028015e-08, 2.050563e-08,
  1.63543e-08, 1.700444e-08, 1.948681e-08, 2.043057e-08, 2.043431e-08, 
    2.001201e-08, 1.779461e-08, 1.58723e-08, 1.537513e-08, 1.657651e-08, 
    1.776036e-08, 1.86503e-08, 1.962901e-08, 1.998168e-08, 2.16734e-08,
  1.826075e-08, 1.757865e-08, 1.998758e-08, 2.007646e-08, 1.915247e-08, 
    1.958309e-08, 1.945016e-08, 1.917103e-08, 1.76738e-08, 1.788048e-08, 
    1.906595e-08, 1.91562e-08, 2.037523e-08, 2.108728e-08, 2.310441e-08,
  1.82617e-08, 1.836143e-08, 1.952677e-08, 1.935436e-08, 1.831436e-08, 
    1.749306e-08, 1.836019e-08, 1.961e-08, 1.860861e-08, 1.822028e-08, 
    1.924004e-08, 1.98445e-08, 2.156084e-08, 2.214018e-08, 2.262629e-08,
  1.796767e-08, 1.806181e-08, 1.958193e-08, 1.819752e-08, 1.79229e-08, 
    1.751877e-08, 1.745345e-08, 1.845471e-08, 1.815532e-08, 1.751354e-08, 
    1.898052e-08, 2.117327e-08, 2.352601e-08, 2.327299e-08, 2.223238e-08,
  1.747881e-08, 1.758479e-08, 1.873554e-08, 1.766727e-08, 1.709262e-08, 
    1.678981e-08, 1.728515e-08, 1.761232e-08, 1.739859e-08, 1.815853e-08, 
    2.035293e-08, 2.147719e-08, 2.315776e-08, 2.382006e-08, 2.183145e-08,
  1.687072e-08, 1.724706e-08, 1.874104e-08, 1.805519e-08, 1.723232e-08, 
    1.707356e-08, 1.678291e-08, 1.73645e-08, 1.802731e-08, 1.92276e-08, 
    2.154907e-08, 2.176256e-08, 2.288666e-08, 2.301407e-08, 2.225158e-08,
  1.700817e-08, 1.718104e-08, 1.884507e-08, 1.852594e-08, 1.779676e-08, 
    1.796581e-08, 1.698369e-08, 1.713627e-08, 1.853968e-08, 2.051316e-08, 
    2.154636e-08, 2.165725e-08, 2.345177e-08, 2.22699e-08, 2.106073e-08,
  1.67818e-08, 1.649133e-08, 1.866225e-08, 1.888078e-08, 1.798965e-08, 
    1.802869e-08, 1.594955e-08, 1.62426e-08, 1.966743e-08, 2.121896e-08, 
    2.153675e-08, 2.170622e-08, 2.231175e-08, 2.173259e-08, 2.082326e-08,
  1.651408e-08, 1.602709e-08, 1.878004e-08, 1.886502e-08, 1.706004e-08, 
    1.678468e-08, 1.521941e-08, 1.738845e-08, 2.115641e-08, 2.166746e-08, 
    2.140176e-08, 2.166326e-08, 2.236092e-08, 2.217472e-08, 2.197083e-08,
  1.108002e-08, 1.207748e-08, 1.302373e-08, 1.402149e-08, 1.622657e-08, 
    1.747048e-08, 1.762321e-08, 1.937683e-08, 1.990016e-08, 2.03215e-08, 
    1.919689e-08, 1.995656e-08, 2.044231e-08, 1.980361e-08, 1.94216e-08,
  1.32354e-08, 1.383349e-08, 1.391723e-08, 1.481268e-08, 1.710422e-08, 
    1.747274e-08, 1.819671e-08, 2.017877e-08, 2.086662e-08, 2.072403e-08, 
    2.046559e-08, 2.080987e-08, 2.010203e-08, 1.93095e-08, 1.92998e-08,
  1.502001e-08, 1.42411e-08, 1.444625e-08, 1.593855e-08, 1.752629e-08, 
    1.738884e-08, 1.885841e-08, 2.057031e-08, 2.09248e-08, 2.107774e-08, 
    2.076277e-08, 2.054463e-08, 1.945693e-08, 1.895038e-08, 1.944824e-08,
  1.392057e-08, 1.33066e-08, 1.438712e-08, 1.559657e-08, 1.689425e-08, 
    1.756562e-08, 1.984136e-08, 2.100505e-08, 2.11249e-08, 2.058945e-08, 
    1.879648e-08, 1.861413e-08, 1.845801e-08, 1.864869e-08, 1.851964e-08,
  1.312159e-08, 1.332424e-08, 1.438131e-08, 1.509526e-08, 1.704492e-08, 
    1.778661e-08, 2.037751e-08, 2.102422e-08, 2.008218e-08, 1.840592e-08, 
    1.862784e-08, 1.958949e-08, 1.953713e-08, 1.884989e-08, 1.850884e-08,
  1.380789e-08, 1.422968e-08, 1.503637e-08, 1.608065e-08, 1.754923e-08, 
    1.846827e-08, 2.062119e-08, 1.998495e-08, 1.916207e-08, 1.923246e-08, 
    1.951498e-08, 1.881754e-08, 1.914595e-08, 1.867984e-08, 1.753635e-08,
  1.420843e-08, 1.500588e-08, 1.578584e-08, 1.711705e-08, 1.793186e-08, 
    1.989149e-08, 2.03989e-08, 1.976852e-08, 1.979684e-08, 1.946194e-08, 
    1.887593e-08, 1.878185e-08, 1.969573e-08, 1.894521e-08, 1.721422e-08,
  1.515475e-08, 1.61092e-08, 1.687102e-08, 1.797437e-08, 1.867693e-08, 
    2.062595e-08, 2.025844e-08, 1.992041e-08, 1.951912e-08, 1.839413e-08, 
    1.819952e-08, 1.846143e-08, 1.994207e-08, 1.80624e-08, 1.653254e-08,
  1.654777e-08, 1.731522e-08, 1.765964e-08, 1.807333e-08, 1.888751e-08, 
    1.929637e-08, 1.87618e-08, 1.902926e-08, 1.917771e-08, 1.820566e-08, 
    1.727413e-08, 1.803363e-08, 1.91108e-08, 1.77549e-08, 1.654424e-08,
  1.744103e-08, 1.742799e-08, 1.756651e-08, 1.775528e-08, 1.808e-08, 
    1.782328e-08, 1.834261e-08, 1.974804e-08, 1.96588e-08, 1.731767e-08, 
    1.676265e-08, 1.816216e-08, 1.91488e-08, 1.822117e-08, 1.75916e-08,
  5.237351e-09, 5.437705e-09, 5.608242e-09, 6.269806e-09, 6.923289e-09, 
    7.431296e-09, 7.796635e-09, 8.383585e-09, 9.11591e-09, 9.605222e-09, 
    9.475887e-09, 1.068585e-08, 1.219301e-08, 1.251854e-08, 1.293684e-08,
  6.711807e-09, 7.006635e-09, 7.107813e-09, 7.215012e-09, 7.860695e-09, 
    8.373388e-09, 8.680077e-09, 9.320173e-09, 1.034268e-08, 1.078669e-08, 
    1.109994e-08, 1.20367e-08, 1.292969e-08, 1.264079e-08, 1.324785e-08,
  9.171679e-09, 9.567327e-09, 9.414873e-09, 9.579005e-09, 9.807378e-09, 
    1.037412e-08, 1.077675e-08, 1.152812e-08, 1.217418e-08, 1.2386e-08, 
    1.275509e-08, 1.363908e-08, 1.439435e-08, 1.416912e-08, 1.572436e-08,
  1.187431e-08, 1.203568e-08, 1.197976e-08, 1.202062e-08, 1.193655e-08, 
    1.216807e-08, 1.274378e-08, 1.33579e-08, 1.342838e-08, 1.357894e-08, 
    1.262077e-08, 1.349695e-08, 1.484046e-08, 1.579842e-08, 1.856452e-08,
  1.314469e-08, 1.330543e-08, 1.328783e-08, 1.310055e-08, 1.335347e-08, 
    1.349562e-08, 1.418991e-08, 1.452376e-08, 1.473721e-08, 1.350897e-08, 
    1.35399e-08, 1.556451e-08, 1.637357e-08, 1.874847e-08, 1.966066e-08,
  1.469497e-08, 1.48066e-08, 1.47709e-08, 1.497819e-08, 1.504569e-08, 
    1.538206e-08, 1.550232e-08, 1.582321e-08, 1.535951e-08, 1.517132e-08, 
    1.720384e-08, 1.734752e-08, 1.786114e-08, 2.11007e-08, 1.968122e-08,
  1.459336e-08, 1.472218e-08, 1.483362e-08, 1.518119e-08, 1.528257e-08, 
    1.588537e-08, 1.610734e-08, 1.675127e-08, 1.653597e-08, 1.75452e-08, 
    1.817997e-08, 1.827585e-08, 2.020232e-08, 2.280414e-08, 1.934891e-08,
  1.486273e-08, 1.511724e-08, 1.551997e-08, 1.59832e-08, 1.647296e-08, 
    1.729567e-08, 1.795419e-08, 1.848639e-08, 1.842237e-08, 1.935527e-08, 
    2.006722e-08, 2.095514e-08, 2.390862e-08, 2.268362e-08, 1.969956e-08,
  1.586696e-08, 1.648508e-08, 1.708464e-08, 1.791478e-08, 1.849916e-08, 
    1.915942e-08, 1.985408e-08, 2.012481e-08, 2.052786e-08, 2.193918e-08, 
    2.369908e-08, 2.485519e-08, 2.641574e-08, 2.490471e-08, 2.392476e-08,
  1.715132e-08, 1.795424e-08, 1.85721e-08, 1.956415e-08, 2.016811e-08, 
    2.070019e-08, 2.119629e-08, 2.221934e-08, 2.404971e-08, 2.602616e-08, 
    2.748286e-08, 2.835278e-08, 2.901126e-08, 2.796574e-08, 2.819043e-08,
  1.149092e-08, 1.152502e-08, 1.14777e-08, 1.102492e-08, 1.070943e-08, 
    1.033456e-08, 9.875994e-09, 9.57196e-09, 8.989065e-09, 8.845633e-09, 
    8.964354e-09, 8.803132e-09, 8.736952e-09, 8.978542e-09, 9.034598e-09,
  1.200602e-08, 1.176717e-08, 1.187669e-08, 1.196615e-08, 1.165252e-08, 
    1.133668e-08, 1.132986e-08, 1.11405e-08, 1.086859e-08, 1.078739e-08, 
    1.095976e-08, 1.098465e-08, 1.112198e-08, 1.132246e-08, 1.129707e-08,
  1.208183e-08, 1.202929e-08, 1.19455e-08, 1.217408e-08, 1.213227e-08, 
    1.228049e-08, 1.241915e-08, 1.238099e-08, 1.251174e-08, 1.258302e-08, 
    1.284545e-08, 1.280935e-08, 1.301753e-08, 1.299709e-08, 1.317491e-08,
  1.225189e-08, 1.234619e-08, 1.223842e-08, 1.215966e-08, 1.232335e-08, 
    1.246683e-08, 1.236327e-08, 1.250124e-08, 1.255888e-08, 1.284912e-08, 
    1.290833e-08, 1.273345e-08, 1.291139e-08, 1.308446e-08, 1.377897e-08,
  1.221217e-08, 1.229404e-08, 1.237364e-08, 1.238495e-08, 1.248139e-08, 
    1.24704e-08, 1.263414e-08, 1.260631e-08, 1.298864e-08, 1.31354e-08, 
    1.307918e-08, 1.397509e-08, 1.458779e-08, 1.526597e-08, 1.6706e-08,
  1.222778e-08, 1.239892e-08, 1.235101e-08, 1.250197e-08, 1.251731e-08, 
    1.283323e-08, 1.304289e-08, 1.402247e-08, 1.459218e-08, 1.591217e-08, 
    1.692592e-08, 1.802314e-08, 1.892074e-08, 2.001628e-08, 2.085398e-08,
  1.309756e-08, 1.313003e-08, 1.346688e-08, 1.380616e-08, 1.460255e-08, 
    1.571188e-08, 1.7406e-08, 1.89264e-08, 2.052838e-08, 2.101568e-08, 
    2.106467e-08, 2.105839e-08, 2.022718e-08, 2.114692e-08, 1.994115e-08,
  1.567459e-08, 1.606979e-08, 1.667444e-08, 1.76936e-08, 1.928525e-08, 
    2.096791e-08, 2.219173e-08, 2.221466e-08, 2.166884e-08, 2.006037e-08, 
    1.89357e-08, 1.707584e-08, 1.723576e-08, 1.638781e-08, 1.377057e-08,
  1.731704e-08, 1.790821e-08, 1.920921e-08, 2.135462e-08, 2.285221e-08, 
    2.318357e-08, 2.141864e-08, 2.075801e-08, 1.923908e-08, 1.657484e-08, 
    1.517028e-08, 1.452267e-08, 1.516168e-08, 1.468558e-08, 1.303265e-08,
  1.888439e-08, 2.014341e-08, 2.32826e-08, 2.440192e-08, 2.370371e-08, 
    2.336033e-08, 2.186321e-08, 1.823101e-08, 1.442073e-08, 1.323137e-08, 
    1.297508e-08, 1.315183e-08, 1.406065e-08, 1.426794e-08, 1.544698e-08,
  1.189469e-08, 1.179945e-08, 1.178367e-08, 1.210152e-08, 1.22606e-08, 
    1.251687e-08, 1.257166e-08, 1.285684e-08, 1.301524e-08, 1.305526e-08, 
    1.290335e-08, 1.288978e-08, 1.324299e-08, 1.290251e-08, 1.303605e-08,
  1.38323e-08, 1.382746e-08, 1.343708e-08, 1.34095e-08, 1.356072e-08, 
    1.358455e-08, 1.351347e-08, 1.369566e-08, 1.37229e-08, 1.361708e-08, 
    1.356594e-08, 1.358861e-08, 1.368099e-08, 1.344304e-08, 1.347984e-08,
  1.454057e-08, 1.443981e-08, 1.421795e-08, 1.394502e-08, 1.380086e-08, 
    1.373294e-08, 1.365267e-08, 1.371581e-08, 1.367831e-08, 1.377552e-08, 
    1.362887e-08, 1.362189e-08, 1.356604e-08, 1.330212e-08, 1.332265e-08,
  1.58054e-08, 1.588023e-08, 1.546574e-08, 1.530635e-08, 1.506751e-08, 
    1.49191e-08, 1.467646e-08, 1.446031e-08, 1.446352e-08, 1.424064e-08, 
    1.449831e-08, 1.424432e-08, 1.405994e-08, 1.370056e-08, 1.34107e-08,
  1.640624e-08, 1.643062e-08, 1.624726e-08, 1.591422e-08, 1.566793e-08, 
    1.538581e-08, 1.526213e-08, 1.497295e-08, 1.516825e-08, 1.529215e-08, 
    1.491963e-08, 1.540787e-08, 1.561302e-08, 1.50653e-08, 1.45456e-08,
  1.770793e-08, 1.767125e-08, 1.734158e-08, 1.715864e-08, 1.662942e-08, 
    1.65099e-08, 1.608488e-08, 1.611629e-08, 1.612687e-08, 1.591365e-08, 
    1.600567e-08, 1.553218e-08, 1.567953e-08, 1.564071e-08, 1.499863e-08,
  1.854607e-08, 1.807646e-08, 1.790432e-08, 1.711534e-08, 1.67795e-08, 
    1.632237e-08, 1.628015e-08, 1.624965e-08, 1.701702e-08, 1.614405e-08, 
    1.563147e-08, 1.520112e-08, 1.501457e-08, 1.754836e-08, 1.410937e-08,
  1.932333e-08, 1.877012e-08, 1.784254e-08, 1.714318e-08, 1.691441e-08, 
    1.644536e-08, 1.698062e-08, 1.707973e-08, 1.694379e-08, 1.600719e-08, 
    1.567212e-08, 1.452883e-08, 1.525632e-08, 1.476498e-08, 1.19157e-08,
  1.862994e-08, 1.834974e-08, 1.777446e-08, 1.774285e-08, 1.776279e-08, 
    1.819804e-08, 1.834206e-08, 1.803873e-08, 1.726462e-08, 1.548515e-08, 
    1.388967e-08, 1.308757e-08, 1.464485e-08, 1.298729e-08, 1.298123e-08,
  1.898592e-08, 1.832542e-08, 1.875453e-08, 1.957597e-08, 1.999698e-08, 
    2.082347e-08, 1.951618e-08, 1.843412e-08, 1.307305e-08, 1.221569e-08, 
    1.261053e-08, 1.411255e-08, 1.549144e-08, 1.601291e-08, 1.683909e-08,
  1.440654e-08, 1.446911e-08, 1.451933e-08, 1.463786e-08, 1.455622e-08, 
    1.423912e-08, 1.392003e-08, 1.362881e-08, 1.345715e-08, 1.284959e-08, 
    1.224649e-08, 1.200452e-08, 1.222276e-08, 1.197133e-08, 1.209893e-08,
  1.82615e-08, 1.848006e-08, 1.825961e-08, 1.798212e-08, 1.800943e-08, 
    1.779894e-08, 1.744683e-08, 1.726346e-08, 1.69621e-08, 1.645286e-08, 
    1.610094e-08, 1.589433e-08, 1.594309e-08, 1.563097e-08, 1.593542e-08,
  1.997236e-08, 2.08711e-08, 2.100182e-08, 2.114012e-08, 2.093443e-08, 
    2.112595e-08, 2.088193e-08, 2.076187e-08, 2.045003e-08, 2.00976e-08, 
    1.983705e-08, 1.952418e-08, 1.951776e-08, 1.920488e-08, 1.955907e-08,
  2.109764e-08, 2.179645e-08, 2.178223e-08, 2.202537e-08, 2.228426e-08, 
    2.237433e-08, 2.218607e-08, 2.207902e-08, 2.190882e-08, 2.161407e-08, 
    2.189194e-08, 2.149326e-08, 2.120939e-08, 2.07463e-08, 2.042708e-08,
  2.101708e-08, 2.147389e-08, 2.199908e-08, 2.203094e-08, 2.200734e-08, 
    2.181866e-08, 2.141281e-08, 2.115977e-08, 2.122587e-08, 2.17072e-08, 
    2.125043e-08, 2.160826e-08, 2.144359e-08, 2.069151e-08, 1.912406e-08,
  2.253687e-08, 2.259736e-08, 2.299825e-08, 2.317836e-08, 2.265576e-08, 
    2.251864e-08, 2.226986e-08, 2.237902e-08, 2.325686e-08, 2.297463e-08, 
    2.119828e-08, 2.026401e-08, 1.943424e-08, 1.875799e-08, 1.756276e-08,
  2.228278e-08, 2.241761e-08, 2.259847e-08, 2.221252e-08, 2.223565e-08, 
    2.197672e-08, 2.172012e-08, 2.09643e-08, 2.06143e-08, 1.803313e-08, 
    1.734643e-08, 1.628145e-08, 1.619339e-08, 1.747066e-08, 1.53138e-08,
  2.286287e-08, 2.219948e-08, 2.135886e-08, 2.090655e-08, 2.016388e-08, 
    1.917911e-08, 1.864127e-08, 1.785718e-08, 1.714383e-08, 1.638943e-08, 
    1.619899e-08, 1.567963e-08, 1.704297e-08, 1.675775e-08, 1.621613e-08,
  2.019124e-08, 2.009304e-08, 1.998502e-08, 1.980527e-08, 1.915963e-08, 
    1.88517e-08, 1.830808e-08, 1.768052e-08, 1.670495e-08, 1.642107e-08, 
    1.623922e-08, 1.66209e-08, 1.780041e-08, 1.78215e-08, 1.864845e-08,
  2.074129e-08, 2.076423e-08, 2.073193e-08, 2.036306e-08, 2.016068e-08, 
    1.995748e-08, 1.856982e-08, 1.658528e-08, 1.623943e-08, 1.647984e-08, 
    1.757595e-08, 1.832544e-08, 1.889279e-08, 1.962742e-08, 2.033097e-08,
  9.995578e-09, 1.043659e-08, 1.062557e-08, 1.098163e-08, 1.124657e-08, 
    1.157428e-08, 1.174493e-08, 1.218346e-08, 1.271215e-08, 1.267224e-08, 
    1.247891e-08, 1.279694e-08, 1.362184e-08, 1.380026e-08, 1.394212e-08,
  1.310916e-08, 1.341313e-08, 1.356548e-08, 1.379917e-08, 1.433532e-08, 
    1.472373e-08, 1.490655e-08, 1.55413e-08, 1.586935e-08, 1.605001e-08, 
    1.621111e-08, 1.647865e-08, 1.700089e-08, 1.710784e-08, 1.745996e-08,
  1.524456e-08, 1.530302e-08, 1.559164e-08, 1.601612e-08, 1.65665e-08, 
    1.689108e-08, 1.713768e-08, 1.765072e-08, 1.817818e-08, 1.846318e-08, 
    1.892939e-08, 1.923991e-08, 1.959688e-08, 1.975573e-08, 2.020837e-08,
  1.658689e-08, 1.650424e-08, 1.666507e-08, 1.698108e-08, 1.720812e-08, 
    1.750541e-08, 1.79289e-08, 1.851987e-08, 1.920241e-08, 1.960234e-08, 
    2.044019e-08, 2.1094e-08, 2.123444e-08, 2.150299e-08, 2.168082e-08,
  1.746746e-08, 1.733751e-08, 1.77756e-08, 1.818587e-08, 1.866309e-08, 
    1.928758e-08, 1.979133e-08, 2.053151e-08, 2.101287e-08, 2.151702e-08, 
    2.179848e-08, 2.248014e-08, 2.293711e-08, 2.262749e-08, 2.155713e-08,
  1.849426e-08, 1.860206e-08, 1.911074e-08, 1.950468e-08, 2.016971e-08, 
    2.059331e-08, 2.103358e-08, 2.114501e-08, 2.154556e-08, 2.15075e-08, 
    2.138483e-08, 2.111914e-08, 2.151627e-08, 2.123965e-08, 2.074198e-08,
  1.845606e-08, 1.886525e-08, 1.939805e-08, 1.980398e-08, 2.044445e-08, 
    2.082768e-08, 2.131363e-08, 2.153163e-08, 2.214823e-08, 2.115524e-08, 
    2.128288e-08, 2.108264e-08, 2.136424e-08, 2.027198e-08, 2.017355e-08,
  2.01012e-08, 2.007774e-08, 2.031223e-08, 2.052373e-08, 2.116631e-08, 
    2.12674e-08, 2.175281e-08, 2.167535e-08, 2.184542e-08, 2.114704e-08, 
    2.168523e-08, 2.131841e-08, 2.131328e-08, 2.018431e-08, 2.009643e-08,
  1.933269e-08, 1.938191e-08, 2.011059e-08, 2.058551e-08, 2.115334e-08, 
    2.146838e-08, 2.168745e-08, 2.217092e-08, 2.13133e-08, 2.194426e-08, 
    2.1956e-08, 2.100922e-08, 2.04901e-08, 1.951793e-08, 1.988555e-08,
  2.018401e-08, 2.01896e-08, 2.111086e-08, 2.135271e-08, 2.200292e-08, 
    2.24308e-08, 2.277024e-08, 2.246897e-08, 2.213853e-08, 2.215695e-08, 
    2.10487e-08, 2.036026e-08, 1.993312e-08, 2.098269e-08, 2.171352e-08,
  6.580434e-09, 6.923285e-09, 7.245577e-09, 7.56609e-09, 7.80468e-09, 
    8.139806e-09, 8.272408e-09, 8.715998e-09, 9.221032e-09, 9.66411e-09, 
    9.939469e-09, 1.051629e-08, 1.154992e-08, 1.202989e-08, 1.262341e-08,
  8.297468e-09, 8.792081e-09, 8.9023e-09, 9.021813e-09, 9.425249e-09, 
    9.505464e-09, 9.710178e-09, 1.034282e-08, 1.103457e-08, 1.146474e-08, 
    1.188186e-08, 1.25814e-08, 1.330564e-08, 1.37993e-08, 1.452771e-08,
  1.033484e-08, 1.047797e-08, 1.054023e-08, 1.075889e-08, 1.103081e-08, 
    1.139945e-08, 1.160706e-08, 1.229344e-08, 1.298853e-08, 1.321335e-08, 
    1.366792e-08, 1.427e-08, 1.476166e-08, 1.529451e-08, 1.608094e-08,
  1.254559e-08, 1.275355e-08, 1.284912e-08, 1.313214e-08, 1.308927e-08, 
    1.328413e-08, 1.357893e-08, 1.404347e-08, 1.43698e-08, 1.458525e-08, 
    1.492507e-08, 1.588523e-08, 1.649647e-08, 1.714715e-08, 1.781291e-08,
  1.473623e-08, 1.474214e-08, 1.484101e-08, 1.481652e-08, 1.499671e-08, 
    1.516269e-08, 1.550991e-08, 1.580575e-08, 1.571093e-08, 1.552482e-08, 
    1.605016e-08, 1.84631e-08, 1.913015e-08, 1.936597e-08, 1.911009e-08,
  1.803107e-08, 1.780854e-08, 1.786686e-08, 1.78947e-08, 1.792394e-08, 
    1.7837e-08, 1.780464e-08, 1.758714e-08, 1.733817e-08, 1.764419e-08, 
    1.883661e-08, 1.857771e-08, 1.974613e-08, 1.97442e-08, 2.012365e-08,
  1.962314e-08, 1.94919e-08, 1.960452e-08, 1.96476e-08, 1.952387e-08, 
    1.948893e-08, 1.922723e-08, 1.89037e-08, 1.91522e-08, 1.927578e-08, 
    1.938801e-08, 1.94516e-08, 2.082766e-08, 2.134995e-08, 2.206303e-08,
  2.244161e-08, 2.224461e-08, 2.221372e-08, 2.207523e-08, 2.196061e-08, 
    2.185386e-08, 2.154237e-08, 2.137963e-08, 2.102374e-08, 2.075802e-08, 
    2.088562e-08, 2.082303e-08, 2.227642e-08, 2.245145e-08, 2.361723e-08,
  2.452392e-08, 2.420499e-08, 2.390146e-08, 2.363859e-08, 2.326934e-08, 
    2.298854e-08, 2.25399e-08, 2.202905e-08, 2.146428e-08, 2.172101e-08, 
    2.180043e-08, 2.200136e-08, 2.256624e-08, 2.358572e-08, 2.358542e-08,
  2.563108e-08, 2.536696e-08, 2.483491e-08, 2.460657e-08, 2.422074e-08, 
    2.399661e-08, 2.35283e-08, 2.321726e-08, 2.344688e-08, 2.332091e-08, 
    2.3294e-08, 2.348255e-08, 2.35196e-08, 2.402979e-08, 2.376943e-08,
  6.036434e-09, 6.56103e-09, 6.980991e-09, 7.284865e-09, 7.56961e-09, 
    7.803991e-09, 7.985181e-09, 8.206786e-09, 8.635275e-09, 8.741168e-09, 
    9.131411e-09, 9.576649e-09, 1.057482e-08, 1.117742e-08, 1.207487e-08,
  1.009606e-08, 1.059814e-08, 1.06897e-08, 1.094064e-08, 1.11391e-08, 
    1.134092e-08, 1.126439e-08, 1.155684e-08, 1.183553e-08, 1.188054e-08, 
    1.231474e-08, 1.273034e-08, 1.371618e-08, 1.429408e-08, 1.518761e-08,
  1.357578e-08, 1.409051e-08, 1.413151e-08, 1.416375e-08, 1.410493e-08, 
    1.449398e-08, 1.438042e-08, 1.483699e-08, 1.505055e-08, 1.542988e-08, 
    1.595606e-08, 1.645653e-08, 1.746348e-08, 1.784454e-08, 1.903782e-08,
  1.680415e-08, 1.750931e-08, 1.728042e-08, 1.720571e-08, 1.738618e-08, 
    1.777335e-08, 1.802574e-08, 1.853179e-08, 1.894961e-08, 1.934784e-08, 
    1.989248e-08, 2.028279e-08, 2.101664e-08, 2.1098e-08, 2.240917e-08,
  1.950247e-08, 1.982805e-08, 2.015335e-08, 2.039079e-08, 2.095034e-08, 
    2.146286e-08, 2.19818e-08, 2.232648e-08, 2.278684e-08, 2.266672e-08, 
    2.220271e-08, 2.372791e-08, 2.449052e-08, 2.465912e-08, 2.477994e-08,
  2.128048e-08, 2.177275e-08, 2.234392e-08, 2.333891e-08, 2.397557e-08, 
    2.452779e-08, 2.50398e-08, 2.545978e-08, 2.535123e-08, 2.53011e-08, 
    2.579861e-08, 2.536361e-08, 2.562565e-08, 2.578449e-08, 2.603051e-08,
  2.22521e-08, 2.355621e-08, 2.403324e-08, 2.470492e-08, 2.491515e-08, 
    2.572849e-08, 2.623904e-08, 2.669187e-08, 2.69219e-08, 2.700691e-08, 
    2.681219e-08, 2.671152e-08, 2.729332e-08, 2.761461e-08, 2.854175e-08,
  2.477008e-08, 2.466972e-08, 2.413323e-08, 2.490506e-08, 2.512137e-08, 
    2.592156e-08, 2.622444e-08, 2.681273e-08, 2.711858e-08, 2.69232e-08, 
    2.709414e-08, 2.694619e-08, 2.7773e-08, 2.826025e-08, 2.998642e-08,
  2.21695e-08, 2.294449e-08, 2.382104e-08, 2.434309e-08, 2.425662e-08, 
    2.48143e-08, 2.479372e-08, 2.585324e-08, 2.566018e-08, 2.662522e-08, 
    2.699174e-08, 2.738438e-08, 2.861536e-08, 3.009951e-08, 3.057248e-08,
  2.267731e-08, 2.372628e-08, 2.374894e-08, 2.254698e-08, 2.231336e-08, 
    2.254967e-08, 2.341521e-08, 2.518448e-08, 2.692211e-08, 2.738502e-08, 
    2.788557e-08, 2.899466e-08, 2.873573e-08, 2.934476e-08, 2.877373e-08,
  3.496958e-09, 3.992793e-09, 4.562559e-09, 5.413475e-09, 6.357168e-09, 
    7.62464e-09, 9.018631e-09, 1.078514e-08, 1.203202e-08, 1.314437e-08, 
    1.532951e-08, 1.619066e-08, 1.738429e-08, 1.768499e-08, 1.804857e-08,
  5.38722e-09, 6.027394e-09, 6.716021e-09, 7.804445e-09, 8.87753e-09, 
    1.05606e-08, 1.211602e-08, 1.355291e-08, 1.443565e-08, 1.606928e-08, 
    1.760213e-08, 1.795645e-08, 1.940874e-08, 1.936938e-08, 2.044234e-08,
  7.624509e-09, 9.001592e-09, 1.006777e-08, 1.139401e-08, 1.256298e-08, 
    1.433481e-08, 1.496038e-08, 1.59559e-08, 1.665076e-08, 1.793131e-08, 
    1.842195e-08, 1.877664e-08, 2.038086e-08, 2.014097e-08, 2.181348e-08,
  1.145621e-08, 1.320255e-08, 1.374395e-08, 1.430057e-08, 1.517233e-08, 
    1.587403e-08, 1.619982e-08, 1.688805e-08, 1.78802e-08, 1.903484e-08, 
    1.975578e-08, 2.117578e-08, 2.188473e-08, 2.188124e-08, 2.244189e-08,
  1.466655e-08, 1.64992e-08, 1.711507e-08, 1.768791e-08, 1.816726e-08, 
    1.842477e-08, 1.852146e-08, 1.898319e-08, 1.991864e-08, 1.977931e-08, 
    2.038069e-08, 2.117603e-08, 2.10987e-08, 2.081065e-08, 2.13524e-08,
  1.771547e-08, 1.817068e-08, 1.814497e-08, 1.830688e-08, 1.809836e-08, 
    1.801429e-08, 1.788819e-08, 1.846094e-08, 1.824232e-08, 1.876874e-08, 
    1.929225e-08, 1.93186e-08, 1.995555e-08, 2.059127e-08, 2.205157e-08,
  1.763268e-08, 1.775082e-08, 1.78833e-08, 1.812243e-08, 1.821594e-08, 
    1.809967e-08, 1.81945e-08, 1.821932e-08, 1.856687e-08, 1.935218e-08, 
    2.008578e-08, 2.048952e-08, 2.165642e-08, 2.231013e-08, 2.362749e-08,
  1.84236e-08, 1.834832e-08, 1.858745e-08, 1.872888e-08, 1.890432e-08, 
    1.92583e-08, 1.938191e-08, 1.947618e-08, 2.048643e-08, 2.114092e-08, 
    2.169678e-08, 2.171412e-08, 2.244149e-08, 2.360954e-08, 2.433558e-08,
  1.780781e-08, 1.865125e-08, 1.927801e-08, 2.052779e-08, 2.137191e-08, 
    2.178281e-08, 2.128835e-08, 2.116028e-08, 2.145476e-08, 2.210757e-08, 
    2.221717e-08, 2.193518e-08, 2.26661e-08, 2.373844e-08, 2.41294e-08,
  2.132143e-08, 2.184093e-08, 2.22422e-08, 2.287168e-08, 2.298249e-08, 
    2.255442e-08, 2.139571e-08, 2.143994e-08, 2.152083e-08, 2.123468e-08, 
    2.113857e-08, 2.150255e-08, 2.207122e-08, 2.307485e-08, 2.433868e-08,
  3.607688e-09, 4.042306e-09, 4.5913e-09, 5.392871e-09, 6.262737e-09, 
    7.165985e-09, 8.286158e-09, 9.601941e-09, 1.049789e-08, 1.161382e-08, 
    1.329951e-08, 1.451718e-08, 1.568415e-08, 1.638595e-08, 1.702005e-08,
  6.202184e-09, 6.853059e-09, 7.566072e-09, 8.500368e-09, 9.342282e-09, 
    1.057391e-08, 1.179826e-08, 1.278621e-08, 1.338485e-08, 1.458297e-08, 
    1.601977e-08, 1.657058e-08, 1.779493e-08, 1.79844e-08, 1.830572e-08,
  9.598152e-09, 1.157937e-08, 1.202698e-08, 1.311184e-08, 1.358682e-08, 
    1.509708e-08, 1.545298e-08, 1.589845e-08, 1.617071e-08, 1.734775e-08, 
    1.789218e-08, 1.761681e-08, 1.881852e-08, 1.813211e-08, 1.900398e-08,
  1.430861e-08, 1.571323e-08, 1.571174e-08, 1.570488e-08, 1.623235e-08, 
    1.666325e-08, 1.678958e-08, 1.69899e-08, 1.740544e-08, 1.835115e-08, 
    1.752866e-08, 1.860968e-08, 1.895094e-08, 1.892578e-08, 2.060064e-08,
  1.717224e-08, 1.840586e-08, 1.8773e-08, 1.891426e-08, 1.916336e-08, 
    1.916223e-08, 1.933468e-08, 1.919063e-08, 1.961252e-08, 1.836191e-08, 
    1.810043e-08, 1.857842e-08, 1.837511e-08, 1.916177e-08, 2.073032e-08,
  1.92291e-08, 1.948491e-08, 1.918685e-08, 1.948411e-08, 1.887358e-08, 
    1.890903e-08, 1.871052e-08, 1.873212e-08, 1.772453e-08, 1.770937e-08, 
    1.86796e-08, 1.89294e-08, 2.039503e-08, 2.239426e-08, 2.594715e-08,
  1.888238e-08, 1.889284e-08, 1.883165e-08, 1.88543e-08, 1.88188e-08, 
    1.893049e-08, 1.87034e-08, 1.83031e-08, 1.757209e-08, 1.915942e-08, 
    2.128331e-08, 2.358206e-08, 2.692912e-08, 2.904975e-08, 2.969699e-08,
  1.909956e-08, 1.903588e-08, 1.891781e-08, 1.88893e-08, 1.869151e-08, 
    1.833923e-08, 1.799815e-08, 1.784692e-08, 1.87879e-08, 2.184403e-08, 
    2.546385e-08, 2.75212e-08, 2.853151e-08, 2.812643e-08, 2.626439e-08,
  1.810371e-08, 1.823544e-08, 1.805386e-08, 1.80026e-08, 1.732927e-08, 
    1.814991e-08, 1.886967e-08, 2.081742e-08, 2.271464e-08, 2.704054e-08, 
    2.892066e-08, 2.867714e-08, 2.781289e-08, 2.560744e-08, 2.472756e-08,
  1.908599e-08, 1.866751e-08, 1.847671e-08, 1.877654e-08, 1.96883e-08, 
    2.179586e-08, 2.333855e-08, 2.632158e-08, 2.956516e-08, 2.979533e-08, 
    2.873588e-08, 2.699393e-08, 2.542228e-08, 2.490924e-08, 2.469751e-08 ;

 sftlf =
  0.0008770345, 0.4596241, 0.9892928, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.01035247, 0.004304647, 0.6546783, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.8534847, 0.8118016, 0.9951549, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9894952, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4452189, 0.3028796, 0.7140614, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9903189, 0.3150955, 0.0007410151, 0, 0.02645395, 
    0.9012984, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.681631, 0, 0, 0, 0.004980796, 0.7708192, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5536854, 0, 0, 0, 0.004666397, 0.9395298, 1,
  1, 1, 1, 1, 1, 1, 1, 0.9995009, 0.3626226, 0, 0, 0, 0, 0.8367797, 1,
  1, 1, 1, 1, 1, 0.8451425, 0.7016711, 0.3953246, 0, 0, 0, 0, 0.006316811, 
    0.8673657, 1 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0.2038203, 25.08469, 362.922, 581.3585, 583.7158, 677.0037, 892.3406, 
    840.3151, 1394.918, 1845.667, 2078.668, 2048.803, 1746.472, 1895.031, 
    903.5963,
  0.04938461, 3.284697, 202.5217, 654.3141, 903.2668, 1076.606, 1196.302, 
    1163.293, 1639.916, 1906.256, 1988.945, 1916.741, 1695.228, 1807.269, 
    774.2457,
  790.1076, 1114.346, 653.3495, 780.126, 1392.106, 1491.591, 1273.753, 
    1344.373, 1825.463, 2046.944, 2142.644, 2067.535, 1930.862, 1770.506, 
    591.146,
  1359.809, 1341.669, 1435.043, 1594.124, 1615.893, 1763.274, 1677.539, 
    1645.991, 1875.931, 2003.645, 2040.039, 1879.801, 1919.839, 1717.029, 
    1138.974,
  1205.389, 1290.31, 1192.454, 1271.409, 1283.839, 1439.06, 1538.882, 
    1587.552, 1685.139, 1482.705, 108.3495, 67.86669, 940.4369, 898.4109, 
    1612.947,
  1168.617, 1342.769, 1106.133, 1029.211, 1110.353, 1151.071, 1218.088, 
    1182.275, 1031.226, 58.02261, 0, 0, 7.641389, 710.6758, 2161.482,
  1244.873, 1316.863, 1112.963, 998.5415, 1017.03, 1014.576, 1020.14, 
    838.6226, 484.287, 0, 0, 0, 0, 1273.715, 2180.106,
  896.0552, 1198.27, 1151.006, 981.8504, 1010.922, 1103.887, 1045.003, 
    880.1057, 498.0692, 0, 0, 0, 0, 1386.297, 1186.975,
  625.923, 1015.673, 1096.604, 994.0698, 1069.039, 1288.357, 1166.806, 
    927.0013, 34.64387, 0, 0, 0, 0, 678.2806, 439.0615,
  346.5426, 755.811, 896.7624, 677.1516, 656.058, 642.5463, 557.833, 
    41.91994, 0, 0, 0, 0, 0, 191.3587, 93.07086 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
