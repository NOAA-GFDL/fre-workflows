netcdf \00010101.river_month.tile3.rv_o_h2o {
dimensions:
	time = UNLIMITED ; // (12 currently)
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float rv_o_h2o(time, grid_yt, grid_xt) ;
		rv_o_h2o:_FillValue = -1.e+08f ;
		rv_o_h2o:missing_value = -1.e+08f ;
		rv_o_h2o:units = "kg/m2/s" ;
		rv_o_h2o:long_name = "river outflow, h2o mass" ;
		rv_o_h2o:cell_methods = "time: mean" ;
		rv_o_h2o:time_avg_info = "average_T1,average_T2,average_DT" ;
		rv_o_h2o:coordinates = "geolon_t geolat_t" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "areacellr: 00010101.river_static_cmip.nc land_area: 00010101.river_static.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Fri Aug 29 14:00:37 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 /work/cew/scratch//00010101.river_month.tile3.nc -O /work/cew/scratch/workflow-test/river_month//ncks_out//00010101.river_month.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31 ;

 average_T1 = 0, 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334 ;

 average_T2 = 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365 ;

 rv_o_h2o =
  0, 0, 0, 2.617788e-05, 8.186758e-05, 6.900839e-12, 4.116433e-06, 
    5.929878e-07, 1.349762e-05, 4.493743e-06, 1.6689e-10, 2.530915e-06, 
    2.021267e-05, 5.420628e-06, 1.002553e-06,
  0, 0, 0, 5.694516e-06, 2.586676e-05, 8.099945e-05, 6.252433e-05, 
    7.424063e-06, 1.49471e-06, 2.339164e-05, 1.741806e-06, 2.068686e-06, 
    1.138043e-05, 1.928165e-11, 2.86131e-14,
  0, 0, 0, 1.816367e-05, 1.993692e-05, 5.029997e-06, 1.026228e-05, 
    5.062478e-05, 3.525908e-05, 5.091795e-06, 1.337564e-06, 4.784417e-06, 
    2.885943e-06, 5.272891e-06, 1.777017e-05,
  1.593423e-05, 1.966898e-13, 2.629285e-09, 9.220214e-06, 1.152539e-05, 
    5.957476e-06, 4.503292e-06, 5.446961e-07, 2.927227e-07, 4.786777e-06, 
    8.812933e-06, 1.398506e-05, 8.988744e-06, 7.394308e-06, 1.104133e-05,
  0, 5.676227e-06, 5.222429e-12, 5.771615e-06, 8.860171e-06, 2.370434e-06, 
    1.323546e-07, 2.958676e-06, 4.235656e-06, 3.577832e-05, 0, 0, 0, 
    2.158154e-06, 5.264946e-07,
  5.941721e-06, 5.34326e-06, 5.45018e-06, 1.429054e-13, 2.08965e-05, 
    1.084888e-06, 2.448143e-06, 5.704496e-07, 0, 0, 0, _, 0, 0, 6.209046e-06,
  4.223536e-06, 3.29576e-06, 1.532907e-05, 4.088094e-06, 1.696128e-05, 
    4.474788e-05, 2.629169e-06, 2.946117e-13, 0, _, _, _, 0, 0, 3.532655e-06,
  7.961248e-14, 5.582266e-06, 6.818887e-06, 1.236927e-05, 5.262688e-06, 
    3.092101e-06, 5.797918e-05, 1.370204e-07, 0, _, _, _, 0, 0, 3.019533e-06,
  3.746007e-13, 3.713347e-06, 9.831861e-07, 8.442126e-06, 8.392013e-07, 
    9.982789e-06, 1.168739e-07, 0, 0, _, _, _, _, 0, 4.781598e-07,
  1.383847e-06, 9.102887e-06, 6.461074e-06, 3.875211e-14, 9.161216e-06, 0, 0, 
    0, _, _, _, _, 0, 0, 1.009807e-05,
  0, 0, 0, 2.469519e-05, 0.0001265501, 5.047449e-12, 3.889873e-06, 
    1.776406e-06, 1.452312e-05, 5.671107e-06, 1.185252e-10, 3.29744e-06, 
    2.517591e-05, 6.185834e-06, 1.80336e-06,
  0, 0, 0, 1.595712e-05, 2.648094e-05, 0.0001275823, 0.0001063644, 
    1.152248e-05, 2.411881e-06, 2.56264e-05, 2.204983e-06, 1.944316e-06, 
    1.271706e-05, 1.625443e-06, 2.622737e-14,
  0, 0, 0, 1.627034e-05, 2.241401e-05, 5.954914e-06, 1.154209e-05, 
    9.033881e-05, 3.744446e-05, 5.248235e-06, 1.400921e-06, 4.814076e-06, 
    2.69315e-06, 5.110899e-06, 1.623482e-05,
  2.416706e-05, 1.807861e-13, 1.820069e-06, 6.955769e-06, 1.083747e-05, 
    3.971957e-06, 4.142009e-06, 1.051165e-06, 6.129151e-07, 4.971618e-06, 
    7.151188e-06, 1.373342e-05, 8.862067e-06, 7.233432e-06, 1.15617e-05,
  0, 1.966492e-06, 1.100307e-06, 9.062911e-06, 1.994331e-05, 9.492059e-06, 
    4.1654e-06, 3.130547e-06, 4.534026e-06, 3.528786e-05, 0, 0, 0, 
    9.068328e-06, 5.352906e-07,
  4.95234e-06, 5.422773e-06, 5.91315e-07, 1.313344e-13, 4.478924e-05, 
    4.226739e-06, 7.173333e-06, 7.078211e-06, 0, 0, 0, _, 0, 0, 5.319757e-06,
  2.216146e-06, 8.165292e-06, 1.691319e-05, 1.61398e-06, 2.609284e-05, 
    9.551698e-05, 2.932414e-06, 2.696491e-13, 0, _, _, _, 0, 0, 3.260584e-06,
  7.311861e-14, 4.030153e-06, 9.104476e-06, 1.992142e-05, 7.37191e-06, 
    2.585918e-06, 0.0001139984, 4.270704e-07, 0, _, _, _, 0, 0, 1.25411e-06,
  3.41487e-13, 3.296346e-06, 1.233126e-06, 1.15025e-05, 4.756208e-07, 
    8.743498e-06, 1.95482e-06, 0, 0, _, _, _, _, 0, 4.709427e-07,
  1.192725e-06, 8.085783e-06, 3.262958e-06, 3.561057e-14, 1.355505e-05, 0, 0, 
    0, _, _, _, _, 0, 0, 8.479298e-06,
  0, 0, 0, 2.530722e-05, 0.0002467867, 3.809845e-12, 3.42831e-06, 
    3.794699e-06, 2.145194e-05, 1.772236e-05, 1.493984e-05, 9.042692e-06, 
    5.582549e-05, 6.504817e-06, 1.336741e-06,
  0, 0, 0, 1.624273e-05, 2.240634e-05, 0.0002529389, 0.0002477323, 
    9.20139e-06, 9.74142e-05, 6.349033e-05, 8.757846e-06, 1.179519e-05, 
    2.63452e-05, 3.475661e-06, 2.410466e-14,
  0, 0, 0, 1.230895e-05, 1.31259e-05, 4.859496e-06, 7.121132e-06, 
    0.0002364442, 7.243914e-05, 6.663633e-06, 5.598437e-06, 8.460404e-06, 
    1.45889e-05, 1.748053e-05, 3.886102e-05,
  2.873782e-05, 1.665642e-13, 6.757332e-08, 6.738964e-06, 5.744504e-06, 
    3.767223e-06, 3.800084e-06, 3.754591e-05, 1.192044e-06, 6.883928e-06, 
    2.429012e-05, 1.358941e-05, 1.133194e-05, 1.275427e-05, 1.236946e-05,
  0, 1.283332e-06, 1.621147e-07, 6.18231e-07, 1.485739e-06, 2.09939e-06, 
    9.228208e-07, 3.0777e-06, 7.000092e-06, 7.945109e-05, 0, 0, 0, 
    2.129334e-05, 2.515845e-06,
  4.82622e-06, 2.512562e-06, 2.358814e-07, 1.209887e-13, 6.86375e-06, 
    3.270574e-07, 3.330241e-06, 2.383704e-06, 0, 0, 0, _, 0, 0, 1.227074e-05,
  4.418622e-07, 1.512934e-06, 3.774576e-06, 1.238319e-06, 6.273865e-06, 
    2.092246e-05, 2.718765e-06, 2.474507e-13, 0, _, _, _, 0, 0, 7.752937e-06,
  6.732555e-14, 1.999205e-06, 4.346489e-06, 3.792169e-06, 1.700166e-06, 
    2.032254e-06, 3.677629e-05, 1.531336e-07, 0, _, _, _, 0, 0, 9.510142e-07,
  3.121957e-13, 3.571673e-06, 7.011393e-07, 5.068442e-06, 5.392116e-07, 
    8.887409e-06, 1.338855e-06, 0, 0, _, _, _, _, 0, 7.815522e-07,
  1.125503e-06, 9.412715e-06, 3.802936e-06, 3.280207e-14, 9.977556e-06, 0, 0, 
    0, _, _, _, _, 0, 0, 8.555058e-06,
  0, 0, 0, 1.597202e-05, 0.0004923114, 2.918487e-12, 3.207608e-06, 
    2.620834e-06, 2.896043e-05, 2.345458e-05, 1.412375e-05, 2.621558e-06, 
    4.265316e-05, 3.383596e-06, 1.002066e-06,
  0, 0, 0, 6.050393e-06, 1.597305e-05, 0.0004784133, 0.0004576303, 
    8.255408e-06, 8.773633e-05, 0.0001016693, 2.365328e-06, 6.337083e-06, 
    2.449281e-05, 2.433265e-06, 2.214274e-14,
  0, 0, 0, 1.07776e-05, 1.105532e-05, 3.668146e-06, 4.752817e-06, 
    0.0004257713, 0.0001758556, 5.626966e-06, 4.60638e-06, 7.324556e-06, 
    1.407241e-05, 5.541348e-06, 2.758153e-05,
  2.985021e-05, 1.533585e-13, 1.398388e-08, 8.776417e-06, 4.953682e-06, 
    3.703187e-06, 4.164657e-06, 2.899519e-05, 9.630784e-05, 6.985602e-06, 
    0.0002077968, 4.970597e-05, 8.908123e-06, 1.052229e-05, 2.894634e-07,
  0, 1.077892e-06, 2.273871e-09, 1.672264e-07, 6.624736e-07, 1.045658e-06, 
    3.295653e-07, 3.681075e-06, 8.970464e-06, 5.528055e-05, 0, 0, 0, 
    1.045283e-05, 7.597749e-05,
  5.586034e-06, 1.769649e-06, 9.875017e-08, 1.113837e-13, 3.201482e-06, 
    9.726502e-08, 2.258181e-06, 5.639213e-07, 0, 0, 0, _, 0, 0, 7.336224e-05,
  2.321672e-07, 1.03069e-06, 2.584989e-06, 1.142112e-06, 4.395613e-06, 
    1.285694e-05, 2.532806e-06, 2.269458e-13, 0, _, _, _, 0, 0, 5.451975e-05,
  6.195829e-14, 1.706403e-06, 4.305748e-06, 2.454221e-06, 1.641676e-06, 
    1.977798e-06, 2.590583e-05, 9.930535e-08, 0, _, _, _, 0, 0, 3.851741e-07,
  6.305489e-08, 3.688714e-06, 6.720907e-07, 5.00535e-06, 5.879588e-07, 
    7.29588e-06, 8.741246e-07, 0, 0, _, _, _, _, 0, 1.132021e-08,
  1.087791e-06, 1.061871e-05, 3.235253e-06, 3.019501e-14, 1.939009e-05, 0, 0, 
    0, _, _, _, _, 0, 0, 4.936197e-06,
  0, 0, 0, 1.456141e-05, 0.0002125845, 2.285908e-12, 3.298163e-06, 
    1.608001e-06, 2.561212e-05, 1.342907e-05, 3.03966e-06, 1.570853e-06, 
    1.537551e-05, 3.02486e-06, 8.753526e-07,
  0, 0, 0, 4.443722e-06, 1.454833e-05, 0.0002032799, 0.0001873525, 
    7.557069e-06, 1.203632e-05, 6.998501e-05, 1.979749e-06, 1.64701e-06, 
    8.027583e-06, 1.876084e-06, 2.038998e-14,
  0, 0, 0, 1.271311e-05, 1.125184e-05, 2.169245e-06, 3.891844e-06, 
    0.0001657795, 0.0001112913, 8.735582e-06, 2.678495e-06, 4.445649e-06, 
    2.624171e-06, 2.513282e-06, 2.748091e-05,
  2.982943e-05, 1.41508e-13, 5.834118e-10, 1.107459e-05, 6.562623e-06, 
    3.456766e-06, 3.900226e-06, 9.124775e-06, 1.578567e-05, 7.403801e-06, 
    6.230763e-05, 5.301007e-05, 1.047997e-05, 8.001629e-06, 2.283517e-07,
  0, 8.497437e-07, 3.223965e-10, 3.68639e-09, 6.033258e-07, 9.707979e-07, 
    3.068943e-07, 3.438523e-06, 8.316944e-06, 2.99345e-05, 0, 0, 0, 
    5.597906e-06, 2.121392e-05,
  6.571906e-06, 1.833733e-06, 3.910399e-08, 1.027657e-13, 2.636456e-06, 
    3.447865e-08, 2.230832e-06, 5.843711e-07, 0, 0, 0, _, 0, 0, 0.000135058,
  4.87621e-09, 1.203379e-06, 2.929931e-06, 1.158544e-06, 5.558775e-06, 
    1.357719e-05, 2.550789e-06, 2.08639e-13, 0, _, _, _, 0, 0, 6.68921e-05,
  5.715179e-14, 2.031931e-06, 4.818882e-06, 3.289427e-06, 1.693514e-06, 
    2.140954e-06, 2.832077e-05, 1.037816e-07, 0, _, _, _, 0, 0, 3.47209e-07,
  1.568045e-07, 4.016868e-06, 7.586781e-07, 5.807705e-06, 1.130879e-06, 
    8.908451e-06, 3.267705e-06, 0, 0, _, _, _, _, 0, 2.641493e-08,
  1.041849e-06, 1.178055e-05, 4.119243e-06, 2.785613e-14, 3.597788e-05, 0, 0, 
    0, _, _, _, _, 0, 0, 2.832879e-06,
  0, 0, 0, 1.215472e-05, 0.000131053, 1.823014e-12, 2.963e-06, 5.715547e-07, 
    1.898331e-05, 2.589239e-06, 1.031151e-07, 1.023268e-06, 1.291275e-05, 
    1.849802e-06, 1.920828e-07,
  0, 0, 0, 1.310939e-06, 1.252349e-05, 0.0001270616, 0.0001174394, 
    5.384097e-06, 4.694662e-06, 3.697798e-05, 2.009297e-06, 1.782183e-06, 
    8.058259e-06, 9.640092e-07, 1.881731e-14,
  0, 0, 0, 1.359805e-05, 1.101685e-05, 7.241014e-07, 2.666778e-06, 
    0.0001055621, 6.803552e-05, 9.015917e-06, 2.809855e-06, 4.577811e-06, 
    2.631568e-06, 2.54253e-06, 1.174112e-05,
  2.942943e-05, 1.308314e-13, 1.244698e-10, 1.202786e-05, 7.472979e-06, 
    3.506899e-06, 4.179195e-06, 5.552299e-06, 1.473229e-05, 7.467484e-06, 
    3.171108e-05, 3.93888e-05, 1.152672e-05, 9.323944e-06, 1.802646e-07,
  0, 7.459383e-07, 1.016449e-10, 7.163954e-10, 5.455199e-07, 9.309438e-07, 
    3.149355e-07, 3.465374e-06, 8.037085e-06, 3.166602e-05, 0, 0, 0, 
    1.280075e-05, 1.191677e-05,
  7.160509e-06, 7.146838e-07, 2.13076e-09, 9.500245e-14, 1.55437e-06, 
    2.308477e-09, 2.177184e-06, 4.879891e-07, 0, 0, 0, _, 0, 0, 3.892368e-05,
  9.9606e-10, 1.067505e-07, 2.948983e-07, 9.296946e-07, 1.146591e-06, 
    7.740258e-06, 2.487982e-06, 1.922245e-13, 0, _, _, _, 0, 0, 2.9327e-05,
  5.282955e-14, 8.192392e-07, 3.461468e-06, 2.821192e-07, 1.562741e-06, 
    1.822467e-06, 1.913594e-05, 1.403351e-07, 0, _, _, _, 0, 0, 4.131388e-07,
  2.560411e-09, 3.823462e-06, 5.126258e-07, 3.940653e-06, 5.071109e-07, 
    5.565277e-06, 2.532408e-07, 0, 0, _, _, _, _, 0, 6.923848e-10,
  5.866406e-07, 1.220642e-05, 8.358329e-07, 2.574951e-14, 9.292492e-06, 0, 0, 
    0, _, _, _, _, 0, 0, 1.85388e-06,
  0, 0, 0, 1.050138e-05, 6.55296e-05, 1.477562e-12, 2.829403e-06, 
    4.106186e-08, 1.403129e-05, 3.743862e-08, 1.071865e-08, 8.646225e-07, 
    1.123883e-05, 1.70149e-07, 1.547322e-08,
  0, 0, 0, 4.149024e-08, 1.128738e-05, 6.481224e-05, 6.104948e-05, 
    4.157121e-06, 1.785198e-06, 2.371533e-05, 1.965328e-06, 1.882725e-06, 
    8.016225e-06, 2.719573e-08, 1.740375e-14,
  0, 0, 0, 1.371931e-05, 1.077471e-05, 7.590111e-08, 1.07451e-06, 
    5.687614e-05, 4.551368e-05, 8.383033e-06, 2.37438e-06, 4.984216e-06, 
    2.267934e-06, 2.350243e-06, 7.106023e-06,
  2.873413e-05, 1.21198e-13, 4.618796e-11, 1.198035e-05, 7.647859e-06, 
    3.549608e-06, 4.405866e-06, 1.037383e-06, 1.651728e-06, 6.987762e-06, 
    1.123097e-05, 3.000286e-05, 1.196183e-05, 8.633877e-06, 5.377062e-08,
  0, 1.418061e-07, 4.480787e-11, 2.564884e-10, 4.822971e-07, 8.717275e-07, 
    2.45031e-07, 3.355695e-06, 5.825153e-06, 2.395731e-05, 0, 0, 0, 
    2.263573e-06, 4.352844e-06,
  7.197377e-06, 1.2906e-08, 3.776569e-10, 8.799865e-14, 7.190619e-07, 
    4.283001e-10, 2.151987e-06, 2.675688e-07, 0, 0, 0, _, 0, 0, 1.40061e-05,
  3.634172e-10, 3.687699e-09, 1.297745e-08, 7.760116e-07, 3.506127e-08, 
    5.105825e-06, 2.475212e-06, 1.774816e-13, 0, _, _, _, 0, 0, 1.078562e-05,
  4.893629e-14, 3.123361e-08, 2.238295e-06, 2.821788e-08, 1.504192e-06, 
    1.773675e-06, 1.50239e-05, 1.33915e-07, 0, _, _, _, 0, 0, 6.992186e-09,
  5.299284e-10, 3.49953e-06, 3.803607e-07, 2.341059e-06, 7.644132e-08, 
    4.778447e-06, 7.369022e-09, 0, 0, _, _, _, _, 0, 1.375361e-10,
  3.59648e-07, 1.25481e-05, 4.118907e-08, 2.384918e-14, 3.489309e-06, 0, 0, 
    0, _, _, _, _, 0, 0, 9.967839e-07,
  0, 0, 0, 1.016807e-05, 4.804608e-05, 1.210149e-12, 3.008789e-06, 
    3.535104e-09, 1.216184e-05, 3.554737e-09, 3.040851e-09, 7.561335e-07, 
    1.108082e-05, 4.637785e-08, 2.054875e-09,
  0, 0, 0, 6.030077e-09, 1.094213e-05, 4.898386e-05, 4.634308e-05, 
    4.090261e-06, 9.522802e-07, 1.952012e-05, 1.936574e-06, 1.974317e-06, 
    8.318734e-06, 1.474079e-09, 1.610869e-14,
  0, 0, 0, 1.365097e-05, 1.061739e-05, 4.084761e-09, 1.320001e-06, 
    4.389382e-05, 3.704692e-05, 7.552902e-06, 1.965188e-06, 5.459471e-06, 
    2.211816e-06, 2.167808e-06, 3.642919e-06,
  2.766839e-05, 1.123405e-13, 2.177051e-11, 1.150707e-05, 7.492901e-06, 
    3.590807e-06, 4.589725e-06, 1.579207e-07, 3.750669e-07, 6.595167e-06, 
    6.843725e-06, 2.271285e-05, 1.186663e-05, 8.583018e-06, 1.690476e-08,
  0, 1.106564e-07, 2.336517e-11, 1.185273e-10, 4.783196e-07, 8.759491e-07, 
    1.867298e-07, 3.32235e-06, 5.099906e-06, 1.810371e-05, 0, 0, 0, 
    5.751747e-07, 2.773124e-06,
  7.232168e-06, 1.615571e-09, 1.270689e-10, 8.155981e-14, 7.05472e-07, 
    1.465892e-10, 2.201662e-06, 1.660126e-07, 0, 0, 0, _, 0, 0, 1.368243e-05,
  1.696941e-10, 6.295089e-10, 2.184172e-09, 7.587507e-07, 4.826971e-09, 
    5.006242e-06, 2.483406e-06, 1.639851e-13, 0, _, _, _, 0, 0, 7.621386e-06,
  4.53622e-14, 4.942963e-09, 1.893455e-06, 6.362152e-09, 1.517887e-06, 
    1.790667e-06, 1.338596e-05, 1.176538e-07, 0, _, _, _, 0, 0, 8.292628e-10,
  1.892666e-10, 3.279406e-06, 3.390257e-07, 1.755655e-06, 2.249683e-09, 
    3.639649e-06, 9.32473e-10, 0, 0, _, _, _, _, 0, 4.832699e-11,
  1.687489e-07, 1.265765e-05, 5.614039e-09, 2.210233e-14, 1.908988e-06, 0, 0, 
    0, _, _, _, _, 0, 0, 4.149943e-07,
  0, 0, 0, 1.051125e-05, 4.609124e-05, 1.006336e-12, 3.285797e-06, 
    9.767721e-10, 1.091327e-05, 1.022296e-09, 1.280637e-09, 9.225828e-07, 
    1.172503e-05, 5.252315e-09, 6.490134e-10,
  0, 0, 0, 1.959073e-09, 1.11567e-05, 4.729876e-05, 4.312547e-05, 
    4.585485e-06, 7.04567e-07, 1.763898e-05, 1.96271e-06, 2.060365e-06, 
    8.615473e-06, 3.744372e-10, 1.495719e-14,
  0, 0, 0, 1.355605e-05, 1.082428e-05, 9.573283e-10, 2.798125e-06, 
    3.97506e-05, 3.325868e-05, 7.12569e-06, 1.774969e-06, 5.782303e-06, 
    2.179944e-06, 2.165048e-06, 2.03229e-06,
  2.618785e-05, 1.044385e-13, 1.205728e-11, 1.082448e-05, 7.102233e-06, 
    3.621022e-06, 4.726998e-06, 9.413192e-08, 1.88184e-07, 6.11629e-06, 
    6.124032e-06, 1.944408e-05, 1.152201e-05, 8.408943e-06, 3.069388e-08,
  0, 5.131062e-07, 1.380564e-11, 6.484655e-11, 5.310446e-07, 9.15878e-07, 
    1.644899e-07, 3.307423e-06, 4.837897e-06, 1.68546e-05, 0, 0, 0, 
    8.991932e-08, 1.359352e-06,
  7.17812e-06, 5.012782e-10, 5.816442e-11, 7.581627e-14, 1.372235e-06, 
    6.769198e-11, 2.280847e-06, 1.690344e-07, 0, 0, 0, _, 0, 0, 1.144549e-05,
  9.343672e-11, 2.158421e-10, 7.452062e-10, 9.106094e-07, 1.541558e-09, 
    5.982934e-06, 2.502932e-06, 1.519944e-13, 0, _, _, _, 0, 0, 7.415434e-06,
  4.217817e-14, 1.6514e-09, 2.595842e-06, 2.423813e-09, 1.671035e-06, 
    1.952701e-06, 1.571438e-05, 1.065732e-07, 0, _, _, _, 0, 0, 2.532865e-10,
  8.937229e-11, 3.296012e-06, 4.654255e-07, 2.730795e-06, 4.085007e-10, 
    4.794161e-06, 2.902553e-10, 0, 0, _, _, _, _, 0, 2.262453e-11,
  1.451439e-07, 1.271688e-05, 1.787387e-09, 2.054429e-14, 2.689589e-06, 0, 0, 
    0, _, _, _, _, 0, 0, 2.763375e-07,
  0, 0, 0, 1.133617e-05, 5.365175e-05, 8.459721e-13, 3.683143e-06, 
    4.044824e-10, 1.093832e-05, 4.312223e-10, 6.593397e-10, 1.531587e-06, 
    1.472186e-05, 1.581382e-06, 2.863545e-10,
  0, 0, 0, 8.765831e-10, 1.130457e-05, 5.391549e-05, 4.610368e-05, 
    5.6323e-06, 6.758479e-07, 1.749306e-05, 2.028039e-06, 2.231285e-06, 
    9.462172e-06, 1.49351e-10, 1.391386e-14,
  0, 0, 0, 1.362992e-05, 1.065886e-05, 3.690032e-10, 4.755944e-06, 
    4.008669e-05, 3.205901e-05, 6.813653e-06, 1.704537e-06, 5.962093e-06, 
    2.612461e-06, 2.557312e-06, 3.883818e-06,
  2.427505e-05, 9.725666e-14, 7.382529e-12, 1.018316e-05, 6.641294e-06, 
    3.643482e-06, 4.82293e-06, 3.351509e-07, 3.930793e-07, 6.179921e-06, 
    8.891666e-06, 1.761918e-05, 1.126628e-05, 9.725782e-06, 2.771912e-07,
  0, 1.453816e-06, 8.844626e-12, 3.937421e-11, 6.464231e-07, 1.014727e-06, 
    1.550616e-07, 3.348276e-06, 5.603927e-06, 2.145925e-05, 0, 0, 0, 
    2.380417e-07, 2.180579e-06,
  7.063832e-06, 3.259301e-08, 3.147438e-11, 7.059677e-14, 2.928008e-06, 
    3.682816e-11, 2.410238e-06, 3.604397e-07, 0, 0, 0, _, 0, 0, 2.378501e-05,
  5.698244e-11, 9.926292e-11, 3.418383e-10, 1.212107e-06, 1.595937e-06, 
    9.619424e-06, 2.543874e-06, 1.411394e-13, 0, _, _, _, 0, 0, 7.903647e-06,
  3.9288e-14, 9.949031e-07, 4.092982e-06, 1.179076e-09, 1.926458e-06, 
    2.245591e-06, 2.158604e-05, 1.019501e-07, 0, _, _, _, 0, 0, 1.099413e-10,
  4.930044e-11, 3.496341e-06, 6.613257e-07, 4.653661e-06, 1.426597e-10, 
    6.936278e-06, 1.271529e-10, 0, 0, _, _, _, _, 0, 1.241371e-11,
  2.829687e-07, 1.282355e-05, 7.917464e-10, 1.912854e-14, 4.470804e-06, 0, 0, 
    0, _, _, _, _, 0, 0, 5.01185e-07,
  0, 0, 0, 1.209215e-05, 7.54293e-05, 7.177593e-13, 4.28046e-06, 
    2.048414e-10, 1.153422e-05, 7.264463e-06, 3.827579e-10, 2.048302e-06, 
    1.698441e-05, 3.025872e-06, 2.587257e-07,
  0, 0, 0, 4.651101e-10, 1.145543e-05, 7.396544e-05, 6.104653e-05, 
    7.30978e-06, 7.848943e-07, 2.549628e-05, 2.144206e-06, 2.417432e-06, 
    9.944202e-06, 7.400232e-11, 1.29653e-14,
  0, 0, 0, 1.302535e-05, 1.04525e-05, 6.656624e-08, 6.793987e-06, 
    5.031624e-05, 4.039057e-05, 7.85817e-06, 2.025e-06, 6.137674e-06, 
    2.892535e-06, 2.64289e-06, 1.03077e-05,
  2.198506e-05, 9.070845e-14, 4.840183e-12, 9.327948e-06, 5.995136e-06, 
    3.813605e-06, 4.869382e-06, 6.097426e-07, 7.556462e-07, 6.368959e-06, 
    2.399294e-05, 1.972987e-05, 1.130807e-05, 9.871059e-06, 2.586128e-07,
  0, 1.598352e-06, 5.998636e-12, 2.565632e-11, 6.921812e-07, 1.040688e-06, 
    3.249311e-07, 3.484632e-06, 6.103945e-06, 4.111583e-05, 0, 0, 0, 
    6.57622e-07, 4.787226e-06,
  6.908341e-06, 3.113743e-06, 1.889746e-11, 6.583827e-14, 3.437733e-06, 
    2.219411e-11, 2.474531e-06, 5.681553e-07, 0, 0, 0, _, 0, 0, 1.999588e-05,
  3.724946e-11, 5.357158e-11, 1.841947e-10, 1.299941e-06, 2.722233e-06, 
    1.206745e-05, 2.578392e-06, 1.312788e-13, 0, _, _, _, 0, 0, 1.016345e-05,
  3.665579e-14, 2.116194e-06, 4.476638e-06, 6.594552e-10, 2.026996e-06, 
    2.402793e-06, 2.623575e-05, 9.792737e-08, 0, _, _, _, 0, 0, 5.726312e-11,
  2.999592e-11, 3.545432e-06, 8.173083e-07, 5.426528e-06, 3.71835e-10, 
    8.319728e-06, 6.659839e-11, 0, 0, _, _, _, _, 0, 7.52489e-12,
  6.31607e-07, 1.267634e-05, 2.530268e-06, 1.783796e-14, 5.409904e-06, 0, 0, 
    0, _, _, _, _, 0, 0, 8.846003e-07,
  0, 0, 0, 1.182119e-05, 8.164552e-05, 6.142635e-13, 3.985951e-06, 
    7.021062e-08, 1.146855e-05, 9.710265e-06, 2.421595e-10, 2.181679e-06, 
    2.209594e-05, 3.308595e-06, 7.612904e-07,
  0, 0, 0, 1.501481e-06, 1.129962e-05, 8.014546e-05, 6.689409e-05, 
    6.694149e-06, 1.722168e-06, 3.017095e-05, 3.29304e-06, 2.908689e-06, 
    1.346346e-05, 4.208429e-11, 1.210182e-14,
  0, 0, 0, 1.265062e-05, 1.028609e-05, 1.509824e-07, 7.44718e-06, 
    5.752066e-05, 4.47979e-05, 6.497828e-06, 2.002406e-06, 6.361643e-06, 
    5.216769e-06, 3.014809e-06, 1.382527e-05,
  1.959407e-05, 8.473158e-14, 3.347832e-12, 8.545213e-06, 5.683377e-06, 
    4.665731e-06, 5.299593e-06, 1.085316e-06, 9.094354e-07, 6.059189e-06, 
    2.530149e-05, 2.329881e-05, 1.108017e-05, 1.287637e-05, 2.662066e-07,
  0, 1.652841e-06, 4.258597e-12, 1.766306e-11, 1.180866e-06, 1.203354e-06, 
    2.469684e-07, 3.425804e-06, 6.184569e-06, 5.899867e-05, 0, 0, 0, 
    1.595345e-05, 1.024484e-05,
  6.689801e-06, 3.280036e-06, 4.753984e-08, 6.149543e-14, 4.543975e-06, 
    1.442157e-11, 2.527114e-06, 4.681212e-07, 0, 0, 0, _, 0, 0, 1.233214e-05,
  2.570698e-11, 3.03149e-06, 2.547617e-06, 1.336447e-06, 2.89121e-06, 
    1.348458e-05, 2.887417e-06, 1.223108e-13, 0, _, _, _, 0, 0, 7.563299e-06,
  3.425571e-14, 2.336902e-06, 4.623937e-06, 2.299132e-07, 2.082628e-06, 
    2.347119e-06, 2.75257e-05, 2.453985e-07, 0, _, _, _, 0, 0, 5.353003e-11,
  1.962662e-11, 3.435223e-06, 7.138174e-07, 5.470481e-06, 2.934681e-07, 
    7.578291e-06, 3.927026e-11, 0, 0, _, _, _, _, 0, 6.122107e-08,
  9.241619e-07, 1.21739e-05, 2.909834e-06, 1.666022e-14, 5.890007e-06, 0, 0, 
    0, _, _, _, _, 0, 0, 1.374491e-06 ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319, 349.5 ;
}
