netcdf atmos_daily.00010101-00010701.ps.tile4 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float ps(time, grid_yt, grid_xt) ;
		ps:_FillValue = 1.e+20f ;
		ps:missing_value = 1.e+20f ;
		ps:units = "Pa" ;
		ps:long_name = "Surface Air Pressure" ;
		ps:cell_methods = "time: mean" ;
		ps:cell_measures = "area: area" ;
		ps:time_avg_info = "average_T1,average_T2,average_DT" ;
		ps:standard_name = "surface_air_pressure" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:03 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile4.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile4.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.2466774, 0.6143242, 0.0668168, 0.2301621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.4924844, 0.2132108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.600569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1560082, 0,
  1, 1, 0.7132517, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02739768, 0,
  0.6230268, 0.6280472, 0.3043983, 0.08344039, 0, 0.3148882, 0.01188002, 0, 
    0, 0, 0, 0.08803581, 0, 0, 0,
  0, 0, 0, 0, 0.01144353, 0.8597386, 0.8205094, 0.5086318, 0.1258651, 
    0.08909279, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.291879, 0.6933324, 1, 0.9996726, 0.6666086, 0.08008575, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.611689, 0.7180831, 0.4623523, 0.2838529, 0.02767258, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0.002817577, 0.8915156, 0.5654301, 0.7485356, 0.3018697, 0, 0, 0, 
    0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 ps =
  102040.9, 102033, 102070.3, 102103, 102157.2, 102227.1, 102279.2, 102321.1, 
    102339.2, 102348.9, 102336.7, 102310.7, 102263.1, 102194.1, 102104.8,
  101909.8, 101904.1, 101952.2, 102005.8, 102035.1, 102099.1, 102153.7, 
    102206.6, 102230.3, 102249.6, 102237.7, 102226.2, 102180.7, 102148.8, 
    102109,
  100148.4, 99891.34, 101856.5, 101984.6, 101971.9, 102014.4, 102047.6, 
    102096.5, 102127.6, 102153.7, 102157.3, 102155.2, 102135.7, 102098.8, 
    102064.9,
  98058.39, 98129.23, 101752.6, 101926.3, 101913.3, 101945.2, 101979.8, 
    102017.2, 102044.5, 102064.2, 102069, 102075.8, 102060.8, 102043, 102041.7,
  98015.91, 98481.62, 100414.6, 101911.1, 101897, 101869, 101914.3, 101944.2, 
    101963, 101989.8, 102004.4, 102018.2, 102000.8, 102010.7, 102013.9,
  97303.56, 98836.88, 101746.2, 101873.2, 101842.9, 101809.2, 101875.1, 
    101909.7, 101923.8, 101944.9, 101927.8, 101917.9, 101967.3, 101980.7, 
    101988.3,
  101737.4, 101762.3, 101833.2, 101853.2, 101807.1, 99985.77, 101533.9, 
    101662.5, 101808.6, 101883.5, 101927.7, 101942.8, 101941.6, 101960.2, 
    101965.3,
  101690.5, 101694.6, 101754.1, 101736.1, 101620.5, 99108.17, 97226.83, 
    96407.77, 99035.68, 101849.5, 101910.3, 101923.2, 101927.8, 101938.3, 
    101943.6,
  101623.2, 101635.1, 101693.1, 101678.4, 96753.35, 98250.14, 99972.99, 
    101553.2, 101775.8, 101847.8, 101881.8, 101892.2, 101902.3, 101919.3, 
    101930.2,
  101743.2, 101634.1, 101645.6, 101598.8, 97255.15, 97520.95, 97035.55, 
    101687.4, 101889.6, 101819.5, 101859.8, 101868.5, 101893.4, 101901.2, 
    101914.2,
  101881.5, 101856.2, 101878.1, 101886.2, 101918.8, 101982.4, 102041.9, 
    102105, 102156.8, 102203.6, 102221.7, 102226.1, 102212.4, 102177.6, 
    102112.2,
  101698.5, 101703.8, 101765.6, 101782.3, 101788, 101818.6, 101878.6, 
    101946.9, 101999.1, 102047.9, 102076.1, 102090.2, 102086.6, 102073.9, 
    102059.5,
  99817.55, 99599.69, 101613.7, 101756.1, 101720.8, 101728.1, 101740.8, 
    101796.5, 101855.8, 101911.9, 101959.3, 101980.6, 101992.6, 101975.9, 
    101957.9,
  97706.83, 97803.58, 101464.8, 101679.3, 101635, 101638.5, 101639.3, 
    101664.6, 101706, 101761.7, 101807.2, 101849.5, 101859.7, 101865, 101872.5,
  97578.34, 98104.56, 100050.6, 101620.3, 101595.4, 101540.5, 101542.6, 
    101560, 101586.4, 101639.8, 101691.9, 101741.2, 101747.6, 101784.8, 
    101795.7,
  96847.7, 98412.94, 101311.3, 101507.4, 101495.9, 101457.8, 101502.9, 
    101512.6, 101516.2, 101554.3, 101569.4, 101587.8, 101659.5, 101690.7, 
    101708.1,
  101173.3, 101255.1, 101359.5, 101426.4, 101403, 99602.24, 101105.6, 
    101216.3, 101329.1, 101417.1, 101479.2, 101535.3, 101575.9, 101605.2, 
    101627,
  101074.3, 101042.7, 101122.2, 101212.3, 101128.8, 98656.71, 96800.1, 
    95955.75, 98515.24, 101348, 101393.5, 101430.1, 101477.2, 101513.2, 
    101545.7,
  101044.9, 100987.1, 100987.6, 101051.8, 96193.46, 97693.62, 99406.49, 
    101009.2, 101245.8, 101304.7, 101308.1, 101337.1, 101385.2, 101428, 
    101457.7,
  101092.3, 100936.4, 100947.4, 100906.2, 96600.02, 96912.02, 96452.68, 
    101090.5, 101302.1, 101199.6, 101231, 101249.4, 101294.6, 101341.9, 
    101387.3,
  101837.1, 101862.7, 101936.3, 101999.3, 102082.9, 102165.8, 102243.7, 
    102314.2, 102355, 102391.1, 102400, 102396.4, 102385.9, 102359.8, 102307.2,
  101655.6, 101696.7, 101790.5, 101871, 101940, 102027.2, 102105.1, 102180.5, 
    102233.8, 102274.6, 102301.6, 102307.9, 102295.1, 102282.6, 102269.5,
  99855.77, 99652.52, 101651.3, 101834.6, 101851.4, 101915.1, 101974, 
    102048.7, 102113.5, 102163.8, 102198.3, 102217.1, 102224.2, 102209.3, 
    102193.1,
  97765.21, 97886.25, 101533.9, 101736.7, 101748.4, 101812.9, 101867, 
    101929.3, 101984.2, 102042.3, 102082.9, 102113.9, 102123.8, 102119.6, 
    102132.5,
  97766.01, 98249.65, 100212, 101727.2, 101713, 101712.9, 101761.8, 101816.3, 
    101861.2, 101917.8, 101972.9, 102018.5, 102020.4, 102054.1, 102064.5,
  96983.62, 98588.28, 101551.6, 101706.9, 101654.1, 101643.8, 101714, 
    101752.8, 101792.3, 101833.8, 101852.3, 101870.4, 101945.3, 101972.5, 
    101988.8,
  101439.8, 101532.6, 101607.3, 101682.3, 101609.9, 99819.76, 101349.4, 
    101463.5, 101584.1, 101688.8, 101768.6, 101821.8, 101870.3, 101894.6, 
    101916.3,
  101360.4, 101382.5, 101453.1, 101510.6, 101378.9, 98893.18, 97043.99, 
    96209.77, 98798.68, 101629, 101681.9, 101725.7, 101777.2, 101815.6, 
    101840.6,
  101159.3, 101203.6, 101293.7, 101384.6, 96456.08, 97978, 99710.35, 
    101325.7, 101552.8, 101601.4, 101603.7, 101644.2, 101690.5, 101735.3, 
    101762.9,
  101154.3, 101141.8, 101125.5, 101169, 96832.36, 97207.52, 96756.88, 
    101441.1, 101636.8, 101539.6, 101550.2, 101567.5, 101611.1, 101653.3, 
    101689.1,
  102056.1, 102087.4, 102123.4, 102169.3, 102227, 102294.9, 102355.1, 
    102416.6, 102459.9, 102501.1, 102515.9, 102527.4, 102519.6, 102488.4, 
    102428.6,
  101893.9, 101944, 102048.2, 102109.6, 102141, 102218.3, 102292.7, 102356.9, 
    102400.8, 102442.9, 102467.2, 102478, 102473.4, 102462.5, 102442.8,
  100024.9, 99867.77, 101896.7, 102087.8, 102093.8, 102150.4, 102208.9, 
    102284.6, 102345.7, 102398.2, 102435.4, 102452.5, 102449.5, 102428.2, 
    102405.2,
  97930.85, 98107.16, 101775, 102021.7, 102028.7, 102094.9, 102155.2, 
    102225.2, 102286.3, 102338.6, 102376.5, 102403.2, 102400.2, 102384.9, 
    102387.1,
  97941.06, 98463.34, 100413.2, 101972.4, 101984.8, 102000.8, 102075.8, 
    102141.2, 102205.9, 102276.2, 102325.7, 102365.7, 102357.4, 102372.6, 
    102363.6,
  97282.22, 98856.1, 101812.8, 101929.9, 101925, 101943.9, 102040.5, 
    102115.5, 102163.1, 102219.9, 102250.1, 102265.2, 102326.4, 102339.5, 
    102334,
  101763.5, 101848.3, 101939.5, 101941.9, 101884.1, 100104.9, 101666.5, 
    101815.5, 101994.3, 102120.6, 102205.4, 102259, 102291.5, 102305.3, 
    102305.2,
  101814, 101809.5, 101865.8, 101845.6, 101716, 99230.52, 97392.27, 96594.94, 
    99211.65, 102072.9, 102139.2, 102192, 102234.8, 102260.9, 102272.6,
  101615.4, 101652.5, 101790, 101793.6, 96792.03, 98337.08, 100081.2, 
    101684.5, 101948.8, 102048.8, 102086, 102132.3, 102178.8, 102211, 102232.1,
  101510.4, 101564, 101694.3, 101695.8, 97303.91, 97598.6, 97150.32, 
    101866.1, 102069.8, 101992.9, 102040.5, 102074.3, 102125.8, 102159.1, 
    102186.8,
  101518.1, 101595.4, 101709.8, 101803.5, 101897.1, 101977.2, 102050.1, 
    102113, 102162.1, 102213.4, 102257.8, 102292.5, 102309.6, 102298.9, 
    102257.2,
  101449, 101519.4, 101675.4, 101786.7, 101874.9, 101970.1, 102048, 102112.2, 
    102156.7, 102200.4, 102238, 102275, 102293.1, 102292.6, 102270,
  99675.08, 99531.15, 101576.3, 101799.6, 101854.5, 101943.4, 102018.2, 
    102085.3, 102135.2, 102186, 102229, 102271.5, 102295.5, 102289.4, 102276.9,
  97630.55, 97850.12, 101490.7, 101779.8, 101840.9, 101944.3, 102022.2, 
    102093.5, 102139.8, 102180.5, 102218.3, 102253.4, 102271.9, 102265.6, 
    102274.5,
  97658.48, 98223.18, 100199, 101768.9, 101840, 101893.6, 101980.2, 102052.8, 
    102107, 102160.9, 102206.1, 102251.3, 102264.8, 102284.9, 102276.8,
  97080.38, 98672.22, 101585.6, 101747.5, 101828.4, 101863.8, 101984.3, 
    102062.5, 102115.6, 102157.6, 102175.9, 102185.9, 102260.8, 102286, 
    102280.4,
  101523.1, 101638.5, 101751, 101790.7, 101830.3, 100123.5, 101646.9, 
    101798.9, 101985.3, 102098.7, 102175.3, 102223.4, 102257.5, 102284.6, 
    102277.7,
  101693.9, 101704.2, 101744.5, 101764.2, 101714.6, 99285.97, 97455.69, 
    96663.6, 99262.65, 102081.2, 102153.4, 102202.8, 102242.7, 102273.1, 
    102271.8,
  101616.7, 101650, 101766.6, 101774.1, 96954.73, 98483.05, 100181.9, 
    101774.2, 102002.2, 102094.1, 102136.3, 102182.5, 102229.7, 102256.4, 
    102262.1,
  101671.8, 101698.6, 101786, 101776.5, 97450.71, 97774.23, 97316.99, 
    101981.8, 102133.5, 102081.2, 102127.1, 102166.6, 102212.4, 102238.9, 
    102251.1,
  101781.3, 101809.5, 101866, 101883.5, 101914.7, 101932.5, 101946.8, 
    101964.3, 101976.2, 101996, 102030.7, 102067.2, 102095.7, 102118.1, 
    102083.5,
  101605.4, 101659.6, 101778.1, 101833.6, 101859.4, 101901.9, 101929.7, 
    101955, 101971.2, 101988.7, 102025.5, 102064.8, 102094.2, 102117.4, 
    102117.4,
  99716.98, 99573.63, 101603.7, 101794.3, 101806.8, 101855, 101884.5, 
    101927.6, 101956.9, 101979, 102019, 102065, 102106.6, 102126.1, 102130.5,
  97543.16, 97771.76, 101430.3, 101719.2, 101756, 101826.4, 101866.7, 
    101909.5, 101947.8, 101975.9, 102014.5, 102059, 102101.5, 102116.9, 
    102139.1,
  97438.09, 98044.46, 100069, 101644.1, 101703.6, 101743.1, 101824, 101874, 
    101915.3, 101959.3, 102008.1, 102055.9, 102094.5, 102139.1, 102150.6,
  96733.72, 98368.35, 101339.5, 101567.7, 101636.1, 101672.9, 101790.2, 
    101862, 101913.6, 101957.2, 101989.5, 102002.7, 102092.2, 102147.2, 
    102158.4,
  101090.4, 101308.7, 101481.4, 101542.1, 101572.5, 99885.92, 101444, 
    101607.9, 101791.5, 101897, 101990.1, 102045.6, 102093.9, 102148.4, 
    102168.5,
  101225, 101278.7, 101391.5, 101429.8, 101389.8, 98993.17, 97228.53, 
    96467.04, 99067.41, 101871.7, 101966.2, 102033.3, 102088.1, 102145.1, 
    102172.5,
  101051.8, 101160.3, 101349.4, 101373.5, 96619.84, 98147.13, 99849.22, 
    101450.9, 101747.4, 101869.3, 101944.9, 102020.2, 102084.2, 102139.1, 
    102176.6,
  101012.4, 101124.5, 101289.5, 101296.4, 97065.4, 97413.23, 97030.59, 
    101623.5, 101853.3, 101852.2, 101934.2, 102008.4, 102080.5, 102133.4, 
    102175.4,
  102042.4, 101997.2, 101963.7, 101923.7, 101886.3, 101879.7, 101891.5, 
    101914.3, 101923.4, 101940.9, 101961, 101970.1, 101970.1, 101952.6, 
    101922.8,
  101924.4, 101920.7, 101963, 101917.3, 101874.6, 101868.2, 101883.1, 
    101909.9, 101925.7, 101937.6, 101953.2, 101970.7, 101984.7, 101982.2, 
    101967.5,
  100091.2, 99870.34, 101842.3, 101946.1, 101859.9, 101845, 101850.6, 
    101882.1, 101912.4, 101932.2, 101961.9, 101988.9, 102001.5, 102003.6, 
    101986,
  97984.07, 98123.57, 101745.5, 101933.6, 101862.8, 101855.7, 101855.6, 
    101884.8, 101917.8, 101938.5, 101964.8, 101996.2, 102019.4, 102012.6, 
    102017.4,
  97977.65, 98484.23, 100428.2, 101921, 101861.5, 101806.5, 101829.2, 
    101860.8, 101898.8, 101938, 101966.8, 102003.6, 102022.8, 102041.5, 
    102046.1,
  97325.98, 98870.32, 101788, 101891.3, 101846.1, 101774.9, 101828.6, 
    101867.8, 101914.7, 101949.1, 101963.8, 101964.2, 102043, 102072, 102073.5,
  101826.5, 101898.8, 101966, 101923.2, 101838.1, 100016, 101496.7, 101626.4, 
    101804.1, 101905.4, 101976.5, 102017.3, 102052.9, 102087.9, 102091,
  101897, 101868.9, 101911.7, 101850.5, 101668.1, 99145.86, 97313.3, 96531.2, 
    99121.36, 101907.6, 101975.2, 102019.5, 102060.4, 102098.8, 102107.8,
  101804.2, 101818, 101918.9, 101838.4, 96895.9, 98325.63, 99972.66, 
    101526.5, 101816.1, 101929.7, 101970.5, 102017.1, 102064.3, 102100, 
    102117.5,
  101811.4, 101812.8, 101888.3, 101785.7, 97367.27, 97606.63, 97148.59, 
    101728.1, 101952.3, 101927, 101976.8, 102017.8, 102065.8, 102102.1, 
    102124.4,
  102726.5, 102679.4, 102626.8, 102563.6, 102486.5, 102406.6, 102303.6, 
    102199.4, 102101.3, 102015.8, 101937.9, 101886.3, 101871.2, 101850.9, 
    101816.9,
  102667.1, 102624.5, 102645.2, 102594.7, 102515.6, 102455.1, 102369.3, 
    102288.1, 102188.2, 102099.7, 102022.9, 101971.6, 101946.9, 101923.2, 
    101896,
  100834.7, 100564.5, 102575, 102618.3, 102540.3, 102487.2, 102401.8, 
    102329.2, 102240.1, 102162.9, 102094.8, 102032.6, 102009.3, 101978.9, 
    101943.7,
  98768.97, 98835.29, 102458.1, 102636.4, 102550.9, 102527, 102452.5, 
    102389.4, 102300.9, 102227.7, 102155.3, 102092.8, 102067.7, 102024.7, 
    102008.3,
  98737.22, 99217.71, 101138.3, 102646.6, 102561.9, 102506.4, 102451.3, 
    102390.6, 102324, 102263.8, 102199.9, 102147.5, 102105.8, 102085.4, 
    102059.2,
  98070.97, 99622.64, 102503.8, 102626.9, 102547.7, 102497.7, 102503.9, 
    102438.9, 102360.1, 102297.9, 102221, 102138.2, 102154.3, 102145.7, 
    102110.7,
  102517.6, 102602.9, 102656.2, 102639.7, 102554.2, 100689.1, 102158.3, 
    102198.4, 102266, 102270.9, 102251.7, 102212.1, 102195.2, 102180.3, 
    102154.5,
  102602.2, 102569.8, 102580.7, 102522.4, 102382.9, 99846.52, 97926.1, 
    97028.27, 99564.57, 102275.1, 102264.4, 102231.4, 102223.4, 102214.1, 
    102195.1,
  102453.2, 102445.5, 102548.5, 102498.7, 97549.74, 98970.83, 100648.4, 
    102167.3, 102322.2, 102303.8, 102279, 102248.2, 102244.3, 102241.6, 
    102223.4,
  102437.5, 102398.3, 102512.2, 102418.3, 98031.02, 98257.98, 97739.75, 
    102278.7, 102437, 102310.7, 102301, 102259.2, 102262.7, 102262.7, 102249.4,
  102653, 102476.8, 102267.6, 101970.8, 101742.1, 101514, 101334.3, 101230.6, 
    101144.6, 101081.2, 101009.5, 101016.1, 101068.1, 101100.7, 101104.9,
  102702.5, 102480.4, 102396.3, 102136.1, 101925.1, 101720.6, 101551.5, 
    101397.7, 101280.1, 101189.4, 101117.9, 101113.1, 101106.3, 101138.7, 
    101173.4,
  100901.2, 100484.9, 102419.8, 102259.7, 102058.3, 101858.6, 101705.9, 
    101572, 101452.9, 101335.2, 101237.9, 101196.4, 101196.1, 101211.9, 
    101234.3,
  98925.09, 98948.03, 102396.1, 102405.6, 102214.1, 102044, 101893.6, 
    101767.3, 101641.5, 101508.4, 101388.2, 101306.3, 101296.1, 101281.3, 
    101311.8,
  98972.02, 99390.29, 101172.6, 102537.9, 102342.4, 102164.6, 102016.1, 
    101894.8, 101783.6, 101667.8, 101530.3, 101436.9, 101372.2, 101377.1, 
    101376.9,
  98423.66, 99903.94, 102653, 102620.9, 102460.1, 102243.9, 102178.8, 
    102039.3, 101931.8, 101788.2, 101651.1, 101517.3, 101495.5, 101496.7, 
    101482.2,
  102980, 102944.8, 102850.6, 102738.5, 102557.8, 100594.8, 101953.3, 101890, 
    101937.2, 101869.1, 101795.1, 101707.5, 101643.5, 101614.3, 101594,
  103099.4, 102993, 102911.4, 102764.4, 102452.8, 99852.77, 97838.03, 
    96926.05, 99429.46, 102032.5, 101925.3, 101849.6, 101786.1, 101750.5, 
    101716.9,
  103072, 102976.2, 102962.5, 102818.1, 97736.25, 99173.84, 100761, 102260.3, 
    102251.4, 102152.6, 102054.8, 101963.7, 101907.6, 101861.9, 101832,
  103101.9, 103011.9, 103013.4, 102850.9, 98364.06, 98533.41, 97866.56, 
    102409.8, 102412.1, 102258.8, 102165.1, 102062.6, 102009, 101957.8, 
    101922.5,
  101116.5, 100711.9, 100354.8, 100265.9, 100335.3, 100455.3, 100569.3, 
    100660.7, 100751, 100841.8, 100910.5, 100941.6, 100960.2, 100964, 100955,
  101175.9, 100758.9, 100494.4, 100335, 100313.8, 100388.8, 100493.1, 100597, 
    100689.5, 100756.8, 100800.5, 100833.1, 100852.8, 100876.2, 100905.5,
  99369.35, 98852.29, 100531.5, 100436.8, 100372.1, 100421.9, 100475.8, 
    100543.5, 100605.6, 100661.6, 100718.4, 100757.6, 100782.8, 100789.6, 
    100791.6,
  97589.66, 97543.7, 100621.4, 100639.7, 100530.3, 100517, 100551.1, 100589, 
    100613.1, 100647.8, 100664.4, 100693.8, 100720.6, 100699.8, 100721,
  97817.23, 98024.59, 99553.23, 100827.6, 100700.6, 100619.1, 100600, 
    100597.9, 100604.4, 100630.8, 100659, 100715.4, 100716.4, 100694.5, 
    100692.4,
  97627.4, 98784, 101181.4, 101030.5, 100870.1, 100673.1, 100708, 100709.2, 
    100727.4, 100721.1, 100706.9, 100686.9, 100730.7, 100713.7, 100698.6,
  102144.9, 101794.1, 101460.4, 101224.7, 100958.9, 99111.77, 100491.8, 
    100556.1, 100702.4, 100746.1, 100784.4, 100791.4, 100785.6, 100770.3, 
    100741.2,
  102296.1, 101963, 101693.2, 101396.3, 100901.4, 98425.45, 96570.7, 95757.1, 
    98276.24, 100883.4, 100876.8, 100878.1, 100851.6, 100827.1, 100805.5,
  102420.9, 102106.1, 101931.1, 101514.6, 96565.16, 97993.76, 99512.9, 
    101015.7, 101053.5, 101040.4, 101013.7, 100980.5, 100946.1, 100916, 
    100885.9,
  102637.1, 102336.9, 102170.1, 101771.3, 97360.33, 97438.41, 96842.9, 
    101311.8, 101317.2, 101232.4, 101155.5, 101101.5, 101058.8, 101024.6, 
    100993.7,
  100714.2, 100651, 100617.7, 100654.9, 100758.3, 100896, 101037.1, 101155.2, 
    101268.4, 101368.3, 101430.1, 101476.4, 101492.6, 101501, 101481.9,
  100467.3, 100371.7, 100418.2, 100419.4, 100479.6, 100613.1, 100781.8, 
    100946, 101078.3, 101178.1, 101268.3, 101344.9, 101389.8, 101422, 101443.5,
  98479.36, 98135.26, 100084, 100213.7, 100254.9, 100366.1, 100521.4, 
    100705.4, 100867.5, 101008, 101120.1, 101211.9, 101278.9, 101322.8, 
    101354.3,
  96369.56, 96398.05, 99775.66, 100033, 100073.1, 100169.8, 100313.1, 
    100497.6, 100676.9, 100839.1, 100969.8, 101080.9, 101163.6, 101219.4, 
    101287,
  96140.14, 96540.56, 98326.32, 99841.58, 99914.94, 99993.66, 100147.9, 
    100320.4, 100496.7, 100672.5, 100823, 100951.7, 101038.6, 101128.9, 101199,
  95418.87, 96786.17, 99511.98, 99682.32, 99781, 99824.02, 100014.6, 
    100183.5, 100365.2, 100539.5, 100683.4, 100783.5, 100938.5, 101037.4, 
    101116.3,
  99537.61, 99474.05, 99516.3, 99584.82, 99671.2, 98050.76, 99633.78, 
    99871.14, 100160.6, 100378.9, 100581.8, 100721.8, 100841.2, 100944.8, 
    101035.6,
  99387.92, 99410.93, 99439.2, 99517.41, 99439.35, 97135.55, 95435.17, 
    94766.48, 97410.12, 100260.5, 100477.2, 100626.7, 100756.6, 100862.1, 
    100961,
  99403.42, 99430.45, 99478.95, 99426.2, 94825.02, 96338.76, 97978.61, 
    99578.84, 99933.32, 100197.8, 100384.3, 100541.1, 100673.5, 100785.1, 
    100885.4,
  99654.49, 99572.99, 99626.82, 99490.62, 95365.83, 95632.64, 95229.04, 
    99741.09, 100030.9, 100149, 100322.2, 100472, 100611.8, 100720.6, 100823.7,
  100681.8, 100776.9, 100936.4, 101062.3, 101191.3, 101307.7, 101402.5, 
    101481.6, 101539.4, 101585.5, 101613, 101622.6, 101623.3, 101609.8, 
    101559.9,
  100378.3, 100471.3, 100692.7, 100862.4, 100987.5, 101140.2, 101260.8, 
    101356.5, 101429.8, 101485.4, 101524.1, 101552.2, 101562.5, 101561.1, 
    101572.2,
  98335, 98254.46, 100343.1, 100663.1, 100780.7, 100932.6, 101064.7, 
    101196.7, 101297.6, 101376.1, 101432.2, 101473.9, 101499.9, 101509.6, 
    101509.5,
  96119.98, 96363.45, 100006.5, 100443.2, 100588.6, 100768.7, 100922.4, 
    101058.1, 101170.5, 101266.5, 101337.8, 101396, 101430.5, 101447, 101478.5,
  95968.34, 96575.18, 98565.86, 100246.7, 100410.9, 100556.1, 100733.2, 
    100891.9, 101018.7, 101135, 101223.9, 101303.6, 101341.2, 101395, 101424.3,
  95178.23, 96831.76, 99743.17, 100072.3, 100219.9, 100372.9, 100597.9, 
    100761.7, 100895.4, 101015.8, 101103.4, 101159.1, 101267.7, 101331.5, 
    101371.5,
  99438.16, 99593.91, 99787.26, 99945.98, 100066.5, 98483.09, 100113.9, 
    100396.2, 100661.7, 100851, 100998.2, 101108.4, 101192, 101257.4, 101310,
  99362.76, 99440.75, 99619.16, 99745.41, 99796.48, 97519.55, 95853.23, 
    95184.22, 97801.86, 100704.3, 100881.9, 101003.7, 101105.3, 101185.6, 
    101250.6,
  99062.47, 99241.02, 99492.79, 99615.69, 94990.56, 96554.26, 98321.2, 
    99970.75, 100385, 100626.2, 100770.5, 100904.9, 101018.3, 101110.3, 
    101185.4,
  98900.14, 99135.07, 99372.6, 99476.38, 95369.62, 95795.67, 95485.05, 
    100135.2, 100468.3, 100524.1, 100687.6, 100817.4, 100942.2, 101039.8, 
    101124.6,
  101447, 101456.4, 101512, 101559, 101604.7, 101657.8, 101701.2, 101733.3, 
    101763.1, 101781.1, 101790.7, 101778.4, 101762.1, 101731.7, 101687.8,
  101249.6, 101253.5, 101377.8, 101436.5, 101477.5, 101537, 101590.5, 
    101646.8, 101683.8, 101709.5, 101727.6, 101740.7, 101729.2, 101720.4, 
    101689.1,
  99313.98, 99096.04, 101115.1, 101313.6, 101334, 101398.9, 101449.3, 
    101506.4, 101565, 101619, 101641.9, 101669, 101670.2, 101665.4, 101652.3,
  97188.89, 97278.32, 100842.9, 101169.9, 101203.7, 101281.8, 101343.9, 
    101410.3, 101459.6, 101523.2, 101569.5, 101612.5, 101622.9, 101617.9, 
    101633.3,
  97039.8, 97562.54, 99443.08, 101006.7, 101057.9, 101103.4, 101182, 
    101266.9, 101333.4, 101403.7, 101464.3, 101522.1, 101542.8, 101569.7, 
    101584.2,
  96232.85, 97842.08, 100677.3, 100885.6, 100892.5, 100944.1, 101070.8, 
    101146.8, 101208.4, 101293.8, 101343.2, 101381.5, 101480.2, 101520.6, 
    101539.5,
  100592.2, 100668.9, 100753.5, 100803.9, 100801.8, 99038.85, 100567.4, 
    100793.3, 100990.4, 101129.8, 101242.1, 101326.1, 101397.9, 101450.7, 
    101484.6,
  100574.9, 100530, 100580, 100582.2, 100504.9, 98131.8, 96319.99, 95541.05, 
    98098.35, 100982, 101115.4, 101217, 101307.2, 101376.4, 101428,
  100367, 100381.5, 100466.4, 100481.1, 95665.86, 97090.2, 98809.25, 
    100406.8, 100735.7, 100895.9, 101001.8, 101110.3, 101204.9, 101291.6, 
    101359.6,
  100165.5, 100204.8, 100316.2, 100298, 96042.55, 96329.77, 95917.72, 
    100491.5, 100794.6, 100776.9, 100909.6, 101004.2, 101109.4, 101201.1, 
    101285.3,
  101886.4, 101850.4, 101835, 101825.8, 101822.5, 101821.6, 101815.6, 
    101803.4, 101789.7, 101771.6, 101755, 101720.7, 101692.5, 101660.2, 
    101606.7,
  101831.1, 101782.9, 101835.4, 101815.4, 101797, 101795.8, 101790.9, 
    101792.7, 101786.7, 101773.7, 101757.8, 101738.3, 101713.8, 101689.4, 
    101662.7,
  99989.05, 99733.2, 101737.5, 101804.5, 101778.9, 101767.1, 101751.8, 
    101750.7, 101751.9, 101751.1, 101754.8, 101730.8, 101717.2, 101696.9, 
    101671.7,
  97983.64, 98082.64, 101590.2, 101790.8, 101755.2, 101756, 101751.3, 
    101742.5, 101744, 101730.9, 101728.8, 101725.8, 101716.4, 101697.6, 101697,
  97960.74, 98453.94, 100294.5, 101786.4, 101739.8, 101706, 101691.2, 
    101696.5, 101703.5, 101703.2, 101707, 101714.3, 101706.8, 101712.1, 
    101706.8,
  97269.26, 98801.46, 101622.3, 101759.2, 101694.6, 101662.2, 101726.4, 
    101706.4, 101670.9, 101668.9, 101666.8, 101644.9, 101697.3, 101703.6, 
    101705.7,
  101771.4, 101773.4, 101768.2, 101741.1, 101692.9, 99822.72, 101309.1, 
    101449.4, 101569.5, 101615.8, 101640.6, 101655.8, 101671.8, 101673.6, 
    101677.1,
  101746.5, 101693.9, 101695.5, 101614.9, 101447.6, 98996.48, 97088.23, 
    96205.61, 98757.46, 101570.7, 101606.4, 101618.9, 101635.4, 101642.6, 
    101655.3,
  101631.6, 101595.1, 101618.8, 101575, 96620.5, 97974.02, 99703.49, 
    101309.5, 101523.7, 101541.4, 101555.9, 101563.4, 101587.2, 101599.5, 
    101618.4,
  101529.6, 101489.5, 101509.6, 101417.7, 97065.1, 97262.52, 96772.52, 
    101306.6, 101575.1, 101471.3, 101519.3, 101505.3, 101536.2, 101554.2, 
    101579.3,
  100910.2, 100962.9, 101041.6, 101137, 101228.8, 101296.1, 101354.8, 
    101397.3, 101385, 101371.2, 101350.9, 101347.6, 101351.2, 101338.7, 
    101305.4,
  100820.9, 100847.7, 100949.9, 101042.7, 101123.8, 101207, 101275.9, 
    101326.5, 101330.9, 101300.7, 101278.8, 101281.8, 101294, 101299.2, 
    101298.2,
  99034.65, 98845.93, 100838.2, 100977.9, 101044.7, 101120.3, 101188.2, 
    101235.9, 101253.4, 101227.4, 101219, 101222.1, 101238.8, 101243, 101231,
  97067.55, 97255.39, 100758.1, 100965.6, 101022.3, 101084.7, 101136.7, 
    101179.6, 101199.7, 101185.1, 101177.6, 101176.5, 101196.1, 101193.4, 
    101190.8,
  97116.54, 97603.19, 99472.77, 100995.3, 101021.9, 101055.3, 101122.6, 
    101145.8, 101144.5, 101136.9, 101134.9, 101148.8, 101149.6, 101163.7, 
    101149.5,
  96653.05, 98127.88, 100882.8, 100982.8, 101010.7, 100992.2, 101105.8, 
    101143.4, 101154.9, 101137.8, 101114, 101087.6, 101140.4, 101151, 101131.4,
  101126.7, 101083.8, 101048.9, 101066.1, 101038.6, 99285.08, 100824.6, 
    100923.9, 101066.5, 101101.3, 101120.9, 101128.1, 101131.6, 101124.9, 
    101108.9,
  101267.6, 101191.9, 101154.6, 101104, 100906.9, 98434.77, 96572.52, 
    95752.71, 98372.32, 101118.2, 101127, 101120.6, 101129.3, 101118.1, 
    101110.8,
  101350.8, 101266.1, 101250, 101123.2, 96225.39, 97729.8, 99409.98, 
    100994.3, 101158.6, 101151.1, 101153, 101131, 101135.7, 101124.3, 101118.7,
  101451.5, 101368.4, 101355.7, 101206, 96844.35, 97059.77, 96498.59, 
    101103.5, 101254.2, 101186.9, 101185.3, 101156, 101145.6, 101147.6, 
    101143.8,
  100676.4, 100827.8, 101036.2, 101247.1, 101450.9, 101616.8, 101761.6, 
    101884.5, 101974.5, 102039.5, 102070, 102077.5, 102059.7, 102034.9, 102004,
  100310.4, 100485.8, 100742, 100970.7, 101166.4, 101384.6, 101540.4, 
    101680.4, 101789, 101886.3, 101939.7, 101974.8, 101977.7, 101979.4, 
    101986.5,
  98177.52, 98148.81, 100287.6, 100689, 100838.9, 101054.5, 101252, 101438.2, 
    101572.6, 101684.6, 101772.3, 101834.7, 101873.2, 101886.8, 101897.1,
  95707.53, 96057.08, 99872.52, 100391.1, 100534.9, 100786.3, 100986.5, 
    101180.7, 101362.8, 101513.3, 101628.5, 101712, 101763.2, 101795.6, 101844,
  95365.86, 96101.83, 98239.35, 100071.2, 100304.3, 100495.4, 100728.8, 
    100959.8, 101140.9, 101314.6, 101441.9, 101559.1, 101620.8, 101693.2, 
    101750.9,
  94369.3, 96143.62, 99305.75, 99777.73, 100015.8, 100245.3, 100519.3, 
    100729.2, 100914.8, 101103.2, 101255.5, 101347.1, 101493.4, 101585.2, 
    101655.2,
  98529.59, 98898.59, 99272.8, 99569.14, 99802.31, 98267.78, 99951.71, 
    100319.4, 100635.3, 100873.4, 101069.1, 101223.2, 101353.1, 101457.8, 
    101546.7,
  98542.33, 98776.5, 99034.6, 99298.64, 99457.21, 97196.45, 95543, 94886.15, 
    97590.11, 100631.8, 100863.1, 101040.9, 101197, 101324.8, 101431.3,
  98460.19, 98635.66, 98906.31, 99133.54, 94521.09, 96151.2, 98014.1, 
    99716.16, 100191.1, 100467.3, 100649.9, 100841.5, 101021.3, 101177.4, 
    101301.7,
  98492.27, 98615.41, 98820.64, 98976.58, 94863.3, 95328.69, 95093.3, 
    99837.61, 100239.9, 100271.2, 100477.3, 100661.6, 100845.9, 101016.6, 
    101164,
  101673.6, 101667.8, 101741.4, 101824.7, 101889.4, 101990.1, 102064, 
    102137.8, 102190.8, 102247.2, 102268.6, 102269.2, 102248.6, 102222.3, 
    102173.4,
  101319.5, 101392.4, 101523, 101620.5, 101674.9, 101746.3, 101857.3, 
    101957.1, 102029.2, 102084.2, 102130.3, 102156.4, 102159.4, 102156.7, 
    102150,
  99244.1, 99070.58, 101127.9, 101418.4, 101412.6, 101506.9, 101576.5, 
    101698.1, 101811.1, 101899.1, 101971.1, 102023, 102054.6, 102063.1, 
    102067.2,
  96844.34, 97023.37, 100627.9, 101130.9, 101170.9, 101306.2, 101394.9, 
    101499.9, 101611.9, 101723.4, 101810.6, 101889, 101932.2, 101959.6, 
    101995.4,
  96499.56, 97087.75, 99052.27, 100814.6, 100927.1, 101025.9, 101154, 101288, 
    101393.4, 101524.2, 101630.7, 101733.8, 101791.8, 101857, 101895.4,
  95377.04, 97093.72, 100126.5, 100541.8, 100676.9, 100832, 100980.7, 
    101104.4, 101195.4, 101327.1, 101429.7, 101517.1, 101659.2, 101743, 
    101794.4,
  99662.82, 99859.31, 100058.6, 100285.1, 100423.9, 98773.66, 100395.6, 
    100701.9, 100920.4, 101097.3, 101243.3, 101380.7, 101509.9, 101602.1, 
    101675.1,
  99447.33, 99573.47, 99761.39, 99911.44, 99988.77, 97702.76, 95952.39, 
    95232.58, 97851.57, 100891.1, 101047.7, 101191.3, 101331.5, 101456.6, 
    101550,
  99114.67, 99155.43, 99423.55, 99644.7, 94917.93, 96440.58, 98308.34, 
    100004.5, 100498.8, 100727.4, 100846.5, 101001.9, 101153.1, 101290.7, 
    101408.9,
  98813.91, 98862.12, 99032.47, 99184.98, 95125.45, 95511.78, 95322.27, 
    99983.71, 100486.8, 100458.5, 100684.8, 100810.3, 100973.2, 101124.4, 
    101258.9,
  102348.6, 102317.6, 102345.1, 102372.3, 102390.2, 102426.3, 102448, 
    102467.8, 102467.3, 102464, 102462.1, 102448.2, 102408.5, 102358.3, 102295,
  102182, 102194, 102268.2, 102293.6, 102289.8, 102328.5, 102350.5, 102376.4, 
    102390.4, 102393.2, 102382.4, 102367.2, 102337.5, 102305, 102275.8,
  100238.1, 100033.9, 102070.8, 102272.8, 102212, 102231.6, 102232.8, 
    102249.3, 102266.6, 102282.5, 102288.3, 102286.4, 102271.4, 102241.1, 
    102205.4,
  98036.27, 98118.12, 101796.7, 102161.8, 102126.2, 102161.6, 102163.8, 
    102181.1, 102176.7, 102186.3, 102186.4, 102195.9, 102178.5, 102162.2, 
    102158,
  97831.98, 98384.11, 100365.3, 102006.8, 102037.9, 102019.6, 102031.9, 
    102052.3, 102055.4, 102073.8, 102079.4, 102101.2, 102088.5, 102095.9, 
    102086.7,
  96908.92, 98600.32, 101562.2, 101836.4, 101851.9, 101892.1, 101958.2, 
    101970.1, 101951.6, 101964.8, 101953.5, 101947.6, 102010.6, 102023, 102017,
  101364.1, 101498.8, 101606.4, 101688, 101690.2, 99886.05, 101431.3, 
    101620.6, 101745.3, 101834.4, 101862.3, 101889.3, 101913.5, 101930.5, 
    101938.1,
  101300.3, 101281.5, 101374.3, 101416, 101326.9, 98885.56, 97012.59, 
    96179.23, 98756.62, 101692.9, 101763.6, 101783.2, 101808.5, 101834.8, 
    101849.6,
  101175.9, 101105.3, 101169.6, 101196.9, 96313.05, 97720.23, 99504.48, 
    101150.7, 101506.4, 101611.2, 101657.5, 101687.5, 101709.6, 101735.8, 
    101755.1,
  101029.1, 100984.1, 101027.6, 100939.9, 96617.09, 96910.43, 96511.38, 
    101169.1, 101530.8, 101431.4, 101532.5, 101559.6, 101602.1, 101627.5, 
    101658.8,
  101816.6, 101845.2, 101924.9, 102003.3, 102080.5, 102151.3, 102208.8, 
    102257.3, 102299.9, 102328, 102338.1, 102333.9, 102308.8, 102284.6, 
    102239.1,
  101613.7, 101699.2, 101834.7, 101928, 101986.1, 102070.4, 102137.6, 102200, 
    102236.5, 102266.8, 102279.5, 102273.8, 102261.6, 102253.2, 102248.7,
  99745.95, 99628.88, 101677.6, 101883.2, 101914.5, 101992.9, 102055, 
    102121.4, 102166.8, 102201.3, 102216.7, 102226.4, 102223.9, 102209.2, 
    102203.7,
  97559.79, 97818.25, 101527.2, 101828.7, 101859, 101943.9, 101997.3, 102062, 
    102101.2, 102138.6, 102149.9, 102169.6, 102165.4, 102164.3, 102180.3,
  97512.55, 98111.52, 100156, 101755.8, 101811.9, 101854.2, 101921.4, 
    101979.3, 102021.4, 102068.9, 102089.7, 102116.3, 102114.4, 102137.6, 
    102140.8,
  96822.14, 98459.02, 101441, 101675, 101739.2, 101783.9, 101883.8, 101940.3, 
    101968.4, 102007.8, 102020.4, 102018.1, 102083.4, 102108.1, 102116.6,
  101241, 101414.6, 101576.3, 101648.1, 101677.7, 99936.8, 101488.2, 
    101655.6, 101832.5, 101928.7, 101993.1, 102022.8, 102045.9, 102069.9, 
    102083.9,
  101341.2, 101384.3, 101477.7, 101515.2, 101477.7, 99035.12, 97199.7, 
    96388.85, 99011.54, 101880.8, 101953.8, 101994.9, 102018.4, 102039, 
    102054.3,
  101260.3, 101315.6, 101453.5, 101453.3, 96622.16, 98123.11, 99872.3, 
    101496.6, 101776.9, 101862.8, 101917.1, 101953, 101990.2, 102017, 102037.5,
  101293.4, 101326.1, 101426.9, 101391.2, 97081.45, 97370.66, 96954.5, 
    101608.3, 101864.2, 101799.5, 101865.6, 101897.9, 101946.7, 101978.7, 
    102003,
  102174.7, 102163.1, 102221.4, 102274.2, 102317.4, 102360, 102385.1, 
    102409.4, 102427.5, 102450.4, 102456.8, 102449.4, 102420.2, 102385.5, 
    102342.1,
  101918.3, 101991.2, 102088.6, 102155.9, 102193.5, 102266.4, 102314.2, 
    102356.6, 102375.2, 102394.3, 102395.8, 102391.7, 102373, 102351.5, 
    102333.8,
  99926.02, 99783.38, 101834.1, 102069.9, 102046.1, 102117.3, 102167.1, 
    102223.6, 102271.6, 102306.9, 102332.5, 102338.3, 102330.3, 102305, 
    102285.3,
  97608.16, 97821.85, 101540.1, 101948.2, 101947.4, 102035.9, 102084.7, 
    102143.9, 102184.6, 102223.5, 102252.8, 102275, 102268.4, 102251.7, 
    102254.6,
  97460.6, 98056.58, 100091.4, 101790.4, 101815.8, 101867.5, 101940.7, 
    102006.2, 102054.9, 102117.9, 102155.8, 102194.1, 102194, 102202, 102200.2,
  96452.42, 98251.24, 101341.5, 101659.8, 101725.2, 101758.2, 101861.9, 
    101927.4, 101960.5, 102012.1, 102040.7, 102048.4, 102121.7, 102134.9, 
    102144.7,
  100856.7, 101175.2, 101385.4, 101538.5, 101565.6, 99810.45, 101392.5, 
    101577, 101740.6, 101862.6, 101945.6, 101999.4, 102041.3, 102055.8, 102078,
  100852, 100962.1, 101146.6, 101281.4, 101294.5, 98823.11, 97007.95, 
    96224.41, 98825.44, 101743.3, 101830, 101890.8, 101944.3, 101972.2, 
    102007.3,
  100473.3, 100674.1, 100965.9, 101099.3, 96207.2, 97734.08, 99540.45, 
    101183.7, 101535.6, 101674.3, 101724.9, 101783.4, 101845.9, 101883, 
    101930.6,
  100307.7, 100485.4, 100724.3, 100823.8, 96540.94, 96942.27, 96621.05, 
    101320, 101628.7, 101548.3, 101638.8, 101676.9, 101747.8, 101790.1, 
    101853.3,
  102071.1, 101977.8, 101891.9, 101840.4, 101789.8, 101802.3, 101832.5, 
    101888.8, 101945, 102013.4, 102082.5, 102121.8, 102148.4, 102177.6, 
    102183.7,
  102016.2, 101969.4, 101984, 101912.9, 101833.2, 101817.6, 101838.4, 
    101893.4, 101945.6, 102005.9, 102045.2, 102087.8, 102132.9, 102172.6, 
    102197.3,
  100114, 99853.89, 101866.3, 101971.4, 101849.5, 101795.3, 101782.2, 
    101830.4, 101887.2, 101953, 102017.3, 102075.3, 102118.7, 102160, 102185.6,
  97974.2, 98011.98, 101695, 101970.6, 101872.8, 101869.9, 101809.9, 101830, 
    101874.2, 101929.2, 101985, 102045.5, 102101.3, 102134.8, 102175.5,
  97829.14, 98353, 100335.1, 101918.3, 101860.3, 101800.5, 101775, 101781.6, 
    101815.8, 101882, 101947.7, 102013.2, 102061.8, 102116, 102151.6,
  96933.9, 98646.9, 101625.7, 101862.4, 101824.8, 101820.9, 101823.1, 
    101779.3, 101788, 101843.6, 101887.6, 101921, 102037.4, 102093.8, 102129.2,
  101413.6, 101561.8, 101694.9, 101795, 101746, 99903.52, 101446.6, 101568.9, 
    101673.2, 101773.6, 101855.7, 101923, 101993.8, 102050.3, 102098.2,
  101378.3, 101438.8, 101546, 101574, 101520.5, 99009.04, 97151.18, 96324.6, 
    98895.38, 101748.4, 101819.2, 101872.5, 101938.2, 102002.7, 102064.7,
  101157.9, 101194, 101396.2, 101442.5, 96496.4, 97954.88, 99740.46, 
    101343.6, 101665.1, 101752, 101791.1, 101828.1, 101890.8, 101954.7, 
    102021.9,
  101150.2, 101101.1, 101204.2, 101222.6, 96882.71, 97208.66, 96841.2, 
    101517.1, 101806.9, 101690.2, 101767, 101783.2, 101845.8, 101902.6, 
    101972.7,
  102384.2, 102267.6, 102244.4, 102202.2, 102194, 102221.8, 102263.4, 
    102296.2, 102317.9, 102339.7, 102338.5, 102311, 102270, 102228.6, 102188.9,
  102163.9, 102160.1, 102203, 102199, 102128.7, 102109.4, 102101.5, 102158.8, 
    102206.2, 102233.1, 102231.7, 102217.3, 102186.9, 102165.5, 102156,
  100201.4, 99974.85, 101948.2, 102123.9, 102012.3, 101989.2, 101956.9, 
    101965.9, 101999.7, 102050.9, 102079.9, 102092.6, 102085.5, 102084, 
    102078.2,
  97934.67, 98053.53, 101725.4, 102066.3, 101961.2, 101957.5, 101909.8, 
    101880.8, 101879.3, 101907.6, 101942.8, 101983.5, 101996.8, 101994.7, 
    102020.3,
  97772.48, 98318.23, 100282.1, 101912.1, 101908.8, 101825.9, 101801.8, 
    101774.6, 101744.8, 101767.5, 101791, 101840.3, 101867.6, 101909.6, 
    101937.2,
  96806.41, 98483.45, 101488.9, 101734.4, 101729.8, 101753.7, 101766.6, 
    101708, 101638.4, 101641.1, 101649.1, 101662.2, 101761.1, 101808.6, 
    101855.5,
  101290, 101430.9, 101493.7, 101584.2, 101554.2, 99726.87, 101278.3, 
    101412.5, 101467.7, 101513, 101527.4, 101583.1, 101643.7, 101701.9, 
    101764.6,
  101145.5, 101160.4, 101258.7, 101278.8, 101210.4, 98721.66, 96837.88, 
    96016.14, 98556.71, 101415.7, 101449.1, 101473, 101523.4, 101592.4, 
    101658.7,
  101033.3, 100942.3, 101022.5, 101073.1, 96133.16, 97599.18, 99379.98, 
    100998.5, 101305, 101372.8, 101368.2, 101382.8, 101424, 101486.6, 101555.6,
  100996.7, 100882.8, 100878.1, 100797.3, 96481.98, 96798.32, 96385.47, 
    101072.1, 101362.3, 101213.2, 101272.4, 101293, 101335.8, 101388.8, 
    101460.7,
  102422.7, 102381.9, 102397.4, 102422.2, 102455.7, 102500.2, 102522.5, 
    102539.8, 102540.8, 102536.2, 102518.2, 102489.2, 102444.9, 102393.1, 
    102329.4,
  102316.8, 102322.5, 102370.7, 102374.2, 102371.5, 102412.8, 102444.1, 
    102480.5, 102485.8, 102476.5, 102454.5, 102418.5, 102377.3, 102343.1, 
    102311.2,
  100412.2, 100186.6, 102224, 102383.3, 102306.3, 102318.3, 102312.3, 
    102339.3, 102361.2, 102379, 102361.5, 102351.3, 102324.6, 102296.1, 
    102263.9,
  98251.49, 98306.92, 102070.8, 102369.6, 102288.8, 102302.8, 102289.9, 
    102299.7, 102291.2, 102295.5, 102284.7, 102283.9, 102259, 102240, 102237.6,
  98082.22, 98641.25, 100672.4, 102298.5, 102272.1, 102206.3, 102194, 
    102200.1, 102192.8, 102210.9, 102201.9, 102214.4, 102192.5, 102193.4, 
    102182.8,
  97150.26, 98913.65, 101939.8, 102199.6, 102172.6, 102192.2, 102209.8, 
    102179.3, 102127.6, 102131.8, 102116.1, 102101, 102145.9, 102146.9, 
    102141.2,
  101692.2, 101849.7, 101970.4, 102076.8, 102038.8, 100192.4, 101752.2, 
    101916, 102008, 102061, 102061.2, 102075.3, 102091.3, 102095.4, 102095.2,
  101614.7, 101673.1, 101776.3, 101801.3, 101715, 99214.74, 97319.82, 
    96483.58, 99098.66, 102020.9, 102046.4, 102033.1, 102034.1, 102041.3, 
    102050.7,
  101384.9, 101374.7, 101559.4, 101610, 96624.98, 98097.43, 99896.45, 
    101565.9, 101888, 101979.4, 102005.3, 101991.4, 101991.5, 101991.9, 
    102000.7,
  101326.1, 101294.5, 101369.9, 101344.2, 96980.87, 97303.97, 96928.62, 
    101661.3, 101979.5, 101863.4, 101935.3, 101928.5, 101946.5, 101946.2, 
    101951.8,
  102497.3, 102437.5, 102428.7, 102453.2, 102499.4, 102564.3, 102614.5, 
    102648.5, 102663.5, 102668.7, 102655.8, 102625.8, 102589.9, 102552.3, 
    102504.6,
  102481.6, 102475.6, 102463.8, 102453.2, 102423.2, 102479.1, 102516.8, 
    102575.4, 102602, 102603.6, 102592.8, 102571.9, 102548.5, 102522.8, 
    102502.6,
  100585.6, 100348.7, 102355.7, 102457.6, 102373.4, 102376.8, 102380, 
    102423.1, 102459.8, 102490.4, 102502, 102502, 102495.4, 102480.4, 102463.2,
  98417, 98513.48, 102234, 102508.3, 102361.6, 102371.6, 102366.2, 102374, 
    102382.2, 102404.9, 102419.5, 102435.4, 102433.9, 102420.1, 102432.6,
  98324.85, 98876.91, 100842.9, 102443.9, 102388.3, 102285.4, 102261.2, 
    102274, 102288.5, 102307.9, 102324.9, 102348.9, 102353.5, 102373.7, 
    102378.5,
  97436.3, 99152.89, 102162.4, 102391, 102308.9, 102327.4, 102302.1, 
    102239.5, 102201.5, 102216.5, 102218.9, 102216.7, 102283.4, 102312.8, 
    102324.7,
  101983.2, 102138.6, 102202, 102305.7, 102228.5, 100342.6, 101885, 102007.8, 
    102082, 102132.1, 102151.5, 102176.6, 102205.8, 102238.5, 102259.4,
  101890, 101928.4, 102010.8, 102043.4, 101962.1, 99414.83, 97486.38, 
    96620.46, 99197.97, 102078.1, 102094.4, 102101.7, 102123.3, 102160.1, 
    102190.2,
  101649.3, 101652.5, 101839.1, 101885.6, 96860.3, 98336.98, 100139.9, 
    101755.6, 102011.9, 102061.3, 102039.5, 102030.4, 102046.3, 102076.2, 
    102113.8,
  101618.3, 101574, 101607.2, 101635.9, 97228.83, 97560.76, 97161.34, 
    101879.3, 102120.7, 101960.2, 101988.7, 101958.9, 101977.6, 101997, 
    102038.6,
  102008.2, 102002.2, 102066.6, 102122.9, 102180.8, 102228.9, 102256.4, 
    102282.6, 102296.1, 102305.8, 102299.3, 102276.6, 102278, 102266.6, 
    102228.6,
  101810.6, 101869.5, 101978.5, 102061.4, 102100.5, 102173.5, 102215.3, 
    102260.4, 102273.3, 102279.3, 102268.4, 102266.9, 102268.9, 102269.1, 
    102260.7,
  99893.89, 99770.89, 101768.7, 102009, 102012.2, 102088.1, 102131.1, 
    102185.6, 102211.1, 102232.7, 102243.8, 102252.8, 102258.2, 102268.5, 
    102257.7,
  97691.52, 97929.96, 101617.5, 101947.1, 101962, 102068.2, 102114.7, 
    102171.1, 102188.2, 102206.1, 102215, 102237.6, 102251.8, 102259.8, 
    102261.8,
  97590.65, 98212.53, 100243.1, 101874.7, 101902.1, 101959.8, 102034.8, 
    102098.4, 102136.5, 102179, 102200.9, 102222.3, 102238.4, 102256.6, 102267,
  96896.08, 98548.02, 101520.5, 101791.2, 101842.6, 101935.5, 102027.2, 
    102103.4, 102121, 102152.9, 102171.4, 102173.8, 102236.5, 102262.7, 
    102271.8,
  101297.6, 101467.5, 101654.6, 101764.8, 101759.3, 100050.9, 101633.3, 
    101831.5, 102014.6, 102117.7, 102183.8, 102222.6, 102238.6, 102260.2, 
    102273.3,
  101328.8, 101370.9, 101521.5, 101564.5, 101577.1, 99113.98, 97331.09, 
    96562.26, 99209.2, 102090.7, 102183.1, 102222.9, 102247.9, 102272.2, 
    102272.3,
  101096.1, 101164.7, 101425.9, 101474.1, 96640.98, 98148.52, 99956.86, 
    101565.9, 101923.9, 102067.4, 102147.1, 102188.6, 102240.3, 102266.7, 
    102270.4,
  101042.3, 101119.7, 101301, 101318.1, 97022.77, 97384.09, 97085.41, 
    101784.9, 102081.6, 102011.9, 102120.3, 102153.1, 102224.5, 102251.5, 
    102265.7,
  103114.3, 103009.2, 102966.4, 102904.6, 102835, 102794.2, 102735.3, 
    102678.1, 102611, 102550.2, 102472, 102387.7, 102291.6, 102229.5, 102171,
  103006.5, 102949.1, 102977.2, 102938.9, 102843.2, 102790.2, 102724.5, 
    102678.5, 102610.9, 102543.7, 102458.5, 102389.2, 102314.1, 102264.3, 
    102213.5,
  101048.1, 100756.8, 102792.7, 102930.5, 102802.9, 102754.6, 102670.9, 
    102616.4, 102565.1, 102509, 102447.6, 102390.2, 102331.1, 102273.7, 
    102222.7,
  98856.69, 98877.74, 102617.5, 102904.1, 102775.6, 102747.4, 102680, 
    102619.7, 102555.8, 102493.7, 102430.1, 102387.3, 102320.2, 102273.1, 
    102237.6,
  98646.37, 99187.88, 101160.7, 102764.5, 102713.8, 102637.9, 102582.4, 
    102533.5, 102482.3, 102450.2, 102403.9, 102369.4, 102307.3, 102275.9, 
    102238.8,
  97805.66, 99508.95, 102436.5, 102654.9, 102569.1, 102573.6, 102594.3, 
    102550.3, 102459.2, 102411.1, 102348.7, 102286.1, 102292, 102265.5, 
    102233.1,
  102355.3, 102483.2, 102517.3, 102580.7, 102455.5, 100565.3, 102072.6, 
    102226.5, 102323.3, 102365.1, 102335.8, 102301.3, 102265.4, 102243.3, 
    102219.7,
  102323, 102262, 102297.4, 102291, 102166.5, 99626.11, 97691.88, 96811.35, 
    99388.05, 102270.9, 102285.6, 102264.3, 102233.5, 102214.2, 102199.2,
  102153.3, 102105, 102144.1, 102139.4, 97082.53, 98480.08, 100267, 101891.5, 
    102164, 102217.3, 102213.6, 102188.6, 102176.4, 102163.9, 102162.5,
  102083.1, 101999.8, 102012.3, 101893.2, 97437.86, 97692.86, 97298.8, 
    101978, 102276.1, 102098, 102144.5, 102107.6, 102121.2, 102108.2, 102117.6,
  102681.3, 102556.5, 102434.8, 102298.9, 102116.4, 101963.3, 101841.7, 
    101760.3, 101719.1, 101704.9, 101694.4, 101702.6, 101716.5, 101726, 
    101711.3,
  102690.3, 102535.6, 102515.1, 102396.7, 102240.1, 102099.8, 101943.1, 
    101842.8, 101784.8, 101756.2, 101749, 101757, 101767.7, 101783.1, 101786.5,
  100771.6, 100402.7, 102476, 102447, 102296.5, 102182.8, 102027.5, 101923.7, 
    101845.8, 101812.6, 101810.9, 101831.3, 101842.6, 101849.4, 101841.2,
  98673.09, 98700.81, 102372.1, 102465.9, 102336.6, 102280.7, 102156.3, 
    102043.3, 101939.4, 101889.6, 101886.2, 101895.9, 101898.9, 101890.2, 
    101898.6,
  98648.45, 99107.98, 100999.9, 102489.9, 102372.5, 102290.9, 102200.1, 
    102124.2, 102032.3, 101986.7, 101968.6, 101965.6, 101954.9, 101963.2, 
    101951.9,
  97971.7, 99558.85, 102425.4, 102477.9, 102373.2, 102326.4, 102309.1, 
    102242.1, 102145.4, 102086.3, 102038.6, 101989.1, 102021.4, 102020.3, 
    102004.9,
  102513.3, 102567.9, 102533.6, 102482.9, 102393, 100470.6, 101982.8, 
    102022.1, 102114, 102124, 102115.8, 102084.1, 102078, 102063.6, 102043.4,
  102632.3, 102530.4, 102533.1, 102391.1, 102251, 99659.07, 97660.16, 
    96745.32, 99344.81, 102146.6, 102143.8, 102113.9, 102109, 102099, 102078.6,
  102586.1, 102494.4, 102532.5, 102439.6, 97311.87, 98765.23, 100513.8, 
    102049.3, 102217.6, 102212.4, 102184.2, 102145.8, 102130.7, 102115.7, 
    102100.6,
  102591.4, 102500.9, 102523.6, 102387.6, 97878.15, 98092.36, 97532.21, 
    102191.2, 102370.8, 102217.6, 102218, 102168.1, 102165.8, 102139, 102126.1,
  101526.1, 101362.4, 101217.8, 101019.8, 100882, 100749, 100678.3, 100686.5, 
    100719.9, 100767.2, 100817.6, 100868.5, 100915, 100945.6, 100968.5,
  101518.3, 101297.8, 101245.1, 101035.7, 100860.2, 100694.3, 100611.5, 
    100615, 100661.2, 100713, 100775.8, 100852.4, 100909.8, 100953, 101009.3,
  99647.73, 99256.45, 101164.8, 101057.6, 100873.4, 100676.2, 100518, 
    100514.8, 100576, 100660.6, 100755.6, 100852.4, 100913.2, 100965.8, 
    101018.8,
  97675.45, 97685.96, 101043.3, 101096.6, 100871.2, 100678, 100485.5, 
    100469.8, 100526.9, 100624.2, 100735, 100842.3, 100909.5, 100969.4, 
    101041.1,
  97728.01, 98106.8, 99785.67, 101143.9, 100885.4, 100651.7, 100466.9, 
    100431.4, 100489.5, 100607, 100727, 100851.1, 100919.8, 101003.8, 101066.1,
  97226.7, 98648.77, 101259.6, 101223.4, 100950.2, 100634.6, 100473, 
    100438.4, 100502.2, 100610.9, 100714.2, 100812.4, 100947.4, 101038.1, 
    101100.7,
  101810.6, 101717.5, 101471.1, 101354.2, 101048.2, 98961.74, 100192, 
    100222.4, 100419.5, 100578.7, 100734.9, 100874.9, 100983.5, 101073.6, 
    101140.4,
  101921, 101778.7, 101584.7, 101416.2, 100950.4, 98247.65, 96216.74, 
    95338.39, 97851.23, 100600, 100744.8, 100898.3, 101012.2, 101108.7, 101180,
  101985.8, 101830.1, 101691.5, 101481.8, 96296.05, 97649.91, 99109.17, 
    100432.2, 100517.8, 100658.1, 100769.5, 100923.6, 101048.9, 101147.6, 
    101223.3,
  102090.8, 101933.2, 101815.4, 101595.5, 97025.76, 97061.3, 96386.3, 
    100787.9, 100782.2, 100705.7, 100812.8, 100954.7, 101092.1, 101187.7, 
    101269.7,
  101800.9, 101755.9, 101715.7, 101661.9, 101661.7, 101685.5, 101696, 
    101698.6, 101694, 101685.3, 101661.4, 101624.8, 101585.7, 101533, 101476.4,
  101775.8, 101702.5, 101724.6, 101675.1, 101602.9, 101567.5, 101562.2, 
    101588.2, 101600.8, 101600.7, 101585.8, 101558.6, 101530.9, 101503.8, 
    101479.8,
  99906.31, 99613.93, 101607.9, 101675.1, 101560.6, 101519, 101451.5, 101443, 
    101465.8, 101483.2, 101491.4, 101493, 101482.6, 101464.9, 101439.8,
  97865.78, 97980.36, 101474.1, 101644.5, 101505, 101452, 101397.6, 101375.5, 
    101358.5, 101370.8, 101386.4, 101406.3, 101414, 101404.2, 101410.9,
  97855.1, 98329.17, 100120.4, 101573.7, 101448.3, 101361.5, 101320.2, 
    101285.1, 101268.8, 101278.8, 101301, 101328.7, 101342.6, 101358.9, 
    101366.9,
  97270.67, 98741.73, 101484.2, 101529.7, 101358, 101265, 101291.5, 101267.6, 
    101234.9, 101224.2, 101212.2, 101204.9, 101274.4, 101303.6, 101323.1,
  101792.9, 101705.6, 101589, 101471.8, 101327.8, 99410.34, 100841.6, 
    100951.6, 101071.8, 101137.6, 101168.8, 101186.4, 101217, 101246.3, 101274,
  101810.1, 101672, 101568.9, 101395.3, 101084.6, 98568.5, 96626.23, 
    95739.72, 98231.1, 101011.7, 101089, 101118.4, 101151, 101187.8, 101224.2,
  101769.9, 101644.9, 101543.6, 101373.9, 96276.32, 97650.34, 99261.55, 
    100798.2, 100950.2, 100975.5, 100998.4, 101037.7, 101079, 101127.8, 
    101171.2,
  101761.7, 101639.7, 101533.8, 101318.9, 96825.74, 96933.3, 96341.16, 
    100811.7, 100986.9, 100858.5, 100901.3, 100936.3, 100998.9, 101057.3, 
    101112.3,
  102263.7, 102222.1, 102176, 102087.9, 102023.9, 101993.2, 101937.4, 
    101897.1, 101848.5, 101806.8, 101772.3, 101698.7, 101642.7, 101601.2, 
    101546.1,
  102178.4, 102138, 102179.3, 102129.9, 102031.4, 101956.8, 101893, 101840, 
    101780.2, 101734.8, 101700.7, 101661.4, 101638.6, 101608.5, 101581.7,
  100340.7, 100081.6, 102082.6, 102152.1, 102045.1, 101970.1, 101875.3, 
    101792.4, 101718.8, 101679.3, 101649.6, 101654.2, 101633, 101612.1, 
    101586.5,
  98275.99, 98355.98, 101953.4, 102149.2, 102051.8, 101998.5, 101917.4, 
    101838.5, 101729.1, 101666.4, 101635.8, 101636.7, 101627.3, 101602, 
    101591.1,
  98228.52, 98718.74, 100610.9, 102112.8, 102044.2, 101984.2, 101916, 
    101854.4, 101797.8, 101740, 101696, 101670.4, 101630.3, 101619.9, 101606,
  97612.11, 99121.12, 101960, 102083.7, 102014.6, 101972.8, 101997.2, 
    101940.9, 101856, 101799.1, 101739.4, 101681.9, 101687.6, 101649.1, 
    101626.3,
  102029, 102080.7, 102092.6, 102085.7, 102006.5, 100159.9, 101644.4, 
    101730.3, 101809.6, 101799.5, 101782.4, 101746.4, 101731.6, 101699.2, 
    101667.7,
  102151.4, 102084, 102069.1, 101976.4, 101813.2, 99328.66, 97407.8, 
    96487.42, 99015.12, 101777.8, 101801.1, 101764.7, 101735.3, 101712.2, 
    101696.1,
  102110.6, 102049, 102067.9, 101973, 96996.47, 98430.73, 100147.2, 101698.6, 
    101853.1, 101845.8, 101828.3, 101776.3, 101748.3, 101718.7, 101695.8,
  102150.8, 102078.6, 102080.4, 101927, 97532.69, 97757.51, 97228.27, 
    101773.8, 101949.6, 101812, 101814.4, 101764.6, 101748.5, 101711.2, 
    101690.3,
  102172.6, 102148.8, 102123.9, 102087.9, 102057.3, 102035.8, 101993.9, 
    101953, 101886.7, 101828.6, 101775.6, 101725.9, 101665.7, 101610.4, 
    101536.2,
  102090.1, 102071.2, 102118.3, 102108.7, 102047.7, 102001.7, 101937.3, 
    101875.5, 101806.9, 101747.6, 101701.1, 101651.5, 101595.8, 101566.6, 
    101529.8,
  100247.1, 99968.83, 101986.3, 102082.2, 102016.8, 101970.5, 101894.9, 
    101816.8, 101709.7, 101639.8, 101599.1, 101568.6, 101531.2, 101503.9, 
    101464,
  98155.57, 98229.84, 101838.1, 102061.5, 101990.3, 101950.9, 101875.5, 
    101789.9, 101657.9, 101565.6, 101516, 101499.5, 101467.4, 101443.5, 
    101432.7,
  98071.53, 98544.62, 100439.1, 101979.9, 101934.9, 101874, 101826.6, 
    101758.7, 101650.1, 101522, 101458.4, 101436.6, 101414.8, 101410.4, 
    101384.2,
  97414.27, 98907.73, 101768.2, 101908.5, 101850.5, 101809.6, 101839.3, 
    101796.2, 101695, 101565.1, 101441.9, 101360.7, 101385.7, 101377.2, 
    101352.9,
  101812.4, 101830.6, 101835, 101850, 101797.6, 99967.48, 101486.8, 101583.7, 
    101615.2, 101557, 101475.9, 101399.1, 101362.7, 101348.9, 101326.7,
  101823, 101799.8, 101769.3, 101720.4, 101591.5, 99106.56, 97197.39, 
    96320.23, 98849.76, 101569.8, 101493.7, 101398.8, 101349.2, 101331.5, 
    101311.5,
  101839.9, 101757.8, 101681.8, 101657.2, 96726.79, 98230.31, 99934.04, 
    101506.3, 101647.7, 101573.2, 101485.2, 101392.2, 101340.4, 101312, 
    101290.6,
  101935.1, 101839.6, 101758.5, 101634.9, 97255.38, 97539.34, 96984.42, 
    101597.5, 101713.3, 101555.5, 101485, 101388.8, 101338.1, 101300.3, 
    101284.1,
  102344.2, 102321.7, 102341.7, 102357.2, 102377.9, 102397.9, 102380.6, 
    102354, 102300, 102250.2, 102198.3, 102115.5, 102029.6, 101975.8, 101914.9,
  102216.6, 102248.3, 102311.2, 102332, 102329.6, 102351.4, 102346.8, 
    102329.9, 102297, 102240, 102193.9, 102128.1, 102057.8, 102001.5, 101954.5,
  100364.3, 100179.4, 102181.6, 102315, 102281.5, 102293.6, 102281.4, 102273, 
    102244.1, 102218.3, 102170.7, 102122.8, 102058.8, 102004, 101956.5,
  98246.07, 98402.06, 102050.9, 102324.2, 102268.2, 102298.3, 102285.3, 
    102276, 102231.8, 102205.4, 102162.8, 102123.1, 102067.2, 102015.7, 
    101983.4,
  98211.09, 98718.83, 100665.2, 102252.2, 102241.4, 102212.9, 102211.6, 
    102209.9, 102194.3, 102172.7, 102147.7, 102108.5, 102071.8, 102036.2, 
    101995.1,
  97479.76, 99042.3, 101953.6, 102174.8, 102163.2, 102186.3, 102230.8, 
    102218.5, 102177.6, 102155.6, 102112.3, 102057.5, 102077.8, 102044.2, 
    102005.7,
  101864.7, 101971.5, 102032, 102107.1, 102082.8, 100290.1, 101819.7, 101972, 
    102081, 102121.6, 102122.1, 102095.7, 102070.7, 102037.7, 101995.3,
  101871.9, 101863.4, 101909.3, 101920.4, 101853.3, 99403.05, 97535.07, 
    96704.98, 99267.74, 102097.1, 102109.5, 102086.8, 102052, 102018.1, 
    101980.1,
  101793.5, 101785.4, 101754.1, 101792.2, 96937.87, 98406.2, 100154, 
    101771.5, 102008.1, 102058.1, 102061.6, 102039.9, 102014.9, 101981.9, 
    101948,
  101772.7, 101769.9, 101696.8, 101631.7, 97338.41, 97681.35, 97249.61, 
    101849.4, 102099.7, 101986.4, 102014.3, 101978.8, 101970.6, 101937.1, 
    101909.4,
  102839.5, 102738.5, 102692.1, 102588.8, 102452, 102345.8, 102244.3, 
    102162.2, 102106.3, 102099.9, 102097.8, 102089.5, 102107.8, 102116, 
    102093.5,
  102826.4, 102730.4, 102748.3, 102652.1, 102556.6, 102452.5, 102336.6, 
    102226.4, 102152.8, 102128.8, 102117.9, 102130.1, 102144.5, 102145.7, 
    102143,
  100954.4, 100625.9, 102668.1, 102712.9, 102585.8, 102502.1, 102393.6, 
    102292.1, 102203.1, 102146.3, 102146.7, 102169.1, 102182.2, 102184.4, 
    102182.6,
  98901.72, 98909.94, 102538.7, 102742.8, 102624.5, 102586.3, 102464.9, 
    102372.1, 102272.5, 102211.6, 102213.1, 102217.2, 102235.9, 102211.9, 
    102234.2,
  98815.6, 99302.77, 101195.9, 102728.8, 102642.8, 102567.6, 102491, 
    102396.6, 102317.6, 102265.6, 102253.1, 102260.3, 102274.3, 102279.6, 
    102278.6,
  98086.98, 99678, 102557.1, 102705.3, 102626.3, 102583.1, 102565.6, 102477, 
    102376.2, 102321.3, 102293.7, 102260.2, 102325.9, 102339.5, 102327.1,
  102567.7, 102632.1, 102682, 102680.6, 102613.8, 100731.6, 102225.6, 
    102259.3, 102334, 102343.4, 102356.6, 102354.5, 102373.3, 102371.8, 
    102352.9,
  102621.1, 102577.7, 102617.9, 102555.4, 102441.7, 99907, 97958.65, 
    97036.75, 99618.16, 102386.6, 102412.8, 102415.3, 102415.9, 102404, 
    102385.1,
  102425.2, 102439.6, 102548.6, 102526.3, 97536.93, 98950.52, 100722, 
    102278.5, 102436.6, 102412.8, 102434.2, 102430.5, 102430.2, 102418.9, 
    102398.7,
  102376.7, 102363.8, 102442.6, 102398.8, 98006.63, 98255.52, 97777.02, 
    102376.2, 102572.9, 102412, 102448.1, 102433.5, 102452.1, 102429.8, 
    102412.9,
  102956.7, 102845.8, 102784.7, 102695.1, 102593.2, 102486.9, 102381.2, 
    102271.5, 102175.1, 102138.8, 102114.4, 102106.8, 102095.7, 102081.4, 
    102061.7,
  102913.9, 102796.9, 102826.5, 102732.5, 102607, 102486.2, 102350.6, 
    102214.4, 102120.5, 102082.2, 102052.2, 102042.4, 102044.7, 102052.9, 
    102058.7,
  101033, 100704.3, 102727.3, 102753.6, 102607.3, 102505.5, 102372.9, 
    102248.4, 102091.4, 102024.8, 102003.6, 102005.2, 102012.9, 102025.8, 
    102033.4,
  98959.83, 99006.64, 102607.9, 102768.7, 102620.9, 102552, 102408.9, 
    102283.3, 102099.4, 102003.4, 101967.8, 101968.3, 101979.3, 101982.6, 
    102017.1,
  98930.58, 99406.08, 101270.6, 102749.1, 102641.3, 102543.5, 102430.3, 
    102279.5, 102082.1, 101983.7, 101938.2, 101937.8, 101939, 101969.1, 
    101996.7,
  98252.95, 99789.05, 102643.9, 102723.3, 102638.4, 102535, 102515.1, 
    102383.7, 102205.3, 102034.5, 101900.9, 101856.4, 101909.9, 101950.6, 
    101979.2,
  102816.5, 102809.4, 102819.1, 102736.9, 102647.9, 100712.1, 102165.2, 
    102102.8, 102109, 102029.6, 101906.2, 101870.3, 101879.9, 101915.2, 
    101952.8,
  102891.4, 102804.2, 102786.6, 102658.6, 102482, 99916.85, 97882.36, 
    96902.59, 99483.09, 102117.1, 101945.3, 101852.5, 101853.2, 101884.8, 
    101930.4,
  102798.2, 102737.3, 102744.6, 102684.2, 97603.16, 99000.08, 100737.7, 
    102274.6, 102326.9, 102156.2, 101997.6, 101850.3, 101832.2, 101852.8, 
    101901.3,
  102833.2, 102751.6, 102743.4, 102619.2, 98147.41, 98346.7, 97762.88, 
    102336.3, 102439.4, 102188.6, 102074.2, 101879, 101830.1, 101831, 101878.5,
  103283.3, 103182.7, 103109.8, 102996.6, 102913.6, 102828.5, 102683.6, 
    102556.4, 102446.7, 102339.4, 102253.2, 102208.4, 102189.4, 102180.4, 
    102140.5,
  103201.4, 103125, 103119.9, 103058.5, 102934.3, 102829.5, 102698.1, 102585, 
    102463.8, 102340.7, 102242.9, 102199.9, 102181, 102176.1, 102156.7,
  101313.1, 100979.1, 102985.5, 103054.5, 102931.1, 102837.3, 102705.8, 
    102583, 102480.7, 102383.9, 102254.6, 102220.9, 102198.4, 102177.5, 
    102160.5,
  99198.22, 99182.24, 102857.7, 103045.2, 102915.9, 102856.2, 102739.7, 
    102630.6, 102504.8, 102412.9, 102290.3, 102232.1, 102205.5, 102170.6, 
    102158.5,
  99100.95, 99570.99, 101480.9, 102999.7, 102899.9, 102809.6, 102727.9, 
    102641, 102542.6, 102439.5, 102332, 102266.8, 102207.4, 102194.8, 102163.4,
  98353.7, 99920.66, 102805.8, 102956, 102846.1, 102797.1, 102790.8, 
    102718.8, 102594.7, 102486.4, 102347.1, 102239.1, 102229, 102211.9, 102177,
  102893, 102922.3, 102926.5, 102930, 102803.3, 100919.8, 102409.9, 102464.1, 
    102501.3, 102457, 102383.6, 102303.2, 102250.8, 102228.2, 102186,
  102886.8, 102819.6, 102830.2, 102750, 102608.3, 100065.3, 98129.36, 
    97189.59, 99720.97, 102464.3, 102407.4, 102327.4, 102267.4, 102239.3, 
    102198.1,
  102777.5, 102725, 102762.8, 102709.1, 97675.52, 99074.52, 100843.3, 
    102395.3, 102540.2, 102496.8, 102406.9, 102334, 102278.9, 102247.9, 
    102201.8,
  102769.5, 102694, 102691.8, 102582.9, 98138.57, 98367.87, 97880.97, 
    102490.1, 102673.5, 102480.2, 102432.1, 102351.4, 102290.5, 102248.3, 
    102208.3,
  103613, 103523.5, 103468.2, 103377.4, 103264.9, 103180.1, 103063.1, 
    102908.2, 102743.5, 102614, 102464.1, 102323.3, 102221.5, 102192.4, 
    102164.8,
  103524.7, 103454.8, 103475.5, 103410.5, 103284, 103183, 103042.1, 102916.4, 
    102773.6, 102628.6, 102462.8, 102332.1, 102229.4, 102183.7, 102182.6,
  101610.1, 101277.2, 103315.8, 103390.1, 103260.5, 103165.7, 103036.8, 
    102908.9, 102759.4, 102630.5, 102487.9, 102355.9, 102259.8, 102195.7, 
    102187,
  99471.95, 99479.9, 103178.4, 103379.5, 103237.5, 103167.7, 103053.4, 
    102936.7, 102788.9, 102665.8, 102520.9, 102389, 102279, 102195.3, 102189.9,
  99367.07, 99856.13, 101750.9, 103304.7, 103203.1, 103111.5, 103029.6, 
    102924.3, 102807.5, 102697, 102545.2, 102429.8, 102303.7, 102233.1, 
    102202.8,
  98615.13, 100208.6, 103117.7, 103245.9, 103140.8, 103080.6, 103073.7, 
    102995.5, 102878.4, 102752.6, 102593.7, 102437.6, 102357.2, 102272.4, 
    102224.5,
  103183.5, 103218.4, 103202.9, 103196.9, 103082.7, 101170.3, 102670, 
    102740.5, 102800, 102741, 102637.3, 102514, 102391.9, 102291.7, 102231.5,
  103170.5, 103110.2, 103120, 103008.7, 102864.3, 100300.4, 98320.24, 
    97382.04, 99959.17, 102743.9, 102669.7, 102547.2, 102419.6, 102306.8, 
    102241.4,
  103077.7, 103034.9, 103065.8, 102988.9, 97904.26, 99326.14, 101090.4, 
    102664.4, 102814.2, 102765.6, 102661.5, 102562.7, 102448.6, 102325.9, 
    102260.7,
  103083.4, 103014.7, 103025.6, 102909.8, 98419.62, 98646.25, 98108.58, 
    102738.9, 102915.8, 102740.6, 102683.5, 102572.9, 102476.8, 102348.4, 
    102265.9,
  103345.3, 103247.2, 103154.1, 103059.4, 102944.2, 102838.3, 102705.4, 
    102552.1, 102401.9, 102283.6, 102136.9, 102049.9, 102036.4, 102049.7, 
    102031.2,
  103328.3, 103202.8, 103205.3, 103100.1, 102961.2, 102856.9, 102714.3, 
    102588.3, 102454.8, 102322.3, 102177.4, 102050.4, 102019.6, 102043.3, 
    102074.3,
  101434.7, 101052.9, 103117.3, 103128.7, 102982.5, 102885.4, 102743, 102613, 
    102463.7, 102347.9, 102226.3, 102096.2, 102053.6, 102061, 102071.1,
  99349.3, 99341.85, 102998.2, 103146.1, 102993.1, 102925.7, 102791, 
    102681.3, 102529.3, 102398.5, 102255.3, 102130.9, 102062.8, 102050.7, 
    102082.4,
  99272.18, 99749.01, 101634.3, 103129.4, 103011.5, 102918.3, 102817.1, 
    102719.8, 102591.8, 102453.6, 102302.2, 102188.2, 102098.2, 102091.7, 
    102093.5,
  98583.61, 100127.9, 103016.2, 103104.1, 103010, 102917.7, 102879.1, 
    102800.2, 102655.2, 102524.4, 102351.4, 102177.8, 102136.2, 102120.5, 
    102108.8,
  103122.3, 103155.5, 103154.2, 103109.2, 103021.9, 101060.1, 102546.5, 
    102580.9, 102589.3, 102534.1, 102413.4, 102275.3, 102176.5, 102148.4, 
    102125.9,
  103152.3, 103094.6, 103102.1, 102994.9, 102845.4, 100254, 98214.78, 
    97227.41, 99836.12, 102582.6, 102462.9, 102323.5, 102211.2, 102169.8, 
    102140.5,
  103065.5, 103022.9, 103049.7, 103000.5, 97914.31, 99344.2, 101083.1, 
    102633.6, 102758.1, 102629.9, 102510.8, 102375.2, 102249.1, 102195.1, 
    102160.6,
  103099.6, 103026.6, 103028.4, 102914.3, 98436.62, 98670.77, 98092.62, 
    102705.3, 102847.2, 102642.6, 102570.4, 102423.3, 102293.2, 102224.3, 
    102179.3,
  102891.1, 102772.6, 102657.8, 102544, 102413.4, 102299.7, 102150.8, 
    102006.1, 101860, 101741.6, 101655, 101559.2, 101514.6, 101528.3, 101533.6,
  102822, 102698, 102677, 102571.3, 102405.2, 102283.3, 102129.6, 101998.9, 
    101839, 101691.9, 101573.1, 101486.1, 101443.3, 101479.2, 101517.9,
  100910.8, 100534.7, 102534.2, 102566.7, 102382.9, 102268.6, 102106.6, 
    101960.6, 101794.5, 101650.7, 101564.1, 101457, 101380.2, 101430.7, 
    101471.1,
  98797.85, 98786.86, 102405.9, 102548.5, 102364.7, 102261.5, 102119.3, 
    101978.2, 101798.6, 101648.5, 101528, 101421.3, 101320.1, 101378.4, 
    101435.4,
  98680.07, 99140.87, 101015.2, 102492.7, 102342.6, 102218.3, 102113.9, 
    101965.3, 101794.2, 101652.5, 101513.7, 101430.2, 101290.9, 101353.3, 
    101399.8,
  97988.19, 99513.92, 102371.8, 102459.2, 102296.2, 102182.6, 102163.7, 
    102037.6, 101869.1, 101700.8, 101521.2, 101402.2, 101298.2, 101334.1, 
    101373.6,
  102492.5, 102506.2, 102467.3, 102415, 102279.4, 100349.7, 101787.1, 
    101769.3, 101758.2, 101668.2, 101539.4, 101416.1, 101305.5, 101314.6, 
    101348.6,
  102577.7, 102463.8, 102420.9, 102293.2, 102072.1, 99504.7, 97480.14, 
    96493.02, 99013.25, 101694.1, 101551.9, 101393.7, 101277.5, 101279.8, 
    101319.6,
  102452.9, 102364, 102367.4, 102278.6, 97181.2, 98566.52, 100274.9, 101816, 
    101887, 101707.5, 101555.9, 101379.4, 101256.5, 101248.3, 101286.6,
  102396.8, 102324.9, 102322.6, 102185.8, 97688.81, 97891.65, 97293.48, 
    101880.7, 101954.3, 101698.6, 101574.8, 101400.3, 101282.9, 101225.7, 
    101263.8,
  102832.3, 102793.4, 102778.3, 102742.9, 102704, 102676.5, 102623.6, 
    102579.4, 102503.7, 102426, 102335.4, 102229, 102116.3, 101990.9, 101861.1,
  102705.7, 102677.3, 102723.1, 102708.2, 102648.5, 102606.2, 102569, 
    102513.5, 102446.7, 102363.4, 102274, 102176.7, 102066.6, 101973.6, 
    101888.5,
  100748.7, 100479.8, 102530.6, 102653.3, 102579.1, 102534.9, 102463.1, 
    102409.1, 102344.5, 102289, 102201.1, 102129.6, 102038.3, 101944.4, 
    101849.4,
  98569.7, 98608.95, 102320.5, 102577.5, 102490.3, 102482.4, 102419.2, 
    102373.4, 102291.5, 102226.1, 102134.5, 102073.1, 101976.5, 101905.8, 
    101828.4,
  98420.95, 98920.58, 100848.9, 102428.5, 102386, 102327.6, 102280.2, 
    102242.3, 102189.9, 102141.5, 102074.2, 102013.8, 101930.6, 101870.8, 
    101791,
  97589.49, 99213.09, 102140.6, 102305.7, 102238, 102219.2, 102236.4, 102196, 
    102122, 102075, 101997.8, 101910.5, 101896.5, 101838.6, 101766.4,
  102065.1, 102161.8, 102158.1, 102184.4, 102115.1, 100242.8, 101750.3, 
    101885.9, 101965, 101994.9, 101956.7, 101895.6, 101839.1, 101784.9, 
    101725.7,
  102062.1, 102017.8, 102005.1, 101947.8, 101811.5, 99289.01, 97337.55, 
    96479.56, 99068.79, 101918.2, 101921.6, 101852.6, 101786.3, 101738.7, 
    101684.3,
  101945.7, 101894.5, 101915.9, 101861.6, 96772.01, 98207.45, 99975.45, 
    101595.2, 101821.4, 101858.8, 101830.6, 101782.4, 101727.9, 101680.9, 
    101629.3,
  101905.9, 101827.4, 101845.2, 101718.4, 97255.08, 97482.98, 96960.59, 
    101630.1, 101857.4, 101721.2, 101734, 101696.9, 101660.6, 101618.2, 
    101573.4,
  102800.9, 102762.5, 102727.5, 102669.8, 102608.9, 102566.5, 102508.7, 
    102441.5, 102366.9, 102293.6, 102223.9, 102143.1, 102088.3, 102037, 
    101981.8,
  102741.8, 102703.3, 102747, 102704.6, 102622, 102578, 102511.4, 102463.8, 
    102404.5, 102334.9, 102260.4, 102189.4, 102135.5, 102095.2, 102058,
  100831.8, 100541.7, 102618.4, 102712.8, 102610.7, 102576.5, 102499.6, 
    102451.8, 102386.5, 102333.5, 102265.2, 102217.2, 102166.6, 102129.8, 
    102077.3,
  98707.6, 98740.24, 102432.1, 102684.1, 102589.5, 102566, 102517.3, 
    102472.1, 102400.9, 102341.5, 102292.1, 102254.6, 102204.6, 102149.9, 
    102121.3,
  98585.52, 99110.59, 101039.1, 102599.7, 102552.1, 102497.6, 102450.5, 
    102419.6, 102374.4, 102341, 102291.6, 102263.5, 102221.5, 102186, 102150.9,
  97761.02, 99420.63, 102327.3, 102532.5, 102454, 102447.2, 102490.8, 
    102457.3, 102374.5, 102341, 102276.9, 102234, 102243.3, 102216.9, 102164.6,
  102269.7, 102386.4, 102432.7, 102464.7, 102409.6, 100519.2, 102051.7, 
    102211.9, 102323.4, 102345.2, 102320.9, 102279.4, 102239.8, 102210.1, 
    102167.4,
  102253.8, 102248.1, 102301.1, 102255.4, 102137, 99642.59, 97702.7, 
    96788.06, 99403.76, 102292.2, 102302.3, 102265.3, 102232.1, 102199, 
    102173.3,
  102087.8, 102094.2, 102173.1, 102175, 97147.52, 98574.34, 100382, 102035.5, 
    102250.1, 102255.6, 102247.9, 102212.4, 102198, 102175.3, 102157.1,
  102026.4, 102019.2, 102064.9, 102010.4, 97566.8, 97837.52, 97370.45, 
    102056.2, 102307.7, 102157.7, 102194.7, 102154.1, 102159.3, 102140.3, 
    102127.7,
  102236.4, 102085.8, 101933.8, 101763.9, 101567.8, 101381.2, 101256.5, 
    101210.5, 101182.9, 101179.6, 101223.3, 101278, 101354.8, 101437.3, 
    101488.6,
  102212.2, 102064.5, 102041.6, 101889.1, 101735, 101557.5, 101386.9, 
    101302.2, 101247.5, 101239, 101256.2, 101305.8, 101386.2, 101462.9, 
    101535.5,
  100369.8, 100038.9, 102034.9, 101971.7, 101835.7, 101685.4, 101516.4, 
    101409, 101329, 101307.6, 101313.7, 101354.1, 101427.1, 101495, 101564.1,
  98346.16, 98427.66, 101971.5, 102073.3, 101958.6, 101845.1, 101687.8, 
    101537.3, 101456.9, 101403.8, 101399.5, 101426.9, 101481, 101528, 101613.2,
  98391.83, 98844.64, 100678.1, 102152.8, 102048.4, 101927.7, 101823.5, 
    101695.1, 101594.7, 101534.9, 101509.7, 101514.9, 101542.9, 101606.1, 
    101679.1,
  97787.6, 99320.83, 102135.4, 102193.7, 102109.8, 101988.4, 101994.3, 
    101873.1, 101749.4, 101681.6, 101618.3, 101571.6, 101637.9, 101687, 
    101736.1,
  102358.6, 102352.3, 102297.9, 102266.8, 102169.1, 100220.3, 101729.6, 
    101720.4, 101803.7, 101769.5, 101739.7, 101713.7, 101728.8, 101758.4, 
    101800.6,
  102442.1, 102358.3, 102332.7, 102240.9, 102037.6, 99443.59, 97451.8, 
    96546.95, 99166.8, 101897, 101855.3, 101811.2, 101817.2, 101833.8, 
    101862.8,
  102429.1, 102357, 102362.2, 102258.8, 97191.33, 98660.68, 100376.7, 
    101924.2, 102063.6, 102010.4, 101957.6, 101903.6, 101896.5, 101899.7, 
    101922.3,
  102436.9, 102376, 102382.6, 102261, 97785.32, 97995.2, 97408.64, 102045.3, 
    102196.7, 102077.8, 102043.3, 101980.3, 101971.3, 101965.5, 101985.9,
  101615.5, 101506.2, 101448.9, 101363.1, 101282.1, 101214.4, 101180.3, 
    101179.7, 101190.2, 101197.8, 101184.3, 101148.6, 101119.8, 101118.1, 
    101108.6,
  101468.2, 101388.9, 101404.8, 101310.9, 101203.4, 101109.6, 101049.8, 
    101050.5, 101076.2, 101103.3, 101113.4, 101095, 101079.2, 101101.4, 
    101126.2,
  99595.66, 99308.39, 101267.1, 101288.1, 101152.2, 101053.1, 100949.8, 
    100931.1, 100956.5, 101002.2, 101041.3, 101047.8, 101055.8, 101086.2, 
    101109.7,
  97523.92, 97602.58, 101112, 101240.4, 101103.4, 101008.5, 100877.3, 
    100839.1, 100858.6, 100906.3, 100964.2, 100998.1, 101023.8, 101056.6, 
    101107.6,
  97530.61, 97972.73, 99785.03, 101218.3, 101087.9, 100948.7, 100828.2, 
    100750.8, 100758.6, 100814.5, 100888.8, 100953.9, 100985.7, 101050.7, 
    101101.3,
  96947.12, 98389.84, 101143.5, 101184.1, 101070.6, 100910.9, 100820.4, 
    100717, 100689.5, 100742.6, 100813.9, 100852.9, 100961.7, 101037.6, 101102,
  101388.2, 101348.9, 101263.1, 101209.6, 101074.2, 99152.32, 100461.7, 
    100471.9, 100565.4, 100636.7, 100755.5, 100838.8, 100927.7, 101013.1, 
    101096,
  101502.7, 101391.9, 101304.8, 101181.9, 100931.5, 98349.27, 96346.2, 
    95452.95, 97896.44, 100576, 100705.1, 100782.2, 100881.6, 100979.2, 
    101082.7,
  101539.6, 101411.2, 101366.6, 101208.1, 96199.8, 97622.07, 99165.88, 
    100599.4, 100604.7, 100600.3, 100667.6, 100735.8, 100840.6, 100945, 
    101062.8,
  101624.8, 101492.5, 101440, 101261.4, 96795.68, 96941.7, 96313.7, 100766.1, 
    100764.1, 100602.5, 100649.6, 100713, 100809.4, 100917.7, 101045.5,
  101910.8, 101880.9, 101891.8, 101902.8, 101913.2, 101929.5, 101938.6, 
    101938.4, 101918.3, 101894.3, 101859.7, 101799.3, 101727.6, 101640.5, 
    101558.2,
  101725.6, 101730.7, 101814.8, 101825.8, 101818.8, 101825.2, 101817.7, 
    101808.9, 101799.1, 101781.6, 101754.1, 101708.1, 101646, 101581.1, 
    101540.6,
  99823.05, 99604.95, 101626.4, 101781.6, 101749, 101744.8, 101719.5, 101700, 
    101678.5, 101658.2, 101637.3, 101611, 101569.6, 101519.9, 101477.7,
  97719.34, 97755.02, 101408.9, 101674.8, 101657.4, 101675.7, 101652.4, 
    101628, 101589.9, 101566.8, 101532.5, 101513.5, 101479.3, 101437.2, 
    101429.7,
  97598.72, 98071.16, 100003.9, 101554.1, 101560, 101539.6, 101540.2, 
    101515.9, 101480.4, 101473.1, 101442.2, 101438.8, 101400.9, 101383.2, 
    101366.4,
  96819.25, 98381.95, 101270.5, 101448.8, 101451.3, 101437.9, 101483.4, 
    101461.6, 101409.6, 101386, 101344.9, 101311.1, 101339.4, 101325.9, 
    101310.3,
  101190.4, 101265, 101340.8, 101373.2, 101346, 99541.49, 101050.9, 101163.7, 
    101272.4, 101299.2, 101294.9, 101275.6, 101273.5, 101264.3, 101251.4,
  101198.1, 101179.7, 101209.9, 101179.4, 101071.1, 98633.09, 96738.75, 
    95886.95, 98422, 101212.7, 101253.8, 101218.7, 101206.3, 101195.9, 101194,
  101071.9, 101056.5, 101130.9, 101104.2, 96200.91, 97649.84, 99373.8, 
    100948.9, 101145.6, 101182.5, 101177.5, 101163.6, 101159.2, 101141.3, 
    101139.5,
  101054.8, 101022.9, 101066.1, 100993.2, 96664.98, 96922.3, 96434.98, 
    100974.2, 101191.2, 101079, 101100.6, 101102.5, 101112.2, 101093.6, 101093,
  102477, 102452.4, 102483.7, 102517.9, 102537.1, 102583.9, 102599.6, 102601, 
    102580.8, 102544.3, 102503.8, 102437.9, 102354.5, 102274.7, 102213,
  102219.2, 102301.9, 102397.7, 102438.2, 102439.5, 102473.3, 102494.2, 
    102519.3, 102513.9, 102491.9, 102459.9, 102397.3, 102325.3, 102273.1, 
    102234.9,
  100294.4, 100162.8, 102187.1, 102393.7, 102366.7, 102395.9, 102401.9, 
    102413.6, 102419.3, 102417.5, 102392.9, 102352, 102298.7, 102253.9, 102215,
  98087.23, 98304.29, 101984.6, 102315.6, 102292.2, 102344.4, 102347.3, 
    102359.9, 102355.2, 102347.7, 102321.5, 102300, 102263.2, 102221.7, 
    102205.5,
  98033.93, 98574, 100583.2, 102218.3, 102224, 102224.9, 102251.3, 102268.8, 
    102263.3, 102277.1, 102268, 102257.2, 102224.7, 102206.5, 102181.9,
  97277.27, 98890.28, 101882.1, 102117.1, 102131.4, 102161.4, 102209.6, 
    102225.5, 102210.5, 102212.6, 102195.7, 102164.5, 102201.8, 102194.2, 
    102165.2,
  101732.6, 101860.3, 101964.1, 102062.8, 102035.1, 100241.3, 101776.3, 
    101925.7, 102053.6, 102131.9, 102155.6, 102165, 102167.7, 102162.3, 
    102146.8,
  101721, 101710.3, 101811.1, 101848.5, 101784.1, 99311.7, 97448.12, 
    96641.78, 99215.02, 102067.3, 102121.1, 102121.6, 102127.2, 102130.2, 
    102121.8,
  101491.1, 101530.8, 101696, 101721.4, 96826.61, 98294.79, 100062.5, 
    101659.6, 101955.3, 102036.9, 102068.9, 102080.6, 102089.1, 102092.5, 
    102092.2,
  101394.6, 101418.3, 101542, 101527.4, 97182.17, 97514.34, 97154.6, 
    101788.6, 102055.3, 101945.4, 102008.2, 102016.1, 102048.8, 102052.8, 
    102060.1,
  103029.9, 103021.2, 103066.8, 103089.8, 103098.4, 103120.1, 103119.9, 
    103102.8, 103054.6, 102992.9, 102915.6, 102818.4, 102696.1, 102566.5, 
    102497,
  102840, 102886.8, 102999, 103031, 103025.4, 103045.9, 103043.7, 103035.9, 
    103003.9, 102953.8, 102887.9, 102797.2, 102704.9, 102620.6, 102544.7,
  100871.6, 100707.1, 102777.9, 102984.8, 102947.7, 102963.6, 102949.4, 
    102944.6, 102926.2, 102898.9, 102851.7, 102784.5, 102707, 102630.9, 
    102563.5,
  98691.47, 98850.39, 102583.7, 102937.5, 102892.8, 102941, 102925.6, 
    102912.8, 102877.8, 102846.9, 102793.8, 102756.7, 102694.1, 102634.4, 
    102585.6,
  98657.82, 99167.28, 101153.5, 102819.9, 102831.4, 102815.6, 102820.1, 
    102817.2, 102801.6, 102786.9, 102755.3, 102724.3, 102676.1, 102632.7, 
    102583.5,
  97839.16, 99506.85, 102503, 102731.2, 102737, 102768.6, 102815.1, 102798.4, 
    102760.3, 102736.3, 102693.6, 102635.2, 102661.7, 102629.3, 102588.9,
  102342.6, 102533.3, 102616.3, 102700.9, 102642.5, 100799.6, 102357.2, 
    102510.2, 102610.3, 102658.8, 102647.2, 102632.2, 102625, 102604.9, 
    102582.2,
  102341.8, 102392.5, 102474.2, 102494.9, 102410.1, 99887.77, 97973.02, 
    97137.24, 99736.7, 102620.7, 102628.5, 102589.8, 102574.6, 102567, 
    102555.8,
  102092.5, 102156.6, 102341.4, 102371.6, 97347.76, 98807.98, 100613.3, 
    102245.8, 102531.8, 102584.2, 102589.6, 102552.5, 102533, 102523.3, 
    102518.3,
  101993, 102034.8, 102165.8, 102157.5, 97742.1, 98042.64, 97656.21, 
    102372.2, 102643.2, 102488, 102520.6, 102498.8, 102492.9, 102478.6, 
    102475.3,
  102973.2, 102959.1, 102950.7, 102933.2, 102903.4, 102877.4, 102826.4, 
    102778.8, 102729.1, 102674.3, 102608.5, 102542.9, 102482.5, 102444.2, 
    102414.3,
  102894, 102901.7, 102966, 102961.2, 102911.8, 102888.3, 102851.7, 102813.7, 
    102761.4, 102695.9, 102621.4, 102558.1, 102523.9, 102504.7, 102465.3,
  101026, 100791.1, 102871.8, 102975.1, 102925.3, 102903.9, 102849.8, 
    102807.9, 102752, 102693, 102633.9, 102572.3, 102552.6, 102527.1, 102495.9,
  98923.95, 99021.55, 102738.6, 102974, 102934, 102942.3, 102892, 102855.8, 
    102781, 102710.2, 102652.3, 102605.5, 102583.1, 102547.2, 102541.4,
  98892.25, 99409.5, 101365.2, 102945.9, 102925.8, 102893.1, 102860.6, 
    102828.2, 102781.2, 102727.2, 102673.5, 102644.4, 102600.3, 102583.3, 
    102562.7,
  98168.02, 99789.52, 102720.2, 102900.4, 102889.5, 102890, 102944.8, 
    102900.2, 102821.3, 102755.8, 102697.6, 102624.4, 102637.9, 102624.5, 
    102590,
  102655, 102770.8, 102844.7, 102887.5, 102868.8, 100987.4, 102537.3, 
    102647.6, 102753.4, 102765, 102733.7, 102690.2, 102667.3, 102637.4, 
    102609.1,
  102714.6, 102711.5, 102768.5, 102737, 102637.8, 100129.4, 98173.02, 
    97249.23, 99891.18, 102743.7, 102740, 102705.3, 102687.6, 102658.7, 
    102629.7,
  102581.6, 102585.2, 102693.3, 102684.4, 97667.27, 99111.37, 100910, 
    102556.6, 102758, 102744, 102730.3, 102694.9, 102683.2, 102661.2, 102635.6,
  102555.2, 102553.9, 102615.3, 102558.5, 98109.4, 98380.62, 97913.85, 
    102596.5, 102841, 102688.2, 102721.1, 102672.4, 102672.2, 102644.8, 
    102627.1,
  102524.6, 102500, 102528.3, 102526.3, 102528.2, 102531.9, 102519.1, 
    102482.4, 102432.9, 102369.4, 102312.8, 102246.4, 102194.6, 102174.1, 
    102151,
  102372.1, 102392.4, 102460.5, 102480.7, 102448.4, 102444.2, 102427.8, 
    102409.9, 102371.8, 102318.9, 102261.9, 102201.3, 102161.3, 102156.8, 
    102152.9,
  100485.8, 100298, 102320.3, 102464, 102405.2, 102387.6, 102345.7, 102321.5, 
    102284, 102237.7, 102184.9, 102148.1, 102127.7, 102122.5, 102128.3,
  98372.75, 98498.65, 102197.3, 102430.4, 102372.1, 102370.7, 102315.2, 
    102293.4, 102242.3, 102196.1, 102138.8, 102105.6, 102089.1, 102083.5, 
    102112.3,
  98339.83, 98839.98, 100823, 102393.6, 102344.6, 102286.2, 102231.2, 
    102196.1, 102154.4, 102121.4, 102083, 102066.8, 102053.5, 102074.5, 
    102093.9,
  97629.38, 99207.27, 102134.5, 102337.1, 102305.8, 102326.4, 102322.7, 
    102244.9, 102145.8, 102086.7, 102029, 101985, 102036, 102068.9, 102086.4,
  102050.6, 102174.3, 102262.5, 102329, 102269.9, 100458.1, 101962.1, 
    102008.4, 102098.6, 102042.6, 102009.9, 102004.9, 102023.9, 102054.6, 
    102086.7,
  102097.8, 102114.7, 102185.2, 102175.7, 102088.4, 99582.74, 97688.7, 
    96824.93, 99402.33, 102096.7, 102028.2, 102004.1, 102013.2, 102050.2, 
    102089,
  101966.6, 102005.6, 102134.2, 102126.6, 97198.13, 98666.53, 100417.2, 
    101930.6, 102151.3, 102122.3, 102046.1, 102009.9, 102016.4, 102047.3, 
    102092.7,
  101924.7, 101961.8, 102061.1, 102032.4, 97651.36, 97958.74, 97487.64, 
    102145.9, 102312.8, 102141.6, 102099.9, 102021.5, 102028, 102054, 102100.6,
  102389, 102470.6, 102556.1, 102624.4, 102671, 102709.8, 102726.9, 102733, 
    102713.2, 102689.5, 102653.4, 102600.2, 102547.7, 102477.1, 102409.9,
  102295.7, 102373.4, 102496.9, 102570.1, 102603.9, 102643.5, 102660.2, 
    102664.6, 102652.7, 102632.2, 102608.3, 102566.1, 102515.1, 102465.8, 
    102423.4,
  100420.2, 100281.7, 102334.1, 102532.8, 102539.4, 102573, 102575.7, 102581, 
    102576.9, 102570.1, 102544.1, 102516, 102472.9, 102432, 102387.7,
  98310.28, 98486.24, 102189, 102495.8, 102497, 102549.4, 102551.4, 102558.8, 
    102539.2, 102522.9, 102489.9, 102475.9, 102434, 102399, 102379.6,
  98284.37, 98826.2, 100811.3, 102431.5, 102459.8, 102458.9, 102472.6, 
    102475.5, 102467.8, 102462.9, 102444.5, 102429.4, 102394.2, 102379.9, 
    102352.5,
  97553.47, 99186.89, 102146.7, 102369.6, 102385.9, 102409.5, 102468.4, 
    102469, 102429.6, 102412.7, 102375.7, 102337, 102369.5, 102354.6, 102333.2,
  102021.6, 102165.2, 102264.6, 102346.1, 102335.4, 100517.8, 102061.7, 
    102207.2, 102324.5, 102363.7, 102361.9, 102332.6, 102326.6, 102315.7, 
    102298.3,
  102084.9, 102090.4, 102187.5, 102195, 102113.1, 99640.28, 97730.04, 
    96879.01, 99474.79, 102326.1, 102343.2, 102308.3, 102285.3, 102274.6, 
    102258.9,
  101926.5, 101966.6, 102117, 102126.5, 97203.8, 98657.57, 100424.6, 
    102033.4, 102252.9, 102277.8, 102276.4, 102252.8, 102238.1, 102226.7, 
    102213.7,
  101863.5, 101901.2, 102020.7, 101998.3, 97640.35, 97915.92, 97469.41, 
    102105.5, 102340.2, 102203.5, 102218.9, 102188.2, 102180.4, 102166.3, 
    102163.1,
  101800.9, 101756.1, 101799.6, 101829.4, 101880, 101912.3, 101952.9, 
    101964.5, 101973, 101977.5, 101975.6, 101991.3, 102021.7, 102039.9, 
    102041.9,
  101681.7, 101679.2, 101788.5, 101821.3, 101866.6, 101919.8, 101961, 
    101990.4, 101986.9, 101983.6, 101995.1, 102017.9, 102046.2, 102070.8, 
    102094.8,
  99839.72, 99645.41, 101639.7, 101815.7, 101834.1, 101886.2, 101926.5, 
    101970.2, 101982.5, 101998.5, 102015.2, 102033.8, 102064.4, 102090.8, 
    102105.6,
  97736.28, 97908.87, 101519, 101789.7, 101820.1, 101902.9, 101932.6, 
    101974.7, 101982.6, 102008.2, 102028.3, 102064.3, 102099.1, 102107.9, 
    102139.2,
  97665.86, 98230.27, 100188.2, 101764.1, 101793.2, 101826.6, 101903.2, 
    101958.9, 101988, 102017.7, 102053, 102096.2, 102122, 102145.9, 102166.7,
  96981.08, 98569.84, 101488.1, 101709.1, 101758.3, 101807.2, 101890.3, 
    101939.8, 101979, 102030.9, 102065.8, 102078, 102157.7, 102186.7, 102206.8,
  101304.5, 101475.3, 101623.7, 101715.1, 101708.7, 99983.99, 101553.1, 
    101734.3, 101915.3, 102002.7, 102082.3, 102137.6, 102182.8, 102222.1, 
    102227.1,
  101403.1, 101416.4, 101546.1, 101583.8, 101534.1, 99122.22, 97328.23, 
    96563.2, 99185.88, 102016.1, 102113.7, 102170.9, 102213.3, 102253, 
    102255.4,
  101223.7, 101292.8, 101500.2, 101544.1, 96739.39, 98242.15, 99995.52, 
    101596.8, 101921.7, 102040.3, 102114, 102174.3, 102233.5, 102271.8, 
    102278.9,
  101166.8, 101249.3, 101425.4, 101439.3, 97160.18, 97529.43, 97147.43, 
    101774.9, 102046.2, 102014.7, 102121.3, 102177.3, 102245.2, 102279.5, 
    102291.4,
  102096.7, 101999.6, 101924.3, 101820.4, 101721.1, 101628.9, 101544.9, 
    101481.4, 101419.9, 101369.4, 101356, 101350.4, 101379, 101424, 101456.2,
  102008.9, 101910.1, 101897.1, 101819.3, 101707.5, 101609, 101509.6, 
    101436.6, 101365, 101316.6, 101311.1, 101308, 101343.5, 101407.4, 101464.6,
  100142.9, 99795.38, 101754.8, 101820.5, 101696.8, 101581.1, 101458.6, 
    101377.7, 101308, 101253.1, 101260, 101280.4, 101315.6, 101382.3, 101451.2,
  98054.43, 98038.12, 101651.2, 101810.1, 101690.7, 101594.6, 101453.5, 
    101351, 101267.7, 101203.1, 101215.1, 101250, 101287.3, 101353.7, 101442.4,
  97969.91, 98433, 100315.7, 101791.7, 101683.7, 101541.3, 101421.7, 
    101305.4, 101219.1, 101157.4, 101173.1, 101214.6, 101261.7, 101344.4, 
    101428.7,
  97215.22, 98785.62, 101680.4, 101768.5, 101658.8, 101508.8, 101418.1, 
    101315.6, 101215.5, 101144.2, 101137.5, 101144.9, 101253.9, 101335.1, 
    101424.7,
  101726.4, 101755.6, 101803.5, 101757.9, 101639.4, 99692.63, 101064.7, 
    101055.8, 101093.5, 101068, 101112.6, 101171.9, 101246.9, 101332.4, 
    101427.5,
  101699.5, 101648.7, 101718.3, 101619.4, 101454.5, 98823.8, 96847.5, 
    95901.34, 98378.89, 101052, 101090.3, 101150.6, 101236.1, 101338.2, 
    101439.7,
  101511.1, 101504, 101639.1, 101578.2, 96574.23, 97903.85, 99551.49, 
    100974.1, 101142.9, 101094.5, 101089.2, 101150.3, 101233.2, 101347.9, 
    101454.4,
  101452.5, 101446.5, 101538.9, 101474.8, 97035.66, 97209.45, 96655.09, 
    101084.1, 101223.8, 101059, 101077.5, 101149.4, 101247.8, 101364.7, 
    101479.6,
  102425.2, 102457, 102493, 102525.9, 102584.4, 102662, 102708.4, 102725.9, 
    102725.5, 102697.7, 102653.5, 102586, 102506.1, 102406, 102291.9,
  102269.4, 102291, 102352.8, 102400.9, 102409.9, 102472, 102533.1, 102582.7, 
    102594.9, 102580.1, 102546.9, 102491.2, 102421.5, 102344.6, 102265.1,
  100367, 100145.2, 102170.1, 102336.1, 102303.3, 102333.2, 102361.5, 
    102399.7, 102430.2, 102440.1, 102423, 102382.1, 102336.4, 102269.1, 
    102196.2,
  98217, 98280.09, 102012.1, 102265.2, 102208.7, 102251.1, 102257, 102287.3, 
    102302.3, 102305.4, 102289.5, 102271.2, 102235.4, 102180.9, 102149.5,
  98155.54, 98625.16, 100613.4, 102198.1, 102166.7, 102121.1, 102131.4, 
    102139.2, 102145.7, 102164.7, 102168.9, 102166, 102137.5, 102114.6, 
    102080.4,
  97299.62, 98957.91, 101966.6, 102148.4, 102086.3, 102064.2, 102091.5, 
    102094, 102070.5, 102061.4, 102040, 102017.8, 102054.9, 102042.3, 102010.6,
  101790.9, 101940.7, 102029.5, 102087.3, 102028.7, 100143.6, 101660.7, 
    101769.5, 101875.2, 101940.5, 101954.7, 101965.7, 101975.4, 101966.5, 
    101945.6,
  101688.8, 101748.5, 101832.9, 101858.3, 101763, 99214.51, 97288.15, 
    96424.55, 99010.98, 101862.9, 101882.2, 101865.2, 101880.7, 101877, 
    101871.4,
  101412.7, 101466.1, 101636.8, 101686.7, 96684.25, 98132.87, 99921.19, 
    101534.1, 101795.8, 101830.8, 101805.6, 101781.4, 101783.4, 101788.6, 
    101788.1,
  101274.7, 101300.5, 101409.2, 101442.5, 97044.58, 97330.59, 96947.11, 
    101645.3, 101897.7, 101731.1, 101737.4, 101706.7, 101707.7, 101704, 
    101710.8,
  102783.2, 102798.7, 102856.1, 102901, 102955.2, 103020.4, 103069.8, 103103, 
    103114.6, 103111.9, 103082.1, 103046.3, 102985, 102919.8, 102832.3,
  102598.4, 102648, 102750.4, 102804.2, 102824.1, 102883.4, 102942.4, 
    103000.9, 103017.9, 103021.7, 102995.9, 102964.4, 102909, 102866, 102822,
  100606.1, 100448.6, 102518.7, 102729.4, 102713.2, 102754.7, 102778.3, 
    102835.3, 102869.4, 102895.1, 102891.2, 102875.4, 102847.4, 102807.2, 
    102770.5,
  98400.59, 98562.78, 102330.8, 102648.5, 102620.6, 102685.1, 102698.6, 
    102738.3, 102754.9, 102772.1, 102767.2, 102775.3, 102764.7, 102738.8, 
    102732.4,
  98356.41, 98867.8, 100903.7, 102551.5, 102561.9, 102545, 102571.1, 102604, 
    102623.6, 102641.2, 102645.8, 102653.8, 102653.2, 102664.3, 102659.6,
  97550.56, 99184.63, 102218.4, 102453.3, 102448.8, 102489.9, 102534.8, 
    102541.6, 102540.3, 102545.8, 102531, 102507.1, 102570.1, 102582.2, 
    102585.6,
  102126.2, 102226.2, 102303.2, 102387.4, 102356.3, 100523.4, 102095.2, 
    102245.5, 102366.7, 102437.7, 102452.3, 102465.2, 102480.7, 102497.2, 
    102511.6,
  102098, 102073.8, 102138.6, 102163.4, 102109.8, 99581.34, 97667.77, 
    96828.72, 99468.31, 102371.5, 102401.4, 102385.5, 102395.2, 102408, 
    102436.4,
  101891.6, 101897.5, 102015.6, 102031.5, 97015.99, 98535.27, 100345.9, 
    101982.9, 102269.6, 102357.4, 102342.6, 102326.1, 102325.2, 102334.2, 
    102359.5,
  101807.6, 101792.2, 101879.1, 101847.9, 97427.37, 97738.46, 97350.22, 
    102124.7, 102372.4, 102247.2, 102281.6, 102261.7, 102267.2, 102269.3, 
    102291.3,
  102676.5, 102775.6, 102863.6, 102937.8, 102988.8, 103029.2, 103046.9, 
    103049.8, 103035.6, 103026.8, 102992.9, 102946.9, 102879.9, 102829.5, 
    102778.9,
  102602.6, 102707.9, 102836.7, 102909.9, 102941.3, 102986.1, 103001.9, 
    103020.1, 102997.8, 102988.3, 102951.9, 102902.1, 102846.8, 102822.9, 
    102797.1,
  100747.4, 100603.3, 102712.8, 102911.2, 102908.3, 102937.3, 102942, 
    102941.6, 102934.1, 102933.4, 102896.8, 102867.2, 102832.8, 102811.6, 
    102782.6,
  98615.73, 98825.3, 102580.6, 102896.7, 102889.4, 102937, 102936.9, 
    102939.5, 102914, 102896.1, 102847.2, 102832.6, 102811.3, 102788.3, 
    102777.5,
  98602.94, 99169.71, 101211.9, 102848.2, 102875.4, 102877.6, 102873.9, 
    102876.2, 102870.2, 102851.5, 102835.2, 102823.5, 102790.5, 102782.1, 
    102762.6,
  97867.24, 99549.78, 102562.7, 102788.6, 102813.5, 102853, 102924.4, 
    102910.2, 102863.3, 102835.5, 102802.5, 102752, 102783.2, 102775.4, 
    102752.4,
  102359, 102553.1, 102689.6, 102773.9, 102779.8, 100953.4, 102525.3, 
    102676.5, 102784.8, 102834, 102821.9, 102797.3, 102772.9, 102760.5, 
    102743.7,
  102453, 102509.4, 102608.3, 102621.8, 102565.5, 100065.9, 98129.48, 
    97250.35, 99890.53, 102795.9, 102809, 102777.2, 102759.9, 102750.9, 
    102732.2,
  102305.1, 102373, 102517.4, 102544.3, 97566.02, 99060.01, 100866.9, 
    102504.1, 102732.8, 102762.8, 102762, 102736.6, 102747.1, 102729.6, 
    102708.6,
  102271.8, 102329.4, 102449.1, 102422.9, 98001.59, 98305.69, 97862.09, 
    102601.9, 102847.6, 102703.5, 102729.5, 102710.4, 102723.5, 102704.7, 
    102682.2,
  102308.1, 102378.7, 102444.9, 102518.7, 102609.1, 102691.3, 102747.6, 
    102789.6, 102805.7, 102811.8, 102795.4, 102771, 102723.6, 102685.9, 
    102653.2,
  102162.6, 102231.8, 102357, 102436.5, 102497.3, 102592.8, 102666.1, 
    102723.2, 102753, 102772, 102763.7, 102733.1, 102693.1, 102682.1, 102664.6,
  100242.7, 100098.6, 102160.1, 102377.7, 102409.9, 102493, 102558.9, 
    102625.3, 102670.1, 102706.2, 102715.5, 102701.6, 102680.8, 102669.3, 
    102655.3,
  98072.13, 98257.83, 101972.8, 102300.3, 102339, 102436, 102497.2, 102560.8, 
    102600.5, 102635.6, 102647.7, 102658, 102647.3, 102647.5, 102651.4,
  97967.23, 98540.93, 100572.5, 102207.6, 102271.4, 102320.2, 102400.5, 
    102461.4, 102508.1, 102561.1, 102585.5, 102616.6, 102610.9, 102636.8, 
    102641.5,
  97187.7, 98861.31, 101871.1, 102124.1, 102191.2, 102247.8, 102353.3, 
    102415.1, 102451.8, 102497.6, 102514.9, 102520.7, 102588.2, 102619.6, 
    102627.1,
  101587, 101814.1, 101968.6, 102075.2, 102121.5, 100400.2, 101976.7, 
    102144.9, 102307.2, 102399.8, 102476.4, 102523.5, 102566.4, 102601, 
    102625.2,
  101637.5, 101720.3, 101845.5, 101921.2, 101907.7, 99470.23, 97663.79, 
    96880.59, 99518.16, 102367.2, 102432.8, 102480.2, 102534.6, 102587.8, 
    102616.8,
  101441.9, 101559.1, 101762.9, 101828.8, 97021.79, 98548.63, 100315.9, 
    101928.2, 102250.9, 102352.6, 102385, 102437.5, 102509.1, 102568.3, 
    102599.3,
  101363.4, 101482.5, 101660.5, 101703.7, 97433.73, 97782.16, 97424.29, 
    102116.6, 102362.5, 102292.6, 102354.2, 102403.1, 102486.4, 102549.8, 
    102584.7,
  102693.1, 102743.6, 102806, 102860.9, 102925.4, 102981.7, 103018.3, 
    103048.7, 103063.7, 103076.3, 103058.6, 103029.8, 102967.5, 102902.3, 
    102847.5,
  102592.1, 102658.7, 102775.5, 102821.5, 102861.3, 102936.4, 102994, 
    103037.1, 103051, 103053.7, 103039.3, 103012.8, 102965.4, 102936.4, 
    102889.7,
  100716, 100560.4, 102629, 102805.6, 102808, 102857.9, 102898.1, 102947.9, 
    102976.4, 103002.8, 102998, 102993.4, 102969.3, 102940, 102893.6,
  98564.48, 98774.83, 102491.4, 102796.2, 102772.8, 102842.5, 102874.5, 
    102918, 102938.2, 102947.9, 102947, 102955, 102939.5, 102917.5, 102910,
  98530.59, 99091.66, 101107.3, 102743.1, 102768.4, 102755.4, 102789.8, 
    102831.3, 102855.2, 102893.4, 102892.8, 102910.7, 102902.2, 102905.9, 
    102895.7,
  97764.05, 99438.57, 102451.5, 102682.7, 102711.5, 102742.9, 102805.5, 
    102809.8, 102804.2, 102823.9, 102828, 102811, 102874.4, 102883.7, 102881.3,
  102231.6, 102415, 102559, 102661.7, 102674, 100837.9, 102397.7, 102553.2, 
    102682.5, 102746.2, 102770.6, 102800.8, 102828, 102847.7, 102858.5,
  102290.7, 102355.6, 102468.1, 102514.2, 102457, 99973.24, 98065.46, 
    97234.59, 99856.26, 102718.8, 102745.4, 102752.3, 102771.3, 102801, 
    102822.2,
  102109.4, 102190.5, 102380.8, 102435.3, 97489.63, 98983.46, 100772.2, 
    102376.1, 102624.4, 102703.4, 102698.2, 102697.3, 102710.6, 102745.1, 
    102772.2,
  102028.3, 102112.2, 102266.5, 102296.3, 97915.2, 98223.12, 97809.91, 
    102533, 102776.6, 102645.8, 102662.4, 102648.9, 102661.1, 102686.9, 
    102718.2,
  102318.2, 102368.8, 102456.4, 102517, 102570.8, 102578.5, 102556.2, 102560, 
    102576.1, 102597.2, 102605.5, 102611.2, 102610.5, 102608.2, 102579.9,
  102215.9, 102299.7, 102425.9, 102509, 102564.4, 102619, 102602.5, 102609.5, 
    102609.1, 102623.9, 102630, 102633.2, 102638.6, 102633.4, 102624.5,
  100379.4, 100259, 102297.8, 102499.4, 102536.8, 102602.8, 102609.3, 
    102609.4, 102618.4, 102636.4, 102656.9, 102661.7, 102672, 102667.6, 
    102647.4,
  98286.11, 98504.23, 102158.1, 102474.6, 102509.8, 102607.5, 102635.8, 
    102630.2, 102633.3, 102650.9, 102660.9, 102683.8, 102688.1, 102681.4, 
    102679.5,
  98249.81, 98817.41, 100817.2, 102427.7, 102485.2, 102518, 102590.4, 
    102608.2, 102617.5, 102648, 102665, 102694.1, 102705.8, 102717.4, 102704.2,
  97563.62, 99166.62, 102121.5, 102361.7, 102445.3, 102500.1, 102584, 
    102615.6, 102617.9, 102639.3, 102651, 102645.3, 102722.4, 102738.8, 102733,
  101909.5, 102107.4, 102258.6, 102371.6, 102387.9, 100642.3, 102216.1, 
    102375.4, 102524, 102594.4, 102651.7, 102683.5, 102723.5, 102749.8, 
    102756.3,
  102040.4, 102069.7, 102197.4, 102236.6, 102225.4, 99791.98, 97943.59, 
    97145.54, 99766.88, 102601.3, 102651.4, 102675.5, 102715.8, 102753.9, 
    102768.7,
  101893.2, 101960.4, 102154.9, 102206.9, 97365.3, 98869.42, 100649.1, 
    102244, 102519.9, 102607.4, 102651.4, 102670.4, 102704.9, 102746.5, 
    102767.4,
  101854.9, 101930.5, 102081.2, 102097.6, 97806.02, 98152.8, 97756.5, 
    102393.8, 102646.9, 102572.2, 102645.5, 102657.4, 102702.5, 102737.4, 
    102767.8,
  102306.4, 102237.3, 102211.3, 102176.7, 102150.3, 102134.8, 102132.9, 
    102107.4, 102091.9, 102084.3, 102070.5, 102080, 102098.4, 102121.6, 
    102118.6,
  102119.6, 102100.8, 102142.4, 102133.1, 102074.5, 102057.6, 102064.3, 
    102068.2, 102059.7, 102058.2, 102046, 102058.5, 102084.7, 102124.1, 
    102154.6,
  100204.2, 99981.81, 101930.9, 102084.9, 102021.6, 102001.5, 101994, 
    102005.8, 102006.3, 102016.8, 102026.4, 102056.5, 102098.3, 102136.1, 
    102168.9,
  98070.92, 98169.84, 101755.3, 101999.8, 101966.4, 101962.9, 101948.6, 
    101966.6, 101967.9, 101982.9, 101998.3, 102040, 102089.5, 102124.6, 
    102183.5,
  97942.13, 98468.62, 100384.4, 101915.8, 101905.4, 101870.6, 101882.3, 
    101900.1, 101912.9, 101946, 101978.5, 102038.2, 102092.2, 102146.7, 
    102196.2,
  97233.76, 98789.33, 101674, 101832.5, 101837.6, 101808.4, 101851.3, 
    101884.5, 101891.7, 101930.6, 101955.2, 101988, 102098.9, 102158.3, 
    102207.1,
  101605, 101706.4, 101771.4, 101799.4, 101766, 99992.74, 101469.1, 101608.6, 
    101765, 101865.2, 101950.4, 102029.9, 102107.9, 102165.7, 102217.4,
  101653.5, 101610.6, 101682, 101646, 101565, 99092.83, 97260.4, 96488.09, 
    99047.03, 101833, 101939.1, 102018.9, 102099.5, 102168.5, 102228.9,
  101497, 101481.6, 101610.3, 101566.4, 96747.79, 98182.41, 99855.74, 
    101393.5, 101700.2, 101833, 101912.5, 102002.1, 102091.9, 102168.5, 
    102233.9,
  101451.1, 101445.2, 101530.5, 101456.5, 97146.43, 97444.73, 97045.88, 
    101589.9, 101838.8, 101801.1, 101903.5, 101983, 102085, 102167.8, 102242.7,
  103469.3, 103428.9, 103432.8, 103408, 103371.4, 103323.9, 103272.6, 
    103203.4, 103119.2, 103009.3, 102893.9, 102763.1, 102614.8, 102467.7, 
    102357.9,
  103315.5, 103293.6, 103380.8, 103381.8, 103323, 103279.2, 103219.9, 
    103158.3, 103084.9, 102983.7, 102871.7, 102719.6, 102589, 102496.2, 
    102409.6,
  101336.7, 101099.9, 103164.5, 103334.7, 103275.2, 103230.6, 103159, 
    103087.8, 103009.8, 102928.2, 102820.5, 102706, 102590, 102487.8, 102400.8,
  99160.23, 99230.77, 102939.3, 103244.2, 103188.1, 103179.8, 103122.3, 
    103058.8, 102979.7, 102887.8, 102785.4, 102687.8, 102579.6, 102483.1, 
    102416.7,
  99032.63, 99553.64, 101532.5, 103144.5, 103117.8, 103063, 103016.9, 
    102955.4, 102894.6, 102828.6, 102760.3, 102671.9, 102579.5, 102491.1, 
    102421.6,
  98203.17, 99854.27, 102839.7, 103053.9, 103012.5, 102993.1, 103007.1, 
    102968.1, 102875.5, 102806.4, 102707.8, 102609.3, 102580.1, 102502.4, 
    102430.6,
  102749, 102871.1, 102932, 102988, 102924.1, 101031, 102531, 102661.1, 
    102743.8, 102774.5, 102732.3, 102651.4, 102560.1, 102486.2, 102419.7,
  102679.2, 102674.6, 102761.9, 102755.3, 102653.3, 100106.4, 98147.38, 
    97238.23, 99798.37, 102667, 102676.5, 102607.1, 102528, 102464.1, 102402.6,
  102512.9, 102514.7, 102630.1, 102629.2, 97591.94, 98988.66, 100771.8, 
    102392.7, 102628.5, 102639.1, 102607.9, 102546.6, 102484.6, 102429.7, 
    102382.8,
  102404, 102407.5, 102468, 102419.2, 97964.51, 98212.09, 97790.87, 102443.1, 
    102718.3, 102545.7, 102547.8, 102490.5, 102453.5, 102398.4, 102359.6,
  103666.2, 103633.4, 103637.4, 103614.8, 103569.3, 103527.5, 103466.9, 
    103401.5, 103290.8, 103199.3, 103064.2, 102888.7, 102730.1, 102629.4, 
    102538.8,
  103526.6, 103505.9, 103589.4, 103585.8, 103532.8, 103500.8, 103435.4, 
    103373.8, 103279.9, 103177.5, 103033.4, 102916.8, 102789.2, 102680.1, 
    102592.4,
  101591.8, 101356.4, 103417.6, 103567.8, 103503.4, 103469.3, 103390.2, 
    103321.4, 103229.9, 103146.8, 103024.8, 102908.4, 102791.1, 102709.7, 
    102622.7,
  99419.84, 99486.09, 103227.7, 103502.7, 103443.6, 103444.2, 103378.1, 
    103311.5, 103212.1, 103110, 103006.6, 102938.7, 102828.2, 102733.6, 
    102660.9,
  99334.94, 99832.34, 101820.3, 103421.2, 103392.2, 103346.6, 103302.1, 
    103235.9, 103165.8, 103099.9, 103015.2, 102956, 102859.9, 102772.2, 
    102696.5,
  98520.41, 100130.3, 103125.5, 103322, 103303.4, 103279.2, 103315, 103266.2, 
    103185.5, 103107.3, 103023.6, 102930.9, 102886.4, 102823.7, 102730.8,
  103060.2, 103157.9, 103222.2, 103281, 103232.3, 101344.8, 102878.2, 
    102992.4, 103098.2, 103104.5, 103065.7, 102973.9, 102897, 102832.9, 
    102766.2,
  103006.8, 103016.4, 103091.1, 103082.1, 102988.8, 100444.9, 98488.74, 
    97568.56, 100184.2, 103030.5, 103037.9, 102954.7, 102901.3, 102849.9, 
    102789.9,
  102900.1, 102902.8, 103015.3, 103001.8, 97971.09, 99436.07, 101236.5, 
    102825.9, 103043.7, 103043.1, 103012.4, 102933.2, 102901.2, 102855.1, 
    102799.6,
  102919.3, 102877.9, 102916.3, 102878, 98429.39, 98702.27, 98201.79, 
    102882.7, 103098.4, 102963.3, 102971.4, 102924.4, 102910.5, 102859.2, 
    102804.9,
  103577.7, 103556.2, 103548.2, 103513.4, 103460.7, 103417.1, 103340.4, 
    103261.7, 103167.3, 103056.4, 102897.4, 102719, 102560, 102401.6, 102298.3,
  103464.1, 103443.8, 103532.3, 103510.7, 103443.9, 103394.9, 103314.8, 
    103239.8, 103145.5, 103044.6, 102903.7, 102750.4, 102629.5, 102475.9, 
    102340.6,
  101553, 101274.4, 103366.5, 103484.3, 103410.8, 103361.8, 103277.2, 103199, 
    103108.6, 103008.5, 102883.9, 102754.7, 102642, 102518.5, 102392.5,
  99397.53, 99455.83, 103168.4, 103431.3, 103363.5, 103345.5, 103274.5, 
    103201.9, 103106.9, 102999.2, 102900.3, 102799.7, 102690.4, 102564.6, 
    102451.9,
  99305.48, 99814.96, 101756.8, 103357.6, 103309.7, 103270.5, 103208.2, 
    103151.5, 103082.8, 102997.3, 102905.8, 102818.6, 102713.7, 102612, 
    102505.8,
  98497.59, 100133.8, 103073.1, 103283.3, 103229.7, 103211.1, 103238, 
    103196.4, 103117, 103026.3, 102932.2, 102809, 102747.9, 102670, 102554.7,
  103009.8, 103125.3, 103183.1, 103230.7, 103178.3, 101290.9, 102818.2, 
    102950.6, 103049.8, 103028.5, 102975, 102873.1, 102776.1, 102693.4, 102603,
  103009.2, 103007.5, 103077.9, 103052.3, 102941.7, 100407, 98448.4, 
    97512.74, 100117.8, 102971.3, 102947.1, 102866.1, 102790.8, 102720.5, 
    102632.7,
  102855, 102859.7, 102980.5, 102983.6, 97955.94, 99383.16, 101183.9, 
    102805.2, 102994.2, 102970.5, 102909.2, 102844.8, 102780.1, 102737.2, 
    102674.5,
  102812.9, 102801.9, 102875.1, 102831.5, 98403.24, 98659.67, 98164.49, 
    102832, 103053.7, 102901.4, 102897, 102833.2, 102785.7, 102750.7, 102699.6,
  103252.5, 103214, 103171.5, 103094.6, 103010.2, 102940.7, 102854.2, 
    102764.6, 102642.3, 102522.7, 102296.2, 102132.4, 101967.3, 101821.9, 
    101713.5,
  103183, 103121.6, 103174, 103116.8, 103014.1, 102933.2, 102831.4, 102738.8, 
    102604, 102471.8, 102302.9, 102152.2, 101990.2, 101825.5, 101713.5,
  101294.4, 100987.4, 103033.6, 103097.3, 102984.2, 102915.7, 102802.4, 
    102703.3, 102576.8, 102447, 102278, 102133.4, 101993, 101837.3, 101697.2,
  99194.51, 99233.95, 102883.3, 103085.5, 102970.2, 102924.7, 102813.7, 
    102716.3, 102576.5, 102464.5, 102341.1, 102186.4, 102026.4, 101868.6, 
    101716.4,
  99138.48, 99617.53, 101514.5, 103040.6, 102953.7, 102876.3, 102801.9, 
    102712.7, 102594.3, 102521.5, 102393.1, 102229.4, 102050.4, 101907.9, 
    101725.5,
  98419.11, 99974.73, 102866.9, 103005.7, 102908.9, 102844.6, 102859.2, 
    102775.8, 102655.1, 102582.9, 102446.8, 102246.5, 102131.7, 101982.5, 
    101767,
  103010.6, 103016.3, 103015.7, 102993.3, 102911.3, 100984.1, 102470.4, 
    102534.2, 102603, 102571.5, 102485.4, 102328.4, 102174.5, 102047.6, 
    101855.3,
  103069.8, 102979.1, 102988.6, 102886.5, 102716.9, 100138.3, 98147.53, 
    97157.77, 99731.7, 102547.8, 102499, 102360.8, 102219.7, 102103.5, 
    101945.1,
  102946.3, 102892.7, 102930.8, 102863.4, 97782.67, 99163.27, 100925.6, 
    102502.7, 102648.1, 102582.5, 102494, 102383, 102250.1, 102141.5, 102010.3,
  102896, 102848.6, 102871.4, 102751.7, 98268.17, 98475.06, 97931.23, 
    102526.1, 102710.5, 102545, 102516.3, 102410.8, 102301.6, 102189.2, 
    102076.8,
  102825.7, 102810, 102791.3, 102747.2, 102706.1, 102672.8, 102627.2, 
    102566.3, 102484, 102409.3, 102304.4, 102192.6, 102060.4, 101928.6, 
    101782.6,
  102759.4, 102696.9, 102767.4, 102739.3, 102678.9, 102626, 102561.3, 102498, 
    102419.4, 102333.8, 102214.6, 102105.3, 101972.2, 101864.6, 101781.5,
  100858.2, 100567.4, 102614.8, 102701.2, 102632.6, 102582.6, 102501, 
    102419.4, 102332.9, 102237, 102133.7, 102037.1, 101925.5, 101826.6, 
    101724.3,
  98721.86, 98806.88, 102452.3, 102654.9, 102583.7, 102552.8, 102468.1, 
    102394.1, 102293.5, 102189.3, 102074.8, 101982.1, 101868.6, 101767.6, 
    101684.5,
  98750.64, 99200.21, 101079, 102618.5, 102561.6, 102486.1, 102413.7, 
    102334.7, 102237.5, 102148.8, 102038.4, 101932.5, 101818.6, 101721.5, 
    101630.3,
  98027.71, 99608.22, 102506.5, 102586.4, 102509.9, 102420.8, 102447.4, 
    102362.4, 102249.6, 102155.7, 102013.8, 101865.8, 101791.7, 101688.1, 
    101588.3,
  102600.5, 102651.4, 102636.9, 102574.3, 102536.6, 100575.9, 102091.7, 
    102094.4, 102145.4, 102098.4, 102033.4, 101898.5, 101769.1, 101665, 
    101560.5,
  102626.7, 102622.3, 102617.1, 102542.8, 102321.5, 99740.06, 97731.23, 
    96736.11, 99353.56, 102127.2, 102042.9, 101896.5, 101757.5, 101643.3, 
    101536.3,
  102580.6, 102579.7, 102599.4, 102532.9, 97384.55, 98862.77, 100548.6, 
    102121.4, 102233.5, 102116.5, 102004.5, 101877.9, 101750.1, 101629.6, 
    101506.1,
  102545.7, 102544.3, 102560.3, 102476.7, 97959.75, 98179.99, 97530.97, 
    102162.1, 102256.1, 102073.7, 101998.8, 101863.3, 101733, 101613.3, 
    101478.1,
  102015.5, 102093.6, 102169.1, 102240.9, 102307.3, 102353.4, 102389.2, 
    102403.5, 102391.6, 102363, 102314.3, 102253.5, 102194.6, 102140.5, 
    102068.6,
  101934.5, 102000.9, 102137.2, 102206, 102252.1, 102313.4, 102336.8, 
    102358.5, 102343.4, 102325.1, 102276.4, 102211.1, 102162.6, 102103.3, 
    102061.2,
  100106.6, 99950.26, 102012.3, 102205.6, 102222.2, 102268.8, 102278, 
    102278.5, 102274.9, 102248.3, 102209.3, 102161.3, 102124.5, 102082.5, 
    102035.7,
  97991.14, 98206.62, 101877.2, 102167.8, 102189.4, 102246.9, 102260.8, 
    102259.6, 102241.7, 102211, 102162.9, 102138.1, 102094.6, 102048.5, 
    102016.6,
  97980.48, 98536.44, 100532.3, 102117.8, 102159.3, 102171.5, 102196.5, 
    102194.6, 102178.7, 102162.8, 102136.7, 102108.3, 102070.9, 102031.3, 
    101992.5,
  97336.16, 98916.42, 101874.2, 102069, 102108.4, 102120.3, 102204.9, 
    102210.5, 102172.6, 102150.4, 102101.5, 102050.2, 102067.7, 102027.6, 
    101974.1,
  101728.8, 101884, 102014.6, 102073.8, 102104.2, 100303, 101838.9, 101968.8, 
    102098.7, 102122.4, 102115.6, 102082, 102045, 102004.7, 101950.4,
  101852, 101899.4, 101983.1, 102003.5, 101922.8, 99453.84, 97545.01, 
    96694.69, 99296.84, 102107.1, 102119.9, 102075.9, 102032.4, 101990.9, 
    101932.3,
  101785.5, 101854.5, 101983.3, 101996.8, 97082.77, 98577.7, 100301.6, 
    101890.1, 102076.9, 102096.6, 102076.1, 102044.1, 102016.1, 101973.5, 
    101918.5,
  101806.1, 101870.9, 101975.8, 101966.9, 97580.55, 97874.42, 97353.74, 
    101998.1, 102178.2, 102071.2, 102073.1, 102034.8, 102011.6, 101952.8, 
    101895.4,
  102160.4, 102195.5, 102221, 102241.5, 102291, 102350.6, 102404.3, 102436.2, 
    102450.9, 102450.6, 102431.6, 102405.4, 102360, 102319.7, 102268.4,
  102003.4, 102024.7, 102140.1, 102165.9, 102187.3, 102231.4, 102287.1, 
    102333.7, 102363.5, 102375.5, 102364.7, 102342.7, 102308.2, 102277, 102255,
  100055.3, 99865.23, 101911, 102089.9, 102083.5, 102131.4, 102169.1, 
    102216.3, 102252.6, 102283.6, 102289.4, 102277.9, 102260.2, 102241.2, 
    102218.5,
  97865.65, 98010.59, 101699.6, 101996.5, 102001.5, 102055.2, 102094, 
    102133.3, 102162.9, 102191.7, 102198.5, 102203.3, 102195.1, 102182.8, 
    102183.7,
  97764.62, 98290.21, 100282, 101874.8, 101918.9, 101933.1, 101984, 102017.6, 
    102054.7, 102092.8, 102118.3, 102134.7, 102129.7, 102147.7, 102142.9,
  96968.59, 98581.77, 101555.4, 101770.8, 101812.9, 101830.5, 101929.5, 
    101972.6, 101989.4, 102016.2, 102028.8, 102027.8, 102091, 102105.9, 
    102104.6,
  101349.5, 101502.1, 101633.5, 101699, 101730.9, 99971.58, 101525.8, 
    101673.7, 101822.4, 101903.1, 101971.5, 102007.7, 102042.4, 102066.8, 
    102075.1,
  101335.6, 101394, 101503.3, 101545.2, 101505.6, 99026.55, 97206.69, 
    96410.95, 99028, 101840.7, 101909.9, 101951.7, 101992.8, 102024.3, 
    102043.6,
  101137.4, 101227.7, 101415.2, 101449.2, 96614.23, 98107.38, 99831.09, 
    101421, 101715.4, 101816.6, 101850, 101897, 101944.4, 101985.5, 102015.8,
  101078.5, 101159.1, 101314.1, 101353.7, 97029.48, 97333.59, 96909.84, 
    101552.7, 101793.5, 101743.3, 101800.7, 101849, 101903.6, 101953.9, 
    101983.4,
  101983.5, 102077.1, 102197.8, 102320, 102417, 102495.3, 102550.5, 102593, 
    102608.4, 102618.5, 102609.5, 102586.7, 102551.1, 102516, 102470.3,
  101876.4, 101972.8, 102142.1, 102271.2, 102360.8, 102453.6, 102509.1, 
    102553.4, 102577.9, 102587, 102572, 102545, 102518, 102500.5, 102482.3,
  100040.9, 99922.94, 101984.2, 102226.5, 102299.3, 102394.5, 102442.6, 
    102478.5, 102502, 102515.2, 102517, 102506, 102491.9, 102468.6, 102455.9,
  97932.16, 98149.02, 101819.7, 102179.5, 102252.5, 102370.1, 102425.3, 
    102463.7, 102470.6, 102470.8, 102460.7, 102459.4, 102431.2, 102421.6, 
    102431.4,
  97929.08, 98475.59, 100468.6, 102109.6, 102197.6, 102267.8, 102337.6, 
    102381.4, 102403.7, 102422.2, 102425.5, 102423.9, 102406.4, 102404.3, 
    102392.9,
  97183.66, 98818.3, 101778.3, 102043.8, 102136, 102209.5, 102340.1, 
    102385.4, 102389.5, 102393.2, 102374.7, 102342.4, 102391.5, 102388.8, 
    102371.3,
  101632.7, 101795.2, 101922.8, 102024.2, 102079.6, 100339.1, 101904.6, 
    102099.2, 102266.1, 102345.1, 102368.1, 102365.7, 102362, 102356.8, 
    102347.9,
  101708.4, 101738.8, 101848.7, 101883.7, 101878.3, 99460.66, 97629.39, 
    96807.71, 99425.73, 102301, 102346.7, 102344.2, 102330.1, 102326.1, 
    102321.2,
  101546.3, 101608.4, 101786.6, 101834.6, 96979.89, 98469.02, 100259, 
    101904.3, 102193.5, 102268, 102291.2, 102290.2, 102286.3, 102289, 102286.5,
  101497.2, 101543.6, 101682.7, 101693, 97380.91, 97726.12, 97347.95, 
    102014.6, 102305.8, 102206.2, 102256, 102234.2, 102247.5, 102248.9, 
    102255.8,
  101957.5, 101914.4, 101906.9, 101909.3, 101939.1, 101967.1, 102000.7, 
    102030.8, 102074.9, 102127.3, 102171.6, 102204.2, 102212.7, 102233.4, 
    102252.8,
  101862.9, 101804.3, 101866.3, 101874.7, 101884.5, 101928.9, 101971.1, 
    102007.3, 102047, 102095, 102134.5, 102163.8, 102181, 102222.4, 102265.8,
  99964.06, 99702.98, 101681.1, 101826, 101820.8, 101862.1, 101903, 101956.2, 
    102006.2, 102060.4, 102108.4, 102141.5, 102172.6, 102203, 102247.1,
  97852.81, 97929.32, 101515.4, 101765.2, 101756.1, 101829.2, 101871.2, 
    101920.8, 101967.9, 102014.8, 102067.9, 102110.6, 102145.3, 102178.2, 
    102243.6,
  97775.79, 98270.53, 100143.2, 101701.2, 101693.7, 101713.1, 101787.5, 
    101849.5, 101912.9, 101971.1, 102028.6, 102085.9, 102114.3, 102178.9, 
    102223.6,
  97038.51, 98617.12, 101449.3, 101620.8, 101617.7, 101642.8, 101736.9, 
    101803.7, 101853.2, 101921.3, 101973.3, 102006, 102108.1, 102177.3, 
    102213.4,
  101465.1, 101530.2, 101579.2, 101609, 101551.6, 99788.07, 101338.5, 
    101518.8, 101714.3, 101834.3, 101940.8, 102021.8, 102096.9, 102162.4, 
    102201.4,
  101556.2, 101506.9, 101524, 101469.1, 101371.6, 98903.75, 97092.69, 
    96335.8, 98933.72, 101777.8, 101892.5, 101988.7, 102068.4, 102140.6, 
    102199.9,
  101381.3, 101398.2, 101489.1, 101451.2, 96558.8, 97978.7, 99675.34, 
    101264.8, 101611.4, 101759.7, 101848.9, 101947, 102033.1, 102116, 102180.6,
  101341.1, 101354.9, 101438.1, 101356.9, 97002.39, 97277.08, 96860.55, 
    101403.6, 101699.2, 101694, 101813.7, 101900.4, 101997.2, 102083, 102160.8,
  102416.5, 102412, 102447.6, 102460.7, 102476.9, 102486.8, 102478.9, 102462, 
    102429.7, 102401.3, 102374.3, 102336.7, 102301.8, 102266.5, 102238,
  102288, 102314.9, 102412.9, 102437.8, 102426.8, 102439.6, 102437.1, 
    102431.1, 102408.1, 102373.2, 102340.1, 102298.5, 102266.3, 102243.4, 
    102241.8,
  100354.9, 100176.8, 102202.4, 102390.7, 102360.3, 102374.8, 102356.8, 
    102345.6, 102332.1, 102315.3, 102288.2, 102262.4, 102234.5, 102213.7, 
    102208.8,
  98196.27, 98332.69, 101999.6, 102331.4, 102306.5, 102350.8, 102345, 
    102332.1, 102301.2, 102273.6, 102240.4, 102226, 102196, 102175.6, 102190.5,
  98138.52, 98648.62, 100599.9, 102213.5, 102244.5, 102232.3, 102239.7, 
    102237.2, 102225.5, 102217.1, 102192.2, 102182.8, 102154.6, 102158.7, 
    102163.2,
  97320.46, 98942.71, 101893, 102107.6, 102128.7, 102156.6, 102219.1, 
    102219.6, 102184.8, 102169.9, 102129.8, 102092.3, 102130.5, 102138.2, 
    102140.9,
  101796.4, 101903.8, 101982.8, 102050, 102035.4, 100221.6, 101746.4, 
    101908.8, 102024.8, 102089.4, 102101.9, 102095.9, 102095.9, 102105, 102115,
  101787, 101785, 101860.1, 101852.4, 101788.1, 99304.41, 97422.92, 96591.78, 
    99164.74, 102025.1, 102059.2, 102063.1, 102059.3, 102069.3, 102086.8,
  101613.7, 101632.9, 101748.9, 101764.1, 96825.27, 98240.7, 99996.4, 
    101600.4, 101880.7, 101949.9, 101978.1, 101991.1, 102005.5, 102022.1, 
    102046.2,
  101585.2, 101547.3, 101621.7, 101595, 97219.58, 97496.59, 97095.09, 
    101698.9, 101976.2, 101860.2, 101910.3, 101906.8, 101934.5, 101956.6, 
    101996,
  102911.9, 102837.6, 102839.2, 102823.4, 102767.8, 102734.1, 102660.5, 
    102605.2, 102572.7, 102543.2, 102516.3, 102481.8, 102463.7, 102440.6, 
    102407.5,
  102777.2, 102773.1, 102860.2, 102849.6, 102799.3, 102760.4, 102711.8, 
    102670.9, 102629.1, 102583.5, 102543.7, 102511.9, 102486, 102463.2, 
    102444.7,
  100872.2, 100642.8, 102667.2, 102822.9, 102763.7, 102752.3, 102701.1, 
    102647.2, 102611.2, 102577, 102542.7, 102516.8, 102492.5, 102473.9, 
    102446.6,
  98723.41, 98835.95, 102484.4, 102794.2, 102738.9, 102759.3, 102728, 102694, 
    102645.3, 102599.8, 102555.9, 102532.7, 102506.2, 102478.6, 102471,
  98646.26, 99164.31, 101100.3, 102692.6, 102689.9, 102664.2, 102650.3, 
    102638.5, 102612.5, 102591, 102561.8, 102548.1, 102507.5, 102490, 102476.4,
  97840.3, 99477.31, 102395.5, 102614.5, 102591, 102606.9, 102665.8, 
    102648.2, 102599.7, 102572.6, 102528.6, 102491.3, 102519.6, 102510.1, 
    102489.4,
  102350.7, 102452.6, 102513.4, 102565.4, 102528.4, 100655.2, 102191.4, 
    102367.2, 102489, 102545.8, 102538.1, 102519.6, 102505.9, 102499, 102483.4,
  102341.4, 102327.4, 102397.9, 102372.8, 102272.5, 99782.89, 97859.74, 
    97016.89, 99609.59, 102495.7, 102525, 102515.6, 102498.4, 102485.2, 
    102480.1,
  102206.1, 102204.9, 102297.1, 102290.1, 97302.91, 98704.75, 100473.3, 
    102092, 102360.6, 102422.4, 102450.7, 102451, 102454.6, 102455.1, 102455.6,
  102132.7, 102143, 102187.5, 102124.1, 97700.59, 97961.16, 97539.48, 
    102179.6, 102454.1, 102331.5, 102397.9, 102383.1, 102403.9, 102408.8, 
    102420.3,
  103014.1, 102950.1, 102887.5, 102847.3, 102801.8, 102665.4, 102484.1, 
    102305.6, 102189.1, 102137, 102173.2, 102221.8, 102271.2, 102296.3, 
    102292.4,
  102909, 102873.6, 102915.7, 102868.7, 102817.3, 102747.7, 102636, 102452.1, 
    102270.2, 102174.5, 102184.2, 102219.4, 102281.5, 102316.5, 102334.8,
  101043.2, 100761.2, 102778.2, 102859.5, 102812.2, 102765, 102650.9, 102505, 
    102421.5, 102225.4, 102190.7, 102247.9, 102303.4, 102340.2, 102352.2,
  98959.31, 98994.24, 102636.7, 102865.2, 102796.8, 102812, 102735.4, 
    102606.8, 102468.7, 102302.2, 102221.9, 102274.6, 102322.4, 102347.4, 
    102388.5,
  98877.7, 99381.35, 101285.3, 102834.2, 102784.6, 102753, 102731.4, 
    102640.9, 102538.4, 102410.7, 102306.5, 102293.7, 102340.2, 102379.5, 
    102416.3,
  98139.38, 99733.58, 102612.6, 102790.5, 102744.7, 102735.9, 102791.3, 
    102754.5, 102616.9, 102489.9, 102346.6, 102300.8, 102379.2, 102415.5, 
    102440.3,
  102637.4, 102706.2, 102757.8, 102788.3, 102709.4, 100843, 102374.1, 
    102495.8, 102557, 102541.4, 102456.3, 102390, 102413.9, 102444.8, 102458.1,
  102646, 102635.4, 102682.9, 102633, 102520.7, 100009.1, 98070.52, 97170.6, 
    99760.52, 102573.8, 102549.3, 102471.6, 102458.9, 102480.9, 102484.3,
  102545.9, 102543, 102621.8, 102602.6, 97600.61, 99003.73, 100791.6, 102393, 
    102592.9, 102569.6, 102566.5, 102523.3, 102497.5, 102507.2, 102510.3,
  102523, 102503.2, 102548.2, 102480, 98046.23, 98293.27, 97838.29, 102484.6, 
    102714.6, 102553.2, 102572.9, 102528.5, 102533.6, 102525.4, 102529.8,
  103086.6, 103087.5, 103111.2, 103093.9, 103076.7, 103036.4, 102984.5, 
    102896.3, 102806.1, 102709.5, 102602.8, 102518.8, 102450.7, 102400.1, 
    102357.6,
  102965.1, 102969, 103067.1, 103066, 103032.2, 102992.5, 102944.1, 102861.1, 
    102777.5, 102676.3, 102568.2, 102473.6, 102407.9, 102372.9, 102364.7,
  101057.7, 100851.2, 102890.8, 103040.7, 102986.7, 102946.7, 102891.9, 
    102793.6, 102719.2, 102632.8, 102522.7, 102441.6, 102383.7, 102355.5, 
    102344.4,
  98926.59, 99040.34, 102707.5, 102987, 102930.9, 102927.4, 102880.4, 
    102796.7, 102704.7, 102589, 102480.5, 102409.8, 102355.2, 102325, 102333.1,
  98854.82, 99394.66, 101327.9, 102909.8, 102884.5, 102833.7, 102811.4, 
    102743.6, 102650.5, 102552.6, 102450.1, 102380.8, 102333.6, 102319.8, 
    102319.7,
  98094.81, 99716.87, 102628.7, 102832.9, 102799.8, 102775.1, 102818.3, 
    102789.1, 102672.6, 102561.6, 102428.3, 102309.2, 102326.8, 102309.8, 
    102311,
  102562.6, 102680, 102754.1, 102805.3, 102742.8, 100879.1, 102380.3, 
    102532.1, 102558.5, 102529.5, 102417.2, 102318.8, 102290.7, 102282.2, 
    102291.6,
  102587, 102598.7, 102662.4, 102634.9, 102515.7, 100000.9, 98077.01, 
    97198.79, 99729.16, 102531.4, 102422.9, 102287.4, 102251.6, 102249.3, 
    102264.5,
  102444.7, 102463.6, 102578, 102574.2, 97593.58, 98995.1, 100772.6, 
    102385.7, 102599.8, 102511.2, 102418.6, 102278, 102213.7, 102213.8, 
    102235.6,
  102393.1, 102415, 102499.7, 102451, 98035.95, 98286.53, 97800.45, 102470.7, 
    102692.2, 102475.4, 102426.1, 102272.3, 102196.5, 102183.3, 102206,
  102787.8, 102849.5, 102923.2, 102998.9, 103054.7, 103090.5, 103091.8, 
    103059.1, 103009, 102954.5, 102904.1, 102807.1, 102727.5, 102660.6, 
    102574.3,
  102695.5, 102750.3, 102881, 102940.6, 102978.9, 103034.6, 103054.8, 
    103053.3, 103005.2, 102954.6, 102882.9, 102808.9, 102744.1, 102697.6, 
    102635.3,
  100838, 100670, 102719, 102914.1, 102925.6, 102975.2, 102981, 102989.7, 
    102958.3, 102933.7, 102873.4, 102824.1, 102759.4, 102706.1, 102648,
  98725.05, 98890.52, 102543.5, 102866.7, 102874.2, 102947.5, 102963.7, 
    102978.2, 102945.2, 102917.6, 102870.1, 102826, 102777.8, 102735.5, 
    102690.3,
  98703.19, 99231.3, 101177.6, 102802.8, 102839.3, 102858.8, 102884.6, 
    102901.7, 102900.5, 102896.8, 102865.9, 102825.3, 102801.9, 102761.1, 
    102719.1,
  97950.86, 99571.02, 102472.8, 102722.3, 102762.2, 102803.1, 102899.9, 
    102916.3, 102887.1, 102876.3, 102837.3, 102795.2, 102822.9, 102798.1, 
    102747.7,
  102394.7, 102518.4, 102621.2, 102711.2, 102727.2, 100926.6, 102474.6, 
    102646.9, 102796.6, 102866.7, 102873.7, 102846.2, 102831.6, 102806, 
    102749.1,
  102473.6, 102484.1, 102560.2, 102557, 102513.1, 100066.7, 98180.54, 
    97347.64, 99947.85, 102825.7, 102864.7, 102842.6, 102825.7, 102792.7, 
    102743.5,
  102320.3, 102365.1, 102499.4, 102523.3, 97620.69, 99073.13, 100853.9, 
    102491, 102732.3, 102789.9, 102802.1, 102782.5, 102776.7, 102759.1, 
    102722.8,
  102269.1, 102308.4, 102408.7, 102394.8, 98047.92, 98349.84, 97922.52, 
    102554.4, 102825.2, 102716.5, 102760.7, 102733.5, 102741.1, 102719.9, 
    102706.4,
  102428.1, 102450.6, 102508.7, 102570.4, 102627.6, 102651.5, 102664.4, 
    102642.3, 102610.2, 102584.2, 102517.9, 102472.3, 102460.9, 102433.7, 
    102416.7,
  102332.7, 102353.2, 102480.9, 102537.6, 102580, 102638.8, 102663.3, 
    102656.6, 102626.6, 102605.5, 102547.5, 102509.7, 102463.2, 102460.9, 
    102455.4,
  100503, 100316.2, 102339.9, 102510.6, 102545.5, 102587.4, 102608.5, 
    102621.9, 102600.2, 102593.4, 102549.1, 102532.4, 102503.7, 102497.2, 
    102487.6,
  98433.15, 98569.41, 102184.6, 102481.2, 102503, 102578, 102602.1, 102616.8, 
    102595.2, 102582.9, 102557.8, 102557.1, 102531, 102513.3, 102527,
  98422.16, 98921.46, 100825.2, 102426.3, 102467.7, 102484, 102528.6, 
    102555.1, 102566.3, 102569.8, 102559.5, 102573.9, 102558.9, 102564.3, 
    102570.3,
  97780.02, 99287.03, 102109.1, 102351.6, 102404.2, 102447.2, 102524.1, 
    102551.6, 102545.3, 102550.1, 102545.2, 102538.7, 102584.7, 102604.2, 
    102605.5,
  102333.7, 102327.9, 102276.2, 102344, 102348.5, 100590.4, 102135, 102292.4, 
    102432, 102499.2, 102538.6, 102577, 102596.9, 102624.7, 102620.6,
  102433.9, 102354.7, 102324.5, 102222.6, 102157.5, 99727.76, 97882.41, 
    97078.56, 99682.91, 102488.6, 102543.4, 102570.4, 102595.6, 102628.4, 
    102634.5,
  102368.4, 102322.1, 102340.4, 102232.6, 97337.84, 98795.63, 100539.1, 
    102125.8, 102381.1, 102478.5, 102522.6, 102551.8, 102588.4, 102618.5, 
    102636.6,
  102396.4, 102353.5, 102349.7, 102225.5, 97787.94, 98091.53, 97660.93, 
    102243.9, 102494.4, 102432.1, 102500.5, 102521, 102565.9, 102591.9, 
    102626.7,
  102556.3, 102541.6, 102516.2, 102482.2, 102475, 102476.1, 102487.8, 
    102487.8, 102474.2, 102457.1, 102427.1, 102380.5, 102328.4, 102299.8, 
    102267.4,
  102494.3, 102431.7, 102497.7, 102473.4, 102440.3, 102438.1, 102452.8, 
    102463.5, 102449.3, 102431.3, 102402.7, 102359, 102321.9, 102284.9, 102267,
  100628.1, 100331.3, 102338.3, 102432.1, 102406.7, 102408, 102403, 102418.7, 
    102414.6, 102402, 102375.1, 102344.5, 102316.3, 102278, 102250.1,
  98551.32, 98650.41, 102187.9, 102448.4, 102420.1, 102429.6, 102401.9, 
    102408.3, 102388.8, 102376.6, 102355.6, 102329.6, 102309.4, 102260.7, 
    102254.1,
  98535.53, 99004.02, 100852.3, 102424.3, 102423.1, 102400.5, 102380.2, 
    102371.4, 102360.6, 102358.3, 102339.6, 102324.3, 102296.5, 102273.3, 
    102253.6,
  97826.3, 99380.03, 102246.5, 102400.6, 102409, 102367.5, 102415.2, 
    102392.4, 102362.4, 102358, 102318.2, 102273.7, 102305.7, 102280.2, 
    102264.9,
  102208.7, 102343.5, 102396.5, 102430.2, 102420.6, 100561.3, 102047, 
    102177.8, 102287, 102331.2, 102324.4, 102312.4, 102304.9, 102281, 102271.8,
  102303.6, 102339.4, 102394.1, 102383.5, 102218.5, 99743.66, 97803.53, 
    96935.52, 99508.35, 102297.2, 102313.8, 102308, 102296.7, 102285.1, 
    102280.1,
  102214.2, 102270.6, 102372.6, 102374, 97376.32, 98851.92, 100557.3, 
    102130.9, 102257.7, 102291, 102285.3, 102287.2, 102293.4, 102291.2, 
    102286.4,
  102162.1, 102243.5, 102344.7, 102320.2, 97910.62, 98158.04, 97619.39, 
    102191, 102373.3, 102288.8, 102296.1, 102281.2, 102295.7, 102292.9, 
    102294.2,
  101492.4, 101532.4, 101591, 101645.7, 101714.7, 101776.9, 101845.2, 
    101896.7, 101954.9, 101999.5, 102034.7, 102057.6, 102074.7, 102091.1, 
    102097.2,
  101373.7, 101442.1, 101564.3, 101633.5, 101695.7, 101760.4, 101824.3, 
    101882.8, 101942.2, 101988.3, 102016.8, 102048.6, 102068.5, 102091, 102111,
  99583.75, 99448.23, 101453.6, 101634.6, 101677.9, 101742.5, 101805.1, 
    101865.3, 101926.7, 101967.3, 102011.1, 102053.7, 102077.3, 102094, 
    102112.4,
  97521.13, 97745.34, 101342, 101608.4, 101670.2, 101744.5, 101800.1, 
    101860.2, 101912.6, 101959.2, 102011.5, 102051.4, 102076.3, 102082.8, 
    102114.4,
  97493.29, 98053.06, 100034.2, 101595, 101670.9, 101714.5, 101783.1, 
    101840.6, 101890.3, 101957.1, 102015.3, 102063.1, 102085, 102103.3, 
    102120.4,
  96870.9, 98423.26, 101331.9, 101561.8, 101662.3, 101685.6, 101808, 
    101865.5, 101917.2, 101976.6, 102015.5, 102018.9, 102090.4, 102115.6, 
    102126.2,
  101160.9, 101317.9, 101504.3, 101589, 101658.7, 99956.55, 101506.8, 
    101661.8, 101856.6, 101952.7, 102045.5, 102067.3, 102102.5, 102122.4, 
    102134.7,
  101349.7, 101382.4, 101494.3, 101540, 101523, 99090.73, 97338.42, 96573.5, 
    99195.45, 101971.7, 102046.1, 102073.1, 102106.3, 102132.8, 102136.3,
  101277.8, 101349.8, 101513.6, 101529.8, 96841.87, 98325.41, 100027.3, 
    101600.5, 101896.3, 101971.3, 102033.4, 102070, 102121, 102135.7, 102136,
  101290.4, 101376.2, 101515.5, 101508.3, 97285.75, 97642.39, 97218.08, 
    101795.4, 102020.4, 101981.2, 102057.2, 102091.8, 102132.4, 102140.4, 
    102139.6,
  101731.5, 101741.2, 101752.7, 101765.1, 101752, 101778.4, 101785.7, 101786, 
    101772, 101749.3, 101725.5, 101706.1, 101683.5, 101664.9, 101661.2,
  101545.3, 101540.1, 101630.5, 101665, 101644.8, 101656.6, 101663.7, 
    101676.2, 101679.7, 101676.7, 101659.4, 101639.6, 101620, 101629.7, 
    101656.2,
  99603.26, 99403.04, 101400.9, 101574.5, 101541.3, 101549.2, 101549.6, 
    101555.8, 101563.2, 101579.5, 101577.4, 101575.4, 101577.1, 101594.4, 
    101623.6,
  97510.62, 97579.79, 101143.9, 101426.4, 101410, 101439.9, 101457, 101470.4, 
    101472.2, 101482.9, 101486.8, 101495.5, 101514.3, 101535.9, 101593.5,
  97468.84, 97945.83, 99785.17, 101314, 101304.8, 101290.5, 101332.7, 
    101362.3, 101369.2, 101393.7, 101416.5, 101438.9, 101461.6, 101508.8, 
    101569.6,
  96827.15, 98346.84, 101125, 101269.4, 101226.3, 101198.5, 101258.7, 
    101297.3, 101306.5, 101325.2, 101332.9, 101329, 101424.6, 101482.1, 
    101544.9,
  101286.4, 101306.9, 101285.9, 101252.2, 101185.3, 99363.27, 100845.5, 
    101001.7, 101154, 101214.6, 101281.6, 101318.6, 101383.9, 101451.4, 
    101526.6,
  101325, 101243.4, 101220.7, 101130, 100948.5, 98479.94, 96608.2, 95826.64, 
    98362.84, 101140.5, 101224.4, 101263.4, 101333.5, 101421.3, 101509,
  101237.6, 101163.3, 101177.6, 101096.6, 96166.53, 97544.2, 99200.99, 
    100725, 101001.3, 101115.3, 101170.1, 101215.4, 101291.7, 101389.4, 
    101492.3,
  101226.3, 101143.2, 101129, 100999, 96610.29, 96827.41, 96369.62, 100830.2, 
    101088.9, 101039, 101121.6, 101169.2, 101254.9, 101359.9, 101477.2,
  101395, 101481.4, 101584.7, 101692.5, 101794.4, 101876.9, 101938.5, 
    101980.5, 102000, 102011.1, 102001.6, 101973.8, 101939.1, 101898.5, 
    101843.9,
  101272.5, 101365.6, 101519.9, 101625.1, 101715.4, 101811.3, 101879.7, 
    101929.4, 101955.9, 101966.6, 101959.6, 101933.8, 101906.4, 101870.2, 
    101846.3,
  99424.55, 99316.52, 101355.8, 101588.7, 101655.3, 101744, 101804.3, 
    101848.3, 101878.4, 101899, 101896, 101883.9, 101862.6, 101835.8, 101817.4,
  97318.14, 97541.76, 101194.8, 101524.3, 101590.4, 101696.3, 101753.8, 
    101807.2, 101828.2, 101842.4, 101840.9, 101838.7, 101816.3, 101800.1, 
    101801.1,
  97246.37, 97838, 99838.11, 101455.9, 101541.7, 101600.1, 101663.5, 
    101699.2, 101727.1, 101763, 101782.2, 101798.1, 101778, 101780.8, 101771.9,
  96602.88, 98169.71, 101115.4, 101380.3, 101472.5, 101527.4, 101659.5, 
    101695.6, 101699.3, 101712.4, 101701.8, 101695.8, 101746.8, 101753.6, 
    101743.8,
  100899.9, 101086.6, 101266.2, 101382.3, 101445.6, 99710.38, 101253.6, 
    101410.8, 101561.3, 101641.3, 101674.7, 101689.5, 101704.7, 101716.5, 
    101710.9,
  101029.7, 101092.6, 101221.3, 101282, 101250.5, 98850.56, 97016.84, 
    96209.54, 98797.77, 101592.4, 101643.5, 101652.2, 101656.9, 101672, 
    101672.9,
  100937.3, 101037.6, 101215.1, 101258, 96471.27, 97957.79, 99686.16, 
    101239.1, 101479.5, 101562.6, 101594.5, 101608.9, 101618.2, 101627.4, 
    101630.2,
  100963, 101058.6, 101199.4, 101207.3, 96915.8, 97239.2, 96812.79, 101373, 
    101598.8, 101509.6, 101549.2, 101561.3, 101577.6, 101585.4, 101592.6,
  102041.3, 102041.4, 102082, 102103.1, 102144.9, 102185.5, 102211.6, 
    102216.4, 102207.7, 102197.7, 102178.5, 102144.8, 102106.2, 102063.5, 
    102019.3,
  101911, 101935.7, 102061.6, 102073.9, 102069.1, 102110.7, 102150.6, 
    102174.7, 102176.5, 102172.5, 102151.5, 102124.3, 102088, 102057.7, 
    102034.4,
  100013.7, 99820.09, 101838.9, 102018.4, 101988.3, 102014.1, 102043.3, 
    102082.7, 102105.2, 102127.4, 102124.7, 102112, 102083.4, 102057.2, 
    102037.5,
  97864.24, 98015.41, 101671.9, 101970.8, 101953.3, 101990.2, 102009, 
    102037.2, 102054.5, 102076.1, 102077.7, 102079.3, 102060.8, 102038.5, 
    102045.1,
  97794.61, 98322.28, 100257.6, 101864, 101889.1, 101877.8, 101918.1, 
    101946.2, 101971.1, 102011, 102031, 102047.6, 102032.3, 102039.7, 102042.8,
  97028.95, 98626.94, 101555.5, 101764.7, 101798.9, 101812.2, 101883.3, 
    101911.9, 101924.7, 101948.4, 101961.1, 101954.6, 102014.9, 102026.4, 
    102034.5,
  101442.1, 101569.3, 101652.6, 101710.6, 101690.7, 99927.1, 101473.1, 
    101615.2, 101769.3, 101855.3, 101919.4, 101953.4, 101986.8, 102006.1, 
    102023,
  101480.6, 101471.8, 101541.2, 101551.2, 101487.5, 99013.87, 97184.37, 
    96394.13, 98978.23, 101791.9, 101866.6, 101904.7, 101942.8, 101975.6, 
    101999.9,
  101326.2, 101362.9, 101491.9, 101481.5, 96586.24, 98056.52, 99773.23, 
    101332.7, 101635.4, 101762.9, 101812.8, 101853.2, 101898.6, 101937.1, 
    101972,
  101240.6, 101286.3, 101400.5, 101370.5, 97030.45, 97325.39, 96906.78, 
    101492, 101745.5, 101694.9, 101760.9, 101797.2, 101856.1, 101895.5, 
    101934.5,
  102287.4, 102270.6, 102270.6, 102271.4, 102247.5, 102215.9, 102164.8, 
    101991, 101902, 101808.6, 101738.2, 101757, 101784.6, 101808.5, 101798.3,
  102196.6, 102199.6, 102274.8, 102280.7, 102269.4, 102254.8, 102219.4, 
    102097.4, 101989.7, 101866.8, 101807.9, 101819.8, 101836.5, 101854.8, 
    101859.4,
  100348.1, 100171.5, 102185.7, 102318.6, 102303.4, 102284.8, 102234.3, 
    102138.9, 102032.2, 101939.5, 101876.2, 101875.7, 101886.5, 101891.6, 
    101891.4,
  98269.79, 98422.45, 102069.6, 102336.2, 102325.8, 102350.9, 102302.5, 
    102238.8, 102110.1, 102021.5, 101951.2, 101935.3, 101935.3, 101928.1, 
    101936.5,
  98238.69, 98763.34, 100741.8, 102321.5, 102339.5, 102327.2, 102313.6, 
    102274.1, 102164.8, 102093, 102024.6, 102000.7, 101980.1, 101984.2, 
    101977.1,
  97567.19, 99132.88, 102068.6, 102286.8, 102329.2, 102328, 102378.9, 102374, 
    102251.2, 102173.8, 102086.2, 102012.7, 102045.2, 102036.2, 102021.7,
  101974.7, 102091.5, 102229.6, 102315.4, 102322.6, 100490, 102033.9, 
    102133.8, 102204.8, 102196, 102163.3, 102115, 102102.9, 102081.6, 102062,
  102079.5, 102068.4, 102191, 102201.8, 102166.6, 99656.5, 97734.74, 96873.4, 
    99462.06, 102226.2, 102236.6, 102183.1, 102156.4, 102128.3, 102101.6,
  101952.1, 101984.1, 102165.9, 102184.4, 97302.25, 98755.45, 100519.4, 
    102092.6, 102270.2, 102286.1, 102282.6, 102229.8, 102203.4, 102166.8, 
    102138,
  101937, 101985.1, 102108.4, 102103.1, 97770.99, 98047.13, 97587.1, 
    102211.8, 102433.7, 102306.3, 102329.7, 102267.6, 102244.2, 102197.1, 
    102172.3,
  102618.4, 102563.7, 102516.5, 102447.4, 102371.3, 102297.5, 102212.9, 
    102124.4, 101995.1, 101907.2, 101857.6, 101816.4, 101774.6, 101728, 
    101677.1,
  102511, 102432, 102473.1, 102422.4, 102332.3, 102256.4, 102159.7, 102066.2, 
    101928, 101832.9, 101778.5, 101736.8, 101706.8, 101687.2, 101669.3,
  100598.4, 100290.9, 102279.9, 102367.3, 102275.1, 102207.7, 102095.7, 
    102006.8, 101848, 101740.3, 101672.7, 101653.1, 101640.4, 101636.6, 
    101630.6,
  98474.83, 98532.7, 102101.4, 102305.1, 102222.6, 102177.5, 102084.3, 
    101998.7, 101845.4, 101701.4, 101604.4, 101594.2, 101582.1, 101585.4, 
    101612,
  98415.3, 98862.46, 100705.6, 102204.4, 102146.6, 102082.7, 102020.5, 
    101926.5, 101784.1, 101639.8, 101540.2, 101537.2, 101529.1, 101563.5, 
    101581.8,
  97787.41, 99251.06, 102079.3, 102201.4, 102106.8, 102041.5, 102034, 
    101974.1, 101814.2, 101634.8, 101469, 101433.1, 101490.7, 101535.7, 
    101556.9,
  102301.4, 102283, 102279.2, 102212.8, 102125.4, 100244.6, 101706.6, 
    101710.4, 101681.7, 101577.6, 101442.2, 101418.9, 101446.5, 101491.8, 
    101523.2,
  102346.2, 102280.1, 102266.7, 102149.9, 101957.6, 99389.7, 97418.56, 
    96460.73, 98985.21, 101562.3, 101435.6, 101365.8, 101404.4, 101453.4, 
    101495.1,
  102273, 102215.9, 102240.3, 102145.7, 97108.55, 98517.2, 100189.5, 101714, 
    101761.7, 101603.3, 101411.3, 101315.4, 101361.2, 101415.7, 101469.1,
  102250.4, 102195.3, 102205.4, 102088.2, 97625.3, 97826.46, 97221.77, 
    101764.5, 101837.5, 101609.6, 101407.2, 101284.4, 101329.7, 101384.7, 
    101450.4,
  102641.4, 102678.9, 102714.6, 102731.9, 102729, 102725.6, 102711, 102682.4, 
    102644.9, 102604.7, 102552.5, 102479.6, 102397.5, 102337, 102263.9,
  102574.5, 102601.9, 102699.5, 102722.7, 102710.3, 102713.1, 102700.2, 
    102681.9, 102644.2, 102605.2, 102542.3, 102473.6, 102406.8, 102354.5, 
    102302.1,
  100733.9, 100529.1, 102566.5, 102713.1, 102683, 102683.6, 102648.8, 
    102627.2, 102590.4, 102573.4, 102516.7, 102463.4, 102403.3, 102344.2, 
    102293.1,
  98638.44, 98764.66, 102391.3, 102685.3, 102647, 102671.7, 102648, 102612.4, 
    102571.9, 102531.4, 102487.1, 102439.3, 102391.2, 102330.2, 102302.6,
  98596.98, 99121.91, 101026.4, 102610.5, 102603.9, 102580.7, 102561.7, 
    102535.5, 102512, 102479.2, 102450.8, 102416.4, 102378, 102339.2, 102299.3,
  97847.86, 99464.16, 102346.4, 102555.9, 102543, 102521.9, 102574.5, 
    102546.1, 102497.9, 102464.9, 102411.9, 102349.6, 102366.3, 102335.6, 
    102296.5,
  102243.7, 102405.9, 102482.6, 102543.8, 102532, 100672.9, 102163.3, 
    102292.4, 102414.5, 102440.3, 102427.8, 102391.9, 102356.9, 102323.4, 
    102290.3,
  102344.2, 102387.6, 102456.6, 102438.1, 102317.9, 99840.7, 97889.09, 
    96993.38, 99553.75, 102370.1, 102392.2, 102364.2, 102333.9, 102309.8, 
    102279.8,
  102239, 102292.4, 102420.6, 102422.4, 97467.77, 98874.41, 100613.3, 
    102190.8, 102356.6, 102367.9, 102352.6, 102325.1, 102301.3, 102279.6, 
    102251.7,
  102202.6, 102265.6, 102378.3, 102339.3, 97934.87, 98166.2, 97658.73, 
    102222, 102441.8, 102313.5, 102320.9, 102285, 102267.6, 102244.1, 102221.7,
  102089.5, 102110.5, 102139.4, 102167.9, 102191.1, 102212.6, 102214.1, 
    102210.4, 102217.2, 102215.4, 102211.5, 102207.8, 102202.1, 102192, 
    102157.4,
  102098.9, 102111.8, 102196, 102235.1, 102258.5, 102279.7, 102292, 102288.3, 
    102284.6, 102270, 102257, 102250.8, 102244.5, 102238, 102212.1,
  100374.2, 100184, 102180.9, 102297, 102303.7, 102320.6, 102327.4, 102324.9, 
    102324.4, 102315.3, 102308.4, 102302.7, 102288.2, 102270.1, 102248.1,
  98363.96, 98567.52, 102116.8, 102339.9, 102360.4, 102383.7, 102393.7, 
    102397.2, 102386.4, 102374.9, 102366.4, 102358.7, 102339.3, 102302.6, 
    102295.7,
  98370.34, 98897.29, 100845.5, 102384.8, 102401.3, 102393.4, 102419.9, 
    102428.3, 102429.9, 102428.8, 102416.9, 102407, 102381.7, 102359.8, 102335,
  97726.95, 99286.49, 102183.9, 102388, 102423.5, 102403.6, 102494.4, 
    102509.6, 102502.5, 102486.7, 102458.9, 102409.2, 102435.1, 102411.2, 
    102382.5,
  101960.3, 102160.7, 102353, 102436.4, 102450.2, 100664.7, 102207.5, 
    102327.2, 102463.5, 102504.8, 102514.6, 102492.9, 102477.6, 102452.1, 
    102422.4,
  102139.8, 102212.9, 102337.9, 102373.5, 102295, 99832.58, 97988.05, 
    97151.13, 99775.53, 102545, 102561.6, 102531.5, 102513.9, 102490.4, 
    102461.5,
  102038.8, 102135.3, 102320, 102356.8, 97561.3, 99017.27, 100757.2, 
    102360.5, 102588.3, 102589.4, 102593.8, 102558.9, 102545.7, 102521.7, 
    102499.2,
  102013.1, 102123.8, 102291.8, 102294.5, 98017.41, 98334.71, 97877.62, 
    102471, 102684.5, 102611.5, 102627.9, 102591, 102578.7, 102551.5, 102536.2,
  100729.9, 100796.9, 100879.9, 100951.7, 101040.3, 101139.2, 101229.6, 
    101311, 101391.2, 101476.5, 101554.2, 101615.9, 101670.6, 101714.6, 101738,
  100661.9, 100727.3, 100868.7, 100963.4, 101055, 101163.5, 101263, 101353.8, 
    101439.2, 101516.5, 101586, 101647.5, 101701.7, 101750.5, 101786.9,
  98942.42, 98824.09, 100783, 100992.4, 101072.3, 101189.7, 101299.2, 
    101396.1, 101484.1, 101557.9, 101627.3, 101690.9, 101744.5, 101786.6, 
    101820.3,
  96990.74, 97229.76, 100697.9, 101000.7, 101101, 101216.8, 101327.1, 101432, 
    101526.2, 101604.7, 101674.1, 101738.5, 101788.7, 101816.7, 101864.9,
  97020.55, 97572.94, 99468.48, 101028.4, 101127.4, 101223.1, 101351.2, 
    101453, 101547.3, 101643, 101724.2, 101792.8, 101832.9, 101874.4, 101905.6,
  96480.88, 97997.16, 100798.1, 101041.2, 101145.5, 101216.1, 101382.7, 
    101500.4, 101604.2, 101696.7, 101767.6, 101796.5, 101890, 101929.8, 
    101947.7,
  100777.8, 100872, 101018, 101104.1, 101163.5, 99571.23, 101143, 101331, 
    101555.5, 101703.4, 101824.4, 101887.3, 101942.4, 101975.1, 101989.7,
  100925.1, 100948.9, 101037.3, 101090, 101067.6, 98735.88, 97075.97, 
    96383.16, 98993.69, 101745.6, 101865, 101934.1, 101990.6, 102022, 102037.5,
  100853.4, 100917.5, 101063.5, 101073.3, 96527.19, 98040.15, 99751.49, 
    101309.8, 101643.7, 101798.3, 101905.8, 101975.1, 102035.7, 102065.7, 
    102083.1,
  100909, 100966.6, 101087.9, 101078, 96999.7, 97387.05, 97041.79, 101565, 
    101809.6, 101837.4, 101944.4, 102013.5, 102078.2, 102107.1, 102127.9,
  101095.5, 101020, 100958.6, 100903.9, 100905.4, 100904.6, 100929.9, 
    100985.8, 101058.2, 101145.4, 101235.6, 101302.6, 101371, 101440.4, 
    101481.9,
  101080, 100990, 101046.8, 100983.9, 100948.6, 100945.2, 100962.8, 101007.5, 
    101071.7, 101157.9, 101234.4, 101314.6, 101388.6, 101456.1, 101510,
  99337.73, 99083.09, 101027.7, 101086.2, 101011.4, 100981.4, 100983.2, 
    101022.8, 101090.2, 101173.1, 101258.5, 101334, 101412.4, 101476.1, 
    101532.5,
  97471.86, 97608.34, 100975.4, 101167.6, 101080.6, 101042.3, 101014.7, 
    101050.8, 101109.4, 101192.3, 101261.9, 101348.5, 101433, 101482, 101557.8,
  97579.84, 98048.49, 99805.56, 101224.1, 101150, 101051.7, 101029.8, 
    101052.1, 101118.6, 101198.4, 101281, 101371.6, 101441.4, 101513, 101579.5,
  97149.15, 98588.09, 101249.2, 101277.7, 101185.8, 101043.7, 101071.2, 
    101075.9, 101134.7, 101194.2, 101278.7, 101329.2, 101463.4, 101537.8, 
    101601.5,
  101578.5, 101511.7, 101418.2, 101338.6, 101229.6, 99350.2, 100756.4, 
    100863.9, 101056.1, 101154.8, 101291.2, 101380.1, 101475.3, 101551.5, 
    101621.6,
  101630.5, 101506.7, 101444.5, 101303, 101024.2, 98588.75, 96719.97, 
    95913.52, 98430.64, 101136.3, 101275.9, 101371.4, 101475.8, 101556.1, 
    101633.2,
  101604.7, 101493.2, 101459.3, 101303.5, 96402.8, 97798.33, 99392.08, 
    100819.3, 101033.8, 101154.7, 101260.6, 101358.9, 101470.3, 101555.8, 
    101638.7,
  101604.5, 101507.8, 101466.8, 101312.3, 96951.13, 97131.4, 96610.76, 
    100998.5, 101174.7, 101143.7, 101245, 101345.7, 101464.2, 101552.8, 
    101641.2,
  100863, 100762.1, 100685, 100612.3, 100555.9, 100542.1, 100539.9, 100574.3, 
    100644.8, 100738.4, 100842.1, 100927.1, 101014.4, 101102.3, 101169.6,
  100802.6, 100686.4, 100707.3, 100635.3, 100555.4, 100530.5, 100541, 
    100582.5, 100636.7, 100718.6, 100821.3, 100916.6, 101017.1, 101117.7, 
    101201.8,
  99020.36, 98687.42, 100586.5, 100671.6, 100589.4, 100531.1, 100531.9, 
    100573.6, 100638.3, 100719.9, 100816.8, 100920.4, 101028.7, 101124.3, 
    101208.3,
  97051.75, 97107.37, 100487.8, 100693.8, 100605.2, 100557.3, 100527, 
    100572.4, 100640, 100721.1, 100812.5, 100921.7, 101033.8, 101122.6, 
    101228.2,
  97035.58, 97494.66, 99237.43, 100677.6, 100594.3, 100528.7, 100508.8, 
    100549.8, 100636.7, 100724.9, 100821.1, 100929.4, 101030, 101139.2, 
    101236.3,
  96440.96, 97909.47, 100578.2, 100667.1, 100570.8, 100490.5, 100518.5, 
    100542.4, 100620.4, 100710.6, 100812.2, 100882.2, 101042.8, 101152, 
    101247.8,
  100820.8, 100810.9, 100731, 100660.7, 100545.5, 98759.45, 100180.3, 
    100321.2, 100533.6, 100659.8, 100818.2, 100933.1, 101049.9, 101156.3, 
    101253.2,
  100874.6, 100767.6, 100702.2, 100568.5, 100340.3, 97926.54, 96135.59, 
    95380.06, 97888.79, 100628.6, 100798.9, 100925.9, 101051, 101156.9, 
    101257.4,
  100833.7, 100729.9, 100699, 100545.8, 95728.11, 97109.89, 98714.07, 
    100173.2, 100448.4, 100621.1, 100768.3, 100907, 101044.5, 101155.1, 
    101254.9,
  100831.9, 100739.2, 100696.9, 100514.4, 96213.98, 96438.77, 95989.91, 
    100360.8, 100567.4, 100576.6, 100736, 100884.5, 101036.4, 101148.5, 101253,
  101454.9, 101372.6, 101300.3, 101227.1, 101168.6, 101106.6, 101050.7, 
    100979.9, 100933.4, 100877.6, 100869.1, 100864.2, 100861.3, 100889.3, 
    100937.7,
  101340.6, 101238, 101258.2, 101193.7, 101123.1, 101072.6, 101029, 100965.1, 
    100927.5, 100878.5, 100847.7, 100843.3, 100846.5, 100890.2, 100964.1,
  99505.47, 99160.96, 101047.3, 101153.6, 101105, 101064.8, 100992, 100930.3, 
    100890.5, 100865, 100832.2, 100838.9, 100836.9, 100883, 100952.4,
  97491.8, 97496.73, 100975.3, 101212, 101115.8, 101064.8, 100971.9, 
    100912.2, 100859.4, 100837.6, 100804, 100818.4, 100827.4, 100857.2, 100957,
  97464.05, 97910.61, 99705.84, 101173.1, 101095.6, 101000.6, 100921.3, 
    100847.6, 100800.3, 100792.2, 100770.2, 100794.4, 100809.5, 100852, 
    100945.4,
  96870.4, 98358.85, 101082.2, 101164.4, 101070.8, 100929.3, 100908.6, 
    100822.1, 100761.9, 100743.1, 100718.5, 100706.6, 100798.2, 100840.2, 
    100930.2,
  101274.1, 101277.3, 101225.6, 101161.4, 101067.4, 99139.43, 100483.3, 
    100511.3, 100598.1, 100637.5, 100674.3, 100700.2, 100769.2, 100821.4, 
    100907.8,
  101309.7, 101219.7, 101188.7, 101089.2, 100831.7, 98324.52, 96365.67, 
    95414.95, 97847.07, 100547.4, 100611.5, 100644.5, 100721.4, 100794.6, 
    100882.2,
  101208.1, 101150.2, 101158, 101086.6, 96116.51, 97417.13, 99039.31, 
    100490.8, 100607.2, 100581.7, 100578.3, 100593.7, 100670.8, 100756.5, 
    100852.1,
  101164.9, 101113.7, 101105.1, 101010.3, 96617.25, 96789.41, 96148.23, 
    100508.2, 100650.1, 100510.7, 100530.3, 100537.5, 100622.7, 100715, 
    100819.8,
  101920.8, 101822.8, 101744, 101649.3, 101556.5, 101477.4, 101405.4, 
    101284.1, 101155.4, 101052.4, 100947.2, 100879.3, 100848, 100826.1, 
    100830.5,
  101847.2, 101729.5, 101759.8, 101664.5, 101550.7, 101487.2, 101410.8, 
    101323.1, 101215, 101109.5, 100978.2, 100876.2, 100844.9, 100830.3, 
    100851.5,
  99982.29, 99630.05, 101602.7, 101638.1, 101568.6, 101528.4, 101411.3, 
    101324.3, 101225, 101112.7, 101002.8, 100910.4, 100846.7, 100821.4, 
    100833.1,
  97937.72, 97965.26, 101452.9, 101668, 101595.5, 101550.4, 101435.4, 
    101339.8, 101248, 101143, 101037.4, 100943.4, 100858.5, 100812.6, 100836.9,
  97873.64, 98328.71, 100136.6, 101650.6, 101605.5, 101523, 101434.9, 
    101337.9, 101242, 101161.4, 101059.5, 100963.5, 100880.9, 100833, 100843.2,
  97179.69, 98694.72, 101517.2, 101662.5, 101601.1, 101489.4, 101476.2, 
    101360.3, 101249.6, 101174.5, 101068.9, 100947.6, 100912, 100852.6, 
    100838.7,
  101635.3, 101675.9, 101705.1, 101675.2, 101618.2, 99694.29, 101107.4, 
    101116.4, 101158.1, 101154, 101093.9, 101009.3, 100932.4, 100874.1, 
    100840.5,
  101687.2, 101644.6, 101674.4, 101589.8, 101418.7, 98907.59, 96945.98, 
    95947.86, 98449.47, 101164.1, 101117.6, 101023.6, 100949.3, 100888, 
    100839.4,
  101535.3, 101550, 101608.2, 101603.4, 96632.97, 97962.77, 99676.11, 
    101195.8, 101308.3, 101220.2, 101132.9, 101042.1, 100966.7, 100902.3, 
    100843.6,
  101489.2, 101509.9, 101557.7, 101506.6, 97117.65, 97312.43, 96747.12, 
    101202.1, 101355.3, 101179, 101156.7, 101062.2, 100991.7, 100913.3, 
    100861.1,
  101766.4, 101720.9, 101664.7, 101614.7, 101536.1, 101458.7, 101380.1, 
    101273.5, 101175.7, 101055.8, 100975.7, 100936.1, 100922.8, 100929, 
    100940.5,
  101693.6, 101612.9, 101653.8, 101605.5, 101500, 101435.1, 101360.1, 
    101260.9, 101145.5, 101014.7, 100916.9, 100860.9, 100847.4, 100868.6, 
    100913.5,
  99802.78, 99491.42, 101492, 101564.5, 101468.8, 101419.7, 101324.6, 
    101217.3, 101092, 100963.6, 100853.3, 100783.5, 100775.8, 100802.8, 
    100851.8,
  97738.53, 97804.02, 101329.6, 101537.2, 101458.4, 101416.2, 101337.6, 
    101233.2, 101086.3, 100938.2, 100790.7, 100713.2, 100705.1, 100724.3, 
    100805.6,
  97667, 98139.08, 99971.22, 101490, 101443.5, 101364.7, 101322.5, 101208.7, 
    101067.6, 100910.1, 100758.8, 100657, 100634, 100672.5, 100749.4,
  96953.88, 98493.2, 101339.9, 101459.1, 101422.6, 101305.6, 101357.2, 
    101247.4, 101115.9, 100922.9, 100743.7, 100570.1, 100580.3, 100616.6, 
    100693.5,
  101369.7, 101446, 101479.8, 101456.1, 101430.4, 99510.98, 101017.9, 
    101011.8, 101021.4, 100904.2, 100769.1, 100597.8, 100537.9, 100566.4, 
    100641.4,
  101431, 101412.9, 101450.3, 101401.9, 101235, 98709.87, 96751.3, 95794.79, 
    98330.11, 100933.4, 100814.3, 100628.7, 100520.4, 100533.5, 100601.9,
  101316.7, 101334.5, 101413.1, 101400.4, 96427.48, 97836.48, 99531.6, 
    101060.3, 101136.3, 100959.3, 100850.5, 100681.5, 100522.3, 100502.6, 
    100571.6,
  101301.1, 101319.8, 101377.8, 101332.8, 96949.17, 97156.52, 96558.62, 
    101094.9, 101188, 100985.6, 100895.3, 100730, 100546.1, 100479.8, 100540.9,
  101987.7, 101963.2, 101951.5, 101914.1, 101858.6, 101828.5, 101773.9, 
    101709, 101593.4, 101474.7, 101374.2, 101295.3, 101249.4, 101246.9, 
    101252.6,
  101895.2, 101859.1, 101936.4, 101924.4, 101858.2, 101827.1, 101789.8, 
    101740.5, 101658.4, 101560.1, 101415.5, 101317.8, 101277, 101273.5, 
    101288.7,
  100047.2, 99765.32, 101767.3, 101881.5, 101834.8, 101810.6, 101755.6, 
    101720.2, 101653.8, 101570, 101448.2, 101377.1, 101314.9, 101287.5, 
    101287.5,
  97988.16, 98039.96, 101574.8, 101852.7, 101804.4, 101816.5, 101762, 
    101728.9, 101670.7, 101595.9, 101502.5, 101412, 101350.2, 101303.3, 
    101317.2,
  97918.42, 98397.29, 100234.6, 101781.8, 101771.6, 101744.8, 101718.1, 
    101695.1, 101660.6, 101599.5, 101527.1, 101460.5, 101389.8, 101343.4, 
    101332.3,
  97167.71, 98718.3, 101529, 101737.9, 101723.5, 101704.9, 101746.9, 
    101699.7, 101669.3, 101626.8, 101547.2, 101445.3, 101436.8, 101387.6, 
    101364.6,
  101555.2, 101617.8, 101688.1, 101719.5, 101706.5, 99864.73, 101349.6, 
    101458.5, 101583.7, 101607.4, 101581, 101515.2, 101451.8, 101416.1, 
    101380.6,
  101597.5, 101583.3, 101645.7, 101598.6, 101505.1, 99043.02, 97130.4, 
    96191.81, 98736.36, 101528.2, 101547.1, 101499.2, 101452.3, 101431.5, 
    101403.2,
  101451.6, 101475.9, 101576.6, 101581, 96705.44, 98080.84, 99838.2, 
    101394.6, 101552, 101532.3, 101533.8, 101488.6, 101450.9, 101421.5, 
    101398.4,
  101432.3, 101435.2, 101490.6, 101468.8, 97153.54, 97388.91, 96888.23, 
    101396.6, 101612.2, 101482.2, 101507.2, 101454.3, 101436.5, 101396.5, 
    101392,
  101891.6, 101809.2, 101758.1, 101670, 101570, 101444.7, 101314.5, 101146.9, 
    100980.5, 100866.1, 100695.1, 100610.3, 100554, 100545.2, 100574.3,
  101833.1, 101727.3, 101775.2, 101705.6, 101613.9, 101516.9, 101362.1, 
    101235.4, 101087, 100977.3, 100832.5, 100717.5, 100583.6, 100546.9, 100590,
  100016.6, 99702.92, 101692.8, 101744, 101654.3, 101559.1, 101404.3, 
    101287.2, 101117.4, 101004.1, 100888.2, 100777.4, 100671.6, 100562.8, 
    100571,
  98019.2, 98073.39, 101571.3, 101786.3, 101695.1, 101629, 101500.8, 
    101374.6, 101224.5, 101099.3, 100998.9, 100853, 100759.4, 100596.7, 
    100589.3,
  98041.72, 98501.61, 100312.6, 101799, 101739, 101629.4, 101535.3, 101425.3, 
    101298.3, 101157.5, 101066.7, 100946.7, 100836.1, 100724.6, 100641.1,
  97405.85, 98908.8, 101701.6, 101812.2, 101755.5, 101627, 101638.1, 
    101525.4, 101406.5, 101250.6, 101135.8, 101024.4, 100949.8, 100858.6, 
    100714.9,
  101910, 101932.5, 101912.5, 101861.4, 101800.8, 99859.24, 101299.2, 101306, 
    101375.2, 101299.7, 101220.8, 101148, 101063.7, 100927.6, 100810.1,
  101937.8, 101896, 101899.2, 101802.7, 101615.7, 99109.35, 97156.88, 
    96184.73, 98732.16, 101384.5, 101321.2, 101238.1, 101192.3, 101054.9, 
    100946.9,
  101865.5, 101841.1, 101879.4, 101836.8, 96856.09, 98238.46, 99918.9, 
    101437.8, 101581, 101490.3, 101404.5, 101311.9, 101273.6, 101169, 101033.9,
  101812.9, 101812.1, 101845.1, 101768, 97377.96, 97585.77, 97022.04, 
    101508.8, 101674.1, 101546.2, 101509.1, 101386.6, 101358.2, 101273.1, 
    101158,
  101897.2, 101837.6, 101787, 101697.4, 101622.4, 101538.6, 101419, 101288.9, 
    101143.1, 101017.7, 100890.9, 100788.3, 100712.8, 100691.1, 100681.3,
  101813.9, 101727.4, 101770.5, 101712.8, 101619.1, 101538, 101422.6, 
    101294.3, 101137.5, 100995.7, 100835.2, 100712.8, 100632.4, 100635.9, 
    100657,
  99976.13, 99669.33, 101673.2, 101737.3, 101621.8, 101528, 101391.4, 
    101257.5, 101103.5, 100955.1, 100786.8, 100655.3, 100556.8, 100558.9, 
    100582.6,
  97960.09, 98083.7, 101581.1, 101747.6, 101625.6, 101534.4, 101417.5, 
    101281.5, 101112.7, 100945.2, 100782.5, 100644, 100519.1, 100494.5, 
    100540.2,
  98040.91, 98492.18, 100280.2, 101730.6, 101625.5, 101501.5, 101396.7, 
    101267.5, 101108.6, 100953.8, 100777.8, 100632.8, 100481.1, 100461.7, 
    100491.5,
  97406.32, 98900.53, 101669.4, 101723.9, 101611.9, 101458.8, 101445.7, 
    101337.5, 101176.4, 100991.6, 100798, 100587.9, 100465.2, 100437.6, 100454,
  101893.4, 101893.9, 101813.6, 101745, 101623, 99687.02, 101106.1, 101090.4, 
    101075.6, 100985.8, 100847.4, 100647.8, 100482.4, 100408.9, 100422.2,
  101913.4, 101853.3, 101809.8, 101713.2, 101409.5, 98907.3, 96913.98, 
    95940.86, 98407.39, 101015.5, 100878.9, 100676.8, 100525.6, 100406.9, 
    100410,
  101896, 101840.4, 101816.4, 101729.1, 96652.95, 98081.7, 99687.04, 
    101213.5, 101217.4, 101056.2, 100906.2, 100703.5, 100543, 100396.1, 
    100396.9,
  101864.6, 101815.3, 101795.8, 101695.1, 97238.95, 97435.32, 96727.98, 
    101241.1, 101285, 101088.2, 100948, 100747.5, 100562.8, 100382.1, 100351.5,
  102216.2, 102188.3, 102181.1, 102143.5, 102105.4, 102066, 102003, 101926.8, 
    101835.2, 101754.9, 101676.5, 101605.4, 101448.2, 101299.9, 101196.8,
  102113.6, 102058.8, 102139.6, 102124, 102071.7, 102030.4, 101982.9, 
    101923.9, 101837.9, 101765.9, 101635, 101536.8, 101442.8, 101353.4, 
    101257.4,
  100267.3, 100005.5, 102000.8, 102088.3, 102044, 102006.8, 101942.1, 
    101876.2, 101793.5, 101720.7, 101618.4, 101540.4, 101431, 101331, 101232.8,
  98182.75, 98287.08, 101824.3, 102081.8, 102029.7, 102018, 101954.3, 
    101875.9, 101781.7, 101697.2, 101595.2, 101528.5, 101441.2, 101350.2, 
    101270.6,
  98244.16, 98681.3, 100518.9, 102064.7, 102027.4, 101964.9, 101907.3, 
    101831.3, 101753.4, 101679, 101587.3, 101521.8, 101428.1, 101360.1, 
    101278.8,
  97603.75, 99132.95, 101948.4, 102049.6, 102013.9, 101921.7, 101929.1, 
    101850.1, 101748.2, 101653, 101564.7, 101461.5, 101436.2, 101379.6, 
    101298.4,
  102119.6, 102130, 102101.4, 102069, 102020.3, 100098.1, 101546.4, 101582, 
    101633.6, 101602.1, 101566, 101493.9, 101430.8, 101376.9, 101307.9,
  102151.7, 102106, 102094.7, 102019.4, 101814.2, 99299.87, 97330.77, 
    96352.36, 98868.37, 101606.8, 101591.6, 101508.6, 101438.7, 101378.9, 
    101326.1,
  102134, 102095.4, 102093, 102036.7, 97014.95, 98377.96, 100066.1, 101617.6, 
    101715.1, 101648, 101570.6, 101486.2, 101439.9, 101378.4, 101329.2,
  102112.5, 102084.2, 102066.8, 101968.6, 97541.48, 97732.73, 97106.88, 
    101592.5, 101741.4, 101589.7, 101559.7, 101489.4, 101452.8, 101382.7, 
    101333.9,
  102310, 102275.8, 102270.9, 102228.2, 102180.8, 102151.9, 102093, 102011.4, 
    101905.4, 101819.1, 101774.8, 101692.1, 101512.4, 101361, 101250.5,
  102211.8, 102153.9, 102229.2, 102209, 102173.9, 102129.9, 102070.6, 
    102003.2, 101918.3, 101831.1, 101714.2, 101601.4, 101503.6, 101397.9, 
    101298.4,
  100374.1, 100095.1, 102089.5, 102178.4, 102137.8, 102095.2, 102039, 
    101976.5, 101892.3, 101801.2, 101695.5, 101610.9, 101500.6, 101362, 
    101240.1,
  98300.67, 98390.81, 101924.4, 102156.6, 102113.5, 102118.2, 102066.6, 
    101989.4, 101903.2, 101779.9, 101680.6, 101601, 101525.4, 101375.6, 101258,
  98324.61, 98753.8, 100591.5, 102113.4, 102104.3, 102072.6, 102044, 
    101965.3, 101902, 101771.5, 101696.3, 101621, 101551.2, 101415.2, 101280.8,
  97658.3, 99175.85, 101994.4, 102110.3, 102107.7, 102044.5, 102070.4, 
    101988.8, 101908.1, 101788.1, 101699.4, 101603.9, 101606.7, 101512, 
    101364.7,
  102156.4, 102174.9, 102159.9, 102158.9, 102115.3, 100228.6, 101718.5, 
    101751.3, 101839, 101800.6, 101744.7, 101660.6, 101636.2, 101567.3, 
    101443.4,
  102197.1, 102188, 102189.5, 102125.2, 101941.8, 99450.17, 97493.18, 
    96541.68, 99098.57, 101826, 101772, 101689.8, 101644.3, 101589.5, 101485.9,
  102191.2, 102190.3, 102211.6, 102164.6, 97148.38, 98571.54, 100271.2, 
    101810.1, 101933, 101871.1, 101786.1, 101710.7, 101667.2, 101599.7, 101518,
  102198.8, 102206, 102219, 102157.3, 97712.22, 97940.22, 97328.72, 101842.9, 
    101991.6, 101867.8, 101831.4, 101740.4, 101687.9, 101615.4, 101562.4,
  102273.1, 102260.5, 102237.3, 102209.5, 102165.8, 102131.8, 102087.5, 
    102028.9, 101961.6, 101896.6, 101803.6, 101740.2, 101673.8, 101634.3, 
    101549.8,
  102214.6, 102157.8, 102222.9, 102201.9, 102155.8, 102123.9, 102086.8, 
    102028.5, 101960.8, 101893.3, 101790.5, 101722.4, 101665.6, 101618.7, 
    101576.1,
  100381.2, 100092.3, 102092.6, 102168.1, 102127.5, 102105.1, 102057.6, 
    101994.3, 101936.5, 101860.3, 101768.1, 101722.3, 101676.5, 101619, 
    101556.6,
  98325.34, 98425.9, 101931, 102154.6, 102112.8, 102110.6, 102062.2, 
    101994.3, 101932, 101845.5, 101778, 101730.3, 101690.2, 101617.9, 101567.1,
  98320.09, 98782.12, 100607.4, 102120.7, 102093.2, 102054.4, 102032, 101993, 
    101936.4, 101852.9, 101780.4, 101738.7, 101695.4, 101627.1, 101575.4,
  97624.66, 99137.25, 101954.1, 102075.5, 102059.9, 102014.6, 102063.5, 
    102001.9, 101934.5, 101856.8, 101776.2, 101692.6, 101706.5, 101656, 
    101591.6,
  102115.2, 102120.5, 102115.9, 102099.9, 102080.2, 100204.1, 101705.4, 
    101767.7, 101845.7, 101820.1, 101787.3, 101725, 101697.9, 101652.4, 
    101604.4,
  102150.6, 102105.8, 102105.3, 102051.5, 101898.1, 99432.34, 97478.95, 
    96548.42, 99093.56, 101849.2, 101818.7, 101737.2, 101709.5, 101664, 
    101619.6,
  102126.8, 102096.3, 102113.8, 102081, 97117.56, 98549.69, 100249.7, 
    101800.8, 101923.9, 101864.4, 101829.7, 101755.8, 101726.8, 101662.8, 
    101629.3,
  102130.5, 102102.9, 102110.7, 102056, 97655.9, 97902.08, 97306.12, 
    101842.7, 102004.1, 101889.7, 101875, 101774, 101733.9, 101669.6, 101636.7,
  102245.9, 102220.7, 102186.2, 102102.8, 102042.2, 102012.7, 101974.3, 
    101924.8, 101879.1, 101834.4, 101762.6, 101691.4, 101646, 101666.9, 
    101639.5,
  102189.3, 102131.9, 102170.6, 102118.3, 102049.9, 102009.9, 101974, 
    101923.1, 101870.4, 101822.1, 101731.4, 101713.2, 101666.5, 101668.4, 
    101659.8,
  100354.4, 100076.6, 102065.8, 102118.4, 102054.2, 101998.6, 101947.7, 
    101905.9, 101860.4, 101799.8, 101740.2, 101705.6, 101667.1, 101686.6, 
    101670.5,
  98291.55, 98396.26, 101948, 102128.6, 102073.6, 102054.5, 101979.7, 
    101932.9, 101854, 101795.1, 101768.5, 101738, 101693.9, 101692.6, 101696.5,
  98313.7, 98748.36, 100608.4, 102122.5, 102076.3, 102024.2, 101987.7, 
    101951.9, 101891.4, 101811.1, 101777.1, 101752.3, 101702.4, 101717.1, 
    101714,
  97642.67, 99134.76, 101986.7, 102086.8, 102079.9, 101984.6, 102007.1, 
    101963.6, 101895.4, 101838.4, 101794.6, 101732.4, 101740.9, 101747, 
    101737.9,
  102058.7, 102097.3, 102126.3, 102134.3, 102092, 100180, 101659.9, 101735.3, 
    101844.7, 101840.6, 101806.8, 101784.6, 101764.7, 101766.3, 101764.8,
  102169.5, 102125.3, 102138.5, 102095.2, 101928.2, 99428.13, 97471.26, 
    96573.76, 99138.09, 101866.2, 101849, 101807.2, 101791.6, 101787.5, 101791,
  102187.5, 102141.1, 102176.8, 102130.1, 97162.61, 98615.65, 100293, 
    101798.8, 101947.1, 101907, 101881.6, 101848.4, 101833.2, 101807, 101815.3,
  102224.3, 102213.1, 102195.8, 102138, 97721.81, 97969.12, 97378.09, 
    101907.4, 102047.9, 101960.5, 101947.2, 101902.3, 101880.3, 101831.6, 
    101842.3,
  102508.9, 102461.6, 102443.4, 102393.7, 102335.6, 102282, 102215.5, 
    102139.6, 102056, 101990.4, 101916.6, 101813.8, 101648.5, 101534.7, 101416,
  102375.6, 102332.7, 102407.1, 102371.4, 102314.7, 102261.2, 102198.8, 
    102133.8, 102053.7, 101980.1, 101892.9, 101809.5, 101709, 101606.2, 
    101512.7,
  100515.4, 100245.7, 102231.4, 102326.6, 102270.9, 102223.7, 102160.3, 
    102089.8, 102015, 101948.1, 101871.2, 101802.2, 101725.6, 101630.8, 
    101546.3,
  98429.08, 98517.58, 102049.3, 102282.6, 102224.8, 102206.9, 102143.2, 
    102077, 102001.6, 101927.2, 101850.6, 101798.3, 101747.1, 101650.7, 
    101600.6,
  98401.72, 98856.09, 100685.4, 102201.6, 102176.6, 102133.7, 102098.4, 
    102045.3, 101974.3, 101907.7, 101836.4, 101797, 101742.8, 101688.3, 
    101628.5,
  97695.12, 99195.38, 102006, 102141.7, 102113.5, 102057.5, 102088.1, 
    102038.5, 101971.5, 101905, 101819.8, 101740.7, 101751.7, 101725.7, 
    101665.5,
  102154.8, 102140.1, 102119.5, 102123.6, 102082.6, 100241.1, 101710, 
    101793.6, 101877.2, 101864.5, 101823, 101772.8, 101751.9, 101736.4, 
    101693.6,
  102157.2, 102098.3, 102069.2, 102031.2, 101898.5, 99406.1, 97475.92, 
    96577.96, 99068.13, 101817.2, 101801.6, 101755.1, 101734, 101739.3, 
    101719.1,
  102165.4, 102103, 102082.2, 102035.1, 97096.41, 98564.69, 100222.3, 
    101752.1, 101874.3, 101834.4, 101770, 101716.9, 101714.2, 101729.2, 
    101727.4,
  102237.9, 102182.9, 102130.2, 102036, 97626.38, 97901.66, 97296.73, 
    101805.5, 101900.1, 101778.6, 101723.1, 101670.6, 101684.8, 101713.8, 
    101727.1,
  102520.3, 102483.2, 102463.9, 102413.1, 102360.6, 102308, 102230, 102134.3, 
    102058.9, 101946.5, 101833.8, 101706.1, 101580, 101519.6, 101409.5,
  102495, 102398.1, 102452.8, 102403.9, 102357.9, 102301.2, 102224.7, 
    102136.1, 102048.8, 101934.1, 101821.8, 101707.6, 101611.5, 101532.4, 
    101423.5,
  100661.8, 100332.1, 102341.9, 102410.2, 102356.8, 102290.6, 102199.4, 
    102111.8, 102032.4, 101934.5, 101814.6, 101711.8, 101632.3, 101538.4, 
    101430.1,
  98656.82, 98721.29, 102228.5, 102420.3, 102362.1, 102311, 102209.9, 
    102117.2, 102027.8, 101933, 101842.1, 101745.4, 101661.7, 101557.8, 
    101461.7,
  98649.16, 99115.21, 100932.9, 102420, 102360.4, 102268.8, 102198.1, 
    102099.6, 102013.8, 101944.2, 101858.3, 101765.2, 101681.2, 101601.7, 
    101487.4,
  98022.71, 99530.41, 102335.9, 102408.3, 102358.5, 102224.6, 102234.2, 
    102129.4, 102031.8, 101961, 101876.3, 101734.7, 101712.3, 101653.1, 
    101532.6,
  102515.7, 102535.7, 102492.4, 102433.6, 102376.1, 100444.2, 101873.4, 
    101898.1, 101955.6, 101946.5, 101895.1, 101791.9, 101736.2, 101678.2, 
    101564.4,
  102562.2, 102514.7, 102478.6, 102390, 102160.9, 99657.34, 97671.96, 
    96710.05, 99214.2, 101938.8, 101909.2, 101813.9, 101751.1, 101703.8, 
    101603.1,
  102517.1, 102479, 102462.5, 102418.6, 97387.28, 98776.24, 100435.6, 
    101964.8, 102038, 101984.3, 101916.2, 101820.9, 101763.9, 101721.2, 
    101630.4,
  102511.7, 102488.8, 102473.5, 102395, 97944.16, 98152.8, 97492.88, 
    101969.8, 102094.1, 101974.4, 101925.2, 101836.4, 101774.2, 101726.7, 
    101661.4,
  102413.9, 102396.2, 102374.9, 102319.1, 102279.4, 102220.7, 102164, 
    102105.4, 102051, 101990.4, 101942.6, 101901.7, 101859.5, 101841.1, 
    101816.6,
  102388.8, 102336, 102401.2, 102339.3, 102303.2, 102240.3, 102172.3, 
    102103.8, 102050.9, 101992.3, 101937.9, 101893.5, 101873.6, 101866.5, 
    101863.7,
  100625.5, 100346.9, 102356.9, 102389.5, 102330.8, 102250.2, 102164.8, 
    102096.9, 102030.6, 101981.9, 101938.3, 101911.9, 101896, 101875.4, 
    101857.5,
  98617.19, 98738.49, 102263.2, 102416.2, 102355.1, 102304.1, 102205.4, 
    102121.7, 102043.1, 101992.4, 101948, 101929.4, 101909.9, 101873.4, 
    101875.6,
  98680.48, 99127.46, 100973.3, 102445.6, 102377.2, 102284.6, 102218.9, 
    102157.8, 102074.2, 102020.8, 101981.1, 101957, 101922.2, 101904.2, 
    101883.1,
  98041.88, 99568.77, 102378.6, 102447.3, 102388.2, 102263, 102248.1, 
    102190.3, 102139, 102071.8, 102006.3, 101931.8, 101952.1, 101928.4, 
    101899.6,
  102465.1, 102531.8, 102519.8, 102514.4, 102421.9, 100493, 101935, 101991.8, 
    102100.1, 102105.6, 102058.1, 102006.2, 101973.6, 101945.9, 101906.2,
  102524, 102542.9, 102544.8, 102491, 102242.4, 99752.73, 97757.86, 96858.31, 
    99407.06, 102141, 102103.7, 102035.4, 101997.2, 101953.6, 101911.8,
  102505.5, 102527.4, 102559.4, 102519, 97479.81, 98943.72, 100597.6, 
    102102.8, 102226.6, 102188.9, 102128.4, 102051.4, 102011.3, 101952, 
    101909.6,
  102518, 102539.4, 102570.6, 102507.6, 98084.45, 98305.7, 97657.21, 
    102190.6, 102311.7, 102201.6, 102156.3, 102066.4, 102017.1, 101949.7, 
    101901.6,
  101911.8, 101905.6, 101874.2, 101806.5, 101763.5, 101722.9, 101683.6, 
    101658.9, 101644.4, 101595.4, 101567.1, 101545.2, 101520.9, 101531, 
    101542.3,
  101849.8, 101792.5, 101842.8, 101788.1, 101732.2, 101655.9, 101602.6, 
    101584.6, 101560.1, 101531.2, 101501.9, 101467.4, 101460.3, 101486.1, 
    101528.9,
  100042.5, 99756.66, 101729.2, 101788.3, 101713.1, 101621.9, 101518.2, 
    101476, 101461.7, 101458.7, 101421.8, 101390.4, 101396.1, 101427, 101479.6,
  98021.04, 98127.26, 101630.9, 101779.9, 101715.5, 101643.2, 101504, 
    101402.8, 101398.7, 101379, 101351.7, 101328.1, 101335.6, 101367.2, 
    101446.7,
  98028.75, 98474.48, 100331.1, 101794.3, 101746.2, 101623.2, 101504, 
    101369.6, 101328.4, 101310.3, 101292.5, 101285.9, 101287.6, 101348.9, 
    101414.4,
  97434.56, 98912.38, 101723.4, 101796.1, 101762.2, 101588.8, 101542.6, 
    101397.2, 101322.1, 101282, 101233.1, 101193.2, 101268.1, 101329.2, 
    101387.9,
  101804, 101840.8, 101872.5, 101852.7, 101787.2, 99863.52, 101275.8, 101205, 
    101251.9, 101239.7, 101221.2, 101230.5, 101263.6, 101320.9, 101377.3,
  101885.4, 101872.4, 101892.1, 101868.2, 101644.7, 99051.82, 97045.01, 
    96129.98, 98614.53, 101270.2, 101242.2, 101247.3, 101275, 101324.7, 
    101380.8,
  101869, 101881.5, 101933.9, 101867.1, 96917.87, 98392.16, 99937.11, 
    101418.1, 101420.2, 101356.1, 101313.5, 101300.7, 101311.6, 101354.9, 
    101400.4,
  101923.6, 101943.1, 101996, 101917, 97532.34, 97712.61, 97044.27, 101583.2, 
    101599.8, 101489.2, 101410.2, 101390.6, 101393.7, 101408.7, 101438.9,
  102142.6, 102133.6, 102157.8, 102152.4, 102150.1, 102163.9, 102178.9, 
    102179.1, 102174.5, 102159.5, 102151.1, 102130.7, 102101.5, 102060.3, 
    102022.8,
  101939.8, 101918.5, 102018.4, 102044.5, 102030.8, 102044.3, 102066.6, 
    102091.5, 102101.3, 102094.9, 102083.2, 102062.5, 102037.4, 102016.9, 
    102006.2,
  99983.55, 99752.33, 101757.2, 101911.9, 101899.1, 101911, 101917.5, 
    101939.7, 101962.9, 101982.7, 101982.8, 101977.8, 101970.2, 101955.8, 
    101948.4,
  97828.95, 97935.15, 101492.3, 101775.3, 101768.1, 101804.8, 101810.9, 
    101827.8, 101844.8, 101869.2, 101877.9, 101881.3, 101880.2, 101871.2, 
    101894,
  97689.93, 98189.5, 100045.9, 101602.4, 101621.7, 101631, 101652.7, 
    101671.5, 101684.6, 101715.5, 101740.3, 101768.5, 101776.8, 101800.4, 
    101818.4,
  96998.73, 98506.95, 101293.9, 101440.1, 101447.4, 101444.2, 101540, 
    101560.9, 101570.8, 101592.3, 101601.5, 101599.6, 101682, 101720, 101744.7,
  101417.4, 101419.6, 101394.1, 101377.7, 101340.9, 99526.89, 101013.1, 
    101167.9, 101330, 101419.7, 101484.8, 101525.1, 101574.8, 101622.4, 
    101662.5,
  101405.8, 101330.6, 101300.2, 101249.5, 101074.5, 98627.15, 96719.04, 
    95875.45, 98385.96, 101224.5, 101335.5, 101398.8, 101459.6, 101522.7, 
    101576.6,
  101277.4, 101221.7, 101234.3, 101191.3, 96251.74, 97624.77, 99236.65, 
    100775.1, 100985, 101094.4, 101171.3, 101254.8, 101335.5, 101414.9, 
    101482.9,
  101176.3, 101134.4, 101151.5, 101099.4, 96722.19, 96891.66, 96277.3, 
    100686.1, 100899.2, 100873.2, 100998.1, 101090.4, 101199.6, 101302.2, 
    101391.2,
  102113.6, 102174.4, 102238.9, 102298.2, 102348.7, 102400.8, 102437.2, 
    102447.7, 102461.5, 102463.8, 102474.1, 102456.7, 102428.8, 102400.5, 
    102369.8,
  101983.7, 102038.6, 102165.9, 102230.1, 102266.1, 102333.4, 102383.1, 
    102427.1, 102438.2, 102448.9, 102443.7, 102434.6, 102417.4, 102397.9, 
    102390.5,
  100098.2, 99930.17, 101961.1, 102163.6, 102174.7, 102235.4, 102276.4, 
    102328.5, 102357.9, 102392.7, 102391.4, 102391.2, 102378.1, 102371.7, 
    102364.8,
  97962.48, 98108.52, 101714.4, 102063.6, 102095.7, 102168.8, 102207.2, 
    102256.8, 102285.2, 102315.6, 102326.8, 102340.2, 102339.1, 102330.8, 
    102346.1,
  97832.94, 98378.07, 100319.9, 101922.7, 101989.5, 102028.1, 102079.9, 
    102134.7, 102173.4, 102215.5, 102237.2, 102261.8, 102268, 102289.4, 
    102299.6,
  96973.8, 98612.93, 101516.8, 101782.8, 101842.6, 101882.8, 102009.3, 
    102051.5, 102077.4, 102117.6, 102136.1, 102132.8, 102211.8, 102243.8, 
    102262.2,
  101275.2, 101433.8, 101579.7, 101680.8, 101739, 99959.09, 101498.2, 
    101715.8, 101888.9, 101990.3, 102045.7, 102088.1, 102132.9, 102175.3, 
    102206.7,
  101293.4, 101338, 101444.7, 101487, 101431.2, 99043.27, 97203.11, 96396.53, 
    98975.66, 101872.7, 101958.5, 101998.1, 102043.6, 102097.3, 102146.3,
  101100.6, 101163.2, 101327.6, 101393.2, 96576.29, 97986.83, 99732.7, 
    101357.6, 101655.2, 101773.9, 101855.2, 101912.9, 101956.2, 102011.4, 
    102068.8,
  100949.7, 101020.4, 101167.5, 101196.5, 96930.51, 97209.17, 96794.96, 
    101389.1, 101698.2, 101644.1, 101749.9, 101795.8, 101869.7, 101926.8, 
    101989.9,
  101361.7, 101413.4, 101503.3, 101589.5, 101674.1, 101755.7, 101828, 
    101896.9, 101967.4, 102014, 102053.7, 102075.5, 102104.5, 102125.7, 
    102123.9,
  101279.2, 101351.3, 101484.8, 101579, 101667, 101763.5, 101842.5, 101915.5, 
    101974.7, 102026.4, 102063.1, 102089.3, 102128.1, 102148.4, 102165,
  99510.64, 99375.38, 101356.1, 101569.9, 101648.3, 101752.7, 101833.5, 
    101911.4, 101977, 102033.5, 102067.6, 102104.5, 102140.1, 102159.9, 
    102176.5,
  97458.46, 97686.34, 101222.5, 101545.6, 101632.1, 101756.9, 101842.5, 
    101923.3, 101985.3, 102035.4, 102070.4, 102112, 102147.9, 102160, 102190.7,
  97403.77, 97970.32, 99903.48, 101511.1, 101611.7, 101694.9, 101803.7, 
    101890.9, 101959.3, 102019.1, 102058.4, 102111.5, 102135.1, 102166.1, 
    102190.2,
  96691.6, 98275.09, 101157.6, 101451.8, 101567.3, 101655.2, 101805.5, 
    101895.6, 101950.5, 102006.3, 102044.7, 102054.8, 102143.9, 102176, 
    102199.4,
  100881.6, 101093.5, 101286, 101441.5, 101535.5, 99861.22, 101443.9, 
    101655.6, 101854.6, 101956.7, 102034.2, 102084.2, 102135.3, 102174.4, 
    102200.1,
  100999.8, 101080.5, 101230.2, 101332.3, 101356.4, 99015.41, 97264.59, 
    96514.71, 99110.3, 101930.8, 102022.8, 102065.7, 102113.7, 102165.2, 
    102198.2,
  100882.5, 100996.1, 101196.2, 101289, 96650.12, 98127.08, 99872.23, 
    101476.2, 101781.1, 101920.9, 101995.6, 102042, 102091.5, 102140.8, 
    102182.2,
  100843.6, 100965.5, 101136.1, 101196, 97055.05, 97411.61, 97038.36, 
    101587.9, 101884, 101871.7, 101968.4, 102009.6, 102078.2, 102119.4, 
    102163.5,
  101814.2, 101767, 101720.1, 101664.1, 101605.9, 101560.6, 101506, 101461, 
    101453.9, 101434.9, 101419, 101426.9, 101442.4, 101478.6, 101525.3,
  101679.6, 101613.7, 101651.4, 101619.9, 101555.2, 101519.5, 101467.1, 
    101414.4, 101410.8, 101399.6, 101379.3, 101380.9, 101388.2, 101442.3, 
    101506.4,
  99774.68, 99479.62, 101433.3, 101539, 101471, 101438.5, 101400.2, 101345.3, 
    101337.1, 101349.6, 101337, 101347.1, 101354.6, 101413.9, 101468,
  97693.35, 97722.12, 101237.6, 101460.4, 101408.6, 101387, 101355.1, 
    101310.9, 101290, 101305.2, 101299, 101316.8, 101324.8, 101371.7, 101448.1,
  97551.45, 98024.43, 99870.74, 101361.5, 101334.9, 101278.4, 101268.7, 
    101239.5, 101223.9, 101253.6, 101256.9, 101289.6, 101301.2, 101357.9, 
    101428.6,
  96779.1, 98338.57, 101125.4, 101263.7, 101230.2, 101165.9, 101214.2, 
    101200.5, 101181.1, 101206.6, 101216.4, 101214.5, 101294.7, 101357.4, 
    101426.3,
  101144.8, 101188.2, 101256.2, 101256.6, 101205, 99361.5, 100804.4, 
    100921.5, 101057.4, 101113, 101181.7, 101231.5, 101282.1, 101349.6, 101423,
  101206.4, 101174, 101208.9, 101148.3, 101002, 98520.05, 96655.93, 95813.27, 
    98317.41, 101077, 101146.5, 101207.5, 101265.7, 101346, 101428.4,
  101003.3, 101028.7, 101148.9, 101128.7, 96298.88, 97627.98, 99271.11, 
    100762.2, 100984.6, 101070.5, 101123.4, 101185.5, 101254.4, 101341.7, 
    101433.6,
  100894.3, 100947.8, 101056.3, 101018.2, 96730.9, 96944.43, 96455.16, 
    100861.3, 101065.3, 101022.2, 101114.8, 101166.5, 101259.8, 101341.6, 
    101444.1,
  101993.1, 102010.5, 102057.5, 102098.7, 102126.1, 102153.1, 102157.7, 
    102149.8, 102132.8, 102110.7, 102088.4, 102050.7, 102007, 101975.7, 
    101929.1,
  101900, 101903.8, 102019.4, 102050.5, 102067.8, 102103.3, 102122.6, 102132, 
    102116.7, 102099, 102063.9, 102024.8, 101986.2, 101961.7, 101932.7,
  100032.9, 99822.45, 101828.5, 102009.1, 101996, 102031.6, 102038.2, 
    102047.3, 102039.6, 102036.3, 102000.2, 101973.6, 101946.2, 101916.2, 
    101888.1,
  97893.26, 98020.21, 101613.2, 101937.1, 101932.4, 101981.6, 101988.4, 
    101998.4, 101985.9, 101969.6, 101948.8, 101929.2, 101905.5, 101872.9, 
    101861.3,
  97801.22, 98336.72, 100244.7, 101816.4, 101852.7, 101854.5, 101870.8, 
    101884.7, 101890.3, 101894.2, 101878.2, 101868.5, 101843, 101834.5, 
    101811.8,
  96974, 98594.2, 101459.7, 101705.1, 101714.1, 101735.9, 101821.8, 101830.2, 
    101815, 101821.2, 101800.5, 101762, 101802.5, 101797.4, 101778.6,
  101373.5, 101497.9, 101570.8, 101624.4, 101630.7, 99812.59, 101316.2, 
    101497.5, 101634.6, 101706.2, 101721.9, 101729.5, 101729.1, 101731.9, 
    101725.8,
  101362.6, 101401.1, 101463, 101454.8, 101363.6, 98940.54, 97061.29, 
    96235.96, 98752.13, 101608.1, 101651.8, 101650.8, 101647.8, 101655.5, 
    101658.9,
  101206.5, 101246.7, 101362.3, 101398.4, 96512.68, 97898.98, 99612.13, 
    101216.5, 101470.2, 101527.2, 101548.8, 101551.3, 101549.8, 101565.4, 
    101578.1,
  101086.2, 101116.1, 101228.9, 101218.2, 96914.52, 97174.02, 96726.38, 
    101255.8, 101531.8, 101419.6, 101463.7, 101442.9, 101456.6, 101469.5, 
    101492.9,
  101292, 101262.7, 101295.2, 101343.8, 101388.8, 101457.8, 101521.5, 
    101580.5, 101631.6, 101683.2, 101727.9, 101766.3, 101808.1, 101830.4, 
    101826.1,
  101324.9, 101271.4, 101358.1, 101390.1, 101447.4, 101510.3, 101564.7, 
    101621.3, 101675.9, 101722.8, 101756.4, 101796.8, 101831.5, 101856.6, 
    101873.3,
  99661.02, 99415.26, 101317, 101448, 101481.8, 101539, 101591.8, 101647.3, 
    101694.2, 101731.4, 101777.8, 101826, 101860.5, 101880.1, 101885.6,
  97699.52, 97797.62, 101299.3, 101514, 101531.1, 101605.5, 101644.2, 
    101691.1, 101722.7, 101761.8, 101807.4, 101854.1, 101886.8, 101890.3, 
    101917.2,
  97787.46, 98238, 100063.3, 101564.1, 101571.7, 101578.9, 101642.3, 
    101691.5, 101727.5, 101778.1, 101822.2, 101873.3, 101902, 101929.6, 101940,
  97091.46, 98632.45, 101450.6, 101601.7, 101592.5, 101613.7, 101701.4, 
    101739.7, 101761.3, 101808.3, 101845.3, 101848.3, 101931.6, 101958.7, 
    101970.9,
  101503.9, 101586.9, 101648.5, 101684, 101633.8, 99842.02, 101364, 101524.9, 
    101706.2, 101794.8, 101859, 101901.4, 101941.7, 101974.6, 101989.5,
  101639.4, 101583.5, 101642.7, 101612.6, 101545.5, 99055.76, 97252.16, 
    96461.55, 99028.41, 101809, 101887.7, 101919.3, 101959.4, 101986.2, 
    102005.3,
  101586.6, 101565.5, 101630.5, 101622.7, 96798.65, 98200.64, 99895.65, 
    101433.9, 101718.8, 101818.9, 101883.9, 101917.5, 101968, 101996.6, 
    102020.3,
  101564.6, 101578.9, 101619.7, 101567.1, 97255.68, 97532.64, 97112.43, 
    101605.6, 101854, 101791.6, 101882, 101901.8, 101965.5, 101994.3, 102023.5,
  100739, 100670.9, 100667.7, 100688.3, 100726.6, 100803.2, 100887, 100963.8, 
    101018.9, 101071.4, 101120.9, 101171.3, 101232.4, 101288.2, 101331,
  100628.8, 100586.1, 100597.7, 100619.2, 100643.5, 100718.9, 100810.8, 
    100905.9, 100987.8, 101047.8, 101099.1, 101159.2, 101227.1, 101295, 
    101365.5,
  98851.42, 98587, 100425.9, 100547.4, 100562.6, 100635.6, 100730.8, 
    100838.1, 100935.1, 101011.1, 101077.6, 101159.7, 101235.9, 101306.6, 
    101375.9,
  96921.41, 97010.29, 100332.3, 100507.9, 100507, 100588.6, 100674.2, 
    100787.4, 100890.4, 100978.1, 101056.7, 101154.3, 101237.5, 101303.5, 
    101394.8,
  96944, 97368.75, 99056.02, 100457.4, 100447.6, 100513.4, 100616.3, 100730, 
    100829.1, 100930.6, 101032.6, 101141.9, 101228.5, 101316.1, 101400.5,
  96465.42, 97849.02, 100451.6, 100440.9, 100403.5, 100448.8, 100579.6, 
    100703.9, 100808.5, 100915.5, 101011.1, 101085.5, 101234.7, 101328.5, 
    101413.7,
  100904, 100772.7, 100603.7, 100437.1, 100336.8, 98680.41, 100229.2, 
    100453.4, 100690, 100848.4, 101009.2, 101126.6, 101244, 101339.8, 101424.8,
  100967.4, 100806.9, 100639.5, 100366.5, 100154, 97790.95, 96129.25, 
    95445.88, 98047.87, 100825.3, 100996.7, 101130.2, 101252.6, 101351.6, 
    101439,
  101000.6, 100849.3, 100713.9, 100410.7, 95567.42, 96999.12, 98683.67, 
    100234.7, 100622.1, 100834.1, 100991.8, 101136.3, 101267.5, 101371.4, 
    101457.5,
  101042.6, 100937, 100836.5, 100525.1, 96113.41, 96351.88, 96011.41, 
    100498.6, 100780.8, 100827.4, 101002.7, 101148.1, 101290.3, 101394, 
    101480.6,
  101782.6, 101758.7, 101807, 101827.5, 101838.7, 101879.8, 101908, 101917.3, 
    101903.6, 101886.9, 101845.8, 101799.9, 101738.4, 101659, 101586.7,
  101548.2, 101544.7, 101681.1, 101713.7, 101714.9, 101756.9, 101790, 
    101817.6, 101817.3, 101804.9, 101777.5, 101737.7, 101682.5, 101623.7, 
    101578.7,
  99649.25, 99452.21, 101414.4, 101589.9, 101579.4, 101614.8, 101639.2, 
    101668.7, 101685.9, 101694.9, 101681.9, 101654.1, 101618.9, 101566.1, 
    101523.9,
  97539.59, 97704.64, 101196.3, 101486.7, 101468.8, 101512.8, 101528.5, 
    101550.7, 101559.3, 101572.4, 101565.2, 101557.2, 101535.2, 101492.8, 
    101478.9,
  97572.19, 98053.69, 99848.3, 101374.5, 101356.1, 101345.8, 101372.6, 
    101393, 101409.8, 101437.4, 101444.8, 101453.8, 101435.5, 101429.1, 
    101411.8,
  96885.46, 98437.7, 101216.2, 101344.6, 101274.5, 101239.9, 101300.4, 
    101309.7, 101304.1, 101321.3, 101318.1, 101300.5, 101356.8, 101364.1, 
    101357.7,
  101344.4, 101364.3, 101314.6, 101312, 101220.8, 99382.47, 100840.9, 
    100983.3, 101113, 101181.6, 101221.2, 101236.9, 101263.5, 101282.6, 
    101294.7,
  101319.9, 101276.8, 101269.4, 101189.7, 100998.3, 98530.91, 96630.12, 
    95780.77, 98278.21, 101068.6, 101131.6, 101137, 101167.3, 101199.8, 
    101229.3,
  101262.2, 101211.3, 101222.2, 101142.9, 96180.74, 97538.62, 99201.45, 
    100735.1, 100937.3, 100996.7, 101026, 101038.2, 101075.5, 101114.1, 
    101157.3,
  101196.5, 101147, 101149.8, 101031.9, 96680.12, 96848.27, 96318.32, 
    100757.6, 100982.5, 100880.6, 100924.6, 100933.7, 100985.7, 101029.2, 
    101085.5,
  101994.5, 102007.3, 102031.6, 102042.9, 102047, 102077.4, 102099, 102113.6, 
    102105.6, 102091, 102062.1, 102024.5, 101980.1, 101931.2, 101873.1,
  101844.1, 101826.7, 101926.9, 101952.8, 101952, 101976.9, 102004.7, 
    102026.2, 102027.3, 102015, 101993.3, 101961.3, 101918.7, 101886.7, 
    101858.9,
  99953.29, 99723.78, 101719.9, 101849.7, 101838.3, 101854.2, 101867.8, 
    101893.4, 101908.3, 101913.5, 101901.5, 101875.4, 101845.6, 101811.8, 
    101787.4,
  97860.8, 97997.9, 101507.7, 101756.6, 101732, 101768.7, 101770.8, 101785.3, 
    101787.5, 101794.9, 101782, 101777.3, 101754.8, 101731, 101731.3,
  97880, 98354.88, 100174.2, 101676.4, 101641.7, 101624.7, 101637.5, 
    101657.3, 101667.9, 101677.1, 101667.1, 101671.1, 101656.1, 101657.9, 
    101648.9,
  97237.98, 98735.47, 101535.7, 101641.5, 101574.2, 101530.5, 101586.4, 
    101578.6, 101574.6, 101578.1, 101557, 101530.1, 101581.1, 101593.2, 
    101591.6,
  101685.2, 101691.2, 101665, 101636, 101575, 99706.15, 101213.6, 101327.8, 
    101442.5, 101482, 101486.5, 101487.3, 101502.5, 101515.9, 101521.9,
  101687.4, 101640.2, 101637.7, 101574.4, 101382.5, 98907.32, 96953.68, 
    96080.09, 98627.76, 101413.8, 101438.9, 101422, 101427.7, 101443.4, 
    101459.3,
  101619, 101592.7, 101600.5, 101556, 96566.93, 97987.94, 99671.7, 101221.2, 
    101365.4, 101373.9, 101375, 101358.1, 101366.5, 101376.1, 101397.1,
  101568.9, 101553.9, 101554.1, 101482, 97098.52, 97311.97, 96725.44, 101248, 
    101424.9, 101320.2, 101333.4, 101304.5, 101314.6, 101318.3, 101337.6,
  101970.1, 101959.5, 101987.1, 102004.6, 102021.7, 102041.5, 102054.3, 
    102057.5, 102052.7, 102047.8, 102029.4, 102016.4, 101995.9, 101970.5, 
    101927.1,
  101856.8, 101835.7, 101938.1, 101949.3, 101943.3, 101964.2, 101982.3, 
    101996.6, 101995, 101989.3, 101980.6, 101968.4, 101943.2, 101930.2, 
    101925.2,
  100013.8, 99781.54, 101779.4, 101903, 101894, 101891.8, 101891.5, 101891.5, 
    101898.5, 101902, 101897.9, 101890.6, 101884.2, 101870.4, 101866.7,
  97950.87, 98100.92, 101605, 101862.8, 101843.6, 101840.9, 101819, 101811.5, 
    101797.8, 101796.9, 101791.8, 101796, 101801.2, 101798.9, 101822.8,
  97957.27, 98433.07, 100271.1, 101821, 101811.2, 101774.2, 101742.8, 
    101711.5, 101701.9, 101689.2, 101686.6, 101700, 101701.8, 101730.2, 101743,
  97290.93, 98812.3, 101672.7, 101800.2, 101788.6, 101703.9, 101743.5, 
    101687.7, 101638.3, 101614.8, 101571, 101557.7, 101629.6, 101660.8, 101682,
  101762.2, 101807.4, 101819.3, 101815.4, 101784.7, 99899.09, 101386.2, 
    101458.8, 101543.5, 101540.6, 101524.5, 101514.7, 101540, 101576.7, 
    101610.5,
  101776.6, 101790.2, 101805.8, 101785.3, 101574.7, 99090.45, 97107.31, 
    96197.94, 98730.3, 101491.3, 101493.1, 101459.7, 101465.8, 101501.1, 
    101543.8,
  101763, 101770.8, 101796.7, 101776, 96741.63, 98210.05, 99852.98, 101419.3, 
    101520.2, 101497.8, 101452.9, 101414.1, 101411, 101436.9, 101475.7,
  101756.8, 101757.5, 101784.8, 101729.3, 97316.4, 97525.24, 96878.16, 
    101424.2, 101550.8, 101461.8, 101412.9, 101372.2, 101361.4, 101384.9, 
    101421.2,
  102198.6, 102210.1, 102225.7, 102241, 102245.1, 102215.6, 102184.3, 
    102187.7, 102212.9, 102215.6, 102202.6, 102179.9, 102136.7, 102125.8, 
    102089.4,
  102107.2, 102091.2, 102188.8, 102195.9, 102199.6, 102216.4, 102218, 
    102215.2, 102204, 102208.7, 102198.3, 102175.8, 102135.6, 102128, 102112.2,
  100260, 100026.9, 102030.3, 102155.8, 102157.5, 102165.6, 102171.7, 
    102175.6, 102179.5, 102178.4, 102166.6, 102139.1, 102120.1, 102104.2, 
    102086.1,
  98183.84, 98315.2, 101838.2, 102103.8, 102102.7, 102120.7, 102123.7, 
    102133.9, 102147.1, 102143.5, 102129.5, 102118.9, 102094.9, 102070.3, 
    102075.5,
  98192.16, 98652.48, 100497, 102036.7, 102055, 102047.5, 102063.6, 102061.4, 
    102070.1, 102076.6, 102066.5, 102064.3, 102044.9, 102040.2, 102035,
  97478.19, 99000.97, 101837.5, 101987, 102006.4, 101978.1, 102060.4, 
    102049.9, 102043.2, 102031.6, 102006.5, 101966.5, 102017.1, 102020.2, 
    102015.9,
  101873.3, 101926.2, 101971.6, 102002.9, 102013.2, 100176.9, 101681.9, 
    101805.2, 101940.7, 101977.1, 101994.2, 101978.5, 101978.3, 101981, 
    101985.2,
  101930.2, 101957.2, 101985.2, 101980.3, 101821.3, 99380.92, 97447.54, 
    96577.31, 99124.94, 101919.1, 101949.9, 101942.7, 101936.9, 101945.9, 
    101954.1,
  101934.7, 101969.7, 102009, 102005.9, 97041.9, 98502.12, 100173.6, 101749, 
    101884.7, 101895.7, 101889.1, 101888.3, 101891, 101899.6, 101913.3,
  101951.6, 101986.2, 102022.3, 101989, 97586.2, 97828.41, 97224.77, 
    101767.9, 101928.8, 101846.4, 101836.4, 101814.9, 101831.4, 101845.8, 
    101868.9,
  102487.3, 102551.2, 102592.5, 102599.4, 102589.6, 102577, 102535, 102479.9, 
    102452.5, 102442.7, 102422.2, 102394.1, 102360.6, 102360.1, 102318.7,
  102395, 102405.8, 102527, 102561.4, 102570.1, 102579.9, 102567.5, 102540, 
    102482, 102458.2, 102431, 102417.1, 102381.8, 102376.4, 102359.1,
  100535, 100341.6, 102375.1, 102522.5, 102526.7, 102534.4, 102529.4, 
    102513.6, 102499.8, 102475.7, 102432.8, 102421.6, 102388.5, 102385.9, 
    102365.4,
  98443.16, 98603.08, 102127.4, 102449.9, 102475, 102504.1, 102504.4, 
    102502.3, 102488.7, 102469.5, 102438.6, 102422.9, 102403.6, 102381.8, 
    102371.3,
  98352.52, 98872.34, 100763.9, 102354.7, 102409.6, 102422.2, 102439.3, 
    102446.6, 102451, 102444.5, 102422.4, 102408.6, 102389.5, 102376.9, 
    102363.2,
  97511.19, 99118.69, 101999.9, 102246.3, 102319.7, 102313, 102420.6, 
    102421.8, 102415.4, 102404.4, 102378.9, 102336.2, 102381.2, 102377.3, 
    102367.8,
  101719.6, 101918.1, 102068.7, 102196.6, 102262.2, 100491, 102014.8, 102171, 
    102319.8, 102357.7, 102362.5, 102353.1, 102353, 102354.2, 102349.3,
  101755.7, 101860.8, 101994.6, 102084.8, 102009.2, 99658.91, 97777.8, 
    96924.04, 99476.91, 102296.8, 102324.7, 102317.6, 102312.8, 102326.1, 
    102329.3,
  101684.1, 101787.2, 101934.2, 102031.6, 97242.5, 98727.02, 100447, 
    102076.2, 102255.2, 102272.4, 102276, 102269, 102272.4, 102284.8, 102296.2,
  101608.9, 101728.3, 101870.1, 101924.6, 97700.83, 98011.77, 97498.23, 
    102045.3, 102271.6, 102212, 102238.7, 102226, 102240.1, 102247.2, 102263.2,
  102375.9, 102427.6, 102453.5, 102471.8, 102473.5, 102466.4, 102451.6, 
    102417.3, 102382.1, 102347.2, 102319.9, 102300, 102278.7, 102263.5, 
    102201.9,
  102332.4, 102341.3, 102438.8, 102471.6, 102492.1, 102503, 102483.6, 
    102457.3, 102431.4, 102387.7, 102342.9, 102327.7, 102311.2, 102302.5, 
    102269.1,
  100541.9, 100344.1, 102349.2, 102473.2, 102481.8, 102498.1, 102482.6, 
    102473, 102451, 102422.2, 102382.5, 102357, 102336.8, 102319.6, 102295.9,
  98487.04, 98625.7, 102149, 102442.1, 102467.3, 102500.4, 102502.4, 
    102495.6, 102470.3, 102441, 102410.8, 102395, 102378.4, 102342.6, 102334,
  98445.34, 98910.69, 100806.9, 102396.2, 102445.9, 102461.7, 102484.5, 
    102491.4, 102484.8, 102465.3, 102437.6, 102420.7, 102392.3, 102371.2, 
    102356.9,
  97631.98, 99210.15, 102032.2, 102288.5, 102383.7, 102379.9, 102485.9, 
    102493.7, 102494.5, 102470.2, 102443.9, 102389.9, 102422, 102407.4, 
    102384.7,
  101863.6, 102002.8, 102129.2, 102259.1, 102339.8, 100592.9, 102128.7, 
    102253.9, 102402.2, 102447.5, 102463.1, 102450.3, 102431.1, 102415.7, 
    102394.3,
  101939.9, 101955.5, 102067, 102157.4, 102105.3, 99743.27, 97882.59, 
    97035.43, 99605.95, 102406.8, 102447.4, 102448.1, 102433.4, 102421.6, 
    102404.7,
  101908.3, 101906.4, 102017.3, 102085.4, 97375.35, 98857.81, 100553.2, 
    102165.8, 102345.5, 102381.6, 102418.1, 102420.5, 102422, 102413.3, 
    102406.1,
  101862.9, 101913.3, 101956.3, 101974, 97816, 98102.74, 97596.38, 102133.7, 
    102350.1, 102321.4, 102375.9, 102388.3, 102409.7, 102406.8, 102405.7,
  101795.3, 101815.8, 101826.8, 101828.7, 101815.7, 101780.8, 101735.7, 
    101677, 101636.3, 101607.6, 101599.9, 101592, 101587.3, 101568, 101527.4,
  101781.3, 101790.1, 101880.7, 101891.8, 101884.9, 101861.4, 101831.4, 
    101797.8, 101763.9, 101729.2, 101708.3, 101699, 101688.3, 101670.8, 
    101650.3,
  100082.5, 99871.88, 101844.4, 101948, 101946.3, 101930.9, 101908.2, 
    101886.2, 101858.7, 101832.4, 101813.5, 101793.1, 101768.4, 101736.4, 
    101712.1,
  98110.2, 98291.59, 101787.4, 101995, 102001.5, 101999.9, 101983, 101970.3, 
    101948.1, 101934, 101914.4, 101895.1, 101873.2, 101823.6, 101806.6,
  98133.82, 98628.19, 100538, 102051.1, 102067.6, 102055.9, 102065.3, 
    102045.3, 102019.1, 102003.2, 101994.3, 101973.5, 101938.7, 101917.7, 
    101889.4,
  97533.71, 99043.11, 101887.7, 102059.7, 102094, 102030.5, 102116.9, 
    102114.9, 102104.4, 102077.3, 102052.4, 101999.9, 102032, 102003, 101970.1,
  101781.2, 101909.7, 102037.1, 102098.4, 102114.9, 100330.6, 101863.4, 
    101947.3, 102075.8, 102098.5, 102120.6, 102104.6, 102096.2, 102076.5, 
    102040.6,
  101921.8, 101958.2, 102051.3, 102096, 101955.4, 99492.36, 97643.98, 
    96821.52, 99407.68, 102149.3, 102165.6, 102159, 102156.3, 102140.4, 102113,
  101883.6, 101938.5, 102076.5, 102063.1, 97278.52, 98796.03, 100448.9, 
    102020.2, 102176.1, 102191.1, 102198.9, 102193.8, 102199.7, 102190, 
    102171.3,
  101910, 101965.4, 102098.1, 102058.5, 97818.88, 98095.05, 97534.88, 
    102072.4, 102236.3, 102198.7, 102208.7, 102216.7, 102234.5, 102231.3, 
    102216.5,
  101242.8, 101258.4, 101199.9, 101195.6, 101149.7, 101002.7, 100843.7, 
    100707.5, 100666.7, 100755.2, 100854.1, 100942.3, 101009.5, 101053.4, 
    101066.5,
  101150.9, 101148.8, 101175, 101190.3, 101125.6, 101007.8, 100836.5, 
    100678.7, 100630.8, 100687.9, 100775.4, 100868.6, 100941.5, 101005.4, 
    101051.1,
  99388.17, 99179.12, 101052.2, 101171.5, 101075, 100988.8, 100785.1, 
    100623.9, 100566.7, 100610.6, 100700, 100808.1, 100901.1, 100974.2, 
    101026.8,
  97401.21, 97569.36, 100931.1, 101159.5, 101074, 100994.2, 100787.4, 
    100625.4, 100555, 100577.4, 100637.6, 100749.3, 100852.9, 100927.7, 
    101011.4,
  97384.75, 97882, 99653.24, 101137.7, 101066, 100949.6, 100772.4, 100628.3, 
    100537.1, 100563.6, 100607, 100719.2, 100818.6, 100928.4, 101009,
  96771.12, 98260.64, 100989.3, 101110.1, 101060.4, 100885.9, 100793.6, 
    100662.6, 100577.9, 100588.1, 100603.7, 100661.5, 100821.9, 100935.1, 
    101015.3,
  101043, 101104.5, 101125.7, 101131.9, 101075.8, 99184.56, 100469.3, 
    100407.4, 100507.7, 100579.1, 100652.2, 100720.7, 100831.2, 100942.8, 
    101030.7,
  101128.9, 101127.3, 101147.3, 101148.6, 100897.9, 98340.91, 96333.62, 
    95439.59, 97956.87, 100623.5, 100704, 100762.7, 100861.8, 100953.2, 
    101049.3,
  101122.2, 101142.6, 101205.3, 101130.1, 96270.2, 97614.57, 99055.73, 
    100463, 100614, 100702, 100765.5, 100821.9, 100909.6, 100986.3, 101087.9,
  101179, 101214, 101228, 101123.2, 96822.7, 96907.58, 96203.91, 100619.5, 
    100764, 100780.3, 100830.7, 100895, 100977.7, 101050.4, 101143.9,
  101586.8, 101604.1, 101643.4, 101690.5, 101722.1, 101764.3, 101778.9, 
    101798.1, 101809.6, 101813.8, 101805.1, 101803.2, 101790.3, 101775.4, 
    101742.9,
  101506.1, 101515.9, 101616.9, 101659, 101696.9, 101746.6, 101775.3, 
    101797.7, 101803.9, 101811.9, 101804.3, 101799.6, 101789.3, 101783.7, 
    101772,
  99738.83, 99522.66, 101464.4, 101622.4, 101633.2, 101693, 101719.8, 
    101751.1, 101773.2, 101793, 101786.8, 101790, 101789.6, 101779.1, 101756.6,
  97726.96, 97841.35, 101278.6, 101573.3, 101589.5, 101650.5, 101685.2, 
    101721.8, 101737.7, 101753.8, 101756.2, 101768.3, 101770.1, 101754, 
    101763.2,
  97664.68, 98145.43, 99946.66, 101471.8, 101521.4, 101548.6, 101595.5, 
    101643.1, 101671.9, 101701.1, 101710.4, 101735.7, 101739.4, 101748.7, 
    101747.5,
  96899.85, 98408.27, 101165.4, 101364.4, 101413.2, 101446.5, 101559.3, 
    101595.9, 101614.8, 101646.7, 101643.9, 101637.2, 101708.4, 101727.6, 
    101733.6,
  101118.8, 101195, 101260.6, 101300.1, 101340.7, 99597.91, 101096.6, 101293, 
    101469.2, 101557.4, 101603.6, 101628.4, 101663, 101690.9, 101708.3,
  101073.2, 101071, 101121.3, 101138.9, 101070.6, 98738.15, 96945.71, 
    96155.44, 98644, 101441.8, 101529.2, 101565.1, 101604.6, 101644.4, 
    101674.9,
  100891.9, 100893.2, 100974, 101021.7, 96318.86, 97690.52, 99384.27, 100972, 
    101263.7, 101359.9, 101440, 101489.7, 101538.2, 101587.8, 101625.9,
  100767.1, 100750.8, 100808.8, 100795.3, 96648.56, 96900.27, 96501.45, 
    100928.2, 101274.7, 101233.4, 101350.9, 101397, 101463.6, 101516.4, 
    101564.5,
  101579.8, 101514, 101493.8, 101445, 101403.3, 101347.5, 101268.3, 101189.3, 
    101125.5, 101091.9, 101077.1, 101072.1, 101072.3, 101098.2, 101130.8,
  101537.1, 101505.3, 101547.5, 101515.6, 101495, 101464.1, 101417.2, 
    101363.1, 101310.1, 101260.3, 101221, 101201.1, 101180.1, 101185.4, 
    101208.4,
  99803.71, 99605.67, 101533.6, 101582.5, 101550, 101530.2, 101504, 101462.2, 
    101416, 101382.9, 101350.1, 101315.5, 101278.6, 101263.9, 101263.4,
  97892.12, 98010.38, 101456.1, 101645.8, 101610.7, 101600.8, 101590.4, 
    101575, 101531.8, 101494.1, 101475.2, 101432.4, 101387.1, 101342.7, 
    101352.4,
  97925.78, 98378.16, 100193.1, 101674.2, 101655, 101613.2, 101610, 101615.3, 
    101610.7, 101582.8, 101563.5, 101547, 101489.2, 101444.3, 101437.4,
  97250.67, 98744.82, 101517.9, 101661.1, 101655.4, 101604.3, 101668.8, 
    101660.5, 101661.9, 101654.2, 101629.3, 101580.3, 101588.1, 101536.7, 
    101523.7,
  101539.6, 101577.7, 101661, 101681.6, 101673.4, 99847.82, 101329.5, 
    101458.8, 101611, 101663.4, 101693.2, 101689, 101667.4, 101612.2, 101594.6,
  101604.9, 101557.6, 101617.4, 101602.5, 101495.8, 99105.34, 97248.97, 
    96411.27, 98928.03, 101670.3, 101732.1, 101736.2, 101727.3, 101676.8, 
    101662.4,
  101537, 101523.9, 101581, 101593.4, 96841.15, 98221.19, 99924.12, 101452.8, 
    101636.6, 101691, 101743.6, 101753.4, 101766.2, 101719.3, 101712.4,
  101489, 101506, 101557.1, 101515.6, 97297.7, 97540.3, 97081.84, 101517.6, 
    101741.3, 101674.6, 101742.6, 101754.9, 101782.5, 101751.5, 101745.5,
  101545.4, 101451.2, 101386.5, 101274.4, 101113.6, 100798.5, 100400.8, 
    100084, 99890.5, 99979.73, 100172.4, 100364.1, 100523.1, 100628, 100695.4,
  101526.3, 101381.4, 101420.5, 101306.9, 101180.9, 100953.5, 100637.4, 
    100224.5, 99904.14, 99826.9, 99941.88, 100142.6, 100335.7, 100489.8, 
    100616.3,
  99732.42, 99457, 101380.4, 101369.1, 101218.9, 101035.4, 100727.2, 
    100382.2, 100036.6, 99801.99, 99787.59, 99941.37, 100149.1, 100335.3, 
    100497,
  97813.58, 97933.45, 101281.8, 101417.9, 101287.3, 101173.4, 100908.6, 
    100591.9, 100239.7, 99948.54, 99785.29, 99833.26, 100009, 100201.5, 
    100411.8,
  97894.41, 98329.46, 100076.4, 101451.1, 101320.4, 101210.9, 101020.5, 
    100729.9, 100448.3, 100155, 99967.77, 99910.66, 99997.41, 100170.2, 
    100358.6,
  97339.93, 98799.86, 101478.1, 101483.9, 101348, 101218.4, 101189.6, 
    100946.2, 100688.7, 100394.9, 100126.7, 100003.6, 100081.1, 100205.8, 
    100359.3,
  101755.5, 101721.9, 101649.8, 101546.5, 101383.2, 99523.23, 100889.5, 
    100709.9, 100667.5, 100566.9, 100363.4, 100196.5, 100171.8, 100269.9, 
    100389.4,
  101800.8, 101698.8, 101661.8, 101546.4, 101229.2, 98767.1, 96866.98, 
    95890.3, 98289.25, 100817.9, 100596, 100389.1, 100283.4, 100335.3, 
    100433.3,
  101734, 101671.9, 101677.7, 101578.8, 96630.18, 97966.04, 99626.05, 
    101117.5, 101118.9, 100995, 100846.1, 100616.2, 100422.8, 100393.9, 
    100493.9,
  101653.8, 101635.2, 101662, 101555.2, 97208.34, 97364.31, 96726.88, 
    101209.2, 101282, 101142.3, 100997.2, 100816.3, 100619.1, 100516.7, 
    100561.3,
  101942.4, 101891.3, 101886.2, 101877.8, 101875.4, 101876.1, 101858.8, 
    101828.2, 101784.5, 101746.6, 101702.5, 101667.8, 101631.1, 101609.4, 
    101592.5,
  101918.2, 101839.2, 101906.5, 101869.5, 101857.6, 101841.7, 101802.8, 
    101769.4, 101720.6, 101676.7, 101621.4, 101575, 101530.9, 101516.9, 
    101518.1,
  100125.3, 99843.48, 101784.8, 101866.7, 101829.6, 101813.1, 101761.3, 
    101718.3, 101655.5, 101605, 101531.2, 101469.7, 101420.2, 101393.7, 
    101394.7,
  98200.5, 98261.32, 101673.2, 101930.2, 101850.8, 101816.7, 101743.1, 
    101679.7, 101603.7, 101528.4, 101435.3, 101358.1, 101287.8, 101243.2, 
    101264,
  98197.55, 98649.35, 100414.2, 101901.3, 101832.6, 101757.7, 101685.5, 
    101614.8, 101542.5, 101463.3, 101355.7, 101262.3, 101168.1, 101120.9, 
    101116,
  97582.97, 99041.88, 101772.5, 101879.1, 101795.6, 101669.7, 101675.2, 
    101588.4, 101492.4, 101398, 101275.1, 101132.9, 101077.5, 101019.7, 
    100990.6,
  102002.9, 101959.7, 101908.3, 101829, 101761.6, 99843.73, 101200.1, 
    101286.6, 101350.2, 101324, 101236.3, 101111.6, 101001.7, 100933.2, 
    100890.1,
  101914.4, 101792.9, 101774, 101675.8, 101473.9, 99002.53, 97078.06, 
    96107.29, 98538.8, 101227.2, 101176.9, 101047.7, 100942.5, 100878.2, 
    100831.5,
  101766.1, 101673.5, 101670.5, 101616.9, 96709.09, 97986.93, 99653.35, 
    101173.6, 101319.6, 101229, 101133.1, 100998.1, 100895.2, 100828.6, 
    100781.6,
  101685, 101586.7, 101572.1, 101468.1, 97152.45, 97326.27, 96747.7, 
    101121.7, 101284.7, 101121, 101069.6, 100929.6, 100813.5, 100741.4, 
    100708.4,
  101921.3, 101910.3, 101899.4, 101865.3, 101856.7, 101828.3, 101794.5, 
    101762.8, 101735.5, 101708.9, 101668.7, 101661.2, 101647.1, 101654.3, 
    101632.7,
  101933, 101886.9, 101958.7, 101919.1, 101901.8, 101875.8, 101840, 101809.2, 
    101777.9, 101751.5, 101700.7, 101678.3, 101655.1, 101657.6, 101651.7,
  100171.6, 99920.69, 101937.5, 101985.6, 101929.7, 101893.8, 101845.7, 
    101811.8, 101778, 101752.5, 101714.3, 101690.5, 101669.1, 101649.6, 
    101646.9,
  98223.27, 98349.59, 101847.1, 102034.1, 101957.7, 101914.8, 101861.8, 
    101820.6, 101782.8, 101747.2, 101717, 101702.6, 101681.2, 101647.9, 
    101656.3,
  98324.22, 98763.69, 100578.3, 102038.3, 101966.9, 101878.8, 101831.4, 
    101780.1, 101750.3, 101732.6, 101711.8, 101699.6, 101677.8, 101669.5, 
    101659.5,
  97748.2, 99234.09, 101994.2, 102036.9, 101956.9, 101818, 101841, 101771, 
    101726, 101706.8, 101682.4, 101637.3, 101674.1, 101669.4, 101654.5,
  102222.8, 102195.9, 102106.6, 102043.8, 101961.6, 100038.7, 101459.7, 
    101532, 101628.8, 101659.6, 101668.4, 101657.9, 101659.5, 101656, 101647.2,
  102242.2, 102166, 102093.3, 102012, 101715.1, 99232.32, 97289.38, 96384.34, 
    98862.96, 101622.1, 101655.9, 101638.9, 101631.6, 101631.4, 101616.8,
  102220.8, 102147.9, 102086.8, 102000.1, 96960.67, 98365.8, 99992.04, 
    101536.6, 101664.8, 101660, 101641.3, 101613.9, 101605.3, 101597.6, 101587,
  102213, 102135.6, 102081.7, 101956.2, 97519.84, 97701.79, 97057.96, 
    101525.7, 101649, 101581.2, 101589.6, 101562.2, 101559, 101543, 101538.8,
  101649.2, 101601.6, 101572.5, 101545.4, 101538.3, 101504.3, 101472.4, 
    101445.1, 101417.5, 101388.7, 101385.5, 101419.5, 101452.5, 101481, 
    101478.7,
  101675, 101623.7, 101647.5, 101601.7, 101593.2, 101568.1, 101538.2, 
    101502.5, 101466.2, 101428.9, 101415.9, 101436.5, 101470.4, 101501, 
    101529.9,
  99967.47, 99702.55, 101662.2, 101670.9, 101632.9, 101613.4, 101571.1, 
    101543.2, 101514.8, 101467.8, 101463.1, 101483.2, 101512.9, 101543.8, 
    101559.6,
  98007.52, 98121.34, 101618.4, 101772.6, 101696.1, 101677.3, 101625.1, 
    101587.5, 101546.5, 101513.6, 101512.8, 101528, 101555.1, 101556.9, 
    101597.6,
  98060.08, 98513.35, 100354.2, 101821, 101751.4, 101694.9, 101669.8, 
    101610.1, 101576.3, 101560.7, 101565.6, 101585.3, 101591.7, 101611.5, 
    101628.8,
  97452.48, 98946.87, 101734.1, 101836.1, 101776.3, 101683.2, 101712.9, 
    101652.2, 101613.6, 101610.5, 101596.3, 101578.6, 101641.1, 101658.1, 
    101658.7,
  101873.7, 101913.7, 101891.3, 101881.8, 101813.2, 99966.5, 101423.4, 
    101484, 101589.5, 101600.6, 101634, 101665.1, 101684.1, 101697.8, 101697,
  101975.5, 101933.6, 101897.7, 101851.5, 101665.9, 99168.42, 97274.8, 
    96429.55, 98950.12, 101653.2, 101673.1, 101695.1, 101716.8, 101724.1, 
    101722.9,
  101975.6, 101922.7, 101924.5, 101841.2, 96941.46, 98399.05, 100021, 
    101529.2, 101692.7, 101694.5, 101699.5, 101725.8, 101738.2, 101741.8, 
    101743.2,
  102011.3, 101949.4, 101953, 101835.5, 97462.98, 97734.42, 97165.88, 
    101660.4, 101780.5, 101714.7, 101730.4, 101745.7, 101760.8, 101765.4, 
    101757.4,
  101594.7, 101580.5, 101584.5, 101563.1, 101533, 101497.8, 101460.6, 
    101469.9, 101432.8, 101400.4, 101393.4, 101430.4, 101457.6, 101490.4, 
    101499.8,
  101582.9, 101552, 101607.6, 101573.1, 101522.8, 101486, 101454.3, 101450.9, 
    101424.4, 101416.4, 101399.4, 101432.9, 101474, 101522.3, 101559,
  99857.73, 99625.5, 101573.7, 101612.3, 101542.3, 101480.9, 101448.3, 
    101415.5, 101400.9, 101394.6, 101402.9, 101464.6, 101510, 101549.3, 
    101582.6,
  97929.62, 98052.58, 101510, 101640.8, 101561.9, 101503.2, 101452.8, 
    101390.5, 101379.4, 101400.3, 101437.3, 101489.7, 101535.7, 101568.3, 
    101622.1,
  98014.13, 98443.77, 100265.3, 101672.7, 101583.2, 101489.5, 101470.2, 
    101394.1, 101377.8, 101420.8, 101469.6, 101521.5, 101559.5, 101615.2, 
    101653.3,
  97475.46, 98925.16, 101650.5, 101681.3, 101609.1, 101460.8, 101515, 
    101452.8, 101443.5, 101477.4, 101510.7, 101513.4, 101620, 101667.8, 
    101697.6,
  101834, 101853.9, 101815.9, 101753.6, 101647, 99774.68, 101245, 101299.8, 
    101425.6, 101487.4, 101566.6, 101607.3, 101674.5, 101715.5, 101736.3,
  101953.2, 101904, 101862.9, 101741, 101522.2, 99034.64, 97127.77, 96294.97, 
    98860.69, 101557.4, 101604.5, 101653.4, 101714.2, 101755.9, 101775.5,
  101981.8, 101933.2, 101920, 101784.3, 96900.15, 98329.48, 99906.02, 101393, 
    101588.6, 101618.4, 101647.4, 101700.3, 101754.2, 101790.3, 101809.8,
  102055.4, 102002.3, 101980.2, 101845.3, 97485.27, 97726.45, 97085.9, 
    101551.5, 101711.5, 101663.6, 101697.4, 101744.2, 101798.4, 101831.3, 
    101853.5,
  101296.2, 101350.8, 101411, 101477.1, 101521.8, 101555, 101564.6, 101551.2, 
    101532.9, 101482.8, 101460.3, 101467.4, 101412.6, 101397.1, 101368.7,
  101227, 101263.2, 101385.3, 101434.4, 101484.9, 101531, 101550.6, 101559.9, 
    101539.7, 101500.4, 101459.2, 101445.7, 101421.5, 101417.7, 101381.9,
  99511.62, 99318.63, 101271.9, 101423.1, 101450.4, 101484.9, 101494.4, 
    101512.4, 101503.6, 101493.5, 101459.1, 101433.4, 101418, 101407.3, 
    101392.7,
  97563.73, 97706.13, 101163.7, 101419.6, 101429.5, 101462.7, 101477.8, 
    101502.1, 101489.5, 101491.5, 101452.2, 101432.5, 101409.3, 101391.6, 
    101414.1,
  97601.81, 98067.28, 99896.26, 101385.6, 101393.9, 101392.1, 101427.4, 
    101450, 101445.4, 101465.6, 101437.7, 101445.4, 101398.9, 101405.4, 
    101436.3,
  97012.36, 98470.45, 101212.4, 101346.7, 101345.3, 101311.6, 101409.2, 
    101441.8, 101426.8, 101450.8, 101407.5, 101396.2, 101412.2, 101425.4, 
    101452.8,
  101333.2, 101350.5, 101351.2, 101337.2, 101334, 99544.2, 101032.2, 
    101181.9, 101297.8, 101377.5, 101394.8, 101433.7, 101414.1, 101441, 101472,
  101444, 101373, 101346.8, 101273.7, 101118.2, 98725.61, 96901.87, 96104.38, 
    98568.6, 101322.7, 101368.6, 101410.6, 101413.1, 101452.5, 101485.6,
  101477, 101404.6, 101387.1, 101277.2, 96467.86, 97861.02, 99471.28, 
    101004.4, 101231.2, 101319.8, 101336.1, 101380.9, 101413.1, 101464.4, 
    101507.2,
  101539.5, 101468.6, 101424.8, 101296.4, 97008.48, 97174.79, 96611.06, 
    101024.9, 101279.4, 101260.2, 101311.6, 101357, 101421, 101479.1, 101533.6,
  101187.2, 101272.9, 101371.3, 101460, 101530.3, 101583.8, 101615.1, 
    101632.8, 101654.2, 101647.4, 101650.4, 101669.1, 101632, 101623.6, 
    101577.8,
  101157.4, 101218.7, 101373.8, 101459.8, 101534.8, 101597.4, 101637.9, 
    101665.8, 101682.4, 101657.6, 101670.3, 101696.3, 101653.6, 101636.6, 
    101611.8,
  99477.2, 99319.76, 101282.7, 101455, 101523, 101589.6, 101624.8, 101654.8, 
    101677, 101661.7, 101676.4, 101717, 101679.8, 101654.7, 101618.5,
  97535.04, 97722.35, 101164.5, 101445.1, 101514.7, 101588.4, 101634.2, 
    101670, 101685.9, 101679.7, 101679.2, 101734.1, 101701.3, 101657.5, 101642,
  97579.47, 98056, 99905.82, 101427.6, 101499.7, 101546.4, 101610.8, 101651, 
    101671.8, 101689.2, 101678.3, 101745.8, 101715.1, 101680.2, 101654.2,
  97014.01, 98427.27, 101183.5, 101384.8, 101467.4, 101494.2, 101625, 
    101663.5, 101679.3, 101688.6, 101665.1, 101705.2, 101734.6, 101700.8, 
    101667.2,
  101309.8, 101308.1, 101339.4, 101395.6, 101449, 99747.86, 101263.2, 
    101432.4, 101598, 101662, 101666.6, 101748.1, 101740.6, 101698.5, 101665,
  101445.9, 101393.2, 101389.7, 101352, 101281.4, 98946.78, 97181.98, 
    96365.88, 98865.22, 101630.4, 101658.3, 101731, 101736.7, 101693.9, 
    101654.7,
  101519.1, 101451.6, 101456.8, 101391.6, 96694.95, 98092.52, 99760.52, 
    101334.1, 101582.2, 101635.6, 101642.6, 101709.6, 101725.6, 101674.5, 
    101634.7,
  101625, 101553.8, 101542.2, 101422.3, 97192.78, 97457.55, 96960.27, 101349, 
    101612.7, 101573.3, 101615, 101675.7, 101705.6, 101649.6, 101616.1,
  100887.2, 100870.5, 100902, 100954.5, 101011.4, 101076.2, 101143.6, 
    101200.2, 101249.1, 101291.7, 101330.9, 101362.1, 101393, 101408.9, 
    101402.2,
  100821.2, 100823.5, 100926.2, 100957.8, 101029.4, 101114.8, 101195.2, 
    101250.2, 101293.3, 101333.3, 101371.7, 101399.9, 101429.5, 101446.9, 
    101451.9,
  99098.77, 98900.27, 100868.5, 100997.9, 101062.6, 101157.7, 101237, 
    101295.3, 101340.2, 101381.1, 101417, 101444.5, 101468.4, 101476.6, 
    101479.3,
  97096.79, 97291.23, 100798.2, 101004.7, 101094.5, 101194.4, 101282.9, 
    101349.5, 101393.9, 101430.7, 101461.9, 101486.9, 101504.8, 101501.9, 
    101524.6,
  97080.54, 97622.3, 99546.42, 101041.9, 101122.9, 101202.8, 101315.7, 
    101378, 101432.6, 101477.8, 101512.3, 101534.3, 101535.9, 101550.5, 
    101561.6,
  96493.72, 98027.4, 100850.6, 101045.8, 101141.7, 101193.1, 101371.9, 
    101453.9, 101503.5, 101535.7, 101553.2, 101536.3, 101598, 101603.4, 
    101598.7,
  100704.5, 100873.9, 101036.9, 101103, 101142.1, 99549.02, 101100.2, 
    101254.5, 101445.8, 101537.7, 101608.3, 101627.3, 101645, 101648.6, 
    101636.4,
  100923.4, 100960.2, 101066.5, 101093.9, 101025, 98709.27, 97031.96, 
    96302.52, 98886.48, 101585.8, 101646, 101672.9, 101687.4, 101688.1, 
    101676.7,
  100912.2, 100986.6, 101120.8, 101068.8, 96517.98, 98003.78, 99698.97, 
    101271.4, 101546.3, 101631.3, 101685.7, 101704.5, 101727.7, 101722.6, 
    101712.7,
  101012.1, 101080.1, 101171.2, 101095.8, 97015.77, 97352.3, 96955.35, 
    101439.9, 101664.5, 101667.2, 101713.6, 101739.4, 101764.3, 101761.5, 
    101749.1,
  100860.8, 100835.6, 100809.1, 100759.6, 100718, 100705.3, 100726.9, 
    100804.5, 100855.7, 100900.5, 100965, 100990, 101034.3, 101089.8, 101136.1,
  100704.9, 100707.2, 100788.1, 100745.4, 100689.1, 100677.2, 100703.3, 
    100782, 100846.9, 100891.7, 100949.1, 100978.8, 101044.6, 101108.3, 
    101168.1,
  98898.7, 98711.18, 100628.6, 100734.7, 100636.4, 100635.2, 100658.6, 
    100735.9, 100811.9, 100874.8, 100940.5, 100989, 101052.7, 101114.8, 
    101180.9,
  96867.22, 97037.88, 100485.2, 100721.3, 100618.1, 100607.3, 100633.7, 
    100703.3, 100792.4, 100864.9, 100940.5, 100989.1, 101050.6, 101106.7, 
    101198.1,
  96795.27, 97339.24, 99185.22, 100656.1, 100591.3, 100522.7, 100585.3, 
    100654.7, 100755.2, 100841.1, 100925.1, 100987.1, 101039.5, 101126.1, 
    101209.4,
  96133.6, 97668.86, 100452.4, 100616.7, 100545.3, 100461.3, 100559.7, 
    100636.7, 100735.4, 100827.4, 100890.9, 100928.6, 101047.3, 101138.3, 
    101226.1,
  100330.3, 100485.7, 100579.4, 100591.6, 100489.4, 98739.31, 100201.2, 
    100388.6, 100616.3, 100756.8, 100880.1, 100964.6, 101055, 101148.6, 
    101240.5,
  100390.5, 100438.6, 100508.2, 100474.6, 100292.1, 97881.45, 96153.05, 
    95431.96, 97958.16, 100711, 100858.5, 100958.8, 101062.4, 101158.4, 
    101254.6,
  100288.2, 100358.9, 100477.8, 100430.9, 95691.54, 97056.8, 98656.12, 
    100193.9, 100534.2, 100716.2, 100841.6, 100952.4, 101066.6, 101169.2, 
    101271.2,
  100288.9, 100333.1, 100442, 100362.1, 96132.67, 96374.53, 95968.22, 
    100366.7, 100657.7, 100703.9, 100839, 100954.3, 101078.3, 101183.9, 
    101289.3,
  101694.7, 101666.5, 101655.7, 101625.2, 101618.2, 101598, 101550.5, 101470, 
    101378.7, 101342.2, 101297.2, 101259.2, 101220, 101224.3, 101241.2,
  101607.9, 101545.6, 101633.1, 101613.6, 101596.7, 101591, 101563.8, 
    101527.4, 101455.1, 101387, 101337.6, 101291.3, 101252.3, 101244.4, 
    101276.4,
  99807.45, 99514, 101495, 101583.8, 101574.9, 101575.2, 101556.9, 101516.4, 
    101467.9, 101398.3, 101382.3, 101315, 101298.2, 101258.1, 101288.6,
  97814.45, 97875.46, 101323.8, 101561.5, 101563.3, 101574.2, 101565.8, 
    101543, 101507.3, 101431.1, 101421.9, 101347.4, 101335.5, 101270.1, 
    101305.5,
  97801.66, 98253.99, 100063.7, 101562, 101550.6, 101522.3, 101517.1, 
    101502.5, 101491.1, 101431.1, 101426.6, 101384.8, 101359.6, 101322.9, 
    101325.1,
  97161.17, 98686.19, 101408.9, 101556.1, 101535.5, 101475.5, 101521.4, 
    101506.8, 101493.5, 101448.3, 101415, 101367.5, 101388.3, 101365.2, 101342,
  101554.9, 101618, 101616.4, 101613.6, 101553.4, 99707.84, 101110.6, 
    101207.5, 101350.2, 101405, 101412.7, 101432.8, 101408.1, 101389.5, 
    101372.5,
  101625.4, 101586.8, 101611.6, 101529.2, 101372.3, 98940.66, 97056.37, 
    96181.27, 98642.22, 101357.7, 101392.9, 101417.3, 101417.3, 101405.6, 
    101397,
  101528.5, 101518.8, 101575.6, 101555.1, 96697.77, 98026.23, 99687.38, 
    101207.5, 101373.8, 101394.6, 101387.3, 101388, 101422.6, 101410.1, 
    101407.8,
  101468, 101464.3, 101517.6, 101460.3, 97173.31, 97367.38, 96853.92, 
    101244.8, 101466.2, 101366.1, 101398, 101367.2, 101411, 101408.7, 101417.3,
  101133.8, 101092.1, 101038.5, 100958.1, 100891.7, 100786.5, 100664.1, 
    100525.8, 100459.8, 100470.2, 100494.6, 100553, 100624.6, 100716.5, 
    100795.9,
  101082.4, 101025.7, 101059.7, 100970.2, 100887.8, 100792.1, 100691.2, 
    100560.1, 100456.5, 100450.2, 100467.5, 100530.4, 100617.7, 100719.1, 
    100815.6,
  99309.8, 99047.58, 100983.2, 101007.1, 100907.9, 100798.9, 100690, 
    100558.6, 100447.7, 100430.1, 100452.6, 100518.4, 100622, 100722.9, 
    100821.2,
  97342.03, 97453.09, 100884.3, 101036, 100937.2, 100845.5, 100740.2, 
    100593.5, 100460.1, 100420.1, 100441.6, 100512.6, 100621.9, 100712.8, 
    100832.7,
  97359.91, 97821.73, 99624.3, 101050.4, 100974.6, 100850.9, 100753.9, 
    100605.6, 100452.3, 100414.2, 100425.3, 100509.5, 100612.3, 100732.6, 
    100846.6,
  96727.9, 98204.57, 100979.5, 101056.3, 100996.8, 100858.1, 100819.4, 
    100686.7, 100507.1, 100428.5, 100408.2, 100450.6, 100612.2, 100741.8, 
    100862.5,
  101006.5, 101103.2, 101123.6, 101106.1, 101029.5, 99167.89, 100526.6, 
    100474.7, 100481.9, 100434.3, 100440.8, 100500.7, 100616.8, 100749.9, 
    100872.6,
  101087.9, 101114.8, 101129.4, 101094.7, 100901.1, 98399.5, 96432.66, 
    95574.09, 97988.27, 100520.2, 100490.3, 100522.1, 100621.4, 100756.5, 
    100880.4,
  101059.7, 101106.7, 101152.7, 101097.9, 96238.24, 97691.16, 99259.04, 
    100714.9, 100723.2, 100585.6, 100516.9, 100558.7, 100637.7, 100760.1, 
    100881.8,
  101097.8, 101137.6, 101181.3, 101112.8, 96820.39, 97034.47, 96408.52, 
    100858.1, 100868.3, 100640, 100563.9, 100588.5, 100661.7, 100769.4, 
    100885.4,
  101207.5, 101227.7, 101285, 101315.2, 101327.2, 101332, 101309.5, 101272.4, 
    101223.6, 101179.2, 101135.2, 101096.3, 101053.6, 101022.8, 100994.6,
  101065, 101083.7, 101211.1, 101249.1, 101261.1, 101277.7, 101263.2, 
    101237.5, 101197.3, 101152, 101101.3, 101065.8, 101037.3, 101024.9, 101013,
  99243.91, 99059.52, 101009.5, 101187.1, 101184.9, 101212.5, 101189.6, 
    101169.9, 101139.3, 101108.5, 101073.9, 101051.5, 101017.1, 101002.2, 
    100992.9,
  97192.81, 97321.8, 100772.4, 101103.3, 101111.7, 101149.9, 101148.2, 
    101136.1, 101105.7, 101072.9, 101040.6, 101019.2, 100995.1, 100973, 
    100981.6,
  97140.15, 97624.1, 99445.1, 100984.3, 101035.2, 101040.4, 101056.1, 
    101051.4, 101032.3, 101010.5, 100996.6, 100978.7, 100958.3, 100957.4, 
    100957.4,
  96390.95, 97896.79, 100655, 100886.5, 100931.2, 100931, 101015.6, 101017.1, 
    100988.7, 100963.5, 100934.2, 100889.5, 100933.6, 100937.3, 100940.6,
  100615.9, 100688.5, 100770.4, 100833.4, 100871.1, 99123.05, 100550.6, 
    100690.2, 100815.8, 100868.7, 100884.8, 100869.1, 100876.2, 100895.9, 
    100914.1,
  100715.2, 100678.9, 100718.1, 100702.7, 100632.8, 98290.7, 96459.91, 
    95606.08, 98063.16, 100788.2, 100830.8, 100811.9, 100816.2, 100840.5, 
    100881.7,
  100608.2, 100608.9, 100674.9, 100682.1, 95965.46, 97329.62, 98993.16, 
    100529.4, 100731, 100765.8, 100747, 100732.9, 100743.4, 100776, 100836.4,
  100552.3, 100581.7, 100635.3, 100598.8, 96400.79, 96648.44, 96164.02, 
    100540.2, 100773.3, 100673.9, 100681, 100663.4, 100687, 100718.3, 100793.2,
  101688.3, 101668.5, 101671.6, 101664.5, 101673.5, 101678.2, 101665.9, 
    101641.2, 101607.1, 101536.8, 101508.2, 101443.1, 101417.1, 101384, 101317,
  101593.4, 101561.2, 101641.7, 101635.3, 101630.6, 101651.4, 101651.9, 
    101639.5, 101614.5, 101570.2, 101530.8, 101482.6, 101442.3, 101419.7, 
    101365.6,
  99784.31, 99530.09, 101484.9, 101604.2, 101578.1, 101598.2, 101598.3, 
    101592.1, 101585, 101559.6, 101529.5, 101495.1, 101453.2, 101433.7, 
    101384.9,
  97784.58, 97857.9, 101287.5, 101555.5, 101536.8, 101561.1, 101574.5, 
    101581.3, 101573.9, 101548.6, 101531, 101496.7, 101471.2, 101427.8, 
    101412.6,
  97719.73, 98207.68, 99988.93, 101465.9, 101476.6, 101474.3, 101497, 
    101513.6, 101527.8, 101520.2, 101508.3, 101489.5, 101467.7, 101447.5, 
    101422.1,
  96996.01, 98502.09, 101264.8, 101424.4, 101402.2, 101396.7, 101494.8, 
    101501.4, 101493.4, 101500.2, 101469.5, 101431.1, 101468.9, 101459, 
    101422.2,
  101366.7, 101410.3, 101444.3, 101437.2, 101421.9, 99606.21, 101050.4, 
    101225.1, 101372.3, 101436.7, 101453.3, 101450.9, 101448.9, 101444.7, 
    101425.1,
  101411.8, 101383.4, 101406, 101331.6, 101211.1, 98840.49, 96985.54, 
    96152.78, 98620.01, 101365.8, 101424.9, 101420.9, 101421.8, 101421.7, 
    101409.3,
  101323.4, 101302.7, 101356.3, 101333.9, 96545.76, 97862.73, 99541.41, 
    101072.3, 101275.7, 101338.2, 101383.5, 101372.6, 101387.2, 101387.4, 
    101380.1,
  101258.9, 101255.9, 101294.1, 101233.1, 96970.87, 97187.85, 96733.21, 
    101122.8, 101366, 101275.2, 101339.8, 101328.2, 101355.6, 101354.7, 
    101362.6,
  101776.8, 101743.9, 101734.7, 101695, 101668.5, 101625.9, 101570.7, 
    101516.6, 101457.2, 101401.1, 101355.6, 101328.8, 101303.1, 101321.4, 
    101263.5,
  101747.8, 101668, 101757.7, 101719.5, 101696.7, 101662.1, 101622.3, 
    101578.5, 101525.5, 101474.2, 101428.3, 101393, 101359.8, 101379.1, 
    101323.3,
  99980.8, 99710.05, 101692.2, 101764.1, 101720.1, 101692.2, 101648.6, 
    101606.1, 101560.7, 101520.7, 101479.2, 101444.6, 101400.1, 101380.7, 
    101395.6,
  98014.45, 98124.77, 101571.6, 101795.7, 101739.6, 101715.4, 101682.8, 
    101653.5, 101604.1, 101561.9, 101528.1, 101497.2, 101464.8, 101409.7, 
    101407,
  98026.5, 98510.77, 100319.5, 101800.3, 101756.3, 101700.1, 101679, 
    101656.1, 101623.1, 101597.5, 101563.7, 101537.2, 101497.4, 101469.8, 
    101445.1,
  97400.88, 98935.22, 101685.5, 101799.2, 101755, 101661.9, 101711.3, 
    101692.6, 101650.8, 101620.1, 101588, 101527.1, 101549.5, 101521, 101485.6,
  101802.4, 101857.6, 101859.7, 101834, 101795, 99917.4, 101321.8, 101441.9, 
    101602.3, 101632.4, 101629.2, 101601.6, 101580.8, 101558, 101518.9,
  101921.3, 101870.1, 101866.5, 101774, 101585.2, 99177.61, 97299.5, 
    96390.67, 98855.3, 101631.8, 101649.5, 101626.1, 101605.7, 101575.5, 
    101547.8,
  101877.4, 101834.1, 101856.3, 101799.8, 96951.72, 98246.48, 99924.02, 
    101452.4, 101654.5, 101670.7, 101675.1, 101641.1, 101630, 101598.2, 101563,
  101879, 101839.9, 101848.2, 101744.5, 97434.58, 97601.47, 97106.31, 
    101472.6, 101710, 101620.9, 101670.8, 101638.9, 101640.5, 101607.4, 101583,
  101963, 101874.5, 101857.3, 101766.4, 101707.9, 101593.9, 101459.3, 
    101420.6, 101331, 101251.1, 101175.9, 101046.2, 100945, 100917.3, 100899.5,
  101971.2, 101841.6, 101924.2, 101832, 101777.5, 101705.7, 101591.8, 
    101482.2, 101434.4, 101379.2, 101330.2, 101255.6, 101142.9, 101048.9, 
    101004.1,
  100221.6, 99925.6, 101912.3, 101929.8, 101836.5, 101770.2, 101686.3, 
    101568.1, 101497.4, 101469.7, 101384.7, 101348, 101280.2, 101177.6, 
    101115.5,
  98365.45, 98421.87, 101832.5, 102009.1, 101894.3, 101829.7, 101753, 
    101698.5, 101574.7, 101530.7, 101515.9, 101434.2, 101390.3, 101308.5, 
    101232.6,
  98462.74, 98875.17, 100624.5, 102056.4, 101949.2, 101845.8, 101770, 
    101715.5, 101664.2, 101587, 101562.4, 101546.9, 101455, 101419.4, 101357.8,
  97938.17, 99367.17, 102058.1, 102102.7, 101980.8, 101805.1, 101835.4, 
    101758.3, 101710.6, 101664.2, 101592.9, 101551.3, 101563.6, 101488.6, 
    101466.8,
  102415.2, 102360.7, 102272.8, 102176.1, 102041.9, 100084.3, 101442.1, 
    101548.4, 101667, 101691.7, 101653.7, 101628.7, 101627.2, 101582.4, 
    101496.3,
  102491.3, 102383.3, 102312.7, 102178, 101846.5, 99383.55, 97427.58, 
    96492.79, 98989.44, 101716.6, 101714.1, 101658.1, 101652.4, 101633.1, 
    101586.2,
  102499.2, 102409.4, 102361.4, 102247.1, 97211.95, 98549.82, 100139.8, 
    101668.9, 101825.3, 101750.6, 101729.2, 101704.6, 101673.2, 101657.3, 
    101635.2,
  102511.1, 102430.1, 102384, 102242.1, 97784.88, 97970.47, 97340.07, 
    101719.2, 101903.1, 101774.4, 101751.3, 101712.7, 101694.4, 101675.4, 
    101668.5,
  102291.9, 102194.9, 102133.3, 101992.6, 101884, 101745.8, 101616.8, 
    101490.5, 101399.3, 101305.9, 101195.2, 101047.8, 100949.8, 100922.9, 
    100914.9,
  102307.6, 102176.4, 102221.5, 102098.1, 101996.9, 101870.4, 101742.6, 
    101609.4, 101496.2, 101418.8, 101345.1, 101260.6, 101119.5, 100977.6, 
    100979.6,
  100552.9, 100255.2, 102223.4, 102204.2, 102070.2, 101951.9, 101833.7, 
    101721.2, 101579.6, 101501, 101421.2, 101366.6, 101297.4, 101139.3, 
    101007.9,
  98666.06, 98765.13, 102145.8, 102292.1, 102147, 102044.8, 101940.9, 101845, 
    101710.8, 101594.5, 101535.3, 101464.8, 101412.7, 101296.5, 101147.5,
  98757.47, 99181.67, 100942.4, 102341, 102193.9, 102069.2, 101995.1, 
    101929.4, 101804.1, 101702.9, 101604.1, 101579.2, 101494.7, 101439.9, 
    101327.2,
  98222.24, 99701.11, 102371.1, 102387.5, 102221.9, 102045.1, 102075.5, 
    102034.9, 101940.1, 101806.4, 101700.6, 101587.1, 101612, 101553.1, 
    101453.5,
  102669.9, 102659.2, 102541.8, 102467, 102268.1, 100348, 101766.3, 101869, 
    101940.1, 101885.3, 101813.2, 101710.6, 101680, 101641.2, 101562.2,
  102750.6, 102678.4, 102605.4, 102492.5, 102099.2, 99666.16, 97697.33, 
    96840.91, 99331.37, 101982.4, 101910.7, 101824.6, 101731.7, 101718, 
    101675.2,
  102768.2, 102695.7, 102660.8, 102540.4, 97450.28, 98903.35, 100457.2, 
    102078.9, 102161.7, 102074.7, 101988.3, 101903.7, 101826.4, 101742.1, 
    101739,
  102783.8, 102731.7, 102705.9, 102564.2, 98101.72, 98306.31, 97600.82, 
    102118.4, 102225.7, 102116.5, 102059.2, 101971.7, 101903.7, 101825.2, 
    101756.4,
  102020.4, 101966.1, 101921.8, 101847.4, 101786.2, 101697.1, 101608.5, 
    101515.2, 101436.2, 101376.7, 101328.7, 101289.1, 101251.1, 101207.6, 
    101180,
  102039.1, 101961.5, 102004.9, 101939.4, 101894.3, 101816.8, 101736.2, 
    101656.3, 101571.4, 101496.9, 101432, 101393.4, 101364.5, 101296.5, 
    101246.7,
  100341.3, 100081.7, 102018.3, 102035.1, 101976.3, 101918.4, 101838.3, 
    101759.9, 101681.2, 101608.8, 101547.5, 101485.4, 101438, 101372, 101326.7,
  98399.7, 98559.57, 101970.7, 102123.1, 102058.2, 102013.6, 101955.1, 
    101884.1, 101807.6, 101729.6, 101658.8, 101587.6, 101529.7, 101433.7, 
    101385.8,
  98451.64, 98904.14, 100754, 102186.8, 102126.5, 102063, 102023.4, 101958.3, 
    101895.1, 101832.6, 101767, 101692.2, 101615.4, 101547.1, 101479.2,
  97887.99, 99365.95, 102140.7, 102209.4, 102162.6, 102042.1, 102118.5, 
    102073.8, 102019.2, 101936.3, 101861.7, 101754.1, 101726.4, 101657.5, 
    101587,
  102157.5, 102255.7, 102281.4, 102267.7, 102192.2, 100397.9, 101850.1, 
    101876.8, 101972.8, 101994.7, 101965.8, 101904.1, 101830.4, 101751.3, 
    101682.1,
  102282.8, 102290.3, 102291.5, 102271.4, 102058.7, 99627.71, 97771.29, 
    96931.98, 99440.91, 102086.8, 102059, 102003.2, 101929.4, 101849.2, 
    101768.1,
  102251, 102265.5, 102315.9, 102244.8, 97449.39, 98963.13, 100551.3, 
    102112.7, 102197.8, 102183.8, 102146.4, 102089.5, 102023.5, 101946.6, 
    101862.7,
  102277.6, 102288.4, 102346.2, 102263.2, 98014.93, 98282.38, 97709.04, 
    102216.5, 102310.3, 102255.8, 102210.5, 102162.4, 102108.5, 102036.3, 
    101956.1,
  101332.6, 101257.5, 101200.8, 101125.6, 101080.2, 101049.5, 101045.3, 
    101056.1, 101090.5, 101136.9, 101189.9, 101230.6, 101275.3, 101311.1, 
    101331.2,
  101409.1, 101321.6, 101332.3, 101255, 101199.8, 101161.3, 101147, 101140.7, 
    101154.5, 101190.7, 101236.9, 101278.4, 101322, 101354.1, 101375.5,
  99794.99, 99526.89, 101399.3, 101391.6, 101324.9, 101271.9, 101246.4, 
    101232.4, 101233.3, 101255.7, 101294.4, 101334.7, 101366.8, 101386.4, 
    101409.4,
  97971.95, 98089.31, 101423.1, 101534.8, 101462.1, 101412.9, 101370.3, 
    101345.6, 101330.9, 101340.2, 101364.5, 101398.2, 101420.5, 101425.3, 
    101466.1,
  98069.06, 98491.8, 100273.7, 101662.5, 101593.7, 101534.5, 101503.8, 
    101469, 101444.2, 101442.5, 101452.8, 101482.2, 101495.3, 101503.4, 
    101516.4,
  97539.46, 98961.13, 101666.5, 101732, 101689.4, 101591.1, 101663.1, 101632, 
    101598.8, 101572.4, 101555.6, 101525.3, 101593.5, 101603, 101599.7,
  101734.8, 101814.1, 101858.3, 101834.5, 101762.5, 99987.99, 101443.2, 
    101519.1, 101644.4, 101667.6, 101688.1, 101676, 101689.5, 101685.8, 
    101682.2,
  101863.4, 101861.8, 101888.5, 101861.2, 101662.8, 99240.03, 97414.85, 
    96616.61, 99159.71, 101809.5, 101800.9, 101784.9, 101779.4, 101776.1, 
    101772.3,
  101793.9, 101835.9, 101922.5, 101880, 97159.73, 98614.97, 100225, 101760.5, 
    101920.2, 101928.4, 101912.6, 101880.1, 101868.4, 101855.9, 101846.8,
  101789.5, 101852.5, 101937.5, 101892.6, 97711.36, 97963.12, 97445.01, 
    101926.1, 102073.6, 102021.1, 102008.2, 101974.4, 101956.8, 101934.4, 
    101919.7,
  100909.8, 100849.5, 100830.1, 100819, 100808.8, 100820.6, 100843.2, 
    100901.7, 100980.1, 101050.8, 101113.2, 101163.4, 101215.5, 101265, 
    101287.5,
  100943.4, 100858, 100907.4, 100882.5, 100872.8, 100872.7, 100893.7, 
    100939.9, 101005.8, 101071.8, 101132.7, 101194.9, 101254.4, 101295.2, 
    101317.3,
  99328.2, 99070.62, 100942.1, 100976.2, 100900.6, 100892.3, 100912.6, 
    100959.5, 101021, 101091.4, 101163.2, 101235.1, 101292.9, 101329.4, 
    101353.9,
  97581.15, 97711.76, 100959, 101065.6, 100946, 100927.4, 100943, 100987.7, 
    101046.4, 101115.7, 101190.5, 101265.5, 101322.2, 101347.9, 101394.8,
  97810.84, 98194.1, 99854.15, 101170, 101013.5, 100924.8, 100950.8, 
    100994.1, 101054.1, 101128.4, 101216.8, 101297.7, 101351.2, 101402.8, 
    101440.8,
  97487.61, 98806.23, 101337.6, 101255.6, 101083.2, 100927.1, 100995.1, 
    101019.4, 101082.7, 101147.8, 101221.9, 101266.4, 101387.6, 101444.3, 
    101483.6,
  101877.9, 101717.2, 101558.5, 101400.9, 101171.1, 99344.43, 100738.2, 
    100839.3, 101017.6, 101137.7, 101257.7, 101342.5, 101424.8, 101484.6, 
    101526.4,
  101955.3, 101804.2, 101673.7, 101468.8, 101078.5, 98635.22, 96814.41, 
    96023.95, 98485.53, 101178.6, 101292, 101387.1, 101463, 101523.6, 101567.4,
  101997.7, 101859.5, 101775.2, 101561.5, 96689.98, 98054.6, 99560.22, 
    101005.2, 101171.1, 101267.3, 101344.3, 101427.3, 101505.3, 101561.8, 
    101607.8,
  102061, 101945.3, 101876.3, 101677.3, 97331.96, 97491.1, 96911.31, 
    101298.1, 101386.7, 101362.4, 101428.7, 101493.7, 101566.5, 101612.6, 
    101658.3,
  100542.2, 100576.8, 100682.5, 100778.5, 100866.7, 100923.8, 100954, 
    100960.2, 100960, 100968.3, 101002.2, 101035.6, 101077.2, 101118.5, 
    101134.1,
  100381.8, 100417.8, 100592.5, 100690.6, 100782.3, 100866.4, 100923.4, 
    100956.4, 100971, 100982, 101010, 101056.9, 101108.2, 101145.8, 101163.9,
  98660.48, 98485.44, 100433.6, 100629.5, 100712.8, 100805.3, 100872.2, 
    100923.5, 100957.2, 100989.9, 101028.4, 101094.4, 101138.3, 101172.6, 
    101191.1,
  96741.8, 96888.74, 100272.9, 100559.2, 100642.3, 100749, 100832.9, 
    100902.6, 100948.3, 100996.8, 101045.8, 101110.9, 101154.6, 101186.4, 
    101232.3,
  96782.53, 97223.27, 99024.12, 100514.5, 100600.8, 100684, 100789.9, 
    100864.4, 100922.1, 100993.7, 101055.6, 101135.1, 101175.8, 101232.4, 
    101267,
  96283.95, 97638.39, 100275.7, 100453.3, 100554.9, 100615.2, 100779.2, 
    100867.6, 100933.6, 100997.1, 101057.7, 101098, 101209.4, 101270.7, 101308,
  100469.8, 100369.4, 100398.5, 100441.2, 100515.5, 98937.05, 100460.7, 
    100640.2, 100841.2, 100957, 101078.1, 101160.9, 101244.7, 101303.3, 
    101345.6,
  100505.1, 100388.2, 100382.3, 100374.1, 100324.6, 98081.45, 96447.69, 
    95737.32, 98249.65, 100942.4, 101084.6, 101184.4, 101275.8, 101338.3, 
    101385.6,
  100491, 100405.7, 100432.4, 100327.3, 95895.6, 97351.34, 98993.14, 
    100486.3, 100787.9, 100959.7, 101077.2, 101192.4, 101290.4, 101360.6, 
    101415.7,
  100581.9, 100492.4, 100501.6, 100344.8, 96349.17, 96723.93, 96328, 
    100686.2, 100903.3, 100951.5, 101074.9, 101200.3, 101310.7, 101390.5, 
    101450.4,
  101200.5, 101208.8, 101224.4, 101211.5, 101209.1, 101194.6, 101188.8, 
    101131.7, 101066.6, 101002.6, 100955.8, 100951.6, 100989.7, 101019.2, 
    101028.6,
  101114.9, 101092.8, 101193.7, 101196.9, 101191.2, 101176.3, 101184, 
    101157.7, 101107.7, 101052.8, 100977.3, 100967.1, 101006.2, 101046.6, 
    101077.3,
  99321.45, 99090.16, 101029.6, 101168.2, 101156.8, 101152.9, 101170.2, 
    101164.8, 101100.8, 101078.6, 101002.8, 100980.9, 101037.8, 101073.5, 
    101104.4,
  97340.15, 97396.45, 100829.5, 101110.2, 101118.7, 101134.3, 101148.9, 
    101174.2, 101119, 101088.3, 101026.4, 100991.9, 101054.2, 101076.3, 
    101141.4,
  97237.18, 97711.77, 99527.25, 101031.2, 101074.8, 101076.7, 101107.1, 
    101139.9, 101120.7, 101073.8, 101039, 101010.1, 101071.7, 101116.8, 
    101173.5,
  96509.27, 98022.05, 100762.1, 100960.9, 101001.9, 100998.9, 101101.7, 
    101132.6, 101142, 101078.7, 101040.2, 100974.9, 101101, 101148.5, 101205.4,
  100687.3, 100791.7, 100884.3, 100937.5, 100970.5, 99254.25, 100713.2, 
    100867.3, 101044.6, 101045.5, 101051.2, 101039.4, 101113.4, 101173, 
    101235.9,
  100749, 100757.6, 100828.5, 100838.9, 100769.6, 98435.34, 96642.65, 
    95828.22, 98341.02, 101033.5, 101046.7, 101060, 101130, 101201.1, 101267.6,
  100624.9, 100678.2, 100796.4, 100816.2, 96196.04, 97566.59, 99169.4, 
    100688.2, 100956.4, 101036.5, 101042.4, 101069.6, 101147.2, 101221.7, 
    101291.1,
  100547.5, 100634.6, 100749.6, 100744.7, 96612.55, 96871.69, 96410.68, 
    100747, 101020.1, 100986.2, 101046.8, 101071.5, 101170.6, 101238.8, 101319,
  101299.2, 101281.7, 101283.9, 101250.8, 101223.6, 101180.8, 101121.9, 
    101022.9, 100912.8, 100822.6, 100819.1, 100863.9, 100915.1, 100952.1, 
    100987.2,
  101246.1, 101189.3, 101287.5, 101255.6, 101216.1, 101188.4, 101135.6, 
    101057.8, 100939.9, 100822.8, 100801.2, 100841.9, 100898.7, 100961.8, 
    101014.1,
  99492.45, 99213.27, 101169.4, 101261.7, 101215.3, 101182.2, 101121, 
    101052.6, 100923, 100800.1, 100776.2, 100827, 100900.2, 100973.5, 101027.9,
  97517.35, 97621.18, 101048, 101266.2, 101213.6, 101192.5, 101134.7, 
    101085.8, 100933.5, 100788.6, 100766.4, 100814.7, 100898.6, 100960.6, 
    101043.6,
  97520.05, 97966.11, 99768.58, 101245.4, 101212.5, 101156.8, 101137.8, 
    101068.9, 100926.6, 100784.9, 100763.9, 100809.1, 100895.8, 100984.8, 
    101066.8,
  96872.27, 98344.73, 101095.6, 101216.2, 101196.1, 101075.6, 101160.7, 
    101099.2, 100995.3, 100834.2, 100756.4, 100761.7, 100911.2, 101000.7, 
    101088.3,
  101078.7, 101171.5, 101226.5, 101237.9, 101194.1, 99355.76, 100815.5, 
    100830.5, 100928, 100842.2, 100809.2, 100826.7, 100926.2, 101014.1, 
    101110.7,
  101141.7, 101169.2, 101224.5, 101198.4, 101009.3, 98608.91, 96766.97, 
    95887.46, 98389.71, 100914.6, 100867.8, 100858.4, 100949.6, 101032.8, 
    101133.6,
  101106.5, 101153.2, 101232.2, 101188.2, 96424.09, 97859.78, 99460.59, 
    100996.1, 101135.7, 100981.6, 100924.3, 100896.8, 100979.5, 101055.3, 
    101159.7,
  101100.7, 101162.7, 101231.6, 101172.1, 96988.57, 97226.43, 96620.85, 
    101065.8, 101199.4, 101032.9, 100979.1, 100938.5, 101016.5, 101082.2, 
    101186.9,
  101322, 101340.1, 101330.2, 101331.1, 101322.3, 101310.3, 101279.8, 
    101228.2, 101142, 101094.5, 101053.3, 101045.5, 101046.2, 101077.6, 
    101097.5,
  101274.9, 101250.8, 101332.7, 101325.8, 101305.4, 101309.2, 101292.4, 
    101280.2, 101216.5, 101132.7, 101085.9, 101079.1, 101085.8, 101110.2, 
    101138.2,
  99543.88, 99278.53, 101205, 101301, 101294.6, 101289, 101279.3, 101268.3, 
    101225.6, 101160.6, 101118.1, 101098.8, 101106.6, 101129.4, 101152.4,
  97594.49, 97686.08, 101054.3, 101283.7, 101281.1, 101276.9, 101268.4, 
    101275.5, 101251.1, 101189.4, 101147.9, 101123.4, 101123.9, 101128, 
    101172.1,
  97578.66, 98014.73, 99769.45, 101257.3, 101253.3, 101230.8, 101234.8, 
    101233.9, 101225.8, 101187.5, 101155.4, 101143.6, 101132.6, 101159.3, 
    101190.3,
  96914.27, 98357.69, 101074.5, 101217.6, 101233.8, 101144.3, 101210.8, 
    101212.8, 101220.7, 101184.9, 101134.4, 101094.1, 101146, 101177.3, 
    101203.7,
  101045.9, 101141.4, 101209.2, 101229.5, 101234.6, 99432.59, 100826.9, 
    100914.8, 101101.1, 101130.4, 101122.8, 101127.2, 101151.6, 101183.6, 
    101216,
  101121.1, 101151, 101199.4, 101208.4, 101045, 98659.52, 96796.23, 95957.75, 
    98461.46, 101106.6, 101105.7, 101111.5, 101148.5, 101188.5, 101229.1,
  101081.5, 101122.9, 101199.5, 101210, 96448.63, 97879.41, 99456.55, 
    100992.2, 101142, 101104.9, 101050.9, 101074.7, 101136.6, 101185.5, 
    101238.5,
  101068.8, 101122.3, 101192.1, 101174.2, 96994.81, 97248.71, 96619.44, 
    101020, 101157.7, 101049.2, 100998.9, 101028.7, 101112.7, 101183.5, 
    101244.4,
  101245.7, 101204.3, 101194.6, 101153.9, 101125, 101090, 101022.6, 100966.6, 
    100904.9, 100887.8, 100900.5, 100934.6, 100978.6, 101025.4, 101058.2,
  101234.3, 101139.1, 101209, 101167.5, 101135.5, 101095.8, 101041.2, 
    100992.6, 100915.9, 100855.5, 100902.6, 100929.6, 100987.7, 101050.9, 
    101088.2,
  99478.68, 99217.57, 101138.1, 101188.2, 101152.6, 101104.3, 101060.3, 
    100988.6, 100921.2, 100847.8, 100893.5, 100932.1, 101007.4, 101070.9, 
    101109.8,
  97603.41, 97725.8, 101043.8, 101206.3, 101170.3, 101127.1, 101080.3, 
    101024, 100935, 100864.6, 100891.8, 100941.2, 101022.1, 101068.4, 101132.1,
  97634.16, 98067.54, 99819.35, 101226.5, 101191.5, 101128.6, 101089.8, 
    101041.1, 100928.5, 100881.4, 100911.2, 100955.4, 101029.9, 101098.7, 
    101162,
  97100.2, 98528.48, 101163.1, 101226.7, 101201.4, 101082.7, 101139, 
    101078.4, 100972.7, 100903, 100914.1, 100925.6, 101052.5, 101125.1, 
    101189.6,
  101323.6, 101331.4, 101300.8, 101286.2, 101224.6, 99411.68, 100837.7, 
    100852.6, 100916.7, 100896, 100948.8, 100997.3, 101080.3, 101153.6, 
    101218.5,
  101377.9, 101366, 101346.2, 101289.5, 101049.9, 98678.55, 96806.82, 
    95991.23, 98407.73, 100963.2, 100992.8, 101045.5, 101117.9, 101190.4, 
    101257.1,
  101409.6, 101372.7, 101391.5, 101282.2, 96555.05, 98012.76, 99554.26, 
    101041.9, 101098.3, 101045.7, 101050.6, 101095, 101161, 101229.6, 101290.9,
  101457.2, 101421.1, 101440.5, 101334.8, 97132.36, 97337.16, 96745.1, 
    101159.2, 101211.2, 101110.6, 101108.9, 101146.7, 101210.9, 101267.3, 
    101322,
  100818, 100795.2, 100789.1, 100752.5, 100732, 100660.3, 100573.9, 100571, 
    100655.4, 100754.3, 100811.1, 100871.2, 100930, 100982.7, 101022.6,
  100760.6, 100718.1, 100788.3, 100748.6, 100727.8, 100689, 100612.8, 
    100593.9, 100662.6, 100741.9, 100811.9, 100877.7, 100941.3, 101010.3, 
    101052.3,
  99055.19, 98811.87, 100702.7, 100764, 100724.9, 100686.8, 100610.5, 
    100585.5, 100658.9, 100741.4, 100817.9, 100889.4, 100982.6, 101041.1, 
    101083.6,
  97173.45, 97286.37, 100594.6, 100763, 100734, 100695.8, 100631.6, 100601.6, 
    100666.9, 100747.1, 100834.9, 100919.4, 101000.7, 101050.2, 101117.6,
  97215.33, 97626.06, 99355.16, 100764.5, 100737, 100659.3, 100637, 100619.3, 
    100668.2, 100757.3, 100849.2, 100935.9, 101018, 101097.5, 101161.1,
  96682.96, 98062.86, 100684.7, 100758, 100736.7, 100604.9, 100640.2, 
    100637.7, 100692.9, 100783, 100850.2, 100906.3, 101046.9, 101129.9, 
    101193.5,
  100890, 100859.5, 100819.3, 100783.8, 100715.5, 98932.95, 100374.8, 
    100465.9, 100637.4, 100757.7, 100886.5, 100987.5, 101088.8, 101163.9, 
    101225.9,
  100972.6, 100897.1, 100857.9, 100784, 100583.2, 98173.88, 96374.22, 
    95630.83, 98120.72, 100796.5, 100917.1, 101028.2, 101125.5, 101201.2, 
    101261.9,
  101022.7, 100959.1, 100936.5, 100799, 96101.62, 97519.8, 99062.52, 
    100540.9, 100717.5, 100844.7, 100947.7, 101068.2, 101167.9, 101243.9, 
    101303.6,
  101095.5, 101051.5, 101028.3, 100888.4, 96687.71, 96890.9, 96352.05, 
    100733.7, 100853.4, 100871.1, 100983.2, 101105.2, 101209.5, 101286.9, 
    101345.9,
  100510.7, 100594.2, 100712.4, 100796.5, 100881.2, 100942.9, 100975.2, 
    100973.7, 100972.9, 100997.5, 100989.7, 100947.2, 100885.5, 100922.7, 
    100919.1,
  100355.9, 100450, 100627.5, 100731.9, 100822.8, 100897.4, 100943.5, 
    100956.7, 100961.7, 100981.9, 100999.4, 100987.6, 100882.1, 100926.3, 
    100939.9,
  98610.3, 98498.41, 100463.9, 100683.9, 100771.1, 100853.1, 100906.3, 
    100929.9, 100941.5, 100954.7, 100983.4, 100984.4, 100907.9, 100923.4, 
    100955.8,
  96597.12, 96812.56, 100292.6, 100618, 100720.2, 100808.5, 100865.2, 
    100898.8, 100919.9, 100938, 100988.6, 100981.7, 100917.3, 100908.9, 
    100983.7,
  96543.88, 97069.2, 98982.28, 100549.3, 100662.9, 100732.8, 100813, 
    100849.8, 100874.8, 100904.4, 100975.2, 100969, 100923.5, 100967.4, 
    101004.6,
  95892.72, 97384.59, 100192, 100470.9, 100590.7, 100635.1, 100763.1, 
    100816.3, 100850.3, 100878.7, 100948.7, 100929.9, 100943.2, 100988.2, 
    101032.4,
  100007.9, 100143.7, 100329.2, 100439.7, 100523.3, 98878.7, 100380.4, 
    100547, 100721.5, 100806.2, 100929.1, 100961.5, 100954.5, 101022.2, 
    101057.4,
  100114.4, 100139.1, 100267.3, 100331.1, 100314, 98011.52, 96297.91, 
    95550.59, 98032.3, 100758.3, 100893.9, 100943.1, 100964.4, 101042.2, 
    101083.7,
  100040.7, 100097.2, 100251, 100276.3, 95753.09, 97157.88, 98762, 100287.2, 
    100573.7, 100759.9, 100853.1, 100935, 100983, 101068.7, 101123.4,
  100073, 100119.1, 100221.8, 100207.9, 96137.66, 96445.48, 96033.8, 100378, 
    100647.5, 100726.4, 100830.9, 100935.7, 101009.9, 101098.6, 101160.6,
  100558.5, 100648.2, 100763.4, 100865.9, 100944.4, 101009.2, 101048.5, 
    101091.9, 101137.4, 101171.1, 101205.4, 101214.8, 101203, 101201.9, 
    101182.3,
  100443.3, 100524.4, 100687.8, 100802.5, 100889.2, 100971.6, 101030, 
    101082.4, 101118.9, 101153.4, 101178.4, 101205.9, 101195.4, 101204.1, 
    101204.4,
  98673.05, 98559.34, 100523.8, 100752, 100839.8, 100929.7, 100987.2, 
    101043.1, 101085.7, 101125, 101152.6, 101177.3, 101180.6, 101196.6, 
    101193.6,
  96648.64, 96861.52, 100350.2, 100701.9, 100794.5, 100905.8, 100975.5, 
    101039.4, 101078, 101112.3, 101125.4, 101152.2, 101162.4, 101161.6, 
    101183.7,
  96561.28, 97119.77, 99051.88, 100634.6, 100749.7, 100827.2, 100918.8, 
    100978.1, 101018.6, 101069.7, 101086.6, 101120, 101128.5, 101149.4, 
    101174.2,
  95831.9, 97405.63, 100246.1, 100561, 100682.8, 100757.5, 100906, 100974.9, 
    101010.2, 101044.4, 101041.8, 101037.6, 101109.8, 101129, 101164.8,
  99906.89, 100142.1, 100367.2, 100531.4, 100634.5, 99003.71, 100519.4, 
    100696.4, 100878.2, 100971.2, 101023.2, 101053.5, 101089.7, 101102.1, 
    101149.8,
  100020.6, 100141.8, 100306.2, 100430.5, 100433.8, 98154.44, 96455.94, 
    95716.56, 98205.32, 100907.9, 100996.4, 101022.4, 101053.5, 101080.3, 
    101135.9,
  99930.49, 100067.7, 100281.1, 100382, 95868.3, 97310.45, 98957.48, 
    100492.1, 100775.2, 100887.1, 100965.6, 100985, 101012.2, 101057.5, 
    101117.9,
  99940.98, 100081.4, 100264, 100322.7, 96286.9, 96618.64, 96226.07, 
    100616.9, 100878.1, 100844.3, 100935, 100942.1, 100975.3, 101041.9, 
    101100.6,
  100597.1, 100685.4, 100794, 100888.5, 100961, 101038.8, 101069.6, 101117.6, 
    101188.1, 101229.6, 101252.8, 101249.4, 101217.1, 101189.7, 101171.8,
  100561.1, 100642.6, 100799.2, 100885.9, 100970.2, 101043.4, 101101.5, 
    101147.3, 101196.4, 101244.5, 101271.7, 101280.7, 101267.2, 101235.6, 
    101216.8,
  98916.11, 98776.38, 100712.3, 100901.9, 100975.9, 101052.2, 101105.2, 
    101147.9, 101188.2, 101242, 101287, 101299, 101289.1, 101261.6, 101236.3,
  97008.57, 97203.54, 100622.9, 100913.2, 100982.7, 101070.1, 101134.7, 
    101183, 101209.4, 101242.3, 101294.8, 101322.1, 101309.9, 101280.5, 
    101268.7,
  97025.74, 97517.57, 99395.54, 100906.6, 100988, 101046, 101124.4, 101174.6, 
    101213.4, 101247.6, 101285.7, 101335, 101325.1, 101310.6, 101296.5,
  96390.6, 97890.24, 100652.5, 100886.3, 100975.9, 101018.4, 101156.9, 
    101205.6, 101228.2, 101260, 101281.2, 101287.4, 101352, 101343.9, 101330.6,
  100514.6, 100636.4, 100788.8, 100907.9, 100982.2, 99319.8, 100825.8, 
    101002.4, 101178, 101246.2, 101298.1, 101327.2, 101372.4, 101367, 101356.5,
  100600.1, 100665.2, 100759.9, 100847.4, 100817.7, 98523.24, 96797.38, 
    96024.81, 98518.16, 101235.2, 101311.2, 101332.7, 101367.7, 101394.5, 
    101374.3,
  100483.7, 100589, 100738.1, 100826.2, 96291.06, 97709.52, 99361.13, 
    100913.4, 101152.8, 101248.8, 101301.5, 101332, 101365.6, 101400.3, 
    101395.4,
  100451, 100561.1, 100717.9, 100761.5, 96734.19, 97039.25, 96600.31, 
    100993.5, 101244.7, 101218.3, 101287.4, 101322.2, 101364.6, 101394.7, 
    101410.8,
  100191.6, 100207.7, 100275.4, 100309.5, 100315.2, 100319.9, 100261.1, 
    100203.5, 100180.8, 100211.1, 100258.4, 100277, 100330.8, 100398.8, 100491,
  100110.2, 100138.6, 100281, 100325.3, 100335.5, 100375.7, 100349.4, 
    100293.5, 100248.4, 100256.7, 100304.9, 100326.7, 100346.4, 100411, 
    100518.1,
  98402.47, 98248.28, 100175.1, 100337.3, 100354.9, 100394, 100391.6, 100367, 
    100297.8, 100277.9, 100329, 100361.9, 100397.5, 100440.1, 100526.5,
  96432.99, 96636.69, 100054.7, 100335.7, 100378.9, 100420.8, 100461, 
    100449.2, 100369.4, 100339.5, 100383.8, 100413.2, 100443.9, 100474.3, 
    100549.3,
  96384.73, 96908.88, 98806.93, 100324.8, 100400.9, 100424.1, 100493.4, 
    100489.1, 100462.6, 100411.5, 100442.3, 100467.2, 100490.8, 100551.3, 
    100596.6,
  95738.06, 97237.66, 100032.1, 100297.7, 100408.4, 100408.2, 100529.9, 
    100560.4, 100539.7, 100498.5, 100473.2, 100486.4, 100545.1, 100609.7, 
    100672.4,
  99786.73, 99949.96, 100168.7, 100313.6, 100409, 98767.04, 100284.8, 
    100397.5, 100523.6, 100551.4, 100539.5, 100582.1, 100602.6, 100642, 100714,
  99928.81, 99978.65, 100148.5, 100270.4, 100266.5, 97974.45, 96248.4, 
    95462.55, 97967.96, 100622.5, 100614.2, 100620.3, 100658.3, 100670.6, 
    100732.7,
  99882.23, 99971.7, 100158.8, 100252.1, 95793.79, 97253.79, 98899.62, 
    100442.7, 100656.9, 100694.5, 100694.6, 100667.8, 100716.9, 100723.7, 
    100764.1,
  99936.62, 100030.9, 100169, 100222.4, 96269.8, 96614.79, 96147.56, 
    100551.5, 100745, 100751.6, 100764, 100737.4, 100763, 100777, 100806.6,
  100325.7, 100310.2, 100337.7, 100334.3, 100335.2, 100341.3, 100340.6, 
    100335.7, 100333.2, 100328.1, 100316, 100319.3, 100343.5, 100363.9, 
    100343.2,
  100201, 100177.5, 100271.7, 100280.5, 100270.5, 100269.5, 100259.9, 
    100265.9, 100262.9, 100258.1, 100258.8, 100265.3, 100298.5, 100331.8, 
    100349,
  98424.05, 98195.32, 100087.3, 100215.1, 100193, 100199.6, 100172.9, 
    100184.2, 100179.7, 100167.3, 100182.5, 100199.1, 100236.2, 100282.9, 
    100315.7,
  96440.38, 96528.73, 99909.97, 100150.9, 100135.4, 100147.4, 100115.5, 
    100129.6, 100094.1, 100062.6, 100082.8, 100126.5, 100175, 100229.1, 
    100293.2,
  96368.21, 96825.09, 98602.55, 100068.8, 100068.8, 100039.6, 100033.2, 
    100046.3, 100013.8, 99972.86, 99981.61, 100049.7, 100099, 100187.2, 
    100259.2,
  95669.77, 97130.89, 99833.96, 99995.68, 99987.7, 99918.12, 99980.23, 
    100002.8, 99970.8, 99901.38, 99865.59, 99915.35, 100036.3, 100138.4, 
    100225.6,
  99836.62, 99892.37, 99950.2, 99958.48, 99952.14, 98158.12, 99573.84, 
    99707.36, 99810.42, 99840.13, 99792.09, 99861.62, 99970.63, 100078.2, 
    100187.3,
  99875.94, 99853.73, 99893.57, 99859.52, 99717.77, 97330.96, 95547.77, 
    94737.32, 97155.6, 99779.24, 99751.88, 99767.57, 99906.84, 100022.8, 
    100155.6,
  99785.13, 99776.19, 99858.49, 99810.92, 95143.02, 96484.65, 98079.45, 
    99571.07, 99777.23, 99739.59, 99688.75, 99679.93, 99841.48, 99967.9, 
    100123.1,
  99783.7, 99763.7, 99825.59, 99745.62, 95601.74, 95792.35, 95295.61, 
    99604.96, 99801.89, 99667.84, 99626.5, 99599.06, 99777.91, 99915.71, 
    100089.1,
  100362.6, 100463.5, 100557.6, 100627.7, 100674.2, 100709.2, 100727, 
    100734.3, 100728.6, 100718.1, 100689.3, 100640.3, 100596, 100552.8, 
    100513.4,
  100327.4, 100417.1, 100551.1, 100630.8, 100690.2, 100733, 100756.9, 100773, 
    100770.8, 100755.1, 100741.1, 100701.6, 100671, 100628.8, 100602.8,
  98643.98, 98521.72, 100460.4, 100633.5, 100680.4, 100733.5, 100756.2, 
    100778, 100781.5, 100778, 100763.8, 100735.8, 100711.8, 100666.3, 100646.7,
  96716.45, 96916.2, 100341.1, 100632.3, 100681.3, 100749.6, 100779.8, 
    100808.9, 100810.3, 100810.2, 100800.3, 100778.9, 100762.8, 100718.9, 
    100710.4,
  96705.58, 97223.14, 99088.98, 100600.5, 100672.2, 100710.2, 100761.4, 
    100793, 100810.9, 100820.6, 100820.5, 100805.6, 100783, 100779.8, 100763.9,
  96037.65, 97561.65, 100313.8, 100561.8, 100638.7, 100664.1, 100785.7, 
    100823.5, 100837.4, 100839.7, 100834, 100786, 100826.3, 100819.2, 100808.3,
  100123, 100284.1, 100440.6, 100550.7, 100618.4, 98929.34, 100405, 100562.7, 
    100747.6, 100811.9, 100852.4, 100845.8, 100852.6, 100856, 100844.5,
  100227.1, 100275.6, 100402, 100456, 100430.7, 98130.42, 96377.77, 95561.47, 
    98052.33, 100770.1, 100841.5, 100852.5, 100864.1, 100876.2, 100870.3,
  100123.5, 100192.8, 100353.7, 100425.6, 95880.59, 97250.12, 98917.93, 
    100466.9, 100706.6, 100764.5, 100819.3, 100841.7, 100870.3, 100880.2, 
    100886.1,
  100093.9, 100155.9, 100291.9, 100328, 96293.23, 96578.19, 96151.07, 
    100499.1, 100761.5, 100722.3, 100812.9, 100827.3, 100870.1, 100878.8, 
    100890.4,
  100127.5, 100154.6, 100235.6, 100308.4, 100359.8, 100397.4, 100416.6, 
    100433.5, 100443.8, 100431.9, 100420.7, 100413.6, 100422.4, 100460.6, 
    100516.1,
  100001, 100073.5, 100219, 100292.2, 100348.5, 100398.4, 100432.3, 100441.1, 
    100453.6, 100440, 100413.4, 100376.3, 100393.5, 100456.1, 100530.9,
  98302.81, 98181.73, 100096.4, 100291.1, 100351.3, 100406.2, 100434, 
    100438.7, 100446.1, 100436.1, 100420.4, 100375.5, 100367.3, 100424.3, 
    100510.2,
  96328.61, 96576.56, 99986.73, 100272.5, 100347.9, 100415, 100453.5, 
    100461.9, 100458.3, 100440, 100412.2, 100347.4, 100338.2, 100390.6, 
    100491.4,
  96283.66, 96852.66, 98748.33, 100257.7, 100349.1, 100405, 100462.7, 
    100461.1, 100450.9, 100430.4, 100401.5, 100336.5, 100319.2, 100400.8, 
    100482.5,
  95677.02, 97197.55, 99984.98, 100229.6, 100339.4, 100360.4, 100488.1, 
    100509.1, 100492, 100446.1, 100388.5, 100295.1, 100326.3, 100418.3, 
    100499.6,
  99741.1, 99927.89, 100144.3, 100254.5, 100317.2, 98711.45, 100201.9, 
    100298.8, 100415.7, 100428.6, 100407.3, 100353.9, 100362.5, 100446.2, 
    100528.1,
  99905.83, 99993, 100147.1, 100215.5, 100158.5, 97869.13, 96163.92, 
    95410.73, 97869.07, 100448.5, 100427, 100384.9, 100409.7, 100485.8, 
    100563.8,
  99856.78, 99980.61, 100169.6, 100181.6, 95723.52, 97190.23, 98834.06, 
    100363.9, 100513.4, 100488.1, 100454.5, 100421, 100461.5, 100532.5, 
    100603.8,
  99907.37, 100027.8, 100190, 100174.5, 96195.95, 96521.45, 96100.37, 
    100489.2, 100609.1, 100526.4, 100486.8, 100470.4, 100522.5, 100592.5, 
    100655.5,
  101045.1, 101048, 101129.2, 101170.1, 101196.4, 101201.6, 101180.3, 101154, 
    101136, 101103.6, 101052.3, 101011.7, 100963.5, 100912.1, 100901.4,
  100840.3, 100870.7, 101025, 101084.3, 101117.5, 101140.6, 101133.2, 
    101120.6, 101112.8, 101099.5, 101053.8, 101003.2, 100967.6, 100925.7, 
    100929.5,
  98980.36, 98826.74, 100762.1, 100983, 101011.4, 101054.1, 101062, 101056.9, 
    101058.4, 101056.4, 101037.6, 100998, 100966.6, 100922.6, 100920.9,
  96855.48, 97047.25, 100500.6, 100861.9, 100918.7, 100985.3, 101013, 
    101011.2, 101016.9, 101014.1, 101012, 100974.6, 100955.2, 100909.7, 100922,
  96716.21, 97254.05, 99120.5, 100708.4, 100807.4, 100852.8, 100913.8, 
    100933.6, 100940.1, 100949.3, 100970.7, 100945.1, 100935.7, 100926, 
    100919.8,
  95899.52, 97448.46, 100263.3, 100564, 100671.9, 100735.1, 100846.1, 100881, 
    100893.9, 100900.8, 100913.4, 100873.7, 100921.5, 100916.9, 100912.9,
  99954.45, 100163, 100324.4, 100469.4, 100563.4, 98919.94, 100402.4, 
    100578.9, 100732.1, 100809.9, 100871.2, 100888.1, 100904.4, 100895.9, 
    100903.2,
  99970.66, 100060.9, 100209.5, 100306.9, 100317.2, 98041.43, 96307.95, 
    95544.18, 97988.45, 100711.7, 100820.7, 100851.2, 100879.6, 100867.3, 
    100892.2,
  99816.98, 99918.44, 100120.7, 100209.2, 95684.55, 97102.25, 98746.65, 
    100267.9, 100537.3, 100664.4, 100748.8, 100804.8, 100847.6, 100841.4, 
    100875.8,
  99741.27, 99854.21, 100022, 100082.5, 96060.8, 96384.7, 95995.1, 100340.2, 
    100607.3, 100565.7, 100673.7, 100743.4, 100812.1, 100817, 100854.9,
  101534.2, 101523.8, 101561.1, 101583.7, 101589.4, 101595.1, 101595.6, 
    101577, 101548.5, 101510.5, 101462.9, 101414.6, 101396, 101348.6, 101277.7,
  101403.2, 101399.8, 101504, 101536.4, 101545.6, 101565.1, 101568.2, 
    101571.7, 101554.8, 101521.8, 101480.7, 101426.6, 101396.4, 101372.4, 
    101331.3,
  99587.85, 99381.59, 101320.9, 101480.8, 101478.7, 101504.9, 101507.2, 
    101512.6, 101512.6, 101498.4, 101467.7, 101435.8, 101389.1, 101363.5, 
    101316.5,
  97571.25, 97671.77, 101107.4, 101395.9, 101403, 101450.5, 101468.1, 
    101483.6, 101482.8, 101476.1, 101458.2, 101430.6, 101398.5, 101356.5, 
    101329.8,
  97481.37, 97975.02, 99787.8, 101287.5, 101323.8, 101340.2, 101380.1, 
    101404.5, 101416.6, 101427.1, 101426.9, 101417.5, 101381.7, 101362.9, 
    101324.8,
  96726.87, 98242.03, 100985.2, 101190, 101225.8, 101241.9, 101348.6, 
    101373.5, 101386.4, 101396.3, 101385.1, 101348.2, 101381.3, 101369.7, 
    101332.2,
  100973.9, 101024, 101092.2, 101131.1, 101156, 99423.89, 100890.1, 101066.5, 
    101230.9, 101315.1, 101358.6, 101366.1, 101363.3, 101360.2, 101331.6,
  101001.2, 100988.4, 101039.7, 101000.8, 100924.7, 98596.49, 96821.72, 
    96003.35, 98473.15, 101216.6, 101306.4, 101322.3, 101333.6, 101337.4, 
    101327.7,
  100837.9, 100865.9, 100973.2, 100984.6, 96297.6, 97626.2, 99309.32, 
    100865.2, 101107.5, 101181.4, 101238.4, 101264.8, 101293.9, 101307.1, 
    101306.8,
  100734.2, 100766.3, 100864.8, 100852.2, 96698.31, 96946.12, 96510.9, 
    100895.6, 101176.1, 101104.1, 101184.6, 101207.8, 101256.6, 101273, 
    101284.7,
  101476.1, 101447.9, 101471.9, 101476.3, 101485.1, 101469.1, 101418, 
    101402.8, 101364.8, 101287.7, 101231.4, 101208.9, 101203.5, 101189.6, 
    101147.6,
  101429.4, 101375.6, 101464.2, 101449.7, 101447.3, 101448.2, 101437.1, 
    101403.7, 101399.9, 101356.4, 101288.7, 101251, 101230.8, 101217.9, 
    101203.6,
  99688.35, 99417.59, 101346.7, 101437.8, 101448.6, 101444.3, 101423.8, 
    101392.8, 101370.8, 101368.1, 101318.6, 101271.8, 101257.9, 101229.1, 
    101218.5,
  97730.53, 97830.37, 101219.9, 101460.7, 101444.8, 101445.2, 101422, 
    101406.4, 101372.1, 101347, 101342.3, 101299.8, 101280, 101241.4, 101245.2,
  97798.31, 98242.33, 100003.5, 101479.7, 101451.2, 101409, 101390.6, 101380, 
    101358.3, 101337, 101322.8, 101308, 101274.8, 101270.6, 101253.3,
  97196.1, 98643.98, 101371.6, 101470.4, 101437.4, 101351.5, 101401.2, 
    101379.2, 101368.8, 101348.1, 101307.5, 101253.3, 101285.7, 101284.4, 
    101269.8,
  101565.5, 101571.5, 101550.6, 101515.5, 101469.4, 99610.31, 101020.6, 
    101128.3, 101288.4, 101318.8, 101323.3, 101300.8, 101296, 101291.5, 
    101274.1,
  101604.8, 101551.2, 101546.8, 101479.3, 101286.8, 98875.22, 97001.9, 
    96103.09, 98562.87, 101292.1, 101320.3, 101298.2, 101290.1, 101286.9, 
    101278,
  101586.3, 101548.9, 101550.1, 101498.2, 96661.06, 98002.24, 99628.12, 
    101149.2, 101302.1, 101313.4, 101310.9, 101284.5, 101281.8, 101276.6, 
    101271.9,
  101567.5, 101543.6, 101533.9, 101446, 97179.77, 97360.64, 96795.09, 
    101155.9, 101356.4, 101274.4, 101307.4, 101282.9, 101281.5, 101266.7, 
    101263.9,
  101690, 101646.6, 101645.3, 101578.2, 101523.8, 101465.9, 101368.3, 
    101266.6, 101170.6, 101048.9, 100988.4, 100992.3, 100990.9, 101010.1, 
    100998.4,
  101667.6, 101597.4, 101687.9, 101623.5, 101594.4, 101527, 101468.3, 
    101398.9, 101304.5, 101216.9, 101108.5, 101062, 101050, 101046.2, 101053.2,
  99946.56, 99678.56, 101660, 101696, 101633.8, 101579.2, 101518.8, 101453.6, 
    101364.1, 101291.7, 101218.4, 101155.5, 101116.7, 101098.8, 101094.8,
  98039.64, 98156.05, 101556.8, 101756.5, 101683.5, 101626.5, 101575.2, 
    101519.8, 101437.6, 101367.8, 101303.8, 101245.6, 101189.2, 101144.5, 
    101150.1,
  98121.47, 98546.09, 100308.7, 101766.9, 101706.2, 101619, 101572.1, 
    101548.7, 101482.9, 101417.7, 101348.7, 101313.3, 101253.1, 101221.4, 
    101204,
  97550.8, 98994.2, 101714.6, 101770.7, 101703.6, 101574.8, 101591, 101561.6, 
    101526.9, 101466.3, 101385.1, 101307.6, 101324.9, 101284.5, 101255.9,
  101911.4, 101922.6, 101850.4, 101799.1, 101707.1, 99824.47, 101273.4, 
    101364.2, 101479.1, 101472.8, 101436.5, 101384.6, 101373.9, 101347.6, 
    101308.9,
  101965.4, 101930.6, 101872.5, 101795.5, 101482.3, 99081.65, 97158.79, 
    96267.71, 98791.06, 101488.7, 101476.7, 101420.9, 101395.6, 101380.6, 
    101356.5,
  101978.8, 101946.5, 101905.7, 101821.1, 96839.84, 98289.26, 99842.72, 
    101396.4, 101544, 101522.3, 101507.2, 101461.3, 101433.8, 101407, 101385,
  101996.4, 101960, 101937.9, 101823.2, 97462.92, 97688.09, 96985.9, 
    101423.4, 101573.6, 101516.1, 101516.1, 101486.3, 101464.9, 101424.9, 
    101411.1,
  101776, 101744.1, 101707.7, 101626.2, 101562.6, 101461.5, 101384, 101271.6, 
    101164.6, 101074.4, 101041, 101038.3, 101021.6, 101052.6, 101087.9,
  101779.5, 101705.6, 101770.7, 101703.8, 101654.4, 101575.2, 101475.8, 
    101388, 101328.6, 101234.3, 101112.5, 101035.8, 101041.4, 101098.9, 
    101114.9,
  100079.5, 99817.49, 101760.2, 101787.8, 101711.5, 101649.7, 101568.6, 
    101472.1, 101383.4, 101357.1, 101325.9, 101254.2, 101165.4, 101139.7, 
    101173.3,
  98159.73, 98308.88, 101675.9, 101847.3, 101779.9, 101730, 101666.9, 
    101592.1, 101505.8, 101413.6, 101392.7, 101380.9, 101285.8, 101224.9, 
    101263.3,
  98236.66, 98660.45, 100467.1, 101880.1, 101821.7, 101758.9, 101726.6, 
    101662.6, 101604.7, 101548.2, 101455.8, 101449.6, 101467.6, 101381, 
    101381.3,
  97675.28, 99140.63, 101834.8, 101873, 101829.6, 101703.8, 101812.7, 
    101767.5, 101701.6, 101625.6, 101573.3, 101476.3, 101473.4, 101502.8, 
    101448.5,
  101941.3, 102009.8, 101963.6, 101921.7, 101844.6, 100031.4, 101487, 
    101582.4, 101697.8, 101697.5, 101658.5, 101640.7, 101597.2, 101552.1, 
    101513.6,
  102039.6, 102040.3, 101989.2, 101937.1, 101669.7, 99310.15, 97441.27, 
    96617.12, 99111.59, 101773.9, 101747.3, 101695.9, 101673.3, 101636.8, 
    101619.5,
  102040.3, 102032.3, 102030.9, 101944.7, 97105.26, 98604.41, 100160.4, 
    101769.4, 101878, 101846.7, 101821.6, 101775.9, 101733.7, 101691.7, 101658,
  102086.6, 102065.6, 102081.6, 101969.1, 97681.36, 97946.76, 97313.12, 
    101788.5, 101935.2, 101886.1, 101863.1, 101819.4, 101789, 101750.3, 
    101724.7,
  101024, 101022.1, 101013.3, 100992.6, 100973.6, 100949.2, 100929.4, 
    100906.8, 100909.1, 100931.5, 100963.2, 101002.5, 101033.6, 101082.6, 
    101093.3,
  101050.5, 101031.9, 101108.2, 101099, 101086.4, 101058.8, 101037, 101007, 
    100974.6, 100966.9, 101001.1, 101050.2, 101093.6, 101123.1, 101131.2,
  99452.35, 99245.03, 101159.1, 101212.5, 101194.1, 101167.8, 101145.5, 
    101130.9, 101122, 101108.7, 101100.9, 101122.7, 101145.1, 101180.3, 
    101195.7,
  97615.22, 97794.88, 101157.6, 101326, 101315.6, 101293.5, 101265.9, 
    101251.5, 101237.9, 101242.8, 101234.5, 101222, 101236.9, 101237.5, 
    101265.7,
  97701.2, 98164.77, 99996.09, 101432.4, 101417.6, 101390.6, 101377.5, 
    101343.2, 101330.7, 101340.7, 101331, 101325.5, 101316.6, 101335.6, 
    101332.3,
  97185.48, 98633.34, 101352, 101459.5, 101474.1, 101403.6, 101500, 101483.5, 
    101458.9, 101438.5, 101407.9, 101404, 101449.2, 101433.1, 101404.3,
  101364.3, 101456.4, 101510.3, 101529.3, 101499.3, 99797.91, 101256.7, 
    101329.7, 101459.8, 101503.2, 101537.9, 101567.6, 101555.9, 101495.6, 
    101499.5,
  101487.9, 101518.7, 101542.6, 101565.4, 101383.5, 99018.87, 97233.14, 
    96454.37, 98984.34, 101615.4, 101604.3, 101601.3, 101583.2, 101598.9, 
    101567.4,
  101456.6, 101517.5, 101584, 101544.2, 96908.97, 98396.8, 99999.04, 
    101545.2, 101693.9, 101716.7, 101720.9, 101705.9, 101690, 101658.6, 
    101624.5,
  101506.3, 101556.3, 101628.3, 101577.8, 97447.45, 97719.46, 97218.41, 
    101670, 101812.8, 101775.4, 101766, 101751.9, 101737.9, 101715.8, 101687.6,
  100059.1, 100079.6, 100160.5, 100235.3, 100322.9, 100400.6, 100456.8, 
    100498.6, 100561.5, 100608.6, 100661.6, 100710, 100759.7, 100801.2, 
    100816.1,
  99944.46, 99972.23, 100102.3, 100193.7, 100284.8, 100380.9, 100469.4, 
    100531.6, 100583, 100638.1, 100699.7, 100755.4, 100804.9, 100834, 100851.1,
  98239.41, 98065.87, 99971.38, 100162.8, 100258.4, 100365.8, 100467.1, 
    100548.3, 100612.1, 100685.6, 100749.3, 100809.1, 100856.8, 100879.7, 
    100900.6,
  96342.27, 96489.39, 99842.38, 100129.5, 100243, 100365.5, 100477, 100574.8, 
    100648.9, 100726.7, 100788.5, 100852.1, 100896, 100910.4, 100949.4,
  96362.41, 96817.39, 98630.52, 100120.8, 100234.8, 100345.5, 100479.4, 
    100585.8, 100674.4, 100761, 100837.2, 100902.3, 100938.6, 100970.2, 
    100990.8,
  95831.46, 97229.45, 99886.47, 100122.6, 100238.3, 100321.6, 100509.4, 
    100634, 100731.8, 100810.2, 100872.8, 100898.1, 100992, 101022.3, 101036.2,
  100025.1, 100006.9, 100088, 100165.4, 100233.9, 98697.84, 100243.5, 100462, 
    100691.5, 100820.7, 100934.7, 100995.7, 101049.8, 101072.9, 101086.5,
  100125, 100084, 100119.9, 100145.2, 100110.1, 97868.98, 96280.41, 95622.75, 
    98204.45, 100876.7, 100989.9, 101050.7, 101102.1, 101129, 101139.5,
  100077.1, 100072.5, 100159.5, 100121.4, 95714.82, 97200.23, 98890.55, 
    100478.2, 100810, 100950.3, 101041.9, 101101.9, 101153.8, 101181.1, 
    101192.6,
  100147.3, 100138.7, 100206.6, 100154, 96196.89, 96574.6, 96271.07, 
    100727.9, 100976.1, 101003.4, 101097.6, 101158, 101211.2, 101234.5, 
    101245.9,
  100853, 100841.4, 100855.9, 100856.4, 100857.5, 100841.8, 100805.1, 
    100748.9, 100692.6, 100676.7, 100676.3, 100706.1, 100701.1, 100749.1, 
    100765.1,
  100767.2, 100734.9, 100836.6, 100851.8, 100840.7, 100845.4, 100823.2, 
    100799.5, 100751.4, 100711.8, 100705.7, 100729.3, 100748.2, 100786.8, 
    100793.8,
  99052.22, 98795.43, 100687.5, 100815.7, 100819, 100835, 100808.5, 100792, 
    100769, 100725.7, 100742.2, 100757.2, 100799.6, 100808.6, 100830.4,
  97127.12, 97199.56, 100519.1, 100796.5, 100806.3, 100827, 100814.7, 100807, 
    100791.5, 100745.7, 100754.9, 100783.6, 100820.1, 100822.8, 100875.1,
  97070.61, 97514.59, 99265.4, 100765, 100786.9, 100780, 100788.5, 100780.6, 
    100776.9, 100760.8, 100765.1, 100810.9, 100838.2, 100870.7, 100899.7,
  96394.39, 97837.7, 100507.8, 100722.8, 100739.6, 100717.5, 100796.4, 
    100794.2, 100789.8, 100770, 100758.8, 100769.8, 100858.4, 100892.3, 
    100916.8,
  100482.6, 100587.9, 100684.2, 100728, 100736.5, 98969.84, 100396, 100551.1, 
    100696.3, 100740.3, 100775.3, 100824.2, 100875.4, 100910.5, 100936.9,
  100552.9, 100572.9, 100651.1, 100638.7, 100525.5, 98202.39, 96411.19, 
    95607.69, 98053.12, 100719.8, 100776.3, 100833.4, 100890.2, 100932.1, 
    100959.4,
  100432.8, 100470.5, 100603, 100619.9, 96031.23, 97355.48, 98919.4, 
    100404.8, 100642.9, 100726.7, 100774.2, 100835, 100904.1, 100949.1, 
    100980.6,
  100370.6, 100412.8, 100546.8, 100533.5, 96457.12, 96685.29, 96194.11, 
    100433, 100696.7, 100689.4, 100769.1, 100832.7, 100917.4, 100964.3, 
    101010.7,
  101231.5, 101198.9, 101179.7, 101098.9, 101032.4, 100950.3, 100889, 
    100786.3, 100733.7, 100722.6, 100725.3, 100757.4, 100795.3, 100833.3, 
    100836.4,
  101251.8, 101162.2, 101234.1, 101165.4, 101109.5, 101044.8, 100980.6, 
    100950.4, 100835.5, 100818, 100799, 100803.5, 100821.3, 100845.6, 100860.2,
  99564.43, 99284.97, 101195, 101240.5, 101156.5, 101087, 101009.7, 100995.5, 
    100935.9, 100898.6, 100872.8, 100856.9, 100877.8, 100888.8, 100903.6,
  97728.58, 97809.13, 101102.8, 101293.3, 101217.7, 101140, 101071.9, 
    101035.1, 101048.7, 100953.8, 100946.9, 100922.1, 100915.3, 100906.9, 
    100945.7,
  97745.44, 98191.02, 99923.98, 101322.3, 101261.7, 101140.4, 101087.2, 
    101044.2, 101031.6, 101014.7, 100989.1, 100987, 100952.1, 100968.8, 
    100978.8,
  97113.95, 98575.53, 101240.7, 101347.5, 101282.2, 101137.2, 101109.9, 
    101090.4, 101063.5, 101111.8, 100984.4, 100973.4, 100988.8, 100999.4, 
    101013.3,
  101344.1, 101391.5, 101402, 101394.4, 101323.5, 99482.3, 100796.1, 
    100853.6, 100978.1, 101047.6, 101021.2, 101025.9, 101034.3, 101016.7, 
    101042.7,
  101339, 101334.8, 101366.4, 101333, 101122.7, 98775.12, 96899.87, 95989.4, 
    98377.77, 101039.8, 101115.6, 101028.8, 101066, 101042.5, 101060,
  101288.5, 101289.2, 101348.1, 101336.6, 96628.92, 97918.37, 99508.29, 
    100950.6, 101126.1, 101068.4, 101080, 101056.4, 101052.9, 101071.7, 
    101078.8,
  101229.9, 101250.4, 101294.9, 101247.9, 97107.94, 97283.3, 96739.41, 
    100960.6, 101155.2, 101059.7, 101077.4, 101088.9, 101049.8, 101085, 
    101085.2,
  101202, 101157.9, 101119.8, 101018, 100913, 100792.6, 100659.3, 100566.3, 
    100539, 100550.4, 100559.4, 100596.1, 100628.9, 100672.9, 100692.1,
  101248.8, 101125.6, 101176.9, 101093.1, 101019.5, 100907.7, 100811.5, 
    100698.4, 100571.2, 100531.4, 100557, 100597.9, 100636.9, 100675.4, 
    100711.6,
  99578.39, 99291.28, 101170.4, 101183.2, 101090.5, 100987.6, 100888, 
    100801.3, 100702.6, 100604.8, 100537, 100586.8, 100638.4, 100672.8, 
    100713.1,
  97694.46, 97816.35, 101103.3, 101250.5, 101172.4, 101097.4, 100993.5, 
    100899.5, 100812.8, 100694.1, 100598.9, 100592.2, 100644.8, 100652.6, 
    100720.4,
  97749.08, 98169.7, 99917.51, 101299.5, 101226.3, 101136.2, 101066.2, 
    100974.4, 100909.8, 100821.9, 100723.7, 100621.1, 100635.3, 100670.2, 
    100724.4,
  97131.4, 98584.9, 101256.5, 101316.1, 101259.8, 101137.8, 101159.9, 
    101049.1, 100996.3, 100923, 100830.2, 100672.3, 100682.2, 100701.1, 100738,
  101375.3, 101379.7, 101385, 101373.9, 101287.2, 99490.7, 100891.6, 
    100896.3, 100944.4, 100965, 100952.9, 100848.3, 100730.6, 100726.1, 
    100752.8,
  101402.3, 101389.7, 101392.5, 101373.3, 101098.6, 98765.04, 96873.11, 
    96017.14, 98442.16, 101008.9, 101032.5, 100957.9, 100842.2, 100761.9, 
    100763.5,
  101421, 101407.8, 101407.5, 101389.1, 96579.44, 97997.12, 99570.32, 
    101088.3, 101168.6, 101103.9, 101066.4, 101042.2, 100939, 100834.5, 
    100797.3,
  101461.2, 101440.5, 101423.5, 101357.4, 97165.41, 97375.52, 96735.15, 
    101123.7, 101241.8, 101154.3, 101110.9, 101094.8, 101020.9, 100924.3, 
    100847.4,
  101133.6, 101085.9, 101043.4, 100951.5, 100869.1, 100759.6, 100637.7, 
    100551, 100483.6, 100500.1, 100531.8, 100576.5, 100599.2, 100644.5, 100643,
  101128.3, 101052.7, 101092.1, 101012, 100949.8, 100864.6, 100740.9, 100624, 
    100519.7, 100509.2, 100520.7, 100556.5, 100582.9, 100638.6, 100670,
  99438.53, 99177.34, 101065.2, 101075.1, 100993.2, 100908.3, 100821.4, 
    100710.8, 100608, 100527.2, 100523.7, 100553.9, 100594.7, 100639.8, 
    100671.9,
  97569.79, 97692.21, 100987.8, 101134.4, 101057, 100987.1, 100911.2, 100815, 
    100722.6, 100613.8, 100538.3, 100559.7, 100610.9, 100630.7, 100681.4,
  97626.43, 98046.25, 99786.55, 101165.6, 101089.8, 101010.4, 100963, 
    100892.4, 100811.1, 100743.8, 100652, 100625.4, 100605.2, 100658.1, 
    100688.7,
  97085.52, 98509.03, 101136.5, 101172.3, 101104, 100965.9, 101023.8, 
    100971.6, 100911.7, 100823.1, 100726.9, 100652.6, 100671, 100679.7, 
    100706.1,
  101317, 101324.8, 101267.3, 101232.5, 101130.5, 99342.65, 100750.1, 
    100778.5, 100855.1, 100885.5, 100846.5, 100770.1, 100732, 100706.1, 
    100716.8,
  101394.8, 101359.5, 101313.8, 101239.1, 100976.5, 98625.52, 96752.48, 
    95939.33, 98371.81, 100944.3, 100921.7, 100857.9, 100802.3, 100746.1, 
    100725.4,
  101438.4, 101390.2, 101359.8, 101253.1, 96469.77, 97940.31, 99480.78, 
    101006.5, 101080.6, 101038.6, 100988, 100922, 100862.1, 100774, 100733.3,
  101484.1, 101450.6, 101429, 101312.2, 97056.69, 97296.12, 96665.53, 
    101078.2, 101177.1, 101107.9, 101048.5, 100982.2, 100923.7, 100850.8, 
    100754.5,
  101071, 101028.7, 101029.5, 100974.9, 100936.1, 100858.8, 100786.3, 
    100706.7, 100654, 100669.4, 100702.9, 100729.6, 100734.4, 100743.9, 
    100729.2,
  101043, 100968.3, 101047.5, 101001.2, 100970, 100911.6, 100831.7, 100742.8, 
    100659.4, 100646.5, 100664.3, 100705.6, 100728, 100754.1, 100747.4,
  99350.59, 99091.42, 100997.4, 101040.9, 100988.7, 100923.3, 100865.1, 
    100765.3, 100675.7, 100625.3, 100633.9, 100674.6, 100702.7, 100745.9, 
    100757.9,
  97455.74, 97583.24, 100903, 101079, 101023.2, 100966.4, 100908.3, 100833.2, 
    100720.6, 100638.3, 100616, 100641.3, 100688.3, 100726, 100759.5,
  97522.54, 97945.98, 99680.29, 101094.8, 101044.1, 100965.9, 100918.3, 
    100863.5, 100750.2, 100668.3, 100600, 100613.8, 100648.5, 100725.3, 
    100758.2,
  96945.45, 98374.42, 101028, 101092.6, 101045.2, 100913.1, 100969.3, 
    100913.1, 100842.6, 100696, 100581.7, 100542.6, 100636.3, 100719.2, 
    100755.6,
  101142.8, 101171.4, 101156.4, 101140.3, 101072.1, 99281.95, 100674.5, 
    100692.8, 100770.7, 100739.6, 100661.1, 100584.7, 100623.2, 100706.5, 
    100754.8,
  101216.9, 101185.4, 101173.8, 101141.5, 100919.4, 98563.66, 96699.38, 
    95865.05, 98253.86, 100810.7, 100705, 100622.2, 100633.5, 100701.5, 
    100755.9,
  101236.3, 101198, 101197.6, 101132.5, 96432.73, 97880.75, 99419.16, 
    100908.2, 100954.5, 100874.5, 100813.9, 100662.5, 100654.1, 100709, 
    100763.8,
  101273.4, 101232.8, 101234.9, 101128.7, 97000.28, 97234.13, 96637.04, 
    100985.6, 101067.5, 100937.6, 100853.5, 100807.8, 100702.3, 100741.3, 
    100778.8,
  101133.3, 101121.7, 101105.1, 101082.3, 101060, 101022.6, 100991.2, 
    100951.6, 100921.4, 100905.6, 100903.6, 100887.5, 100877.8, 100874.2, 
    100865.1,
  101124.5, 101078.9, 101153.2, 101138.9, 101126.8, 101089.3, 101052.1, 
    101004.3, 100969.8, 100939.5, 100927.4, 100919.6, 100913.1, 100905, 
    100903.1,
  99468.5, 99230.67, 101130.2, 101188.3, 101172.1, 101141.2, 101104.4, 
    101061, 101015, 100976.2, 100959.2, 100955.2, 100949.7, 100943.9, 100941.7,
  97584.42, 97727.3, 101064.7, 101240.1, 101224.6, 101203.5, 101173.4, 
    101130.2, 101078.9, 101021.2, 100985.1, 100980.5, 100980, 100955.9, 100984,
  97624.98, 98061.59, 99855.72, 101274.7, 101266.3, 101225.1, 101215.9, 
    101178.9, 101146, 101085.7, 101033.4, 101010.7, 101003.8, 101004.7, 
    101014.6,
  97042.97, 98468.75, 101176, 101270.6, 101283.5, 101180.3, 101273.4, 
    101238.7, 101216.4, 101154.5, 101083, 101000.3, 101036.8, 101033.9, 
    101038.5,
  101183.1, 101257.3, 101315.6, 101308, 101274.8, 99512.43, 100981, 101056.6, 
    101166.7, 101181, 101153.9, 101106.3, 101076.3, 101070.4, 101063.2,
  101271.9, 101290.2, 101319, 101311.8, 101140.7, 98820.3, 96995.42, 
    96170.55, 98646.98, 101243.9, 101213, 101157.8, 101108.9, 101087.7, 
    101085.5,
  101250.8, 101291.6, 101336.3, 101316.8, 96647.29, 98124.91, 99712.52, 
    101248.2, 101349.3, 101315.2, 101266.1, 101211.8, 101154.2, 101107, 
    101106.8,
  101284.4, 101320.8, 101353.5, 101315, 97196.91, 97478.13, 96895.18, 
    101293.7, 101416.1, 101360.6, 101313, 101247.5, 101195.3, 101137.8, 
    101120.9,
  101052.8, 100996, 100879.9, 100837.6, 100797.6, 100748.1, 100673.6, 100600, 
    100576.2, 100603.2, 100635.1, 100669.5, 100689.9, 100713, 100711.4,
  101104.9, 101067.1, 101079, 101008.2, 100928.3, 100830.5, 100767.1, 100708, 
    100675.4, 100683.4, 100722.6, 100772.7, 100797.4, 100817.3, 100811.5,
  99473.13, 99218.54, 101077.8, 101086.9, 101049.1, 100968.8, 100894.3, 
    100801.7, 100771.5, 100762.1, 100790.6, 100842.9, 100891.2, 100890.5, 
    100882.6,
  97657.75, 97765.73, 101061.8, 101206.7, 101145.7, 101076.8, 101028.2, 
    100929.8, 100868.7, 100843.8, 100869.9, 100906, 100960.8, 100974.8, 100975,
  97714.03, 98132.91, 99886.96, 101263, 101254.2, 101175.6, 101136.4, 
    101062.5, 100988.7, 100949.8, 100962.3, 100990.5, 101028.9, 101069.5, 
    101060.7,
  97140.19, 98573.48, 101251.8, 101307.6, 101298.9, 101184.1, 101240.9, 
    101180.6, 101140.1, 101063.8, 101040.1, 101022.4, 101104.6, 101131.2, 
    101143.3,
  101273.1, 101338, 101402.8, 101381.4, 101339.8, 99589.85, 101031.3, 
    101044.7, 101142, 101145.4, 101140.5, 101131.9, 101166.9, 101189.4, 
    101193.3,
  101353, 101385.6, 101453.5, 101442.8, 101259.1, 98872.45, 97053.79, 
    96239.73, 98699.17, 101264.7, 101252.6, 101226.9, 101233.2, 101233.4, 
    101246.4,
  101334.9, 101385, 101477.3, 101439.8, 96799.37, 98262.25, 99829.38, 
    101356.5, 101426.6, 101386.1, 101348.8, 101321.7, 101305.5, 101292.5, 
    101289.9,
  101352.2, 101410.9, 101503.5, 101466.9, 97363.71, 97603.4, 97048.45, 
    101458.2, 101559.8, 101494.9, 101440.4, 101400.9, 101375.7, 101353.5, 
    101344.4,
  100784.1, 100694, 100597.8, 100471.3, 100367.8, 100275, 100199.6, 100189, 
    100228.9, 100295.1, 100350, 100407.1, 100424.4, 100469.7, 100490.6,
  100776.1, 100655.7, 100642.1, 100498.4, 100353.5, 100212.5, 100084.8, 
    100067.2, 100111.5, 100188, 100261.6, 100342.9, 100378.6, 100456.5, 
    100493.6,
  99097.39, 98793.1, 100595.1, 100555.4, 100379.2, 100224.2, 100033.8, 
    99948.04, 99979.34, 100070.4, 100156.7, 100263.1, 100336.6, 100413.8, 
    100468,
  97270.29, 97355.2, 100496.5, 100594.8, 100439, 100253.9, 100085, 99924.77, 
    99893.15, 99966.96, 100063.8, 100181.7, 100283.4, 100361, 100458.2,
  97333.12, 97701.14, 99358.44, 100606.1, 100484.6, 100253.6, 100102.6, 
    99927.8, 99833.11, 99877.11, 99987.2, 100116.1, 100232.3, 100344.4, 
    100448.2,
  96826.39, 98178.69, 100721.9, 100631.3, 100519.3, 100249.1, 100132.8, 
    99959.66, 99833.52, 99831.88, 99928.7, 100037.2, 100222.6, 100348.2, 
    100453.8,
  100996.1, 100946.9, 100875.4, 100712.9, 100561.3, 98664.89, 99858.69, 
    99723.57, 99760.15, 99795.3, 99915.23, 100061.6, 100212.6, 100351.9, 
    100464,
  101078.8, 100995.4, 100951.7, 100773.8, 100387.2, 97983.59, 95997.67, 
    95008.83, 97332.3, 99865.62, 99943.53, 100070.7, 100221.1, 100368.5, 
    100482.6,
  101114.6, 101034.1, 101018.7, 100804.1, 96024.32, 97395.77, 98767.6, 
    100070.4, 100002, 99997.29, 100022.3, 100129.4, 100255.5, 100400.5, 
    100521.9,
  101165.8, 101097.3, 101109.2, 100881.2, 96705.71, 96824.15, 96081.76, 
    100295.8, 100248.8, 100158.5, 100156.7, 100238.2, 100333.6, 100459.4, 
    100572.2,
  100178.8, 100212.7, 100255.5, 100290, 100321.4, 100351.1, 100376.9, 
    100400.7, 100426.8, 100458.1, 100477, 100502.5, 100510.7, 100523.5, 
    100533.8,
  100131.9, 100119.7, 100233.4, 100263.3, 100289.2, 100320.7, 100347.4, 
    100375.8, 100406, 100435.2, 100457.5, 100479.8, 100502.6, 100530.7, 
    100550.6,
  98447.94, 98220.97, 100102.3, 100226.6, 100243, 100272.8, 100290.1, 
    100315.2, 100342.1, 100379.7, 100415.2, 100447.4, 100479.6, 100506.4, 
    100537,
  96563.8, 96715.43, 99981.49, 100222.4, 100213.9, 100229.8, 100234.8, 
    100256.3, 100284.9, 100320, 100358.3, 100398.4, 100446.6, 100468.6, 
    100525.2,
  96622.66, 97062.79, 98784.12, 100183.3, 100169, 100132.5, 100131.8, 
    100137.6, 100171, 100225, 100281.8, 100332.3, 100387.1, 100443, 100494.6,
  96087.73, 97475.01, 100060.8, 100133.3, 100085.1, 99972.73, 100037, 
    100037.3, 100062.1, 100115.4, 100175.3, 100202, 100322.3, 100398, 100459,
  100202.8, 100225.6, 100172.6, 100110.1, 100031.4, 98226, 99533.05, 
    99652.29, 99826.67, 99947.03, 100063, 100146.4, 100244, 100333.1, 100413.5,
  100266.8, 100216.2, 100147.4, 100042.9, 99703.34, 97376.09, 95556.27, 
    94692.2, 97047.34, 99742.75, 99923.13, 100032.4, 100146.7, 100257.9, 
    100357.8,
  100267.2, 100191.6, 100151.3, 100021.7, 95247.4, 96530.97, 97968.14, 
    99427.38, 99599.91, 99681.73, 99783.28, 99909.03, 100044.9, 100174.1, 
    100292.8,
  100287.2, 100188.1, 100161.5, 99976.6, 95779.69, 95884.8, 95192.39, 
    99352.12, 99542.07, 99557.84, 99678.8, 99804.69, 99952.15, 100092.3, 
    100228.4,
  99531.5, 99601.41, 99710.88, 99805.33, 99887.31, 99957.27, 100012.5, 
    100068.9, 100114.1, 100171.4, 100231.4, 100288.3, 100332.8, 100397.5, 
    100461.4,
  99421.34, 99519.31, 99676.55, 99778.82, 99865.43, 99950.04, 100022.6, 
    100075.9, 100124.8, 100175.3, 100227.4, 100281.9, 100348.3, 100430.7, 
    100493.2,
  97781.84, 97674.45, 99567.46, 99773.14, 99851.08, 99946.41, 100021.2, 
    100082.8, 100125.9, 100175, 100234.1, 100291, 100373.2, 100443, 100509.1,
  95877.34, 96105.2, 99466.15, 99752.74, 99837.85, 99943.63, 100026.4, 
    100095.6, 100133.6, 100175.3, 100241.9, 100309.3, 100389.9, 100441.6, 
    100533.6,
  95883.21, 96414.45, 98266.47, 99743.57, 99835.45, 99912.7, 100009.6, 
    100069.8, 100119.2, 100179.7, 100252.4, 100327.3, 100394.1, 100468.8, 
    100552.4,
  95320.97, 96779.92, 99504.21, 99729.65, 99827.02, 99867.31, 100012.6, 
    100080.8, 100133.4, 100190.4, 100249.8, 100292.9, 100414.2, 100491.3, 
    100566.1,
  99357.72, 99509.94, 99679.06, 99756.34, 99806.01, 98202.07, 99694.63, 
    99858.15, 100055.1, 100158.3, 100270.4, 100344.4, 100432.5, 100507.7, 
    100579.1,
  99503.7, 99558.97, 99665.6, 99709.89, 99658.39, 97393.83, 95730.3, 
    95008.64, 97472.84, 100146.3, 100275, 100353.6, 100443.4, 100521.4, 
    100593.5,
  99465.16, 99546.85, 99686.03, 99695.2, 95234.91, 96624.68, 98211.89, 
    99713.03, 99995.09, 100157.2, 100262.7, 100349.4, 100445.3, 100532.2, 
    100606.2,
  99534.35, 99589.09, 99695.89, 99671.25, 95673.27, 95978.66, 95555.05, 
    99834.37, 100103.9, 100139.6, 100254.3, 100346.2, 100443.7, 100532.6, 
    100612.7,
  99565.38, 99665.12, 99780.76, 99913.84, 100033.3, 100148.2, 100244.6, 
    100347, 100422.6, 100468, 100480.5, 100517.6, 100546.6, 100502.9, 100515.6,
  99420.85, 99515.41, 99706.94, 99863.52, 99999.77, 100127.9, 100231.4, 
    100347.5, 100414.5, 100456.8, 100472, 100503.1, 100524.6, 100514, 100531.4,
  97757.17, 97645.33, 99570.98, 99830.34, 99969.34, 100112.4, 100232.4, 
    100331.5, 100394.9, 100435.5, 100454.6, 100479.2, 100508.3, 100501.5, 
    100521,
  95795.55, 96032.91, 99436.85, 99782.36, 99940.06, 100099.5, 100229.7, 
    100330.6, 100389, 100421.4, 100432.9, 100457.3, 100491.7, 100478.8, 
    100522.9,
  95758.75, 96320.75, 98221.26, 99762.96, 99928.59, 100072.7, 100217.1, 
    100305, 100356.5, 100393.3, 100411.1, 100443, 100460.1, 100482.4, 100535.6,
  95148.95, 96645.38, 99444.43, 99735.85, 99896.47, 100024.7, 100222.5, 
    100323.3, 100364.2, 100383.9, 100384, 100385.1, 100461.8, 100492.9, 
    100539.2,
  99165.02, 99378.44, 99615.14, 99742.95, 99869.74, 98371.03, 99911.74, 
    100090.1, 100256.7, 100333.4, 100380.2, 100419.8, 100454.8, 100495.4, 
    100549.5,
  99316.84, 99400.55, 99579.78, 99659.55, 99719.12, 97545.38, 95920.54, 
    95186.88, 97636.36, 100295.4, 100357.7, 100412, 100449.8, 100496.7, 
    100561.7,
  99250.07, 99374.37, 99576.84, 99626.94, 95315.41, 96771.23, 98440.52, 
    99958.46, 100223.4, 100307.9, 100340.9, 100406.4, 100446.6, 100493.5, 
    100575.3,
  99278.98, 99406.66, 99571.59, 99603.2, 95757.35, 96106.42, 95750.04, 
    100081.8, 100305.3, 100278.9, 100333.3, 100405, 100449.3, 100491.5, 
    100590.3,
  100086.5, 100159.6, 100229.4, 100309.3, 100391.2, 100464.4, 100544.8, 
    100625.6, 100700.5, 100775.9, 100816.4, 100854.6, 100898.3, 100855.2, 
    100803.8,
  99977.44, 100032.1, 100169, 100267.5, 100364.2, 100450.2, 100531.2, 100620, 
    100694.9, 100786.4, 100815.2, 100854.4, 100958.9, 100910.5, 100869.2,
  98272.05, 98131.68, 100035.5, 100231.7, 100326.5, 100426.1, 100513.1, 
    100606.5, 100685.8, 100778.9, 100816.5, 100862.7, 100957.3, 100927.9, 
    100890.4,
  96299.31, 96507.88, 99874.28, 100186, 100291.8, 100416.7, 100508.4, 
    100609.3, 100691.6, 100774.9, 100824.3, 100866.7, 100967.8, 100927.3, 
    100899.3,
  96245.97, 96765.7, 98612.05, 100141.7, 100259, 100367.7, 100486.8, 
    100586.5, 100674.6, 100763.7, 100833.8, 100862.7, 100972.7, 100936.2, 
    100894.9,
  95577.2, 97064.03, 99795.59, 100076.8, 100210.3, 100310.5, 100485.1, 
    100592.2, 100692.5, 100776.4, 100823.7, 100828.6, 100977.2, 100947.6, 
    100899.1,
  99557.19, 99741.54, 99921.17, 100062.4, 100175.6, 98637.34, 100185.8, 
    100392.4, 100630.6, 100748.2, 100840.8, 100888.5, 100979.5, 100954.1, 
    100900.6,
  99642.48, 99739.51, 99868.67, 99980.71, 99999.27, 97803.73, 96213.69, 
    95531.5, 98057.65, 100738.7, 100847.8, 100900.8, 100975.9, 100966.4, 
    100909.3,
  99558.59, 99669.11, 99850.46, 99935.57, 95555.84, 97018.19, 98693.22, 
    100253.6, 100616, 100751.9, 100845.3, 100906.2, 100968, 100971.3, 100912.4,
  99543.5, 99664.41, 99829.23, 99882.52, 95974.86, 96351.73, 96052.38, 
    100416.1, 100733.1, 100736.5, 100864.1, 100907.4, 100979.8, 100978.7, 
    100914,
  100656.7, 100670.1, 100699.9, 100733.4, 100772.6, 100799.2, 100833.9, 
    100855.8, 100845.4, 100818.8, 100753.5, 100691.7, 100650.9, 100601.9, 
    100660.9,
  100621.4, 100606.8, 100699.5, 100728.8, 100771.1, 100818.1, 100860.3, 
    100890.9, 100890.8, 100864.8, 100815.9, 100748.1, 100762.7, 100741.9, 
    100735.2,
  98950.13, 98728.16, 100607.1, 100731.9, 100767.1, 100813.2, 100857.3, 
    100900.1, 100916.6, 100909.7, 100885.5, 100816.4, 100801.5, 100793.2, 
    100799.1,
  97030.36, 97166.78, 100492.5, 100736.3, 100763.4, 100827.4, 100875.7, 
    100932, 100959.6, 100963.3, 100961.9, 100925.9, 100886.4, 100875.2, 
    100890.4,
  97041.45, 97482.58, 99268.2, 100730.6, 100765.4, 100797.8, 100865.6, 
    100923.5, 100968, 100988, 101012.7, 101003.3, 100960.8, 100976.4, 100974.8,
  96434.8, 97857.19, 100520.5, 100707, 100753.5, 100768.9, 100896.6, 
    100955.9, 101009.5, 101029.9, 101052.8, 101022.4, 101049.5, 101063.1, 
    101050,
  100619.3, 100623.9, 100667.6, 100730.4, 100751, 99084.05, 100585.4, 
    100759.8, 100946.2, 101022.2, 101095.2, 101101.1, 101104.6, 101105.9, 
    101108.3,
  100715.9, 100656.5, 100665.1, 100687, 100592, 98306.73, 96619.95, 95879.09, 
    98368.68, 101040.6, 101122.2, 101140, 101149.6, 101151.4, 101156.5,
  100664.1, 100643.1, 100687.4, 100688.7, 96144.34, 97531.32, 99144.52, 
    100666.1, 100943.3, 101068.7, 101133.1, 101162, 101178.7, 101179.6, 101178,
  100655.1, 100656.8, 100701.7, 100659, 96603.23, 96888.01, 96450.69, 
    100782.8, 101050, 101065.5, 101148.5, 101182.9, 101214.7, 101214.6, 
    101201.1,
  100569, 100587.9, 100588.1, 100577.2, 100548, 100496.3, 100457.4, 100425.4, 
    100415.1, 100433.6, 100473, 100544.8, 100593.4, 100652.9, 100708.3,
  100539, 100543.2, 100615.9, 100596, 100558, 100512.5, 100461.1, 100420.2, 
    100394.7, 100403.1, 100450.4, 100524, 100596.5, 100679.7, 100739.7,
  98921.03, 98714.7, 100577.5, 100642.3, 100587.5, 100506.9, 100419.4, 
    100394.9, 100406, 100423.6, 100453.4, 100524.8, 100612.8, 100684.1, 
    100764.8,
  97071.1, 97230.21, 100511.1, 100680.7, 100610.8, 100521.9, 100472.4, 
    100412.8, 100390.7, 100419.4, 100468.2, 100527.6, 100630.1, 100696.3, 
    100814.5,
  97110.84, 97567.42, 99329.2, 100725, 100640.8, 100571, 100488, 100417.4, 
    100445.9, 100493.4, 100541.9, 100598.7, 100675.9, 100779.3, 100881.6,
  96606.74, 98003.87, 100655.2, 100732.7, 100666.1, 100563.5, 100560.9, 
    100542.2, 100538.9, 100570.2, 100597.6, 100632.4, 100758.5, 100860.7, 
    100944.8,
  100760.1, 100799.6, 100821.4, 100782.8, 100700.4, 98957.56, 100340.9, 
    100389.4, 100517.6, 100622.8, 100706.4, 100764.9, 100850.2, 100932.8, 
    100994.3,
  100904.7, 100865.8, 100864.8, 100793.9, 100609, 98246.35, 96428.32, 
    95624.98, 98095.91, 100730.3, 100798.4, 100867.7, 100943, 101004.3, 
    101055.1,
  100938.5, 100912.8, 100929.9, 100818.6, 96242.4, 97636.27, 99173.89, 
    100620.3, 100777.8, 100839.9, 100902.3, 100958.3, 101031.2, 101088.7, 
    101125.8,
  101028.2, 101005.2, 101005.5, 100867.9, 96812.21, 97052.26, 96520.77, 
    100841.7, 100958.4, 100953.6, 101003.8, 101062.8, 101128.9, 101166.1, 
    101197.4,
  100511.7, 100467.6, 100439.8, 100354.8, 100342.8, 100245, 100181.4, 
    100111.6, 100129, 100251.3, 100352.6, 100468.3, 100553.9, 100639.2, 
    100703.8,
  100440.9, 100371.5, 100444.4, 100375.5, 100337.7, 100336.6, 100232.6, 
    100163.6, 100172.2, 100254.7, 100361, 100478.1, 100584.3, 100676.5, 
    100746.9,
  98736.28, 98462.24, 100318.8, 100405.8, 100323.5, 100356.6, 100251.3, 
    100200.5, 100182.1, 100282.2, 100364.7, 100487.3, 100611.7, 100696.7, 
    100767.7,
  96824.75, 96925.65, 100179.7, 100418.3, 100320.6, 100370, 100262.3, 
    100243.8, 100188.1, 100301.9, 100378.8, 100521.8, 100625.4, 100700.3, 
    100796,
  96800.47, 97233.44, 98950.35, 100394.4, 100311.3, 100310.7, 100238.5, 
    100253.1, 100213.8, 100309.9, 100391.9, 100542.8, 100632.3, 100732.5, 
    100822.1,
  96201.25, 97616.22, 100251.9, 100369, 100289, 100242.7, 100258.2, 100249.6, 
    100228.4, 100319.4, 100397.6, 100504.7, 100657.5, 100755.2, 100845.6,
  100324.9, 100389.2, 100378.7, 100372.8, 100299.8, 98554.88, 99926.02, 
    100083.1, 100196.4, 100316.3, 100425.1, 100564.8, 100682.4, 100778.4, 
    100871.6,
  100389, 100387, 100370.6, 100317.9, 100091.1, 97776.35, 96005.01, 95229.06, 
    97669.71, 100348.9, 100433.7, 100588.5, 100706.1, 100805.6, 100899.5,
  100387.9, 100389.7, 100383.3, 100302.2, 95623.87, 96944.48, 98511.09, 
    99982.78, 100253.7, 100388.3, 100460.2, 100610.1, 100737.9, 100836.6, 
    100934.8,
  100437.2, 100416.7, 100381.7, 100268.7, 96120.47, 96286.07, 95759.53, 
    100096.4, 100353.4, 100394.3, 100498.1, 100641.6, 100785.6, 100875.2, 
    100971.4,
  100748.4, 100720.9, 100700.5, 100677.3, 100669.1, 100639.8, 100618.3, 
    100595, 100587.7, 100592.3, 100612.7, 100630.6, 100664.8, 100720.9, 
    100770.4,
  100673.4, 100605.6, 100678.6, 100666.3, 100645.5, 100622, 100597.7, 
    100594.5, 100596, 100600.2, 100632, 100641.1, 100689.5, 100737.9, 100799.9,
  98947.49, 98669.77, 100543.9, 100628.3, 100619.6, 100594.7, 100560.9, 
    100548.5, 100565.7, 100588.9, 100628, 100636, 100713, 100750.7, 100819.7,
  97049.8, 97137.96, 100409.4, 100606.4, 100605.7, 100578.1, 100543.8, 
    100516.2, 100507.2, 100569.6, 100600.6, 100634.6, 100717.5, 100744, 
    100841.4,
  97049.78, 97458.1, 99170.61, 100592.3, 100592.7, 100524.7, 100497.6, 
    100438, 100413.1, 100494.1, 100555.4, 100627.7, 100705.3, 100764.3, 
    100858.9,
  96447.38, 97846.09, 100475.2, 100584.1, 100568.9, 100442.9, 100465.8, 
    100403.6, 100345.9, 100405.1, 100501.4, 100530.9, 100695, 100774.8, 
    100870.8,
  100625.3, 100642.4, 100639.1, 100606.1, 100571.5, 98772.58, 100134.9, 
    100209.3, 100234.4, 100275.5, 100471.6, 100539.2, 100688.8, 100780.3, 
    100882.9,
  100666, 100628.4, 100625.8, 100586.7, 100372.4, 98040.03, 96239.75, 
    95409.39, 97735.02, 100280.8, 100439.3, 100508.5, 100692, 100784, 100897.1,
  100614.3, 100614.6, 100646.7, 100611.9, 95921.03, 97268.25, 98824.52, 
    100369.2, 100416.8, 100355.9, 100431.2, 100515.5, 100698.8, 100797.8, 
    100916.7,
  100621.2, 100629.6, 100659, 100581.3, 96446.25, 96662.71, 96033.12, 
    100372.6, 100447.6, 100356.1, 100431.1, 100521.3, 100706.1, 100815.5, 
    100934.8,
  100840.8, 100803.6, 100770.6, 100713.5, 100603.8, 100512.4, 100382.5, 
    100250.5, 100202.6, 100256.2, 100378.2, 100499.6, 100616.8, 100712.7, 
    100783.2,
  100794.4, 100743.2, 100794.6, 100747.3, 100674.8, 100566.2, 100512.6, 
    100352, 100277.3, 100316.1, 100409.8, 100525.5, 100631, 100729, 100813.4,
  99144.67, 98901.35, 100754.9, 100788.8, 100708.5, 100589.8, 100509.2, 
    100415, 100337.8, 100369.6, 100449.8, 100541.2, 100646.4, 100741.2, 
    100832.8,
  97306.92, 97422.78, 100698, 100843.4, 100762.5, 100688.5, 100574.8, 100493, 
    100404.3, 100437, 100495.5, 100566.2, 100670.6, 100749.9, 100861.7,
  97380.83, 97798.93, 99520.71, 100893.7, 100793.1, 100723.2, 100634.5, 
    100524.8, 100456.9, 100490.5, 100539.7, 100601.1, 100696.8, 100788.4, 
    100893.9,
  96906.52, 98291.87, 100879.8, 100924.1, 100828.7, 100698.8, 100739.1, 
    100624.7, 100574.4, 100552.3, 100583.4, 100596.7, 100736.9, 100827.3, 
    100926,
  101125.6, 101094.7, 101030.4, 100981, 100862.5, 99052.26, 100500.1, 
    100492.9, 100595.1, 100614.5, 100667.5, 100712.9, 100780.6, 100869.3, 
    100957.4,
  101156.6, 101086.4, 101042.4, 100975.6, 100698.7, 98333.82, 96509.98, 
    95672.18, 98136.14, 100738.3, 100762, 100780.9, 100830.2, 100914.1, 
    100990.2,
  101140.1, 101084.4, 101072.7, 100998.5, 96213.02, 97622.02, 99183.71, 
    100689.2, 100818.7, 100831.1, 100847.7, 100857.8, 100875.5, 100962, 
    101021.6,
  101154.2, 101101.8, 101085.7, 101009.4, 96776.25, 96998.26, 96403.44, 
    100750.8, 100911.9, 100882.3, 100903.4, 100903.3, 100917, 101000.6, 101058,
  101027.9, 101020.7, 101008, 100998.9, 101008.6, 100992.9, 100976.4, 
    100967.8, 100964, 100955.8, 100941.9, 100941, 100941.3, 100926.3, 100963.5,
  101018.6, 100937.8, 101018.8, 100991.7, 100974.7, 100962.8, 100945.3, 
    100936.6, 100930.3, 100930.5, 100931.7, 100931.3, 100930.4, 100932.3, 
    100963.8,
  99317.52, 99038.68, 100931.1, 101032.7, 100973.7, 100938.7, 100897.7, 
    100881.1, 100877.2, 100879.7, 100883.4, 100898.4, 100909.6, 100925.5, 
    100942.7,
  97479.18, 97589.48, 100841.9, 101035.6, 100953.5, 100901.6, 100855.2, 
    100828.2, 100814, 100819.1, 100831.9, 100860.1, 100887.3, 100897.9, 
    100939.2,
  97514.28, 97934.78, 99623.67, 101012.9, 100924.6, 100827.6, 100774.9, 
    100736.7, 100703.4, 100730.9, 100760.1, 100809.7, 100846.4, 100889.6, 
    100933.4,
  97021.56, 98390.82, 100966.4, 100997, 100870.1, 100718.8, 100725.3, 
    100662.6, 100607.2, 100623.5, 100667.5, 100701.6, 100814.7, 100875.5, 
    100930.7,
  101271.7, 101186.7, 101076.5, 100992.5, 100830.6, 99020.34, 100315.2, 
    100353.6, 100416.5, 100470.6, 100573.6, 100662.9, 100764.9, 100848.4, 
    100920.6,
  101283.7, 101180, 101086, 100961.6, 100580.3, 98256.29, 96349.46, 95503.33, 
    97792.75, 100385.1, 100511.9, 100604.3, 100714.4, 100820.4, 100909.3,
  101295.6, 101179.8, 101100.3, 100951.9, 96086.25, 97489.76, 98936.34, 
    100404.9, 100410.1, 100366.8, 100458.4, 100553.9, 100672.8, 100796.4, 
    100896.2,
  101302.1, 101185, 101118, 100947.7, 96651.98, 96859.16, 96169.38, 100413, 
    100454.8, 100312, 100411.6, 100516.8, 100643.6, 100776.6, 100889.8,
  101430.6, 101420.7, 101397.2, 101356.6, 101328.5, 101288.8, 101248.6, 
    101233.8, 101169.2, 101101.2, 101026.6, 100984.9, 100942.5, 100948.2, 
    100939.4,
  101454.1, 101373, 101449, 101393.7, 101366.2, 101320.1, 101266.6, 101274.4, 
    101234, 101166.6, 101109.4, 101052.5, 100991.8, 100981.6, 100963.8,
  99759.84, 99469.63, 101415.2, 101447.5, 101390.9, 101339.1, 101282.7, 
    101270.8, 101251.2, 101194.7, 101134.3, 101099.2, 101033.6, 101001.2, 
    100987.3,
  97864.45, 97998.91, 101312, 101478.6, 101407.4, 101348.7, 101304, 101268.1, 
    101279.8, 101241.2, 101175.4, 101144.1, 101086.2, 101027.2, 101012.6,
  97950.41, 98361.02, 100098, 101494.9, 101415.3, 101317.1, 101291.9, 
    101256.7, 101271.1, 101249.9, 101193.2, 101170.5, 101120.2, 101092, 
    101057.8,
  97382.84, 98821.4, 101470, 101502, 101416.1, 101240.8, 101263.6, 101253.5, 
    101266.6, 101262.5, 101209.5, 101139.9, 101158, 101124.8, 101087.7,
  101671.4, 101665.4, 101597, 101543, 101432.8, 99556.7, 100947.4, 101032, 
    101182.5, 101216, 101223.9, 101192, 101179, 101153.4, 101122.7,
  101705.7, 101659, 101614.4, 101535.1, 101239.8, 98835.38, 96958.62, 
    96109.12, 98556.05, 101225.9, 101241.9, 101208.8, 101199.6, 101178.3, 
    101151.9,
  101697.2, 101651.9, 101626.8, 101552, 96689.72, 98089.68, 99616.59, 
    101141.1, 101295.8, 101263.9, 101250, 101225.6, 101217.1, 101199.7, 
    101177.3,
  101690.8, 101645.1, 101629.8, 101542.4, 97263.73, 97479.34, 96807.86, 
    101154.7, 101319, 101263.8, 101266.4, 101245.8, 101250.7, 101226.2, 101207,
  101502.2, 101459.2, 101426.6, 101349.9, 101302.4, 101241.6, 101158.9, 
    101084.4, 100992.5, 100954, 100908, 100895.4, 100893.6, 100953, 100960.4,
  101517, 101427.6, 101470.5, 101388.6, 101332, 101312.2, 101229.1, 101152.8, 
    101059.1, 101021.3, 100972, 100936.7, 100940, 100986.6, 100978.9,
  99824.24, 99544.55, 101446.3, 101469.4, 101364.8, 101333.8, 101266.7, 
    101205.7, 101102.9, 101063.1, 101012, 101010.1, 100947.3, 101010.6, 
    100998.5,
  97954.47, 98074.72, 101361.3, 101507.5, 101410.9, 101372, 101340.5, 
    101262.9, 101167.3, 101107.8, 101052.3, 101026.2, 100998.8, 101003.4, 
    101032.6,
  98030.46, 98436.83, 100176.9, 101540.1, 101447.5, 101386, 101363.7, 
    101289.6, 101220.6, 101149.2, 101083.8, 101032.3, 101015.1, 101044, 
    101062.4,
  97494.02, 98932.84, 101539.7, 101548.4, 101470.1, 101345.6, 101432, 
    101365.4, 101296.2, 101215.5, 101115.8, 101018.6, 101053, 101069.5, 
    101088.1,
  101753.1, 101749.2, 101665.5, 101604.8, 101502, 99717.93, 101143.8, 
    101148.8, 101241.1, 101241.6, 101182.4, 101111.7, 101114, 101101.2, 
    101122.9,
  101827.3, 101775.8, 101715.1, 101631.8, 101362.8, 98988.51, 97121.09, 
    96281.96, 98723.36, 101307.1, 101231.5, 101186.4, 101163.4, 101141.7, 
    101160.4,
  101867.5, 101796.3, 101768.5, 101627.7, 96878.62, 98343.81, 99880.79, 
    101384.3, 101422, 101368.4, 101279.3, 101230.2, 101210.8, 101197.6, 
    101202.4,
  101914.2, 101851.1, 101851.9, 101687.2, 97481.14, 97698.54, 97073.42, 
    101479.6, 101527.8, 101461.4, 101361.7, 101299.4, 101293.5, 101252.5, 
    101245,
  101336.9, 101270.7, 101241.7, 101140.3, 101049.8, 100932.6, 100803.9, 
    100726, 100754.1, 100837.5, 100915.9, 100977, 101023.3, 101050.6, 101051.1,
  101329.2, 101223, 101272.5, 101180.7, 101095.1, 101011.2, 100871.2, 100772, 
    100815, 100873.7, 100947.5, 101015, 101047.3, 101078.2, 101087.9,
  99627.1, 99345.38, 101227.4, 101240.1, 101132.5, 101028.1, 100939.1, 
    100830.7, 100841.3, 100913.3, 100969.5, 101036.6, 101063.2, 101101.1, 
    101115.1,
  97776.71, 97875.41, 101126, 101280.1, 101189.6, 101089.5, 101017.8, 
    100904.4, 100894.2, 100951.8, 101008.3, 101059.1, 101101.3, 101111.6, 
    101152.7,
  97833.02, 98229.08, 99930.34, 101302.3, 101219.1, 101104.5, 101032.4, 
    100963.6, 100952.5, 100999.2, 101039.1, 101085.7, 101111.7, 101157.4, 
    101178.3,
  97312.95, 98709.78, 101275.2, 101302.6, 101217.9, 101085.3, 101101.7, 
    101043.9, 101016.1, 101048.4, 101069.8, 101050.3, 101156, 101193.2, 
    101210.3,
  101504.8, 101479, 101397.2, 101347, 101228.1, 99450.1, 100814, 100888, 
    100991.4, 101053.6, 101110.6, 101132.6, 101194.4, 101217.8, 101243.1,
  101564.9, 101501, 101430.7, 101337.9, 101008, 98695.75, 96829.32, 95997.02, 
    98448.09, 101100.8, 101148.2, 101164, 101229.2, 101252.1, 101283.9,
  101593.9, 101506.2, 101463.2, 101333.1, 96560.5, 97939.41, 99455.14, 
    100931.3, 101082.5, 101149.6, 101174.4, 101208.2, 101266.2, 101290, 101318,
  101636.9, 101542.2, 101512.8, 101342.3, 97136.8, 97267.12, 96641.56, 
    100963.1, 101116.1, 101153.2, 101193.9, 101258.5, 101312, 101334.4, 101360,
  101152.2, 101123.1, 101139.6, 101114.4, 101114.9, 101110.7, 101118.5, 
    101131, 101162.2, 101196.1, 101226.6, 101255.2, 101273.6, 101258.9, 101245,
  101135.4, 101068.6, 101155.6, 101133.9, 101135.2, 101127.9, 101131.8, 
    101143.6, 101184, 101219.6, 101251.2, 101284.5, 101304.3, 101305.8, 
    101296.8,
  99459.81, 99215.09, 101100.8, 101168.5, 101142.3, 101118.2, 101130.3, 
    101132.6, 101178.4, 101224.6, 101264.7, 101318, 101338.6, 101331.9, 
    101328.4,
  97602.44, 97742.91, 100991.7, 101178.9, 101134.3, 101111.2, 101114.4, 
    101124.5, 101176.7, 101228.8, 101286.2, 101348.1, 101373.5, 101352.5, 
    101377.5,
  97657.69, 98081.16, 99803.31, 101174.7, 101116.6, 101059, 101063.4, 
    101078.7, 101160.8, 101224.6, 101298.4, 101367.9, 101386.1, 101400.8, 
    101401.8,
  97138.89, 98556.43, 101119.7, 101156.9, 101083.1, 100948.8, 101036.2, 
    101051.3, 101154.9, 101220.3, 101303.8, 101333.1, 101411.5, 101435.9, 
    101429.5,
  101308.2, 101323.3, 101253, 101194.9, 101054.1, 99300.77, 100739, 100866.5, 
    101084.3, 101199, 101335.4, 101397.1, 101440.6, 101462.1, 101456.6,
  101378.8, 101336.7, 101288.8, 101181.2, 100867.9, 98567.69, 96760.84, 
    96010.3, 98532.35, 101218.4, 101359.3, 101426.2, 101475.1, 101491.1, 
    101490.1,
  101384, 101334.4, 101321.4, 101200.9, 96456.08, 97875.56, 99373.57, 
    100856.2, 101133.6, 101285, 101387.6, 101461.9, 101491.5, 101524.4, 
    101522.8,
  101397.5, 101352.4, 101335.8, 101229.1, 97027.88, 97238.6, 96656.88, 
    101018.7, 101256.4, 101315.7, 101413, 101491.6, 101536.1, 101555.1, 
    101556.5,
  100517.5, 100525.4, 100573.1, 100637.5, 100708.5, 100785.1, 100867.3, 
    100953.3, 101021.1, 101078.8, 101121, 101176, 101207.9, 101234, 101242.2,
  100471.1, 100488.2, 100603.4, 100678.8, 100751, 100832.3, 100918.4, 
    101002.9, 101073.1, 101123.5, 101166.5, 101208.2, 101238.9, 101270.5, 
    101278.9,
  98830.44, 98657.7, 100552.1, 100711.8, 100788.6, 100878.2, 100962.1, 
    101040.6, 101108.7, 101164.4, 101211.8, 101250.3, 101286.9, 101302.4, 
    101318.4,
  96955.7, 97166.26, 100499.2, 100750.9, 100837.9, 100926.1, 101004.9, 
    101083.4, 101154.7, 101206.2, 101247.5, 101293.1, 101327.9, 101328.3, 
    101364.9,
  97002.26, 97495, 99308.23, 100801.1, 100875.7, 100950.8, 101050.8, 101125, 
    101190.2, 101246.7, 101292.1, 101338.1, 101355.2, 101384.1, 101396.9,
  96516.44, 97968.16, 100620, 100812.9, 100903.9, 100932.2, 101092.4, 
    101168.9, 101245.3, 101290.8, 101325.6, 101321.9, 101408.5, 101422.3, 
    101431.4,
  100658.6, 100734.7, 100793.3, 100872, 100918.8, 99323.27, 100856.8, 
    101022.2, 101215.8, 101300.5, 101373.8, 101405.5, 101443.9, 101461.7, 
    101470.5,
  100788.2, 100833.2, 100859, 100897.8, 100803, 98521.72, 96846.06, 96116.63, 
    98652.81, 101339, 101407.1, 101441.6, 101479.7, 101501.7, 101508.1,
  100857.8, 100895.4, 100942.8, 100878.5, 96375.62, 97846.97, 99461.09, 
    100993.2, 101279.2, 101390.2, 101443.1, 101478.4, 101518.6, 101541.2, 
    101545.7,
  100993, 100992.7, 101030.7, 100936.1, 96903.13, 97218.71, 96727.41, 
    101138.6, 101365.7, 101408.3, 101473.7, 101516.4, 101555.4, 101581.9, 
    101570.1,
  100896.5, 100915.2, 101005.4, 100964.6, 101042.7, 101036.5, 101058.4, 
    101068.4, 101110.2, 101131.5, 101160.7, 101199.3, 101229.3, 101255.1, 
    101255.3,
  100834.8, 100837.6, 101004.9, 101015.3, 101053.1, 101065.4, 101080.3, 
    101076.6, 101136, 101166.8, 101179.7, 101221.8, 101253.7, 101278, 101289.8,
  99156.53, 98972.2, 100884.7, 101020.8, 101026.2, 101102.1, 101126.5, 
    101159.9, 101174.4, 101208.8, 101222.9, 101261.7, 101286.9, 101305.4, 
    101319.2,
  97234.88, 97380.38, 100742.9, 101014.4, 101035.7, 101082.1, 101159.4, 
    101170.4, 101212.3, 101250.5, 101256.7, 101291, 101317.7, 101323, 101354.7,
  97204.09, 97669.57, 99474.71, 100971.9, 101045.4, 101046.5, 101152.1, 
    101178.5, 101232.6, 101277.7, 101286.9, 101323.2, 101343.9, 101361.8, 
    101382.9,
  96554.88, 97988.73, 100670.4, 100911.3, 101033.1, 101005.1, 101181.3, 
    101190.7, 101238, 101311.2, 101309, 101300.2, 101380.8, 101395.5, 101407.1,
  100612, 100667.8, 100798.6, 100896.2, 101008.5, 99343.22, 100884.8, 
    101008.7, 101189.6, 101285.1, 101350.7, 101373, 101415.4, 101425.7, 
    101433.7,
  100719.2, 100715.5, 100788.5, 100841.1, 100844.2, 98556.76, 96882.55, 
    96135.42, 98594.58, 101301, 101384.4, 101405, 101441.2, 101452.3, 101457.8,
  100613.2, 100655, 100791.6, 100827.3, 96401.31, 97786.22, 99411.25, 
    100944.6, 101207.4, 101331.9, 101409.2, 101441.2, 101468.1, 101482.9, 
    101486.2,
  100591.3, 100656.8, 100777, 100782.3, 96832.33, 97145.4, 96707.49, 101064, 
    101302.7, 101316.6, 101424.8, 101480.7, 101488, 101508.9, 101508.8,
  100975.6, 100907.3, 100784.3, 100740.2, 100629.6, 100590.7, 100653.4, 
    100671.9, 100739.2, 100821.8, 100900.7, 100969.5, 101021.1, 101054.3, 
    101068,
  100976.1, 100889.7, 100909.6, 100838.9, 100708.9, 100626.1, 100658.6, 
    100704.5, 100762, 100833.8, 100917.3, 100983.5, 101040, 101072.7, 101094.4,
  99328.59, 99034.12, 100882.9, 100893.5, 100861.2, 100799.5, 100705.6, 
    100734.9, 100806.3, 100856.9, 100938.5, 101005.3, 101063.7, 101095.5, 
    101119.6,
  97437.92, 97532.23, 100833.7, 100987.9, 100964.6, 100930.4, 100869.6, 
    100834.2, 100883.9, 100892.4, 100973.1, 101027.6, 101084.8, 101105.9, 
    101152.2,
  97443.62, 97847.73, 99613.02, 101028.7, 101014.8, 100980.9, 101039.2, 
    100952, 100967, 100945, 101006.9, 101057.4, 101102.9, 101149.3, 101180.5,
  96784.8, 98204.97, 100861.1, 101031.7, 101059, 100994.1, 101062.3, 101045, 
    101025.1, 101034.4, 101028, 101042.9, 101137.6, 101181.5, 101199.9,
  100859.7, 100886.9, 100952.6, 101042.7, 101063.1, 99347.3, 100824.8, 
    100945.3, 101011.8, 101058.6, 101074, 101127.1, 101164.6, 101211, 101223.8,
  100954.3, 100919.8, 100939.4, 101001.2, 100910.5, 98592.33, 96818.54, 
    96016.73, 98471.14, 101085.2, 101126.2, 101149.5, 101192, 101230.2, 
    101253.4,
  100892.3, 100899.3, 100944, 101000.2, 96455.77, 97859.16, 99479.12, 
    101025.1, 101156.2, 101164.6, 101185.9, 101177.9, 101225, 101250.6, 
    101272.5,
  100869.9, 100889.2, 100935, 100953.3, 96933.91, 97227.55, 96673.52, 101059, 
    101233.5, 101212, 101237.7, 101222.3, 101251.4, 101280.2, 101291.1,
  100574.8, 100494.4, 100455.6, 100396.6, 100327.5, 100247.1, 100226.6, 
    100245.8, 100279.6, 100334.4, 100421.4, 100486.4, 100548.5, 100598.4, 
    100645.6,
  100548.6, 100411.3, 100447.7, 100367.6, 100268, 100193.1, 100169.4, 
    100188.4, 100237.5, 100289.9, 100385.2, 100458.8, 100534.8, 100597.2, 
    100651.4,
  98836.66, 98549.6, 100369.6, 100373.9, 100251.1, 100100.3, 100052.1, 
    100089.9, 100164.5, 100240.8, 100351.3, 100448.4, 100534.2, 100591.2, 
    100651.5,
  97022.22, 97097.95, 100249.5, 100371.5, 100248.6, 100073.2, 99980.6, 
    100008.7, 100095.5, 100189, 100306.6, 100414.7, 100515.9, 100570.1, 
    100652.4,
  97052.13, 97416.59, 99070.48, 100367.7, 100248.9, 100027.6, 99897.02, 
    99900.02, 100014.5, 100129.4, 100264.4, 100390.9, 100491.4, 100575.5, 
    100657.2,
  96555.39, 97887.3, 100389.5, 100372.1, 100257.4, 100026.7, 99913.27, 
    99859.1, 99947.86, 100070.5, 100205, 100308.2, 100478.5, 100576.3, 
    100657.9,
  100716.6, 100640.4, 100517.3, 100430.1, 100284.6, 98465.51, 99666.64, 
    99704.84, 99859.2, 100011.8, 100180.4, 100328.6, 100472.4, 100577.4, 
    100659.6,
  100745.5, 100658.5, 100548.3, 100454.6, 100058.6, 97782.5, 95840.77, 
    94974.82, 97339.49, 100012.5, 100186.3, 100319.6, 100470.4, 100577.3, 
    100665.9,
  100744.8, 100661.6, 100577.9, 100472, 95679.59, 97048.18, 98511.09, 
    99862.91, 99937.91, 100071, 100201, 100331, 100470.6, 100582.4, 100675.7,
  100749.1, 100673.6, 100614.3, 100480.1, 96249.16, 96411.27, 95775.25, 
    100025.4, 100087.6, 100092.4, 100223.7, 100354.5, 100482, 100597, 100687.1,
  100800.6, 100754.1, 100744.5, 100738.5, 100744.2, 100749, 100753.2, 
    100735.9, 100716.1, 100689, 100660.8, 100655.7, 100635.8, 100576.9, 
    100560.1,
  100775.4, 100675.2, 100733.8, 100721.2, 100723.2, 100727.4, 100719.2, 
    100703.8, 100689.6, 100670.3, 100641.5, 100630.5, 100622.6, 100591.5, 
    100571.3,
  99057.16, 98759.33, 100606.9, 100703.5, 100707.3, 100698.1, 100670.8, 
    100653.8, 100632.4, 100619.1, 100599.2, 100593.9, 100587.8, 100583.5, 
    100557.9,
  97207.24, 97275.67, 100514.4, 100743.1, 100695.9, 100673.2, 100634.1, 
    100607.6, 100578.2, 100565, 100549.8, 100559.1, 100553.2, 100559.6, 
    100552.4,
  97184.3, 97588.48, 99287.06, 100696.6, 100656.3, 100596.1, 100556.2, 
    100517.1, 100488.7, 100487.3, 100479.8, 100502.5, 100504.7, 100544.7, 
    100541.6,
  96604.16, 97992.37, 100588.4, 100658.6, 100591.4, 100465, 100483.7, 100439, 
    100406.5, 100403.1, 100397.6, 100391.3, 100461.8, 100515.4, 100525.8,
  100801.5, 100736.4, 100662, 100598.7, 100530.7, 98729.34, 100045.2, 
    100108.7, 100208, 100262.8, 100313.2, 100357.7, 100403.5, 100471.5, 
    100505.1,
  100751.2, 100645.3, 100580.7, 100508.6, 100254.9, 97909.95, 96042.79, 
    95171.09, 97531.9, 100144.1, 100215.7, 100270, 100333.1, 100421.9, 
    100476.7,
  100661.6, 100570.6, 100518, 100451.9, 95721.12, 96995.08, 98524.08, 
    100011.6, 100173.5, 100171.7, 100176.2, 100209.8, 100273.3, 100370.5, 
    100445.2,
  100608, 100505.4, 100455.8, 100357.4, 96191.62, 96343.02, 95718.78, 
    99911.25, 100114.5, 100072.8, 100117.3, 100154.4, 100229.1, 100328.2, 
    100416.4,
  101155, 101117.2, 101107.7, 101108.4, 101139.9, 101145.8, 101131.7, 
    101103.4, 101066.1, 101020, 100953.6, 100978.1, 100926.7, 100801.2, 
    100768.9,
  101115.9, 101045.1, 101135.9, 101109, 101118.4, 101117.5, 101116, 101104.1, 
    101078.3, 101039.7, 100991.2, 100961.6, 101018.8, 100885.7, 100847,
  99383.3, 99111.59, 101049.5, 101160.2, 101136.2, 101132.3, 101108.9, 
    101084.8, 101061.1, 101026.9, 101000.6, 100954.3, 101034.9, 100903.7, 
    100885.1,
  97456.49, 97574.57, 100922.5, 101167.6, 101125.7, 101118.1, 101088.7, 
    101073.3, 101052.3, 101031.4, 101009.9, 100980, 101052.1, 100946.9, 
    100923.2,
  97495.16, 97959.48, 99700.61, 101148.3, 101111.4, 101062.9, 101040, 
    101012.8, 100998.1, 100986.6, 100995.7, 100968.3, 101015.6, 100994.7, 
    100949.4,
  96925.74, 98359.92, 101025.4, 101116.4, 101073.1, 100960.9, 101005.5, 
    100977.4, 100966, 100949.4, 100956.1, 100912, 101010, 101003.1, 100988.6,
  101164.2, 101167.4, 101145.3, 101097.5, 101052.9, 99242.3, 100607, 
    100675.9, 100802.2, 100867.5, 100916.3, 100924.2, 100982.2, 100984.5, 
    101007,
  101168.4, 101110.7, 101087.9, 101034.1, 100810.7, 98439.49, 96583.28, 
    95737.46, 98128.41, 100802.7, 100883, 100893.4, 100948.4, 100970.6, 
    101014.3,
  101102.8, 101061.2, 101054.1, 101007.9, 96251.85, 97593.65, 99151.52, 
    100662.5, 100813.1, 100841, 100860.2, 100859.3, 100904, 100953.1, 101007.1,
  101063.5, 101018.3, 101008.9, 100941.2, 96764.28, 96951.78, 96342.77, 
    100630.1, 100820.5, 100814.5, 100841, 100831.1, 100875.6, 100942.5, 
    100998.7 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.2466774, 0.6143242, 0.0668168, 0.2301621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.4924844, 0.2132108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.600569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1560082, 0,
  1, 1, 0.7132517, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02739768, 0,
  0.6230268, 0.6280472, 0.3043983, 0.08344039, 0, 0.3148882, 0.01188002, 0, 
    0, 0, 0, 0.08803581, 0, 0, 0,
  0, 0, 0, 0, 0.01144353, 0.8597386, 0.8205094, 0.5086318, 0.1258651, 
    0.08909279, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.291879, 0.6933324, 1, 0.9996726, 0.6666086, 0.08008575, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.611689, 0.7180831, 0.4623523, 0.2838529, 0.02767258, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0.002817577, 0.8915156, 0.5654301, 0.7485356, 0.3018697, 0, 0, 0, 
    0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0.04916316, 0.5638732, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3486554,
  2.316188, 6.745579, 0.5592819, 0.3199724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  147.4583, 171.3604, 6.513342, 0.3383408, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03840884, 0.4204801, 0,
  316.1323, 305.6766, 15.46485, 0.007546596, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1807817, 1.695307, 0,
  309.9182, 276.4409, 123.1236, 0.0108671, 0, 1.460928, 0.05467265, 0, 0, 0, 
    0.009753421, 0.03281464, 0.7768181, 0.4781904, 0,
  365.1592, 241.1036, 8.988194, 1.559117, 0.4356286, 6.775464, 0.2077458, 
    1.032432, 0.002793631, 0.1432027, 0.862155, 4.338077, 0.2366837, 0, 0,
  0, 0, 0, 0, 0.1289662, 151.094, 22.45284, 14.93281, 5.254983, 2.574013, 
    0.002986824, 0.1528066, 0.0002596498, 0, 0,
  0, 0, 0, 0, 13.93511, 217.993, 380.8379, 455.4515, 234.498, 2.407733, 0, 0, 
    0, 0, 0,
  0, 0.0003258124, 0, 0, 414.0298, 282.8423, 143.9435, 10.21257, 0.1187258, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 1.536109, 363.0271, 340.0019, 397.2344, 11.61882, 0, 0, 0, 0, 0, 
    0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
