netcdf \00010101.atmos_daily.tile5.pv350K {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pv350K(time, grid_yt, grid_xt) ;
		pv350K:_FillValue = -1.e+10f ;
		pv350K:missing_value = -1.e+10f ;
		pv350K:units = "(K m**2) / (kg s)" ;
		pv350K:long_name = "350-K potential vorticity; needs x350 scaling" ;
		pv350K:cell_methods = "time: mean" ;
		pv350K:time_avg_info = "average_T1,average_T2,average_DT" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:07 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile5.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile5.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pv350K =
  1.077065e-08, 1.114623e-08, 1.136199e-08, 1.162456e-08, 1.214554e-08, 
    1.225421e-08, 1.185387e-08, 1.204939e-08, 1.286765e-08, 1.455854e-08, 
    1.453603e-08, 1.360528e-08, 1.243845e-08, 1.153944e-08, 1.081346e-08,
  1.055041e-08, 1.099809e-08, 1.086566e-08, 1.080498e-08, 1.094127e-08, 
    1.100735e-08, 1.098444e-08, 1.109374e-08, 1.162859e-08, 1.182201e-08, 
    1.191837e-08, 1.21684e-08, 1.168439e-08, 1.0998e-08, 1.029028e-08,
  1.007313e-08, 1.038926e-08, 1.060879e-08, 1.060983e-08, 1.041678e-08, 
    1.018566e-08, 1.000124e-08, 9.84196e-09, 1.03594e-08, 1.078498e-08, 
    1.112211e-08, 1.093262e-08, 1.058033e-08, 1.007447e-08, 9.734066e-09,
  9.625282e-09, 9.934295e-09, 1.038893e-08, 1.0561e-08, 1.03295e-08, 
    9.815206e-09, 9.18982e-09, 9.322907e-09, 9.680473e-09, 1.01443e-08, 
    1.037776e-08, 1.045307e-08, 1.016155e-08, 9.75322e-09, 9.413911e-09,
  9.015888e-09, 9.082238e-09, 9.600978e-09, 1.012446e-08, 1.042128e-08, 
    9.926807e-09, 9.132613e-09, 9.041591e-09, 9.192716e-09, 9.501803e-09, 
    9.988168e-09, 9.970814e-09, 9.665446e-09, 9.291607e-09, 9.001242e-09,
  8.692938e-09, 9.062582e-09, 8.934681e-09, 8.946779e-09, 9.815182e-09, 
    9.930666e-09, 9.806392e-09, 9.376428e-09, 8.933441e-09, 8.964181e-09, 
    9.135223e-09, 9.237795e-09, 9.337667e-09, 9.056492e-09, 8.792031e-09,
  8.607887e-09, 8.576743e-09, 8.884525e-09, 9.099584e-09, 8.740129e-09, 
    9.079596e-09, 9.490757e-09, 9.633938e-09, 9.760279e-09, 9.023769e-09, 
    8.73175e-09, 8.529407e-09, 8.31785e-09, 8.563333e-09, 8.535355e-09,
  1.027698e-08, 8.844641e-09, 8.526656e-09, 8.760428e-09, 8.951129e-09, 
    9.024562e-09, 8.710558e-09, 9.008783e-09, 9.475812e-09, 9.554944e-09, 
    9.277049e-09, 8.403863e-09, 8.035793e-09, 7.827961e-09, 7.96329e-09,
  1.377155e-08, 1.141117e-08, 9.599258e-09, 8.747882e-09, 8.597522e-09, 
    8.782045e-09, 9.013406e-09, 8.885174e-09, 8.66129e-09, 9.064359e-09, 
    9.239213e-09, 8.946264e-09, 8.130666e-09, 7.578271e-09, 7.337832e-09,
  1.718522e-08, 1.56732e-08, 1.307816e-08, 1.065425e-08, 9.140617e-09, 
    8.623088e-09, 8.583498e-09, 8.826181e-09, 8.944205e-09, 8.85406e-09, 
    8.841702e-09, 8.836732e-09, 8.621551e-09, 8.005579e-09, 7.325271e-09,
  1.22358e-08, 1.232517e-08, 1.287451e-08, 1.301622e-08, 1.489208e-08, 
    1.885528e-08, 2.307798e-08, 2.562338e-08, 2.826058e-08, 2.861358e-08, 
    2.86514e-08, 2.62968e-08, 2.512976e-08, 2.436967e-08, 2.391433e-08,
  1.124958e-08, 1.181817e-08, 1.215875e-08, 1.21346e-08, 1.232693e-08, 
    1.437828e-08, 1.889441e-08, 2.287401e-08, 2.428556e-08, 2.704217e-08, 
    2.828111e-08, 2.75279e-08, 2.587243e-08, 2.444884e-08, 2.319005e-08,
  1.076454e-08, 1.158715e-08, 1.209425e-08, 1.233176e-08, 1.224045e-08, 
    1.248808e-08, 1.471297e-08, 1.868534e-08, 2.209345e-08, 2.416165e-08, 
    2.672111e-08, 2.755645e-08, 2.658359e-08, 2.520484e-08, 2.394197e-08,
  1.048201e-08, 1.055626e-08, 1.090695e-08, 1.139569e-08, 1.190007e-08, 
    1.197113e-08, 1.322305e-08, 1.46242e-08, 1.689887e-08, 2.006261e-08, 
    2.329652e-08, 2.5031e-08, 2.524672e-08, 2.470151e-08, 2.333034e-08,
  1.108692e-08, 1.063539e-08, 1.070005e-08, 1.125021e-08, 1.154781e-08, 
    1.203606e-08, 1.222082e-08, 1.356421e-08, 1.469606e-08, 1.66817e-08, 
    1.984277e-08, 2.22352e-08, 2.282699e-08, 2.311288e-08, 2.265939e-08,
  1.25835e-08, 1.172565e-08, 1.125334e-08, 1.084565e-08, 1.092526e-08, 
    1.131362e-08, 1.125441e-08, 1.135814e-08, 1.263628e-08, 1.366946e-08, 
    1.580948e-08, 1.795284e-08, 1.95951e-08, 2.183374e-08, 2.220383e-08,
  1.445256e-08, 1.337211e-08, 1.227646e-08, 1.155741e-08, 1.090811e-08, 
    1.073474e-08, 1.105528e-08, 1.024445e-08, 1.029556e-08, 1.126342e-08, 
    1.223803e-08, 1.40665e-08, 1.655157e-08, 1.977522e-08, 2.086765e-08,
  1.625058e-08, 1.535762e-08, 1.422371e-08, 1.276109e-08, 1.179469e-08, 
    1.076011e-08, 1.061831e-08, 1.054584e-08, 9.741319e-09, 9.635023e-09, 
    1.013481e-08, 1.140745e-08, 1.235798e-08, 1.472914e-08, 1.76815e-08,
  1.628493e-08, 1.657098e-08, 1.602279e-08, 1.489487e-08, 1.321224e-08, 
    1.181081e-08, 1.058241e-08, 1.058408e-08, 1.032081e-08, 9.149045e-09, 
    9.250105e-09, 1.007203e-08, 1.140096e-08, 1.145486e-08, 1.266125e-08,
  1.611819e-08, 1.654671e-08, 1.687382e-08, 1.661459e-08, 1.550021e-08, 
    1.379785e-08, 1.179013e-08, 1.049488e-08, 1.04111e-08, 1.007109e-08, 
    8.901529e-09, 9.246845e-09, 1.006812e-08, 1.111573e-08, 1.14682e-08,
  1.352782e-08, 1.334315e-08, 1.370189e-08, 1.567782e-08, 1.588992e-08, 
    1.488912e-08, 1.558284e-08, 1.708639e-08, 1.800803e-08, 1.70973e-08, 
    1.507638e-08, 1.321676e-08, 1.164891e-08, 9.961733e-09, 8.470929e-09,
  1.298248e-08, 1.343857e-08, 1.47643e-08, 1.637992e-08, 1.515253e-08, 
    1.479068e-08, 1.652923e-08, 1.91507e-08, 1.960353e-08, 1.968791e-08, 
    1.784666e-08, 1.552909e-08, 1.358058e-08, 1.200097e-08, 1.040285e-08,
  1.311804e-08, 1.404468e-08, 1.46217e-08, 1.564775e-08, 1.709895e-08, 
    1.768686e-08, 1.816137e-08, 1.902974e-08, 2.148065e-08, 2.193346e-08, 
    2.097252e-08, 1.840117e-08, 1.574538e-08, 1.377184e-08, 1.219944e-08,
  1.40997e-08, 1.446328e-08, 1.551564e-08, 1.729212e-08, 1.658102e-08, 
    1.791285e-08, 1.920183e-08, 1.846651e-08, 2.065461e-08, 2.327249e-08, 
    2.36221e-08, 2.16784e-08, 1.885603e-08, 1.639675e-08, 1.429774e-08,
  1.433672e-08, 1.494251e-08, 1.545641e-08, 1.610284e-08, 1.604031e-08, 
    1.713246e-08, 1.971417e-08, 1.856697e-08, 1.900782e-08, 2.282526e-08, 
    2.451094e-08, 2.301167e-08, 2.061392e-08, 1.743662e-08, 1.543073e-08,
  1.48507e-08, 1.521428e-08, 1.564894e-08, 1.611735e-08, 1.599342e-08, 
    1.662535e-08, 1.94128e-08, 1.746705e-08, 1.755835e-08, 2.085645e-08, 
    2.397661e-08, 2.388156e-08, 2.221724e-08, 1.945103e-08, 1.691224e-08,
  1.463265e-08, 1.531549e-08, 1.570856e-08, 1.610844e-08, 1.613184e-08, 
    1.629235e-08, 1.860643e-08, 1.875794e-08, 1.639066e-08, 1.804308e-08, 
    2.198572e-08, 2.45911e-08, 2.486594e-08, 2.234752e-08, 1.795944e-08,
  1.399309e-08, 1.45909e-08, 1.55093e-08, 1.585392e-08, 1.638273e-08, 
    1.640857e-08, 1.820976e-08, 1.834015e-08, 1.562199e-08, 1.485313e-08, 
    1.715408e-08, 2.237953e-08, 2.558812e-08, 2.460127e-08, 2.011265e-08,
  1.367932e-08, 1.402589e-08, 1.479333e-08, 1.527094e-08, 1.61008e-08, 
    1.658463e-08, 1.795855e-08, 1.798395e-08, 1.525895e-08, 1.355645e-08, 
    1.488084e-08, 1.891005e-08, 2.310697e-08, 2.4621e-08, 2.236025e-08,
  1.345182e-08, 1.368666e-08, 1.442875e-08, 1.480135e-08, 1.567514e-08, 
    1.630898e-08, 1.766951e-08, 1.832674e-08, 1.557957e-08, 1.324147e-08, 
    1.331729e-08, 1.578585e-08, 2.124961e-08, 2.209834e-08, 2.225188e-08,
  1.107435e-08, 1.080493e-08, 1.046846e-08, 9.530004e-09, 8.885659e-09, 
    8.412453e-09, 8.13902e-09, 7.689329e-09, 7.394605e-09, 6.748282e-09, 
    5.933173e-09, 5.403697e-09, 5.010456e-09, 4.447189e-09, 3.792338e-09,
  1.185251e-08, 1.151527e-08, 1.156564e-08, 1.099651e-08, 1.015252e-08, 
    9.253841e-09, 8.608432e-09, 8.07552e-09, 7.678793e-09, 7.138776e-09, 
    6.401156e-09, 5.665793e-09, 5.173455e-09, 4.693445e-09, 4.081342e-09,
  1.233136e-08, 1.21885e-08, 1.19851e-08, 1.176531e-08, 1.135064e-08, 
    1.043411e-08, 9.411158e-09, 8.616533e-09, 8.130144e-09, 7.6275e-09, 
    6.854236e-09, 6.092287e-09, 5.423015e-09, 5.021864e-09, 4.473051e-09,
  1.256854e-08, 1.283666e-08, 1.296432e-08, 1.331173e-08, 1.265694e-08, 
    1.19299e-08, 1.082812e-08, 9.410286e-09, 8.749804e-09, 8.259211e-09, 
    7.591701e-09, 6.750985e-09, 6.043246e-09, 5.447348e-09, 4.937871e-09,
  1.313893e-08, 1.324726e-08, 1.36287e-08, 1.376695e-08, 1.411344e-08, 
    1.330507e-08, 1.269607e-08, 1.135805e-08, 9.864255e-09, 9.072469e-09, 
    8.374043e-09, 7.645927e-09, 6.937783e-09, 6.223378e-09, 5.55695e-09,
  1.308403e-08, 1.341356e-08, 1.378524e-08, 1.431032e-08, 1.471822e-08, 
    1.480483e-08, 1.420738e-08, 1.303505e-08, 1.142377e-08, 1.025772e-08, 
    9.288855e-09, 8.487902e-09, 7.816602e-09, 7.031226e-09, 6.26726e-09,
  1.269766e-08, 1.32797e-08, 1.399496e-08, 1.505292e-08, 1.5245e-08, 
    1.525016e-08, 1.562148e-08, 1.487353e-08, 1.330919e-08, 1.172169e-08, 
    1.03147e-08, 9.219556e-09, 8.601817e-09, 7.864236e-09, 6.993671e-09,
  1.237967e-08, 1.277724e-08, 1.371152e-08, 1.517595e-08, 1.503853e-08, 
    1.526798e-08, 1.66357e-08, 1.649899e-08, 1.516582e-08, 1.324303e-08, 
    1.148682e-08, 1.012959e-08, 9.208645e-09, 8.631718e-09, 7.90585e-09,
  1.2167e-08, 1.238959e-08, 1.339609e-08, 1.465125e-08, 1.49521e-08, 
    1.522571e-08, 1.735006e-08, 1.739522e-08, 1.679112e-08, 1.491035e-08, 
    1.289976e-08, 1.10845e-08, 9.848542e-09, 9.07039e-09, 8.463767e-09,
  1.192979e-08, 1.203842e-08, 1.280875e-08, 1.418001e-08, 1.467799e-08, 
    1.506893e-08, 1.712682e-08, 1.801457e-08, 1.758125e-08, 1.610244e-08, 
    1.432862e-08, 1.236622e-08, 1.06181e-08, 9.780125e-09, 9.099809e-09,
  1.524232e-08, 1.5427e-08, 1.59667e-08, 1.654355e-08, 1.565059e-08, 
    1.455039e-08, 1.3199e-08, 1.23618e-08, 1.174528e-08, 1.10267e-08, 
    1.016752e-08, 9.572625e-09, 8.824729e-09, 8.069773e-09, 7.475284e-09,
  1.482629e-08, 1.447651e-08, 1.493422e-08, 1.537489e-08, 1.514301e-08, 
    1.409772e-08, 1.309166e-08, 1.214225e-08, 1.145006e-08, 1.087383e-08, 
    1.019548e-08, 9.654388e-09, 8.9712e-09, 8.247055e-09, 7.692069e-09,
  1.438531e-08, 1.341104e-08, 1.394128e-08, 1.419982e-08, 1.406023e-08, 
    1.353197e-08, 1.26382e-08, 1.177619e-08, 1.116883e-08, 1.066065e-08, 
    1.006289e-08, 9.622011e-09, 8.986939e-09, 8.426908e-09, 7.700329e-09,
  1.383671e-08, 1.288739e-08, 1.320062e-08, 1.329351e-08, 1.312116e-08, 
    1.26688e-08, 1.221952e-08, 1.153702e-08, 1.079217e-08, 1.022594e-08, 
    9.639565e-09, 9.226269e-09, 8.753307e-09, 8.127989e-09, 7.567235e-09,
  1.327181e-08, 1.256681e-08, 1.277741e-08, 1.257095e-08, 1.236667e-08, 
    1.194641e-08, 1.161765e-08, 1.105145e-08, 1.051593e-08, 9.981955e-09, 
    9.340033e-09, 8.876393e-09, 8.405998e-09, 8.060765e-09, 7.640171e-09,
  1.288831e-08, 1.243837e-08, 1.241859e-08, 1.210871e-08, 1.172046e-08, 
    1.124767e-08, 1.098956e-08, 1.071143e-08, 1.023974e-08, 9.755557e-09, 
    9.115747e-09, 8.628145e-09, 8.202102e-09, 7.90217e-09, 7.356145e-09,
  1.285662e-08, 1.275248e-08, 1.234559e-08, 1.190386e-08, 1.126505e-08, 
    1.086941e-08, 1.054759e-08, 1.033699e-08, 1.003888e-08, 9.539425e-09, 
    8.883629e-09, 8.373839e-09, 7.843615e-09, 7.402595e-09, 6.837134e-09,
  1.279764e-08, 1.285716e-08, 1.281e-08, 1.209817e-08, 1.112639e-08, 
    1.065852e-08, 1.035582e-08, 1.005599e-08, 9.710226e-09, 9.313162e-09, 
    8.644308e-09, 8.044077e-09, 7.509856e-09, 6.967969e-09, 6.36661e-09,
  1.287398e-08, 1.27663e-08, 1.301187e-08, 1.265657e-08, 1.138949e-08, 
    1.071943e-08, 1.03189e-08, 1.008309e-08, 9.413981e-09, 8.909104e-09, 
    8.4653e-09, 7.946498e-09, 7.352726e-09, 6.784542e-09, 6.10428e-09,
  1.328112e-08, 1.308289e-08, 1.297685e-08, 1.296527e-08, 1.192858e-08, 
    1.117603e-08, 1.044568e-08, 1.016553e-08, 9.594288e-09, 8.81696e-09, 
    8.273314e-09, 7.775353e-09, 7.345544e-09, 6.787296e-09, 6.109852e-09,
  1.239105e-08, 1.117215e-08, 1.007119e-08, 8.749908e-09, 7.596477e-09, 
    6.815514e-09, 6.293052e-09, 5.877877e-09, 5.320964e-09, 4.765899e-09, 
    4.205917e-09, 3.5794e-09, 3.008924e-09, 2.481943e-09, 1.981488e-09,
  1.318189e-08, 1.231367e-08, 1.1303e-08, 1.010799e-08, 8.811598e-09, 
    7.735255e-09, 6.99321e-09, 6.365782e-09, 5.685147e-09, 5.131899e-09, 
    4.578272e-09, 3.975144e-09, 3.367214e-09, 2.847154e-09, 2.344258e-09,
  1.3723e-08, 1.324492e-08, 1.248616e-08, 1.131398e-08, 1.023357e-08, 
    8.839655e-09, 7.809071e-09, 7.026293e-09, 6.269936e-09, 5.56895e-09, 
    5.011055e-09, 4.421359e-09, 3.790738e-09, 3.209349e-09, 2.7106e-09,
  1.402727e-08, 1.40121e-08, 1.349246e-08, 1.271445e-08, 1.151786e-08, 
    1.030809e-08, 8.857294e-09, 7.791155e-09, 6.97675e-09, 6.124604e-09, 
    5.528793e-09, 4.934417e-09, 4.284338e-09, 3.665266e-09, 3.129809e-09,
  1.386513e-08, 1.425415e-08, 1.417403e-08, 1.370486e-08, 1.278965e-08, 
    1.142428e-08, 1.016923e-08, 8.812499e-09, 7.772121e-09, 6.826486e-09, 
    6.152296e-09, 5.522543e-09, 4.833733e-09, 4.18929e-09, 3.637344e-09,
  1.37849e-08, 1.431468e-08, 1.480132e-08, 1.446045e-08, 1.394342e-08, 
    1.259164e-08, 1.119338e-08, 9.957459e-09, 8.623014e-09, 7.742382e-09, 
    6.922218e-09, 6.181825e-09, 5.500503e-09, 4.809992e-09, 4.216972e-09,
  1.359433e-08, 1.390639e-08, 1.486559e-08, 1.500837e-08, 1.463459e-08, 
    1.374553e-08, 1.211372e-08, 1.085469e-08, 9.334439e-09, 8.551907e-09, 
    7.709652e-09, 6.914884e-09, 6.205989e-09, 5.535113e-09, 4.85827e-09,
  1.366552e-08, 1.360614e-08, 1.448337e-08, 1.538239e-08, 1.510022e-08, 
    1.474463e-08, 1.298894e-08, 1.176515e-08, 1.002872e-08, 9.240989e-09, 
    8.506455e-09, 7.680897e-09, 6.964476e-09, 6.280884e-09, 5.570064e-09,
  1.357181e-08, 1.350782e-08, 1.400907e-08, 1.537275e-08, 1.543437e-08, 
    1.551266e-08, 1.397287e-08, 1.264071e-08, 1.08975e-08, 9.868805e-09, 
    9.187028e-09, 8.387802e-09, 7.683094e-09, 6.967969e-09, 6.269589e-09,
  1.366662e-08, 1.33463e-08, 1.382598e-08, 1.5041e-08, 1.564065e-08, 
    1.602394e-08, 1.484637e-08, 1.353764e-08, 1.184103e-08, 1.045637e-08, 
    9.786421e-09, 9.001595e-09, 8.26661e-09, 7.577143e-09, 6.855275e-09,
  1.093067e-08, 9.878891e-09, 9.027786e-09, 8.059205e-09, 7.168938e-09, 
    6.304557e-09, 5.704877e-09, 5.101345e-09, 4.472861e-09, 3.857426e-09, 
    3.418264e-09, 3.302334e-09, 3.186788e-09, 2.899185e-09, 2.347676e-09,
  1.060835e-08, 9.579818e-09, 8.810093e-09, 7.868606e-09, 7.048538e-09, 
    6.251231e-09, 5.593997e-09, 5.042173e-09, 4.490719e-09, 3.957892e-09, 
    3.409861e-09, 3.174579e-09, 3.201602e-09, 3.083201e-09, 2.625591e-09,
  1.044388e-08, 9.284312e-09, 8.527085e-09, 7.68633e-09, 6.933298e-09, 
    6.212554e-09, 5.574596e-09, 4.973363e-09, 4.489578e-09, 4.059881e-09, 
    3.483799e-09, 3.148732e-09, 3.223571e-09, 3.218884e-09, 2.89375e-09,
  1.024015e-08, 9.018126e-09, 8.285546e-09, 7.437328e-09, 6.837384e-09, 
    6.143225e-09, 5.540881e-09, 4.94806e-09, 4.49992e-09, 4.156886e-09, 
    3.643885e-09, 3.234585e-09, 3.212676e-09, 3.23871e-09, 3.056529e-09,
  1.004212e-08, 8.984729e-09, 8.108975e-09, 7.19664e-09, 6.654925e-09, 
    6.064945e-09, 5.519767e-09, 4.943754e-09, 4.55263e-09, 4.215056e-09, 
    3.796978e-09, 3.395327e-09, 3.219698e-09, 3.178152e-09, 3.102083e-09,
  9.879821e-09, 8.964494e-09, 8.094781e-09, 7.194589e-09, 6.512472e-09, 
    5.974229e-09, 5.518077e-09, 4.961447e-09, 4.585081e-09, 4.258919e-09, 
    3.908731e-09, 3.545485e-09, 3.259895e-09, 3.142267e-09, 3.072762e-09,
  9.701555e-09, 8.922473e-09, 8.162417e-09, 7.325882e-09, 6.581426e-09, 
    5.900715e-09, 5.472062e-09, 4.982843e-09, 4.606205e-09, 4.262638e-09, 
    3.969973e-09, 3.681924e-09, 3.331477e-09, 3.166613e-09, 3.087138e-09,
  9.506182e-09, 8.916118e-09, 8.176642e-09, 7.396288e-09, 6.682265e-09, 
    5.998984e-09, 5.45681e-09, 5.006544e-09, 4.655657e-09, 4.291282e-09, 
    3.992781e-09, 3.777559e-09, 3.461549e-09, 3.274768e-09, 3.131626e-09,
  9.514698e-09, 8.809589e-09, 8.148271e-09, 7.380534e-09, 6.702809e-09, 
    6.208054e-09, 5.52951e-09, 5.085671e-09, 4.747177e-09, 4.371295e-09, 
    4.065028e-09, 3.90212e-09, 3.593087e-09, 3.416857e-09, 3.23437e-09,
  9.739518e-09, 8.89244e-09, 8.088186e-09, 7.362507e-09, 6.666904e-09, 
    6.339262e-09, 5.675308e-09, 5.228239e-09, 4.922065e-09, 4.512596e-09, 
    4.129665e-09, 3.959087e-09, 3.735174e-09, 3.537783e-09, 3.361479e-09,
  1.198233e-08, 1.040903e-08, 9.091969e-09, 7.682718e-09, 6.593491e-09, 
    5.672553e-09, 4.702269e-09, 3.815905e-09, 3.129168e-09, 2.716614e-09, 
    2.219892e-09, 1.63216e-09, 1.360945e-09, 1.274909e-09, 1.165737e-09,
  1.191335e-08, 1.036638e-08, 9.13518e-09, 7.76305e-09, 6.681328e-09, 
    5.747121e-09, 4.777015e-09, 3.861277e-09, 3.189508e-09, 2.861385e-09, 
    2.454268e-09, 1.860319e-09, 1.502435e-09, 1.395193e-09, 1.282842e-09,
  1.196536e-08, 1.044022e-08, 9.197449e-09, 7.782933e-09, 6.771016e-09, 
    5.861675e-09, 4.87378e-09, 3.970699e-09, 3.286224e-09, 2.941392e-09, 
    2.677682e-09, 2.173307e-09, 1.669527e-09, 1.520442e-09, 1.38707e-09,
  1.210222e-08, 1.058602e-08, 9.281128e-09, 7.845409e-09, 6.834167e-09, 
    5.981677e-09, 5.034229e-09, 4.17082e-09, 3.422602e-09, 2.950556e-09, 
    2.737024e-09, 2.432374e-09, 1.916713e-09, 1.664668e-09, 1.515312e-09,
  1.224299e-08, 1.081826e-08, 9.431446e-09, 7.895191e-09, 6.888679e-09, 
    6.078084e-09, 5.202762e-09, 4.402208e-09, 3.626355e-09, 3.00439e-09, 
    2.714841e-09, 2.54512e-09, 2.148047e-09, 1.831965e-09, 1.608506e-09,
  1.241311e-08, 1.112811e-08, 9.602113e-09, 7.964066e-09, 6.886912e-09, 
    6.148929e-09, 5.34747e-09, 4.633434e-09, 3.876588e-09, 3.120999e-09, 
    2.713533e-09, 2.623592e-09, 2.367449e-09, 2.00478e-09, 1.737031e-09,
  1.263737e-08, 1.143821e-08, 9.801685e-09, 8.044987e-09, 6.891185e-09, 
    6.203215e-09, 5.473458e-09, 4.805003e-09, 4.129302e-09, 3.314654e-09, 
    2.819502e-09, 2.661283e-09, 2.486772e-09, 2.183905e-09, 1.892521e-09,
  1.29006e-08, 1.171525e-08, 1.001033e-08, 8.171728e-09, 6.919446e-09, 
    6.262336e-09, 5.565902e-09, 4.923673e-09, 4.344198e-09, 3.563888e-09, 
    2.991642e-09, 2.725899e-09, 2.580717e-09, 2.336427e-09, 2.084403e-09,
  1.308934e-08, 1.195577e-08, 1.02448e-08, 8.348072e-09, 7.024955e-09, 
    6.319485e-09, 5.640469e-09, 4.979978e-09, 4.456315e-09, 3.834979e-09, 
    3.214873e-09, 2.795071e-09, 2.667215e-09, 2.438652e-09, 2.243871e-09,
  1.325208e-08, 1.208871e-08, 1.04533e-08, 8.610917e-09, 7.189153e-09, 
    6.381454e-09, 5.683203e-09, 5.000476e-09, 4.486636e-09, 4.022076e-09, 
    3.442528e-09, 2.958724e-09, 2.742749e-09, 2.511784e-09, 2.339067e-09,
  1.770753e-08, 1.616102e-08, 1.398192e-08, 1.201903e-08, 1.053569e-08, 
    9.206845e-09, 8.160315e-09, 7.291053e-09, 6.568573e-09, 6.077579e-09, 
    5.320093e-09, 4.585261e-09, 4.013059e-09, 3.48139e-09, 2.996136e-09,
  1.778617e-08, 1.642738e-08, 1.430262e-08, 1.227315e-08, 1.063141e-08, 
    9.317207e-09, 8.204781e-09, 7.331582e-09, 6.498652e-09, 6.102072e-09, 
    5.548679e-09, 4.741767e-09, 4.10014e-09, 3.533872e-09, 3.051351e-09,
  1.789376e-08, 1.678642e-08, 1.470056e-08, 1.254658e-08, 1.075027e-08, 
    9.367217e-09, 8.241545e-09, 7.34994e-09, 6.475623e-09, 5.965241e-09, 
    5.650503e-09, 4.957792e-09, 4.223454e-09, 3.643161e-09, 3.140574e-09,
  1.796678e-08, 1.690946e-08, 1.515529e-08, 1.28671e-08, 1.092845e-08, 
    9.417282e-09, 8.300268e-09, 7.388043e-09, 6.48108e-09, 5.869334e-09, 
    5.616965e-09, 5.155419e-09, 4.42383e-09, 3.780291e-09, 3.26046e-09,
  1.805184e-08, 1.702808e-08, 1.558725e-08, 1.330428e-08, 1.116755e-08, 
    9.465057e-09, 8.374746e-09, 7.43551e-09, 6.497984e-09, 5.793922e-09, 
    5.486607e-09, 5.223127e-09, 4.57714e-09, 3.912336e-09, 3.384989e-09,
  1.815611e-08, 1.723613e-08, 1.597259e-08, 1.384182e-08, 1.153179e-08, 
    9.581846e-09, 8.471605e-09, 7.504733e-09, 6.489529e-09, 5.73356e-09, 
    5.363265e-09, 5.140382e-09, 4.65486e-09, 4.014016e-09, 3.482505e-09,
  1.851349e-08, 1.732533e-08, 1.628179e-08, 1.44274e-08, 1.195067e-08, 
    9.812603e-09, 8.668023e-09, 7.564682e-09, 6.511487e-09, 5.709788e-09, 
    5.216948e-09, 4.975286e-09, 4.61482e-09, 4.066817e-09, 3.558329e-09,
  1.885588e-08, 1.734269e-08, 1.661006e-08, 1.515392e-08, 1.239671e-08, 
    1.022261e-08, 8.904403e-09, 7.672293e-09, 6.514697e-09, 5.712157e-09, 
    5.144717e-09, 4.821908e-09, 4.527196e-09, 4.05846e-09, 3.596057e-09,
  1.903195e-08, 1.728784e-08, 1.663678e-08, 1.581258e-08, 1.285808e-08, 
    1.063893e-08, 9.148409e-09, 7.856668e-09, 6.575897e-09, 5.72235e-09, 
    5.088129e-09, 4.680695e-09, 4.412595e-09, 4.020297e-09, 3.610061e-09,
  1.918069e-08, 1.729024e-08, 1.722564e-08, 1.638914e-08, 1.348697e-08, 
    1.103752e-08, 9.422843e-09, 8.08868e-09, 6.683984e-09, 5.754153e-09, 
    5.13195e-09, 4.599058e-09, 4.307807e-09, 3.960274e-09, 3.584977e-09,
  1.420207e-08, 1.236706e-08, 1.068955e-08, 9.402856e-09, 8.354625e-09, 
    7.39113e-09, 6.666289e-09, 5.808473e-09, 4.670903e-09, 3.725084e-09, 
    3.261599e-09, 2.757462e-09, 2.308219e-09, 1.815015e-09, 1.402614e-09,
  1.53825e-08, 1.356756e-08, 1.15283e-08, 1.004383e-08, 8.936435e-09, 
    8.023302e-09, 7.244057e-09, 6.419104e-09, 5.393348e-09, 4.276931e-09, 
    3.533962e-09, 3.047179e-09, 2.667483e-09, 2.242767e-09, 1.767661e-09,
  1.666075e-08, 1.493854e-08, 1.256407e-08, 1.077196e-08, 9.498745e-09, 
    8.568034e-09, 7.846556e-09, 7.042081e-09, 6.046496e-09, 4.99024e-09, 
    3.987453e-09, 3.356789e-09, 2.935695e-09, 2.623308e-09, 2.182455e-09,
  1.774873e-08, 1.615571e-08, 1.373641e-08, 1.166838e-08, 1.007524e-08, 
    9.089596e-09, 8.410404e-09, 7.636177e-09, 6.660646e-09, 5.713852e-09, 
    4.680099e-09, 3.812873e-09, 3.181643e-09, 2.925521e-09, 2.624795e-09,
  1.862214e-08, 1.723219e-08, 1.501465e-08, 1.270701e-08, 1.081934e-08, 
    9.55741e-09, 8.883012e-09, 8.147725e-09, 7.216671e-09, 6.33405e-09, 
    5.474877e-09, 4.435739e-09, 3.593737e-09, 3.123348e-09, 2.912299e-09,
  1.944695e-08, 1.807262e-08, 1.631117e-08, 1.382381e-08, 1.174087e-08, 
    1.00743e-08, 9.286637e-09, 8.633974e-09, 7.728775e-09, 6.880126e-09, 
    6.168421e-09, 5.204383e-09, 4.200195e-09, 3.456946e-09, 3.127164e-09,
  2.019187e-08, 1.889785e-08, 1.738626e-08, 1.495401e-08, 1.272954e-08, 
    1.074049e-08, 9.63924e-09, 9.099126e-09, 8.232513e-09, 7.337849e-09, 
    6.727724e-09, 5.903961e-09, 4.92974e-09, 3.968147e-09, 3.448158e-09,
  2.082718e-08, 1.970277e-08, 1.829017e-08, 1.60623e-08, 1.371727e-08, 
    1.145146e-08, 1.00377e-08, 9.523153e-09, 8.729753e-09, 7.792257e-09, 
    7.167373e-09, 6.511121e-09, 5.64078e-09, 4.62206e-09, 3.876981e-09,
  2.138735e-08, 2.039245e-08, 1.905705e-08, 1.706991e-08, 1.465638e-08, 
    1.225785e-08, 1.047735e-08, 9.904054e-09, 9.254993e-09, 8.232894e-09, 
    7.492284e-09, 6.995226e-09, 6.217223e-09, 5.32089e-09, 4.421048e-09,
  2.178742e-08, 2.096614e-08, 1.973123e-08, 1.790855e-08, 1.5558e-08, 
    1.308482e-08, 1.105054e-08, 1.024666e-08, 9.724415e-09, 8.705982e-09, 
    7.850947e-09, 7.382257e-09, 6.724017e-09, 5.925372e-09, 5.015957e-09,
  1.552531e-08, 1.45223e-08, 1.389522e-08, 1.266564e-08, 1.125843e-08, 
    9.604863e-09, 7.833083e-09, 6.172534e-09, 4.939549e-09, 4.085994e-09, 
    3.418248e-09, 2.862939e-09, 2.502046e-09, 2.35945e-09, 2.192188e-09,
  1.564379e-08, 1.465863e-08, 1.40987e-08, 1.304027e-08, 1.174367e-08, 
    1.026196e-08, 8.46465e-09, 6.852869e-09, 5.395212e-09, 4.472712e-09, 
    3.728911e-09, 3.158712e-09, 2.663751e-09, 2.423427e-09, 2.256512e-09,
  1.574636e-08, 1.480882e-08, 1.425053e-08, 1.335257e-08, 1.218572e-08, 
    1.079774e-08, 9.099652e-09, 7.466229e-09, 5.941678e-09, 4.838181e-09, 
    4.019183e-09, 3.425207e-09, 2.901297e-09, 2.525481e-09, 2.320793e-09,
  1.587909e-08, 1.493789e-08, 1.434584e-08, 1.360428e-08, 1.254003e-08, 
    1.123741e-08, 9.633993e-09, 8.000008e-09, 6.503054e-09, 5.205326e-09, 
    4.317834e-09, 3.678255e-09, 3.144177e-09, 2.688374e-09, 2.391318e-09,
  1.59479e-08, 1.507991e-08, 1.441223e-08, 1.377125e-08, 1.279696e-08, 
    1.157569e-08, 1.008442e-08, 8.468148e-09, 7.014701e-09, 5.639475e-09, 
    4.622792e-09, 3.919548e-09, 3.350165e-09, 2.881312e-09, 2.460786e-09,
  1.605037e-08, 1.517867e-08, 1.445311e-08, 1.386908e-08, 1.294617e-08, 
    1.177286e-08, 1.044329e-08, 8.882453e-09, 7.498965e-09, 6.1328e-09, 
    4.933064e-09, 4.159507e-09, 3.528018e-09, 3.060124e-09, 2.592224e-09,
  1.608859e-08, 1.52614e-08, 1.446006e-08, 1.390582e-08, 1.304949e-08, 
    1.189305e-08, 1.072238e-08, 9.273991e-09, 7.917368e-09, 6.608586e-09, 
    5.25778e-09, 4.386049e-09, 3.699412e-09, 3.21095e-09, 2.75878e-09,
  1.612618e-08, 1.530253e-08, 1.447299e-08, 1.392326e-08, 1.31547e-08, 
    1.194143e-08, 1.093583e-08, 9.637501e-09, 8.273302e-09, 7.021271e-09, 
    5.64369e-09, 4.612125e-09, 3.883402e-09, 3.349831e-09, 2.897816e-09,
  1.615632e-08, 1.534385e-08, 1.45541e-08, 1.397822e-08, 1.322018e-08, 
    1.242731e-08, 1.106799e-08, 9.921739e-09, 8.569357e-09, 7.371511e-09, 
    6.037854e-09, 4.852478e-09, 4.06705e-09, 3.485858e-09, 3.017438e-09,
  1.623688e-08, 1.540778e-08, 1.468064e-08, 1.406035e-08, 1.317518e-08, 
    1.248315e-08, 1.124124e-08, 1.018972e-08, 8.823238e-09, 7.646167e-09, 
    6.408564e-09, 5.154037e-09, 4.262813e-09, 3.624484e-09, 3.10671e-09,
  1.838086e-08, 1.736816e-08, 1.656864e-08, 1.544949e-08, 1.370137e-08, 
    1.231216e-08, 1.163287e-08, 1.010134e-08, 7.105599e-09, 5.9479e-09, 
    5.062774e-09, 4.188042e-09, 3.449453e-09, 2.933214e-09, 2.472212e-09,
  1.861142e-08, 1.797519e-08, 1.693385e-08, 1.616606e-08, 1.46838e-08, 
    1.292331e-08, 1.181366e-08, 1.062085e-08, 8.002202e-09, 6.126918e-09, 
    5.358251e-09, 4.717384e-09, 3.899774e-09, 3.167455e-09, 2.548282e-09,
  1.887284e-08, 1.843473e-08, 1.725432e-08, 1.645108e-08, 1.537635e-08, 
    1.366221e-08, 1.212949e-08, 1.094578e-08, 8.867183e-09, 6.541681e-09, 
    5.490842e-09, 5.028832e-09, 4.343821e-09, 3.532836e-09, 2.763026e-09,
  1.900703e-08, 1.858386e-08, 1.761475e-08, 1.664757e-08, 1.584828e-08, 
    1.435912e-08, 1.26983e-08, 1.138763e-08, 9.546336e-09, 7.151406e-09, 
    5.66938e-09, 5.098617e-09, 4.673379e-09, 3.938989e-09, 3.106032e-09,
  1.911708e-08, 1.860481e-08, 1.785681e-08, 1.691984e-08, 1.615454e-08, 
    1.491599e-08, 1.337906e-08, 1.187335e-08, 1.011485e-08, 7.74531e-09, 
    5.828539e-09, 5.10472e-09, 4.722223e-09, 4.249229e-09, 3.509853e-09,
  1.91716e-08, 1.862034e-08, 1.797597e-08, 1.721331e-08, 1.637093e-08, 
    1.530079e-08, 1.39431e-08, 1.23934e-08, 1.070764e-08, 8.378563e-09, 
    6.253974e-09, 5.177063e-09, 4.747891e-09, 4.374697e-09, 3.848691e-09,
  1.920543e-08, 1.865135e-08, 1.804426e-08, 1.745783e-08, 1.655249e-08, 
    1.56073e-08, 1.424718e-08, 1.282929e-08, 1.119577e-08, 8.994225e-09, 
    6.87807e-09, 5.36091e-09, 4.771511e-09, 4.452116e-09, 4.071472e-09,
  1.925431e-08, 1.872013e-08, 1.808428e-08, 1.761576e-08, 1.67508e-08, 
    1.585456e-08, 1.444639e-08, 1.314261e-08, 1.162803e-08, 9.532219e-09, 
    7.556692e-09, 5.779279e-09, 4.846749e-09, 4.484606e-09, 4.226883e-09,
  1.929575e-08, 1.880359e-08, 1.814377e-08, 1.770449e-08, 1.695867e-08, 
    1.604898e-08, 1.463426e-08, 1.328817e-08, 1.198527e-08, 9.973602e-09, 
    8.209866e-09, 6.347292e-09, 5.034088e-09, 4.552199e-09, 4.337934e-09,
  1.937324e-08, 1.890506e-08, 1.821427e-08, 1.778487e-08, 1.712514e-08, 
    1.6245e-08, 1.481287e-08, 1.336601e-08, 1.219859e-08, 1.041675e-08, 
    8.703079e-09, 7.001308e-09, 5.366959e-09, 4.705383e-09, 4.451361e-09,
  1.845351e-08, 1.716488e-08, 1.648989e-08, 1.468854e-08, 1.173251e-08, 
    9.313846e-09, 7.895897e-09, 7.133356e-09, 6.594715e-09, 5.980892e-09, 
    4.659862e-09, 3.980721e-09, 3.639592e-09, 3.383216e-09, 3.162291e-09,
  2.094659e-08, 1.827377e-08, 1.6652e-08, 1.523342e-08, 1.309905e-08, 
    1.074773e-08, 9.041976e-09, 7.845053e-09, 6.948087e-09, 6.374767e-09, 
    5.668203e-09, 4.466527e-09, 3.846339e-09, 3.572942e-09, 3.389213e-09,
  2.155533e-08, 2.013693e-08, 1.806039e-08, 1.644641e-08, 1.452598e-08, 
    1.214606e-08, 1.00945e-08, 8.657559e-09, 7.623383e-09, 6.82178e-09, 
    6.220731e-09, 5.39805e-09, 4.277309e-09, 3.762592e-09, 3.555241e-09,
  2.113658e-08, 2.107351e-08, 1.946284e-08, 1.809802e-08, 1.564175e-08, 
    1.330752e-08, 1.115654e-08, 9.575976e-09, 8.429296e-09, 7.455481e-09, 
    6.633524e-09, 6.050893e-09, 5.181218e-09, 4.241214e-09, 3.764992e-09,
  2.171969e-08, 2.128697e-08, 2.002708e-08, 1.889986e-08, 1.708832e-08, 
    1.426245e-08, 1.201019e-08, 1.047731e-08, 9.287543e-09, 8.321473e-09, 
    7.28948e-09, 6.464336e-09, 5.97261e-09, 5.094737e-09, 4.309272e-09,
  2.213341e-08, 2.147531e-08, 2.02632e-08, 1.916713e-08, 1.823832e-08, 
    1.582634e-08, 1.29282e-08, 1.110464e-08, 9.853477e-09, 8.785768e-09, 
    8.014961e-09, 7.098242e-09, 6.404915e-09, 5.866753e-09, 5.081349e-09,
  2.237797e-08, 2.176701e-08, 2.034224e-08, 1.911954e-08, 1.841061e-08, 
    1.713108e-08, 1.430943e-08, 1.183397e-08, 1.051127e-08, 9.211385e-09, 
    8.455488e-09, 7.737579e-09, 6.981751e-09, 6.354329e-09, 5.807617e-09,
  2.261203e-08, 2.244094e-08, 2.108064e-08, 1.932378e-08, 1.821523e-08, 
    1.753808e-08, 1.560665e-08, 1.293954e-08, 1.111615e-08, 9.971235e-09, 
    8.785221e-09, 8.327156e-09, 7.622353e-09, 6.820445e-09, 6.371141e-09,
  2.292459e-08, 2.292339e-08, 2.223624e-08, 2.067621e-08, 1.850758e-08, 
    1.772281e-08, 1.647419e-08, 1.421785e-08, 1.192421e-08, 1.056252e-08, 
    9.454597e-09, 8.588962e-09, 8.206408e-09, 7.278863e-09, 6.741327e-09,
  2.286282e-08, 2.305019e-08, 2.291677e-08, 2.214102e-08, 2.007699e-08, 
    1.838505e-08, 1.726499e-08, 1.528343e-08, 1.298387e-08, 1.124642e-08, 
    9.905833e-09, 9.014039e-09, 8.520351e-09, 7.872774e-09, 7.08803e-09,
  1.23983e-08, 1.249827e-08, 1.192243e-08, 9.91178e-09, 8.394141e-09, 
    7.466531e-09, 6.597559e-09, 5.752854e-09, 5.081811e-09, 4.4188e-09, 
    3.636286e-09, 2.919117e-09, 2.276143e-09, 1.842288e-09, 1.633922e-09,
  1.184576e-08, 1.206783e-08, 1.199228e-08, 1.07152e-08, 8.890116e-09, 
    7.766504e-09, 6.931225e-09, 6.067486e-09, 5.370903e-09, 4.779284e-09, 
    4.071762e-09, 3.367426e-09, 2.648309e-09, 2.115723e-09, 1.807818e-09,
  1.293895e-08, 1.206027e-08, 1.188624e-08, 1.124283e-08, 9.476511e-09, 
    8.125625e-09, 7.281857e-09, 6.421736e-09, 5.603644e-09, 5.066577e-09, 
    4.451874e-09, 3.803858e-09, 3.139726e-09, 2.533665e-09, 2.110153e-09,
  1.436813e-08, 1.287069e-08, 1.20013e-08, 1.129756e-08, 1.038836e-08, 
    8.720777e-09, 7.608519e-09, 6.819798e-09, 5.903706e-09, 5.268165e-09, 
    4.701955e-09, 4.145591e-09, 3.53641e-09, 2.997747e-09, 2.573743e-09,
  1.578061e-08, 1.404661e-08, 1.255278e-08, 1.168962e-08, 1.081955e-08, 
    9.598166e-09, 8.214821e-09, 7.211114e-09, 6.303072e-09, 5.520668e-09, 
    4.95251e-09, 4.344114e-09, 3.75234e-09, 3.252916e-09, 2.81594e-09,
  1.76121e-08, 1.567831e-08, 1.362741e-08, 1.233205e-08, 1.141421e-08, 
    1.036517e-08, 9.003615e-09, 7.885639e-09, 6.909705e-09, 5.867111e-09, 
    5.160169e-09, 4.550924e-09, 3.930107e-09, 3.38114e-09, 2.879828e-09,
  2.024503e-08, 1.786058e-08, 1.54237e-08, 1.360397e-08, 1.233376e-08, 
    1.112025e-08, 9.942989e-09, 8.555504e-09, 7.577106e-09, 6.568312e-09, 
    5.568499e-09, 4.786519e-09, 4.114163e-09, 3.509669e-09, 2.982822e-09,
  2.142414e-08, 2.025398e-08, 1.753924e-08, 1.528654e-08, 1.364183e-08, 
    1.225662e-08, 1.087514e-08, 9.57999e-09, 8.299474e-09, 7.257859e-09, 
    6.233795e-09, 5.284444e-09, 4.473269e-09, 3.834034e-09, 3.290352e-09,
  1.941752e-08, 2.072903e-08, 1.956237e-08, 1.71316e-08, 1.503938e-08, 
    1.342573e-08, 1.203819e-08, 1.058765e-08, 9.349104e-09, 8.071448e-09, 
    7.001919e-09, 6.001644e-09, 5.110146e-09, 4.394314e-09, 3.825925e-09,
  1.813931e-08, 1.886406e-08, 1.917968e-08, 1.835694e-08, 1.648704e-08, 
    1.440235e-08, 1.292774e-08, 1.173107e-08, 1.029645e-08, 9.081499e-09, 
    7.878915e-09, 6.848481e-09, 5.880266e-09, 5.084297e-09, 4.426264e-09,
  1.91728e-08, 1.704021e-08, 1.541747e-08, 1.283112e-08, 1.097465e-08, 
    9.692467e-09, 8.936345e-09, 8.252142e-09, 7.752571e-09, 7.340029e-09, 
    6.833667e-09, 5.909364e-09, 4.867063e-09, 3.972629e-09, 3.242622e-09,
  1.72511e-08, 1.538589e-08, 1.459363e-08, 1.257734e-08, 1.12346e-08, 
    1.010928e-08, 9.232619e-09, 8.46373e-09, 7.772301e-09, 7.265897e-09, 
    6.834857e-09, 5.976109e-09, 4.946726e-09, 4.061392e-09, 3.310344e-09,
  1.643575e-08, 1.443374e-08, 1.385114e-08, 1.26051e-08, 1.159044e-08, 
    1.060674e-08, 9.65904e-09, 8.626608e-09, 7.679802e-09, 7.159869e-09, 
    6.76697e-09, 6.066347e-09, 5.063369e-09, 4.165204e-09, 3.41051e-09,
  1.653253e-08, 1.397307e-08, 1.354607e-08, 1.286974e-08, 1.20281e-08, 
    1.112185e-08, 9.869712e-09, 8.645082e-09, 7.571773e-09, 7.029811e-09, 
    6.70997e-09, 6.121275e-09, 5.203277e-09, 4.284001e-09, 3.514656e-09,
  1.687494e-08, 1.419514e-08, 1.349394e-08, 1.28767e-08, 1.213669e-08, 
    1.123938e-08, 9.893962e-09, 8.600155e-09, 7.524518e-09, 6.904091e-09, 
    6.595954e-09, 6.153614e-09, 5.3556e-09, 4.437782e-09, 3.648995e-09,
  1.708969e-08, 1.453377e-08, 1.331832e-08, 1.255722e-08, 1.200123e-08, 
    1.126178e-08, 9.992191e-09, 8.675406e-09, 7.607802e-09, 6.871957e-09, 
    6.456591e-09, 6.155106e-09, 5.515321e-09, 4.606296e-09, 3.794375e-09,
  1.679005e-08, 1.476795e-08, 1.318119e-08, 1.231391e-08, 1.183753e-08, 
    1.120193e-08, 1.009988e-08, 8.833131e-09, 7.851939e-09, 6.982243e-09, 
    6.344458e-09, 6.115321e-09, 5.640174e-09, 4.803461e-09, 3.966475e-09,
  1.621389e-08, 1.483682e-08, 1.312557e-08, 1.234545e-08, 1.186793e-08, 
    1.1119e-08, 1.013407e-08, 9.055592e-09, 8.128223e-09, 7.212415e-09, 
    6.367781e-09, 6.050362e-09, 5.760837e-09, 5.03039e-09, 4.190412e-09,
  1.581317e-08, 1.478068e-08, 1.344975e-08, 1.280206e-08, 1.195743e-08, 
    1.100602e-08, 1.006145e-08, 9.240464e-09, 8.416746e-09, 7.400649e-09, 
    6.486129e-09, 6.023189e-09, 5.861331e-09, 5.246692e-09, 4.467923e-09,
  1.557219e-08, 1.486175e-08, 1.414264e-08, 1.345154e-08, 1.229348e-08, 
    1.107823e-08, 1.002084e-08, 9.341084e-09, 8.652767e-09, 7.653705e-09, 
    6.679913e-09, 6.033953e-09, 5.878213e-09, 5.487256e-09, 4.733498e-09,
  2.517931e-08, 2.58782e-08, 2.618176e-08, 2.597479e-08, 2.531906e-08, 
    2.488728e-08, 2.405497e-08, 2.33098e-08, 2.127107e-08, 1.84254e-08, 
    1.651919e-08, 1.402152e-08, 1.253425e-08, 1.064853e-08, 9.331501e-09,
  2.440363e-08, 2.560171e-08, 2.547596e-08, 2.490941e-08, 2.444609e-08, 
    2.416607e-08, 2.367333e-08, 2.319725e-08, 2.145956e-08, 1.841859e-08, 
    1.660542e-08, 1.398571e-08, 1.221125e-08, 1.042829e-08, 9.185531e-09,
  2.506042e-08, 2.575188e-08, 2.516454e-08, 2.458389e-08, 2.41745e-08, 
    2.398568e-08, 2.360922e-08, 2.311083e-08, 2.163046e-08, 1.848907e-08, 
    1.660983e-08, 1.397653e-08, 1.205922e-08, 1.02291e-08, 9.051839e-09,
  2.59472e-08, 2.550723e-08, 2.440163e-08, 2.406986e-08, 2.377554e-08, 
    2.366525e-08, 2.345435e-08, 2.28643e-08, 2.171588e-08, 1.862743e-08, 
    1.663682e-08, 1.400088e-08, 1.183419e-08, 1.000951e-08, 8.986057e-09,
  2.598877e-08, 2.480266e-08, 2.341348e-08, 2.339624e-08, 2.316531e-08, 
    2.318211e-08, 2.310003e-08, 2.234644e-08, 2.151232e-08, 1.86524e-08, 
    1.65206e-08, 1.385063e-08, 1.153874e-08, 9.769402e-09, 8.905955e-09,
  2.567159e-08, 2.425748e-08, 2.260366e-08, 2.260145e-08, 2.244863e-08, 
    2.266356e-08, 2.255977e-08, 2.171585e-08, 2.10776e-08, 1.836403e-08, 
    1.622596e-08, 1.363126e-08, 1.124304e-08, 9.570907e-09, 8.820013e-09,
  2.513629e-08, 2.366363e-08, 2.165184e-08, 2.1801e-08, 2.184257e-08, 
    2.198752e-08, 2.186083e-08, 2.096245e-08, 2.023958e-08, 1.781406e-08, 
    1.572101e-08, 1.326843e-08, 1.087487e-08, 9.366184e-09, 8.681569e-09,
  2.431181e-08, 2.282057e-08, 2.065917e-08, 2.132191e-08, 2.140142e-08, 
    2.13134e-08, 2.096555e-08, 2.009137e-08, 1.927194e-08, 1.699781e-08, 
    1.505063e-08, 1.27827e-08, 1.05439e-08, 9.182912e-09, 8.518879e-09,
  2.316934e-08, 2.182823e-08, 1.997576e-08, 2.090962e-08, 2.112207e-08, 
    2.057423e-08, 1.993313e-08, 1.895373e-08, 1.814316e-08, 1.608306e-08, 
    1.430919e-08, 1.227936e-08, 1.020517e-08, 9.015559e-09, 8.300473e-09,
  2.19633e-08, 2.104277e-08, 1.94961e-08, 2.062451e-08, 2.051111e-08, 
    1.962322e-08, 1.876245e-08, 1.776914e-08, 1.703249e-08, 1.516753e-08, 
    1.360259e-08, 1.176699e-08, 9.962716e-09, 8.897185e-09, 8.030796e-09,
  2.054086e-08, 2.011887e-08, 1.980226e-08, 1.937794e-08, 1.91582e-08, 
    1.8991e-08, 1.884832e-08, 1.885256e-08, 1.891399e-08, 1.855587e-08, 
    1.787332e-08, 1.680498e-08, 1.558959e-08, 1.470932e-08, 1.380156e-08,
  2.20121e-08, 2.111472e-08, 2.038502e-08, 1.986806e-08, 1.924371e-08, 
    1.919422e-08, 1.924752e-08, 1.931912e-08, 1.938321e-08, 1.900167e-08, 
    1.815001e-08, 1.719967e-08, 1.583236e-08, 1.484086e-08, 1.398304e-08,
  2.301781e-08, 2.236696e-08, 2.13381e-08, 2.075111e-08, 1.98562e-08, 
    1.939038e-08, 1.956988e-08, 1.989665e-08, 1.992396e-08, 1.952661e-08, 
    1.841795e-08, 1.749333e-08, 1.609243e-08, 1.494809e-08, 1.409569e-08,
  2.373424e-08, 2.35277e-08, 2.243424e-08, 2.168048e-08, 2.097872e-08, 
    2.004607e-08, 1.996615e-08, 2.046315e-08, 2.063572e-08, 2.013001e-08, 
    1.870676e-08, 1.77168e-08, 1.628983e-08, 1.501839e-08, 1.411067e-08,
  2.419959e-08, 2.44232e-08, 2.396677e-08, 2.290375e-08, 2.21947e-08, 
    2.095002e-08, 2.057684e-08, 2.106633e-08, 2.128955e-08, 2.072807e-08, 
    1.903103e-08, 1.791876e-08, 1.645604e-08, 1.506502e-08, 1.408459e-08,
  2.485838e-08, 2.494465e-08, 2.509956e-08, 2.428527e-08, 2.350004e-08, 
    2.231575e-08, 2.131976e-08, 2.174463e-08, 2.198028e-08, 2.137323e-08, 
    1.941031e-08, 1.813375e-08, 1.659627e-08, 1.505389e-08, 1.394103e-08,
  2.544841e-08, 2.545323e-08, 2.575314e-08, 2.584835e-08, 2.46791e-08, 
    2.390468e-08, 2.238469e-08, 2.270544e-08, 2.272129e-08, 2.200182e-08, 
    1.981466e-08, 1.833114e-08, 1.674304e-08, 1.49786e-08, 1.379357e-08,
  2.561823e-08, 2.574159e-08, 2.608528e-08, 2.679873e-08, 2.596223e-08, 
    2.505631e-08, 2.356873e-08, 2.359543e-08, 2.342056e-08, 2.252184e-08, 
    2.011361e-08, 1.848163e-08, 1.69232e-08, 1.494263e-08, 1.367711e-08,
  2.543119e-08, 2.569858e-08, 2.608794e-08, 2.720576e-08, 2.750186e-08, 
    2.617413e-08, 2.472442e-08, 2.471441e-08, 2.411728e-08, 2.286069e-08, 
    2.040831e-08, 1.862979e-08, 1.709808e-08, 1.501008e-08, 1.372204e-08,
  2.525725e-08, 2.560136e-08, 2.603124e-08, 2.711252e-08, 2.821692e-08, 
    2.756782e-08, 2.565063e-08, 2.567903e-08, 2.490421e-08, 2.295594e-08, 
    2.055581e-08, 1.884566e-08, 1.726659e-08, 1.51272e-08, 1.388591e-08,
  1.745893e-08, 1.694666e-08, 1.646206e-08, 1.607747e-08, 1.589308e-08, 
    1.559985e-08, 1.52257e-08, 1.472266e-08, 1.404358e-08, 1.340602e-08, 
    1.265995e-08, 1.174141e-08, 1.082821e-08, 9.832174e-09, 8.938108e-09,
  1.777763e-08, 1.730497e-08, 1.678804e-08, 1.619287e-08, 1.587658e-08, 
    1.564396e-08, 1.531839e-08, 1.485632e-08, 1.4282e-08, 1.360983e-08, 
    1.290814e-08, 1.205093e-08, 1.113562e-08, 1.010351e-08, 9.097794e-09,
  1.807752e-08, 1.763034e-08, 1.713183e-08, 1.640149e-08, 1.590803e-08, 
    1.569542e-08, 1.539909e-08, 1.498272e-08, 1.443474e-08, 1.383615e-08, 
    1.317334e-08, 1.230414e-08, 1.142004e-08, 1.040346e-08, 9.307485e-09,
  1.932578e-08, 1.797702e-08, 1.744855e-08, 1.68746e-08, 1.613354e-08, 
    1.568769e-08, 1.54462e-08, 1.503862e-08, 1.452193e-08, 1.39208e-08, 
    1.334457e-08, 1.254965e-08, 1.1701e-08, 1.072281e-08, 9.600119e-09,
  2.003056e-08, 1.915836e-08, 1.780974e-08, 1.724831e-08, 1.662705e-08, 
    1.598661e-08, 1.55214e-08, 1.515453e-08, 1.463359e-08, 1.40743e-08, 
    1.349797e-08, 1.274813e-08, 1.196038e-08, 1.100845e-08, 9.908534e-09,
  2.021288e-08, 1.985768e-08, 1.878795e-08, 1.761565e-08, 1.706323e-08, 
    1.640401e-08, 1.58038e-08, 1.532225e-08, 1.476747e-08, 1.418346e-08, 
    1.365532e-08, 1.293754e-08, 1.220915e-08, 1.133715e-08, 1.022955e-08,
  2.040673e-08, 2.001153e-08, 1.942444e-08, 1.842722e-08, 1.736918e-08, 
    1.704887e-08, 1.629591e-08, 1.561918e-08, 1.507873e-08, 1.435398e-08, 
    1.378809e-08, 1.310847e-08, 1.242705e-08, 1.161567e-08, 1.054657e-08,
  2.09799e-08, 2.054721e-08, 1.971669e-08, 1.911837e-08, 1.799311e-08, 
    1.714023e-08, 1.706353e-08, 1.615731e-08, 1.535412e-08, 1.46622e-08, 
    1.402263e-08, 1.331392e-08, 1.265925e-08, 1.194504e-08, 1.084279e-08,
  2.187667e-08, 2.12201e-08, 2.03869e-08, 1.949067e-08, 1.876466e-08, 
    1.756244e-08, 1.718834e-08, 1.693729e-08, 1.60025e-08, 1.500353e-08, 
    1.426739e-08, 1.35533e-08, 1.286647e-08, 1.223666e-08, 1.118639e-08,
  2.250425e-08, 2.215872e-08, 2.116175e-08, 2.013189e-08, 1.922537e-08, 
    1.82894e-08, 1.740169e-08, 1.71884e-08, 1.667729e-08, 1.56393e-08, 
    1.464522e-08, 1.382653e-08, 1.311291e-08, 1.249357e-08, 1.150504e-08,
  1.987194e-08, 1.976354e-08, 1.953039e-08, 1.937192e-08, 1.903585e-08, 
    1.895335e-08, 1.879853e-08, 1.844951e-08, 1.795717e-08, 1.737949e-08, 
    1.668765e-08, 1.613303e-08, 1.549754e-08, 1.479763e-08, 1.387634e-08,
  1.992577e-08, 1.966821e-08, 1.95245e-08, 1.940041e-08, 1.903985e-08, 
    1.876506e-08, 1.864488e-08, 1.836101e-08, 1.785758e-08, 1.730932e-08, 
    1.659712e-08, 1.602203e-08, 1.54055e-08, 1.470782e-08, 1.379415e-08,
  1.998362e-08, 1.971392e-08, 1.958125e-08, 1.945936e-08, 1.909446e-08, 
    1.86609e-08, 1.838095e-08, 1.820854e-08, 1.776077e-08, 1.721429e-08, 
    1.649886e-08, 1.590067e-08, 1.528905e-08, 1.460258e-08, 1.368536e-08,
  2.010382e-08, 1.975166e-08, 1.951923e-08, 1.936399e-08, 1.89893e-08, 
    1.859974e-08, 1.830366e-08, 1.802439e-08, 1.763012e-08, 1.709796e-08, 
    1.641219e-08, 1.577272e-08, 1.5159e-08, 1.448534e-08, 1.362673e-08,
  2.015677e-08, 1.985097e-08, 1.949211e-08, 1.92272e-08, 1.887188e-08, 
    1.847362e-08, 1.819554e-08, 1.796082e-08, 1.760488e-08, 1.69972e-08, 
    1.62653e-08, 1.565856e-08, 1.505832e-08, 1.439721e-08, 1.35501e-08,
  2.030639e-08, 1.98369e-08, 1.939326e-08, 1.903453e-08, 1.868355e-08, 
    1.831703e-08, 1.810689e-08, 1.78269e-08, 1.747805e-08, 1.694689e-08, 
    1.619934e-08, 1.552479e-08, 1.494788e-08, 1.434038e-08, 1.353602e-08,
  2.052539e-08, 2.004696e-08, 1.931691e-08, 1.884177e-08, 1.850137e-08, 
    1.813092e-08, 1.797389e-08, 1.772107e-08, 1.735374e-08, 1.689711e-08, 
    1.618356e-08, 1.542801e-08, 1.482066e-08, 1.426371e-08, 1.349004e-08,
  2.041427e-08, 1.993377e-08, 1.925885e-08, 1.869038e-08, 1.831318e-08, 
    1.800703e-08, 1.780504e-08, 1.762646e-08, 1.722205e-08, 1.676472e-08, 
    1.620451e-08, 1.543576e-08, 1.4679e-08, 1.414205e-08, 1.345101e-08,
  2.005724e-08, 1.968784e-08, 1.901646e-08, 1.854509e-08, 1.826271e-08, 
    1.793135e-08, 1.769139e-08, 1.745955e-08, 1.711538e-08, 1.665803e-08, 
    1.61435e-08, 1.54516e-08, 1.464933e-08, 1.397727e-08, 1.336555e-08,
  1.981991e-08, 1.941807e-08, 1.882928e-08, 1.827116e-08, 1.810881e-08, 
    1.790098e-08, 1.761903e-08, 1.747078e-08, 1.697489e-08, 1.653239e-08, 
    1.606147e-08, 1.550273e-08, 1.46442e-08, 1.389119e-08, 1.324721e-08,
  2.035561e-08, 2.068025e-08, 2.078762e-08, 2.083198e-08, 2.077513e-08, 
    2.069686e-08, 2.061918e-08, 2.043583e-08, 2.004695e-08, 1.960385e-08, 
    1.910318e-08, 1.857819e-08, 1.803293e-08, 1.714613e-08, 1.656778e-08,
  2.087369e-08, 2.113411e-08, 2.138222e-08, 2.159409e-08, 2.17362e-08, 
    2.169273e-08, 2.152009e-08, 2.12637e-08, 2.091217e-08, 2.043316e-08, 
    1.984859e-08, 1.926794e-08, 1.878106e-08, 1.817736e-08, 1.74607e-08,
  2.107148e-08, 2.123049e-08, 2.13234e-08, 2.172713e-08, 2.222262e-08, 
    2.24744e-08, 2.248482e-08, 2.217262e-08, 2.186109e-08, 2.129794e-08, 
    2.071696e-08, 1.998909e-08, 1.937256e-08, 1.880657e-08, 1.809348e-08,
  2.146482e-08, 2.148901e-08, 2.153987e-08, 2.182528e-08, 2.253465e-08, 
    2.284728e-08, 2.28615e-08, 2.25315e-08, 2.228438e-08, 2.178446e-08, 
    2.124654e-08, 2.058048e-08, 1.989697e-08, 1.929872e-08, 1.855321e-08,
  2.224778e-08, 2.220122e-08, 2.210801e-08, 2.227827e-08, 2.282381e-08, 
    2.313247e-08, 2.295956e-08, 2.259718e-08, 2.22895e-08, 2.195238e-08, 
    2.145722e-08, 2.095162e-08, 2.028131e-08, 1.96099e-08, 1.891986e-08,
  2.318316e-08, 2.294041e-08, 2.276619e-08, 2.280433e-08, 2.310112e-08, 
    2.31402e-08, 2.278069e-08, 2.240703e-08, 2.207904e-08, 2.179795e-08, 
    2.140401e-08, 2.10298e-08, 2.037112e-08, 1.973457e-08, 1.913763e-08,
  2.43889e-08, 2.404368e-08, 2.364175e-08, 2.352985e-08, 2.345174e-08, 
    2.322022e-08, 2.259459e-08, 2.212339e-08, 2.175069e-08, 2.153e-08, 
    2.121434e-08, 2.098051e-08, 2.036021e-08, 1.973038e-08, 1.927367e-08,
  2.49253e-08, 2.472393e-08, 2.437492e-08, 2.406535e-08, 2.369275e-08, 
    2.314894e-08, 2.243598e-08, 2.183184e-08, 2.145853e-08, 2.116795e-08, 
    2.097187e-08, 2.080255e-08, 2.024376e-08, 1.963352e-08, 1.922677e-08,
  2.453655e-08, 2.454964e-08, 2.432499e-08, 2.411457e-08, 2.367885e-08, 
    2.30296e-08, 2.226124e-08, 2.166017e-08, 2.125921e-08, 2.097847e-08, 
    2.073717e-08, 2.056238e-08, 2.003419e-08, 1.941642e-08, 1.906048e-08,
  2.413537e-08, 2.403549e-08, 2.398878e-08, 2.373443e-08, 2.333717e-08, 
    2.274173e-08, 2.211843e-08, 2.146841e-08, 2.112408e-08, 2.081632e-08, 
    2.059186e-08, 2.032596e-08, 1.980802e-08, 1.921555e-08, 1.890684e-08,
  1.546325e-08, 1.492434e-08, 1.467658e-08, 1.469599e-08, 1.462674e-08, 
    1.455118e-08, 1.439178e-08, 1.424888e-08, 1.403882e-08, 1.368265e-08, 
    1.344846e-08, 1.286316e-08, 1.220274e-08, 1.145884e-08, 1.067228e-08,
  1.752084e-08, 1.669766e-08, 1.596429e-08, 1.556625e-08, 1.536077e-08, 
    1.51934e-08, 1.506517e-08, 1.486743e-08, 1.478655e-08, 1.45111e-08, 
    1.446057e-08, 1.420526e-08, 1.379497e-08, 1.316161e-08, 1.229193e-08,
  1.892899e-08, 1.883109e-08, 1.796588e-08, 1.729873e-08, 1.692028e-08, 
    1.670304e-08, 1.655801e-08, 1.61833e-08, 1.596898e-08, 1.557395e-08, 
    1.526901e-08, 1.503858e-08, 1.474994e-08, 1.436642e-08, 1.373722e-08,
  1.95298e-08, 1.960888e-08, 1.945329e-08, 1.883213e-08, 1.819696e-08, 
    1.789594e-08, 1.787638e-08, 1.774466e-08, 1.75628e-08, 1.721432e-08, 
    1.687093e-08, 1.623476e-08, 1.582012e-08, 1.521717e-08, 1.483317e-08,
  2.01784e-08, 2.022894e-08, 2.019938e-08, 1.99316e-08, 1.955108e-08, 
    1.909303e-08, 1.890769e-08, 1.887341e-08, 1.879125e-08, 1.868164e-08, 
    1.839282e-08, 1.779906e-08, 1.696883e-08, 1.634594e-08, 1.555689e-08,
  2.075914e-08, 2.067811e-08, 2.064614e-08, 2.0632e-08, 2.042214e-08, 
    2.017397e-08, 1.995353e-08, 1.996752e-08, 1.986018e-08, 2.001816e-08, 
    1.977021e-08, 1.919638e-08, 1.828002e-08, 1.730439e-08, 1.655982e-08,
  2.167002e-08, 2.141605e-08, 2.153753e-08, 2.141649e-08, 2.119921e-08, 
    2.102949e-08, 2.058268e-08, 2.054367e-08, 2.067855e-08, 2.083432e-08, 
    2.073901e-08, 2.021032e-08, 1.930797e-08, 1.837688e-08, 1.722169e-08,
  2.174788e-08, 2.218211e-08, 2.21485e-08, 2.238366e-08, 2.238311e-08, 
    2.220776e-08, 2.176668e-08, 2.131046e-08, 2.144811e-08, 2.160646e-08, 
    2.147397e-08, 2.092952e-08, 1.99746e-08, 1.896766e-08, 1.797363e-08,
  2.227415e-08, 2.297893e-08, 2.312522e-08, 2.330267e-08, 2.325299e-08, 
    2.315245e-08, 2.26842e-08, 2.214956e-08, 2.183394e-08, 2.200486e-08, 
    2.186194e-08, 2.133644e-08, 2.045964e-08, 1.944749e-08, 1.820215e-08,
  2.327608e-08, 2.387376e-08, 2.426313e-08, 2.428425e-08, 2.431255e-08, 
    2.430281e-08, 2.415494e-08, 2.363546e-08, 2.310581e-08, 2.260047e-08, 
    2.214348e-08, 2.166169e-08, 2.077713e-08, 1.966955e-08, 1.841988e-08,
  1.420914e-08, 1.39201e-08, 1.362164e-08, 1.357955e-08, 1.336354e-08, 
    1.314311e-08, 1.259304e-08, 1.209967e-08, 1.152174e-08, 1.0863e-08, 
    1.024406e-08, 9.593835e-09, 8.671973e-09, 7.60302e-09, 6.574993e-09,
  1.487755e-08, 1.439393e-08, 1.394691e-08, 1.372686e-08, 1.345895e-08, 
    1.3331e-08, 1.322234e-08, 1.281481e-08, 1.237537e-08, 1.186275e-08, 
    1.119732e-08, 1.050448e-08, 9.883237e-09, 9.052645e-09, 8.11016e-09,
  1.670815e-08, 1.56495e-08, 1.481627e-08, 1.415245e-08, 1.378884e-08, 
    1.348343e-08, 1.328706e-08, 1.310806e-08, 1.292616e-08, 1.264428e-08, 
    1.228605e-08, 1.171434e-08, 1.10223e-08, 1.034218e-08, 9.500539e-09,
  2.010659e-08, 1.875352e-08, 1.723388e-08, 1.580077e-08, 1.460835e-08, 
    1.390355e-08, 1.357931e-08, 1.330562e-08, 1.307696e-08, 1.281391e-08, 
    1.27024e-08, 1.247394e-08, 1.215263e-08, 1.156928e-08, 1.085556e-08,
  2.336924e-08, 2.21962e-08, 2.102058e-08, 1.940437e-08, 1.771308e-08, 
    1.574802e-08, 1.449817e-08, 1.391107e-08, 1.354807e-08, 1.321533e-08, 
    1.290892e-08, 1.271512e-08, 1.253274e-08, 1.237852e-08, 1.199068e-08,
  2.365177e-08, 2.376763e-08, 2.289414e-08, 2.201092e-08, 2.089994e-08, 
    1.9276e-08, 1.698104e-08, 1.52313e-08, 1.437076e-08, 1.403159e-08, 
    1.367764e-08, 1.334446e-08, 1.301046e-08, 1.280797e-08, 1.267406e-08,
  2.412724e-08, 2.416901e-08, 2.392443e-08, 2.321866e-08, 2.25266e-08, 
    2.195965e-08, 2.055187e-08, 1.833535e-08, 1.595961e-08, 1.483186e-08, 
    1.449458e-08, 1.421845e-08, 1.393776e-08, 1.343011e-08, 1.326929e-08,
  2.391548e-08, 2.414951e-08, 2.357845e-08, 2.344495e-08, 2.268367e-08, 
    2.224377e-08, 2.227738e-08, 2.125117e-08, 1.949e-08, 1.680428e-08, 
    1.55371e-08, 1.517559e-08, 1.497081e-08, 1.462411e-08, 1.412298e-08,
  2.479254e-08, 2.428719e-08, 2.395979e-08, 2.359068e-08, 2.319192e-08, 
    2.242375e-08, 2.199144e-08, 2.19235e-08, 2.118403e-08, 1.952036e-08, 
    1.723959e-08, 1.62245e-08, 1.584457e-08, 1.567799e-08, 1.523151e-08,
  2.421707e-08, 2.391814e-08, 2.413982e-08, 2.418144e-08, 2.409802e-08, 
    2.363618e-08, 2.264017e-08, 2.251767e-08, 2.19406e-08, 2.119182e-08, 
    1.950111e-08, 1.76152e-08, 1.675095e-08, 1.64158e-08, 1.609559e-08,
  1.724229e-08, 1.693927e-08, 1.653816e-08, 1.633449e-08, 1.661595e-08, 
    1.648799e-08, 1.67968e-08, 1.678969e-08, 1.65628e-08, 1.602078e-08, 
    1.521915e-08, 1.419079e-08, 1.289783e-08, 1.186883e-08, 1.075515e-08,
  1.773238e-08, 1.741127e-08, 1.700112e-08, 1.649123e-08, 1.648957e-08, 
    1.642809e-08, 1.653823e-08, 1.652117e-08, 1.626625e-08, 1.604429e-08, 
    1.558785e-08, 1.491027e-08, 1.37804e-08, 1.252169e-08, 1.156235e-08,
  2.13551e-08, 1.911617e-08, 1.786248e-08, 1.693717e-08, 1.653802e-08, 
    1.648608e-08, 1.640184e-08, 1.651629e-08, 1.632515e-08, 1.5995e-08, 
    1.576039e-08, 1.539454e-08, 1.472293e-08, 1.38676e-08, 1.250484e-08,
  2.529634e-08, 2.313153e-08, 2.055157e-08, 1.855997e-08, 1.705579e-08, 
    1.656715e-08, 1.644344e-08, 1.641408e-08, 1.642256e-08, 1.617881e-08, 
    1.58268e-08, 1.554475e-08, 1.513416e-08, 1.47143e-08, 1.390872e-08,
  2.58793e-08, 2.567048e-08, 2.430111e-08, 2.18643e-08, 1.934897e-08, 
    1.736432e-08, 1.652634e-08, 1.647046e-08, 1.648684e-08, 1.625679e-08, 
    1.597222e-08, 1.567646e-08, 1.537799e-08, 1.495219e-08, 1.471472e-08,
  2.588097e-08, 2.599456e-08, 2.554643e-08, 2.473359e-08, 2.251969e-08, 
    2.007019e-08, 1.769132e-08, 1.663089e-08, 1.653252e-08, 1.655592e-08, 
    1.610665e-08, 1.583724e-08, 1.549163e-08, 1.520265e-08, 1.49459e-08,
  2.539846e-08, 2.595428e-08, 2.598594e-08, 2.554451e-08, 2.461396e-08, 
    2.283098e-08, 2.049042e-08, 1.809579e-08, 1.675613e-08, 1.656782e-08, 
    1.647173e-08, 1.601072e-08, 1.568551e-08, 1.535417e-08, 1.504345e-08,
  2.509871e-08, 2.58001e-08, 2.605387e-08, 2.622107e-08, 2.559695e-08, 
    2.466471e-08, 2.295238e-08, 2.069291e-08, 1.849103e-08, 1.693931e-08, 
    1.649016e-08, 1.631493e-08, 1.584796e-08, 1.557129e-08, 1.519983e-08,
  2.507061e-08, 2.472621e-08, 2.541294e-08, 2.562957e-08, 2.60282e-08, 
    2.558926e-08, 2.460307e-08, 2.29086e-08, 2.073596e-08, 1.872514e-08, 
    1.700034e-08, 1.643296e-08, 1.610946e-08, 1.566057e-08, 1.532275e-08,
  2.42092e-08, 2.387138e-08, 2.454318e-08, 2.515651e-08, 2.537559e-08, 
    2.55088e-08, 2.52618e-08, 2.427512e-08, 2.247291e-08, 2.068604e-08, 
    1.857983e-08, 1.681451e-08, 1.624816e-08, 1.586567e-08, 1.539352e-08,
  1.830698e-08, 1.860941e-08, 1.873226e-08, 1.878571e-08, 1.848369e-08, 
    1.820322e-08, 1.808501e-08, 1.772259e-08, 1.714697e-08, 1.645611e-08, 
    1.52389e-08, 1.386313e-08, 1.215869e-08, 1.029183e-08, 8.187115e-09,
  1.853541e-08, 1.869022e-08, 1.867857e-08, 1.875309e-08, 1.861052e-08, 
    1.823981e-08, 1.811247e-08, 1.766989e-08, 1.721447e-08, 1.641476e-08, 
    1.548866e-08, 1.410827e-08, 1.240273e-08, 1.059503e-08, 8.720762e-09,
  1.887112e-08, 1.884699e-08, 1.849458e-08, 1.843562e-08, 1.858821e-08, 
    1.837936e-08, 1.802996e-08, 1.74984e-08, 1.693862e-08, 1.63517e-08, 
    1.554056e-08, 1.421735e-08, 1.260162e-08, 1.082891e-08, 9.107672e-09,
  1.910648e-08, 1.864368e-08, 1.82091e-08, 1.806135e-08, 1.808345e-08, 
    1.80929e-08, 1.805545e-08, 1.755937e-08, 1.696746e-08, 1.627613e-08, 
    1.541848e-08, 1.430821e-08, 1.273909e-08, 1.107908e-08, 9.372167e-09,
  1.965748e-08, 1.878321e-08, 1.818458e-08, 1.801712e-08, 1.769882e-08, 
    1.773385e-08, 1.798392e-08, 1.765509e-08, 1.700149e-08, 1.611494e-08, 
    1.515486e-08, 1.410373e-08, 1.281166e-08, 1.124241e-08, 9.622875e-09,
  2.048651e-08, 1.939392e-08, 1.825197e-08, 1.802881e-08, 1.746331e-08, 
    1.752445e-08, 1.776833e-08, 1.77838e-08, 1.724073e-08, 1.611996e-08, 
    1.504223e-08, 1.389414e-08, 1.270979e-08, 1.138056e-08, 9.905356e-09,
  2.098536e-08, 1.987002e-08, 1.879072e-08, 1.818562e-08, 1.744172e-08, 
    1.729741e-08, 1.734672e-08, 1.752469e-08, 1.728704e-08, 1.644659e-08, 
    1.506241e-08, 1.383958e-08, 1.268494e-08, 1.15383e-08, 1.020089e-08,
  2.141165e-08, 2.051723e-08, 1.956327e-08, 1.8646e-08, 1.768605e-08, 
    1.723081e-08, 1.706478e-08, 1.71449e-08, 1.719233e-08, 1.643082e-08, 
    1.522614e-08, 1.392305e-08, 1.26466e-08, 1.168988e-08, 1.054833e-08,
  2.191102e-08, 2.076391e-08, 2.039672e-08, 1.943203e-08, 1.797821e-08, 
    1.707802e-08, 1.666982e-08, 1.670298e-08, 1.674126e-08, 1.642875e-08, 
    1.545769e-08, 1.42054e-08, 1.296709e-08, 1.193463e-08, 1.089376e-08,
  2.230916e-08, 2.114241e-08, 2.081598e-08, 2.028668e-08, 1.891426e-08, 
    1.73672e-08, 1.662924e-08, 1.654859e-08, 1.645727e-08, 1.63143e-08, 
    1.561202e-08, 1.436459e-08, 1.328492e-08, 1.245296e-08, 1.129501e-08,
  1.851916e-08, 1.893051e-08, 1.906266e-08, 1.908199e-08, 1.915095e-08, 
    1.91156e-08, 1.87309e-08, 1.811419e-08, 1.761755e-08, 1.753073e-08, 
    1.742e-08, 1.708284e-08, 1.618622e-08, 1.492932e-08, 1.346543e-08,
  1.900646e-08, 1.921712e-08, 1.925231e-08, 1.929233e-08, 1.921822e-08, 
    1.895304e-08, 1.853421e-08, 1.787119e-08, 1.746477e-08, 1.742481e-08, 
    1.730785e-08, 1.690081e-08, 1.609506e-08, 1.487896e-08, 1.34212e-08,
  1.924769e-08, 1.916752e-08, 1.929263e-08, 1.91835e-08, 1.904094e-08, 
    1.867396e-08, 1.823385e-08, 1.763194e-08, 1.728882e-08, 1.724145e-08, 
    1.714148e-08, 1.672902e-08, 1.593228e-08, 1.472435e-08, 1.325978e-08,
  1.96432e-08, 1.934501e-08, 1.935324e-08, 1.904418e-08, 1.889187e-08, 
    1.834866e-08, 1.791978e-08, 1.741403e-08, 1.730191e-08, 1.733182e-08, 
    1.708618e-08, 1.651943e-08, 1.563077e-08, 1.440782e-08, 1.297477e-08,
  1.973447e-08, 1.9199e-08, 1.90516e-08, 1.839879e-08, 1.822906e-08, 
    1.762379e-08, 1.742028e-08, 1.70993e-08, 1.71524e-08, 1.706294e-08, 
    1.67187e-08, 1.615732e-08, 1.516894e-08, 1.394754e-08, 1.256579e-08,
  1.946554e-08, 1.896632e-08, 1.890125e-08, 1.831712e-08, 1.809715e-08, 
    1.762793e-08, 1.754375e-08, 1.734512e-08, 1.736044e-08, 1.700327e-08, 
    1.657997e-08, 1.583334e-08, 1.484291e-08, 1.360542e-08, 1.221438e-08,
  1.887506e-08, 1.831921e-08, 1.828806e-08, 1.791421e-08, 1.790975e-08, 
    1.762231e-08, 1.750848e-08, 1.728871e-08, 1.701431e-08, 1.643355e-08, 
    1.583909e-08, 1.501778e-08, 1.409869e-08, 1.28685e-08, 1.151736e-08,
  1.800818e-08, 1.784812e-08, 1.817158e-08, 1.816379e-08, 1.816111e-08, 
    1.789089e-08, 1.768346e-08, 1.736973e-08, 1.690893e-08, 1.629222e-08, 
    1.56111e-08, 1.466721e-08, 1.371405e-08, 1.252805e-08, 1.129831e-08,
  1.798463e-08, 1.786017e-08, 1.809548e-08, 1.836483e-08, 1.847954e-08, 
    1.840319e-08, 1.813019e-08, 1.76335e-08, 1.699627e-08, 1.626729e-08, 
    1.542284e-08, 1.444522e-08, 1.328555e-08, 1.183308e-08, 1.061165e-08,
  1.856514e-08, 1.848682e-08, 1.884903e-08, 1.886376e-08, 1.901944e-08, 
    1.904657e-08, 1.849432e-08, 1.77091e-08, 1.683691e-08, 1.592552e-08, 
    1.484873e-08, 1.363233e-08, 1.225956e-08, 1.083229e-08, 9.591467e-09,
  1.974347e-08, 1.971758e-08, 1.954235e-08, 1.921515e-08, 1.887148e-08, 
    1.817906e-08, 1.741969e-08, 1.674938e-08, 1.588439e-08, 1.48486e-08, 
    1.361747e-08, 1.201889e-08, 1.044652e-08, 8.777456e-09, 7.297723e-09,
  2.000711e-08, 1.985476e-08, 1.969897e-08, 1.941131e-08, 1.91692e-08, 
    1.873517e-08, 1.807109e-08, 1.743211e-08, 1.677312e-08, 1.589489e-08, 
    1.486037e-08, 1.35328e-08, 1.204811e-08, 1.047749e-08, 8.821256e-09,
  1.999516e-08, 1.996742e-08, 1.987617e-08, 1.965715e-08, 1.944577e-08, 
    1.915318e-08, 1.867775e-08, 1.808292e-08, 1.750208e-08, 1.683883e-08, 
    1.591095e-08, 1.478749e-08, 1.340355e-08, 1.191884e-08, 1.033707e-08,
  2.014191e-08, 1.993789e-08, 1.981293e-08, 1.975459e-08, 1.96596e-08, 
    1.943732e-08, 1.903976e-08, 1.852522e-08, 1.801612e-08, 1.744986e-08, 
    1.668445e-08, 1.573942e-08, 1.459221e-08, 1.321983e-08, 1.173154e-08,
  2.0171e-08, 1.99153e-08, 1.981246e-08, 1.970415e-08, 1.968906e-08, 
    1.958611e-08, 1.936536e-08, 1.901035e-08, 1.850316e-08, 1.801177e-08, 
    1.743537e-08, 1.652585e-08, 1.551565e-08, 1.421178e-08, 1.284394e-08,
  2.022457e-08, 1.995392e-08, 1.986075e-08, 1.987844e-08, 1.970399e-08, 
    1.964816e-08, 1.939968e-08, 1.910118e-08, 1.875037e-08, 1.831642e-08, 
    1.778554e-08, 1.704401e-08, 1.612432e-08, 1.50818e-08, 1.376367e-08,
  2.025813e-08, 1.982319e-08, 1.998558e-08, 1.977042e-08, 1.966177e-08, 
    1.966809e-08, 1.956373e-08, 1.943145e-08, 1.913406e-08, 1.871399e-08, 
    1.823857e-08, 1.750894e-08, 1.66575e-08, 1.56336e-08, 1.44554e-08,
  2.065924e-08, 2.00356e-08, 2.038729e-08, 1.994695e-08, 1.993755e-08, 
    1.976657e-08, 1.95987e-08, 1.945516e-08, 1.921162e-08, 1.893546e-08, 
    1.848904e-08, 1.793792e-08, 1.717112e-08, 1.623063e-08, 1.511856e-08,
  2.03813e-08, 1.982921e-08, 2.016533e-08, 1.973218e-08, 2.016409e-08, 
    1.991143e-08, 1.968747e-08, 1.946088e-08, 1.930803e-08, 1.922941e-08, 
    1.883881e-08, 1.828128e-08, 1.747772e-08, 1.648996e-08, 1.552974e-08,
  2.0394e-08, 1.996289e-08, 2.04491e-08, 2.044325e-08, 2.061029e-08, 
    2.006859e-08, 1.977159e-08, 1.943566e-08, 1.929368e-08, 1.914041e-08, 
    1.879659e-08, 1.832704e-08, 1.75295e-08, 1.665688e-08, 1.58244e-08,
  1.818401e-08, 1.735783e-08, 1.605687e-08, 1.441126e-08, 1.293315e-08, 
    1.134489e-08, 1.011662e-08, 8.919813e-09, 7.569142e-09, 6.085894e-09, 
    4.559247e-09, 3.635067e-09, 2.840573e-09, 2.030065e-09, 1.560356e-09,
  1.859055e-08, 1.804449e-08, 1.716155e-08, 1.567562e-08, 1.415254e-08, 
    1.273751e-08, 1.138591e-08, 9.98614e-09, 8.815856e-09, 7.374722e-09, 
    5.821976e-09, 4.466981e-09, 3.588069e-09, 2.666394e-09, 1.953024e-09,
  1.883628e-08, 1.841751e-08, 1.781794e-08, 1.67878e-08, 1.534028e-08, 
    1.387485e-08, 1.256333e-08, 1.114607e-08, 9.795129e-09, 8.590831e-09, 
    7.082148e-09, 5.593011e-09, 4.366837e-09, 3.459248e-09, 2.520148e-09,
  1.929848e-08, 1.873021e-08, 1.830318e-08, 1.763602e-08, 1.645438e-08, 
    1.506003e-08, 1.366385e-08, 1.241856e-08, 1.096029e-08, 9.655374e-09, 
    8.35517e-09, 6.806352e-09, 5.406787e-09, 4.249071e-09, 3.304504e-09,
  1.956137e-08, 1.910812e-08, 1.861404e-08, 1.814001e-08, 1.742818e-08, 
    1.616544e-08, 1.48136e-08, 1.347812e-08, 1.220443e-08, 1.082443e-08, 
    9.534745e-09, 8.143672e-09, 6.596677e-09, 5.227188e-09, 4.038153e-09,
  1.994253e-08, 1.938694e-08, 1.892587e-08, 1.852846e-08, 1.795154e-08, 
    1.713955e-08, 1.588293e-08, 1.457182e-08, 1.33015e-08, 1.197385e-08, 
    1.059383e-08, 9.359933e-09, 7.902509e-09, 6.361588e-09, 5.004295e-09,
  2.016536e-08, 1.99074e-08, 1.938841e-08, 1.894082e-08, 1.841834e-08, 
    1.772741e-08, 1.682008e-08, 1.559889e-08, 1.435841e-08, 1.307872e-08, 
    1.168291e-08, 1.041732e-08, 9.144167e-09, 7.647745e-09, 6.074248e-09,
  2.026163e-08, 1.994107e-08, 1.959562e-08, 1.931553e-08, 1.889097e-08, 
    1.83364e-08, 1.749905e-08, 1.648269e-08, 1.534886e-08, 1.418083e-08, 
    1.277279e-08, 1.148327e-08, 1.020303e-08, 8.922873e-09, 7.34907e-09,
  2.01204e-08, 1.989882e-08, 1.993376e-08, 1.96954e-08, 1.924863e-08, 
    1.875966e-08, 1.810085e-08, 1.719934e-08, 1.617489e-08, 1.506526e-08, 
    1.373079e-08, 1.243468e-08, 1.116335e-08, 9.964579e-09, 8.620449e-09,
  1.981786e-08, 2.006677e-08, 2.004106e-08, 1.970146e-08, 1.958693e-08, 
    1.914328e-08, 1.857997e-08, 1.785135e-08, 1.691892e-08, 1.59513e-08, 
    1.473363e-08, 1.342351e-08, 1.20827e-08, 1.089521e-08, 9.703398e-09,
  2.381129e-08, 2.31144e-08, 2.267007e-08, 2.129521e-08, 1.956746e-08, 
    1.644024e-08, 1.34288e-08, 1.083365e-08, 8.96874e-09, 7.346834e-09, 
    5.553442e-09, 3.80473e-09, 2.744154e-09, 2.184312e-09, 1.828818e-09,
  2.424594e-08, 2.336431e-08, 2.296438e-08, 2.191634e-08, 2.057885e-08, 
    1.829151e-08, 1.533845e-08, 1.233752e-08, 9.962129e-09, 8.281906e-09, 
    6.573389e-09, 4.805048e-09, 3.340069e-09, 2.44093e-09, 1.96224e-09,
  2.428599e-08, 2.344327e-08, 2.313191e-08, 2.222844e-08, 2.109882e-08, 
    1.952805e-08, 1.705195e-08, 1.401905e-08, 1.115855e-08, 9.067171e-09, 
    7.444725e-09, 5.675251e-09, 4.063154e-09, 2.861249e-09, 2.129932e-09,
  2.428464e-08, 2.342314e-08, 2.325185e-08, 2.243412e-08, 2.126284e-08, 
    1.999102e-08, 1.821061e-08, 1.555783e-08, 1.254365e-08, 1.002857e-08, 
    8.21796e-09, 6.563567e-09, 4.912237e-09, 3.470791e-09, 2.463715e-09,
  2.396554e-08, 2.333686e-08, 2.325217e-08, 2.251773e-08, 2.157802e-08, 
    2.014629e-08, 1.890458e-08, 1.673787e-08, 1.389532e-08, 1.104203e-08, 
    9.039686e-09, 7.338988e-09, 5.707056e-09, 4.173768e-09, 2.896203e-09,
  2.3716e-08, 2.307616e-08, 2.317397e-08, 2.256285e-08, 2.176333e-08, 
    2.043438e-08, 1.912173e-08, 1.750051e-08, 1.507999e-08, 1.213247e-08, 
    9.847653e-09, 8.073216e-09, 6.404533e-09, 4.863279e-09, 3.436587e-09,
  2.326804e-08, 2.284618e-08, 2.302888e-08, 2.247823e-08, 2.175266e-08, 
    2.057786e-08, 1.933557e-08, 1.7907e-08, 1.590581e-08, 1.311581e-08, 
    1.0639e-08, 8.749211e-09, 7.069966e-09, 5.504455e-09, 4.000779e-09,
  2.274987e-08, 2.281153e-08, 2.280337e-08, 2.231845e-08, 2.169087e-08, 
    2.064636e-08, 1.944928e-08, 1.816185e-08, 1.649016e-08, 1.394093e-08, 
    1.141245e-08, 9.402376e-09, 7.678573e-09, 6.110546e-09, 4.567893e-09,
  2.236699e-08, 2.256346e-08, 2.255872e-08, 2.216168e-08, 2.15807e-08, 
    2.067781e-08, 1.950346e-08, 1.820467e-08, 1.680066e-08, 1.461937e-08, 
    1.207252e-08, 1.001586e-08, 8.275769e-09, 6.673822e-09, 5.102455e-09,
  2.196654e-08, 2.223744e-08, 2.229827e-08, 2.198236e-08, 2.138513e-08, 
    2.065338e-08, 1.960573e-08, 1.831971e-08, 1.694645e-08, 1.507494e-08, 
    1.269926e-08, 1.055488e-08, 8.810932e-09, 7.222616e-09, 5.623151e-09,
  2.051644e-08, 1.865281e-08, 1.561091e-08, 1.340115e-08, 1.118865e-08, 
    8.765492e-09, 6.869236e-09, 5.656681e-09, 4.696141e-09, 3.854677e-09, 
    2.938917e-09, 2.267504e-09, 1.951655e-09, 1.753762e-09, 1.580359e-09,
  2.105065e-08, 2.047942e-08, 1.861859e-08, 1.592347e-08, 1.337718e-08, 
    1.103256e-08, 8.803774e-09, 7.048142e-09, 5.727873e-09, 4.698538e-09, 
    3.82157e-09, 2.945583e-09, 2.299647e-09, 1.981566e-09, 1.785538e-09,
  2.168585e-08, 2.127589e-08, 2.031142e-08, 1.867517e-08, 1.603179e-08, 
    1.330519e-08, 1.083855e-08, 8.773307e-09, 7.100831e-09, 5.76354e-09, 
    4.631151e-09, 3.728677e-09, 2.88869e-09, 2.301901e-09, 2.00794e-09,
  2.210913e-08, 2.172827e-08, 2.13347e-08, 2.039274e-08, 1.870225e-08, 
    1.609179e-08, 1.324212e-08, 1.060293e-08, 8.672508e-09, 7.080373e-09, 
    5.696865e-09, 4.578286e-09, 3.675515e-09, 2.872334e-09, 2.320817e-09,
  2.201295e-08, 2.190326e-08, 2.177022e-08, 2.148549e-08, 2.052742e-08, 
    1.860492e-08, 1.600585e-08, 1.303514e-08, 1.035484e-08, 8.528553e-09, 
    6.978021e-09, 5.572671e-09, 4.492724e-09, 3.600818e-09, 2.826587e-09,
  2.242923e-08, 2.212776e-08, 2.191564e-08, 2.192049e-08, 2.163368e-08, 
    2.061378e-08, 1.850949e-08, 1.571933e-08, 1.261463e-08, 1.012722e-08, 
    8.334045e-09, 6.804433e-09, 5.416839e-09, 4.354233e-09, 3.468193e-09,
  2.260884e-08, 2.250216e-08, 2.212655e-08, 2.199991e-08, 2.20342e-08, 
    2.181107e-08, 2.054906e-08, 1.838887e-08, 1.513653e-08, 1.213707e-08, 
    9.831457e-09, 8.079942e-09, 6.586878e-09, 5.226784e-09, 4.169489e-09,
  2.230753e-08, 2.260598e-08, 2.246517e-08, 2.241708e-08, 2.227072e-08, 
    2.232432e-08, 2.186169e-08, 2.046089e-08, 1.784392e-08, 1.446579e-08, 
    1.158334e-08, 9.477395e-09, 7.757389e-09, 6.305547e-09, 4.964374e-09,
  2.213562e-08, 2.231873e-08, 2.245547e-08, 2.247505e-08, 2.258496e-08, 
    2.255267e-08, 2.257512e-08, 2.186993e-08, 2.011655e-08, 1.698867e-08, 
    1.364826e-08, 1.098337e-08, 9.051726e-09, 7.371885e-09, 5.952984e-09,
  2.225424e-08, 2.220514e-08, 2.226562e-08, 2.250581e-08, 2.260976e-08, 
    2.284046e-08, 2.284846e-08, 2.263653e-08, 2.161602e-08, 1.939863e-08, 
    1.59479e-08, 1.27633e-08, 1.035702e-08, 8.5429e-09, 6.934562e-09,
  1.293996e-08, 1.180478e-08, 1.083228e-08, 9.655745e-09, 8.579732e-09, 
    7.727982e-09, 6.997809e-09, 6.371811e-09, 5.623091e-09, 4.677538e-09, 
    3.563935e-09, 2.632485e-09, 2.123055e-09, 1.754443e-09, 1.446877e-09,
  1.3021e-08, 1.215841e-08, 1.117983e-08, 1.009647e-08, 8.944065e-09, 
    8.034389e-09, 7.232219e-09, 6.527589e-09, 5.849133e-09, 4.998787e-09, 
    3.977061e-09, 2.973968e-09, 2.281849e-09, 1.837337e-09, 1.491898e-09,
  1.334641e-08, 1.245075e-08, 1.147297e-08, 1.046957e-08, 9.371746e-09, 
    8.382091e-09, 7.545895e-09, 6.760708e-09, 6.043571e-09, 5.273749e-09, 
    4.343395e-09, 3.33851e-09, 2.526264e-09, 1.992014e-09, 1.601705e-09,
  1.372531e-08, 1.286113e-08, 1.188849e-08, 1.083479e-08, 9.764896e-09, 
    8.793571e-09, 7.903708e-09, 7.114361e-09, 6.372713e-09, 5.633776e-09, 
    4.720828e-09, 3.776905e-09, 2.852898e-09, 2.190267e-09, 1.731057e-09,
  1.392585e-08, 1.331673e-08, 1.242625e-08, 1.135689e-08, 1.020814e-08, 
    9.196699e-09, 8.327652e-09, 7.48249e-09, 6.720008e-09, 6.023004e-09, 
    5.138394e-09, 4.189457e-09, 3.269276e-09, 2.478612e-09, 1.899432e-09,
  1.414728e-08, 1.360479e-08, 1.294081e-08, 1.209859e-08, 1.084747e-08, 
    9.70185e-09, 8.773159e-09, 7.954044e-09, 7.10931e-09, 6.377518e-09, 
    5.609307e-09, 4.654411e-09, 3.722012e-09, 2.87772e-09, 2.157981e-09,
  1.459621e-08, 1.37336e-08, 1.32938e-08, 1.271386e-08, 1.166196e-08, 
    1.038999e-08, 9.320928e-09, 8.44161e-09, 7.582907e-09, 6.751026e-09, 
    5.973601e-09, 5.143195e-09, 4.214254e-09, 3.33689e-09, 2.537992e-09,
  1.553123e-08, 1.434846e-08, 1.354397e-08, 1.311394e-08, 1.243155e-08, 
    1.123369e-08, 1.003343e-08, 9.000025e-09, 8.08371e-09, 7.219179e-09, 
    6.399164e-09, 5.550552e-09, 4.703279e-09, 3.828157e-09, 3.003071e-09,
  1.653996e-08, 1.52295e-08, 1.416614e-08, 1.341054e-08, 1.298261e-08, 
    1.203584e-08, 1.092822e-08, 9.751155e-09, 8.706733e-09, 7.762283e-09, 
    6.911613e-09, 6.034045e-09, 5.157827e-09, 4.322565e-09, 3.471315e-09,
  1.734282e-08, 1.632009e-08, 1.505856e-08, 1.406256e-08, 1.338664e-08, 
    1.280641e-08, 1.172055e-08, 1.071181e-08, 9.499388e-09, 8.460866e-09, 
    7.534292e-09, 6.62096e-09, 5.656072e-09, 4.800615e-09, 3.973315e-09,
  1.828657e-08, 1.649838e-08, 1.475033e-08, 1.353736e-08, 1.242676e-08, 
    1.122433e-08, 9.959648e-09, 8.938823e-09, 8.115807e-09, 7.514927e-09, 
    6.849819e-09, 5.999699e-09, 5.073742e-09, 4.298319e-09, 3.637161e-09,
  1.890388e-08, 1.729769e-08, 1.558508e-08, 1.421881e-08, 1.307008e-08, 
    1.197973e-08, 1.06882e-08, 9.562775e-09, 8.656534e-09, 7.970897e-09, 
    7.37195e-09, 6.662766e-09, 5.731058e-09, 4.876452e-09, 4.186623e-09,
  1.964806e-08, 1.802342e-08, 1.631277e-08, 1.488649e-08, 1.368453e-08, 
    1.262333e-08, 1.143689e-08, 1.020367e-08, 9.198033e-09, 8.431769e-09, 
    7.805399e-09, 7.182198e-09, 6.361176e-09, 5.431002e-09, 4.685545e-09,
  2.047712e-08, 1.87674e-08, 1.700103e-08, 1.550066e-08, 1.422519e-08, 
    1.320415e-08, 1.209078e-08, 1.089393e-08, 9.792807e-09, 8.908871e-09, 
    8.205886e-09, 7.589835e-09, 6.93788e-09, 6.006609e-09, 5.184797e-09,
  2.13272e-08, 1.948729e-08, 1.763071e-08, 1.607022e-08, 1.473636e-08, 
    1.368355e-08, 1.267132e-08, 1.153741e-08, 1.038329e-08, 9.429167e-09, 
    8.655815e-09, 7.963898e-09, 7.346033e-09, 6.568804e-09, 5.680876e-09,
  2.189843e-08, 2.017978e-08, 1.827346e-08, 1.667561e-08, 1.523966e-08, 
    1.409268e-08, 1.313236e-08, 1.208565e-08, 1.100619e-08, 9.947895e-09, 
    9.150197e-09, 8.348351e-09, 7.705594e-09, 6.982182e-09, 6.174854e-09,
  2.223791e-08, 2.068165e-08, 1.884795e-08, 1.718197e-08, 1.575186e-08, 
    1.448995e-08, 1.350585e-08, 1.251613e-08, 1.151226e-08, 1.047361e-08, 
    9.592549e-09, 8.766871e-09, 8.010946e-09, 7.336397e-09, 6.587209e-09,
  2.25913e-08, 2.106896e-08, 1.936398e-08, 1.764346e-08, 1.619639e-08, 
    1.484932e-08, 1.37709e-08, 1.286019e-08, 1.193501e-08, 1.092007e-08, 
    1.000248e-08, 9.171577e-09, 8.356816e-09, 7.645557e-09, 6.90504e-09,
  2.275363e-08, 2.129191e-08, 1.969344e-08, 1.80613e-08, 1.663773e-08, 
    1.519414e-08, 1.408132e-08, 1.308257e-08, 1.223652e-08, 1.128509e-08, 
    1.037059e-08, 9.535214e-09, 8.710025e-09, 7.938516e-09, 7.20103e-09,
  2.29615e-08, 2.150046e-08, 2.001321e-08, 1.862897e-08, 1.710491e-08, 
    1.552059e-08, 1.435251e-08, 1.340737e-08, 1.250788e-08, 1.161236e-08, 
    1.072376e-08, 9.897752e-09, 9.053267e-09, 8.23584e-09, 7.466166e-09,
  1.073415e-08, 9.261208e-09, 8.041351e-09, 7.013871e-09, 6.080088e-09, 
    5.252662e-09, 4.523147e-09, 3.919421e-09, 3.394237e-09, 2.8138e-09, 
    2.22734e-09, 1.846243e-09, 1.672744e-09, 1.575409e-09, 1.397331e-09,
  1.138709e-08, 1.019073e-08, 8.856194e-09, 7.709892e-09, 6.775638e-09, 
    5.932855e-09, 5.17856e-09, 4.494451e-09, 3.939981e-09, 3.393163e-09, 
    2.858135e-09, 2.321354e-09, 1.915697e-09, 1.71338e-09, 1.615695e-09,
  1.205173e-08, 1.097465e-08, 9.793737e-09, 8.49037e-09, 7.458686e-09, 
    6.585701e-09, 5.836755e-09, 5.10633e-09, 4.494932e-09, 3.969259e-09, 
    3.457613e-09, 2.948287e-09, 2.443256e-09, 2.032637e-09, 1.793288e-09,
  1.270073e-08, 1.169933e-08, 1.061163e-08, 9.454025e-09, 8.260797e-09, 
    7.282586e-09, 6.50745e-09, 5.786527e-09, 5.127957e-09, 4.564981e-09, 
    4.058077e-09, 3.570412e-09, 3.107849e-09, 2.636387e-09, 2.235549e-09,
  1.329132e-08, 1.233994e-08, 1.134749e-08, 1.031163e-08, 9.26569e-09, 
    8.114803e-09, 7.207038e-09, 6.461662e-09, 5.771487e-09, 5.197373e-09, 
    4.667262e-09, 4.172636e-09, 3.730625e-09, 3.300761e-09, 2.854116e-09,
  1.393425e-08, 1.293527e-08, 1.202995e-08, 1.106628e-08, 1.011771e-08, 
    9.097683e-09, 8.021046e-09, 7.213988e-09, 6.458096e-09, 5.827242e-09, 
    5.276795e-09, 4.786837e-09, 4.33148e-09, 3.928356e-09, 3.500827e-09,
  1.453158e-08, 1.361492e-08, 1.272216e-08, 1.179199e-08, 1.086697e-08, 
    9.903506e-09, 8.932965e-09, 8.018326e-09, 7.224352e-09, 6.504741e-09, 
    5.900936e-09, 5.384996e-09, 4.918426e-09, 4.501878e-09, 4.10988e-09,
  1.508281e-08, 1.42946e-08, 1.34454e-08, 1.256513e-08, 1.166536e-08, 
    1.073568e-08, 9.780464e-09, 8.913329e-09, 8.068975e-09, 7.288401e-09, 
    6.600598e-09, 6.031721e-09, 5.542808e-09, 5.091498e-09, 4.697878e-09,
  1.569817e-08, 1.491222e-08, 1.416747e-08, 1.332639e-08, 1.24629e-08, 
    1.156293e-08, 1.064926e-08, 9.741654e-09, 8.944903e-09, 8.158555e-09, 
    7.396405e-09, 6.742303e-09, 6.190093e-09, 5.69692e-09, 5.268042e-09,
  1.643728e-08, 1.555549e-08, 1.477628e-08, 1.403215e-08, 1.323761e-08, 
    1.238333e-08, 1.151462e-08, 1.063433e-08, 9.743098e-09, 8.999105e-09, 
    8.260257e-09, 7.524556e-09, 6.892654e-09, 6.342574e-09, 5.864325e-09,
  1.1549e-08, 9.444501e-09, 7.769154e-09, 6.082141e-09, 4.800697e-09, 
    3.677845e-09, 2.804967e-09, 2.196357e-09, 1.640347e-09, 1.268757e-09, 
    1.065318e-09, 9.145142e-10, 7.538501e-10, 6.460393e-10, 5.770887e-10,
  1.208416e-08, 1.034253e-08, 8.539154e-09, 6.884501e-09, 5.493842e-09, 
    4.347942e-09, 3.35642e-09, 2.603477e-09, 2.024098e-09, 1.546342e-09, 
    1.199778e-09, 1.019727e-09, 8.613336e-10, 7.408864e-10, 6.316891e-10,
  1.262877e-08, 1.106529e-08, 9.375303e-09, 7.638417e-09, 6.195806e-09, 
    4.977105e-09, 3.991645e-09, 3.123544e-09, 2.441881e-09, 1.919504e-09, 
    1.483514e-09, 1.16185e-09, 9.801691e-10, 8.376176e-10, 7.312914e-10,
  1.315636e-08, 1.170926e-08, 1.016444e-08, 8.508178e-09, 6.965504e-09, 
    5.656265e-09, 4.58971e-09, 3.719145e-09, 2.953094e-09, 2.351896e-09, 
    1.871189e-09, 1.4597e-09, 1.157376e-09, 9.787985e-10, 8.516201e-10,
  1.376821e-08, 1.235081e-08, 1.086834e-08, 9.27887e-09, 7.76328e-09, 
    6.411911e-09, 5.236934e-09, 4.31627e-09, 3.523826e-09, 2.848086e-09, 
    2.288313e-09, 1.848938e-09, 1.460502e-09, 1.194049e-09, 1.008895e-09,
  1.430794e-08, 1.286583e-08, 1.145494e-08, 1.006044e-08, 8.498244e-09, 
    7.17139e-09, 5.921901e-09, 4.918611e-09, 4.116411e-09, 3.409844e-09, 
    2.78724e-09, 2.266307e-09, 1.852463e-09, 1.519071e-09, 1.26477e-09,
  1.484861e-08, 1.340778e-08, 1.19703e-08, 1.072135e-08, 9.276858e-09, 
    7.947101e-09, 6.625774e-09, 5.573523e-09, 4.716116e-09, 4.006345e-09, 
    3.354295e-09, 2.784613e-09, 2.286253e-09, 1.894181e-09, 1.587254e-09,
  1.51097e-08, 1.377983e-08, 1.251804e-08, 1.132833e-08, 1.00131e-08, 
    8.771841e-09, 7.332205e-09, 6.214964e-09, 5.331344e-09, 4.616681e-09, 
    3.962621e-09, 3.367512e-09, 2.850209e-09, 2.355674e-09, 1.975011e-09,
  1.518571e-08, 1.414809e-08, 1.296975e-08, 1.180054e-08, 1.06776e-08, 
    9.578686e-09, 8.125334e-09, 6.895426e-09, 5.974023e-09, 5.209672e-09, 
    4.554924e-09, 3.954323e-09, 3.426445e-09, 2.937496e-09, 2.485246e-09,
  1.515095e-08, 1.432258e-08, 1.320488e-08, 1.212197e-08, 1.114419e-08, 
    1.024752e-08, 8.940581e-09, 7.641153e-09, 6.668672e-09, 5.849625e-09, 
    5.14413e-09, 4.54241e-09, 4.025624e-09, 3.542898e-09, 3.089858e-09,
  1.899355e-08, 1.759601e-08, 1.630402e-08, 1.449718e-08, 1.237958e-08, 
    1.008132e-08, 7.304134e-09, 5.503791e-09, 4.373152e-09, 3.61455e-09, 
    3.067619e-09, 2.724548e-09, 2.525187e-09, 2.122022e-09, 1.78871e-09,
  1.918642e-08, 1.80472e-08, 1.69208e-08, 1.534194e-08, 1.341419e-08, 
    1.125109e-08, 8.697757e-09, 6.464402e-09, 5.103168e-09, 4.161125e-09, 
    3.455808e-09, 2.9264e-09, 2.647259e-09, 2.364435e-09, 2.02849e-09,
  1.934632e-08, 1.847411e-08, 1.735626e-08, 1.604477e-08, 1.437852e-08, 
    1.236665e-08, 1.00233e-08, 7.65641e-09, 5.883006e-09, 4.765619e-09, 
    3.950089e-09, 3.279959e-09, 2.871126e-09, 2.52353e-09, 2.248449e-09,
  1.957761e-08, 1.867033e-08, 1.767981e-08, 1.644703e-08, 1.511578e-08, 
    1.331877e-08, 1.120712e-08, 8.828756e-09, 6.813709e-09, 5.416072e-09, 
    4.475785e-09, 3.735003e-09, 3.185448e-09, 2.766632e-09, 2.446405e-09,
  1.964639e-08, 1.890724e-08, 1.801444e-08, 1.68907e-08, 1.57065e-08, 
    1.417976e-08, 1.229083e-08, 1.005095e-08, 7.880002e-09, 6.148735e-09, 
    5.064237e-09, 4.230638e-09, 3.559118e-09, 3.06228e-09, 2.622842e-09,
  1.967572e-08, 1.896575e-08, 1.820269e-08, 1.720708e-08, 1.618765e-08, 
    1.501839e-08, 1.320679e-08, 1.106749e-08, 8.898033e-09, 7.060012e-09, 
    5.639333e-09, 4.752793e-09, 3.987483e-09, 3.405571e-09, 2.907113e-09,
  1.973986e-08, 1.923141e-08, 1.852259e-08, 1.756012e-08, 1.669691e-08, 
    1.579287e-08, 1.421728e-08, 1.214665e-08, 9.820996e-09, 7.920718e-09, 
    6.425951e-09, 5.311657e-09, 4.471399e-09, 3.790793e-09, 3.26922e-09,
  1.963461e-08, 1.909156e-08, 1.863394e-08, 1.772971e-08, 1.684008e-08, 
    1.592632e-08, 1.463334e-08, 1.308045e-08, 1.093176e-08, 8.8165e-09, 
    7.206969e-09, 5.998686e-09, 5.049549e-09, 4.231703e-09, 3.626782e-09,
  1.918078e-08, 1.901129e-08, 1.87849e-08, 1.75507e-08, 1.672175e-08, 
    1.58532e-08, 1.460671e-08, 1.357311e-08, 1.171406e-08, 9.71975e-09, 
    8.022877e-09, 6.652668e-09, 5.681476e-09, 4.813812e-09, 4.006614e-09,
  1.903061e-08, 1.890447e-08, 1.871074e-08, 1.743025e-08, 1.669859e-08, 
    1.568677e-08, 1.499833e-08, 1.399561e-08, 1.236285e-08, 1.032837e-08, 
    8.749483e-09, 7.250948e-09, 6.152706e-09, 5.314537e-09, 4.501951e-09,
  1.252577e-08, 1.105044e-08, 9.482317e-09, 7.734244e-09, 6.651649e-09, 
    5.892204e-09, 5.221487e-09, 4.530554e-09, 3.815804e-09, 3.38228e-09, 
    2.83898e-09, 2.275155e-09, 1.967282e-09, 1.815816e-09, 1.70282e-09,
  1.353681e-08, 1.197571e-08, 1.068198e-08, 9.06802e-09, 7.591721e-09, 
    6.610349e-09, 5.894723e-09, 5.263712e-09, 4.600054e-09, 3.953315e-09, 
    3.413682e-09, 2.904866e-09, 2.436194e-09, 2.132401e-09, 1.896376e-09,
  1.508035e-08, 1.338415e-08, 1.19035e-08, 1.039921e-08, 8.859921e-09, 
    7.548873e-09, 6.574244e-09, 5.829981e-09, 5.194075e-09, 4.648288e-09, 
    3.992753e-09, 3.440422e-09, 2.959218e-09, 2.537269e-09, 2.219344e-09,
  1.604044e-08, 1.496152e-08, 1.340608e-08, 1.183652e-08, 1.033248e-08, 
    8.877206e-09, 7.532007e-09, 6.531392e-09, 5.769661e-09, 5.205237e-09, 
    4.702426e-09, 4.071722e-09, 3.517655e-09, 3.079161e-09, 2.675299e-09,
  1.704171e-08, 1.639647e-08, 1.499201e-08, 1.340322e-08, 1.183329e-08, 
    1.035832e-08, 8.879063e-09, 7.492711e-09, 6.48192e-09, 5.781655e-09, 
    5.251449e-09, 4.789074e-09, 4.171686e-09, 3.617216e-09, 3.199471e-09,
  1.742146e-08, 1.71974e-08, 1.641126e-08, 1.496093e-08, 1.344528e-08, 
    1.176465e-08, 1.03113e-08, 8.833217e-09, 7.502544e-09, 6.541829e-09, 
    5.881881e-09, 5.358956e-09, 4.914967e-09, 4.328666e-09, 3.781779e-09,
  1.783229e-08, 1.762154e-08, 1.724307e-08, 1.637247e-08, 1.513119e-08, 
    1.358397e-08, 1.187767e-08, 1.034723e-08, 8.938331e-09, 7.744173e-09, 
    6.773918e-09, 6.048344e-09, 5.567275e-09, 5.147919e-09, 4.615072e-09,
  1.881941e-08, 1.817367e-08, 1.786414e-08, 1.719673e-08, 1.63282e-08, 
    1.522008e-08, 1.374229e-08, 1.208795e-08, 1.047067e-08, 9.135124e-09, 
    8.076391e-09, 7.125439e-09, 6.367378e-09, 5.856332e-09, 5.437522e-09,
  1.980322e-08, 1.899349e-08, 1.863133e-08, 1.816724e-08, 1.755745e-08, 
    1.661186e-08, 1.54554e-08, 1.38914e-08, 1.222122e-08, 1.056672e-08, 
    9.266766e-09, 8.406277e-09, 7.555007e-09, 6.870533e-09, 6.300893e-09,
  2.129679e-08, 2.058576e-08, 1.94743e-08, 1.895467e-08, 1.830873e-08, 
    1.782843e-08, 1.707231e-08, 1.565507e-08, 1.403096e-08, 1.234129e-08, 
    1.075412e-08, 9.57237e-09, 8.766595e-09, 8.043845e-09, 7.345449e-09,
  1.103682e-08, 8.636e-09, 6.671418e-09, 5.208119e-09, 4.031464e-09, 
    3.001103e-09, 2.252891e-09, 1.730426e-09, 1.434864e-09, 1.223343e-09, 
    9.635683e-10, 8.139682e-10, 6.844273e-10, 6.117269e-10, 5.547461e-10,
  1.183212e-08, 9.929528e-09, 7.862923e-09, 6.131611e-09, 4.839249e-09, 
    3.74848e-09, 2.867404e-09, 2.183498e-09, 1.704957e-09, 1.465635e-09, 
    1.245275e-09, 9.842961e-10, 8.111596e-10, 6.81766e-10, 5.82891e-10,
  1.26405e-08, 1.092771e-08, 9.162393e-09, 7.24942e-09, 5.679081e-09, 
    4.504066e-09, 3.498625e-09, 2.698727e-09, 2.078584e-09, 1.652124e-09, 
    1.442145e-09, 1.225719e-09, 9.875494e-10, 8.057311e-10, 6.95462e-10,
  1.347988e-08, 1.189156e-08, 1.024417e-08, 8.388936e-09, 6.65394e-09, 
    5.322719e-09, 4.2578e-09, 3.347343e-09, 2.617723e-09, 2.036509e-09, 
    1.659139e-09, 1.443182e-09, 1.252204e-09, 1.036994e-09, 8.677686e-10,
  1.42645e-08, 1.279601e-08, 1.125559e-08, 9.374125e-09, 7.657571e-09, 
    6.20104e-09, 5.049878e-09, 4.053677e-09, 3.256918e-09, 2.577887e-09, 
    2.056364e-09, 1.701879e-09, 1.482605e-09, 1.301828e-09, 1.129845e-09,
  1.495454e-08, 1.35293e-08, 1.21276e-08, 1.037788e-08, 8.67918e-09, 
    7.19885e-09, 5.920676e-09, 4.832196e-09, 3.927573e-09, 3.209548e-09, 
    2.593501e-09, 2.110136e-09, 1.778779e-09, 1.540652e-09, 1.364383e-09,
  1.54507e-08, 1.424016e-08, 1.300519e-08, 1.138972e-08, 9.698356e-09, 
    8.262697e-09, 6.885609e-09, 5.718325e-09, 4.724605e-09, 3.901649e-09, 
    3.223666e-09, 2.64949e-09, 2.191464e-09, 1.847812e-09, 1.599002e-09,
  1.576123e-08, 1.481791e-08, 1.377603e-08, 1.24157e-08, 1.077217e-08, 
    9.330043e-09, 7.93404e-09, 6.703959e-09, 5.612977e-09, 4.708231e-09, 
    3.963278e-09, 3.297359e-09, 2.761692e-09, 2.321831e-09, 1.978484e-09,
  1.590209e-08, 1.528455e-08, 1.444777e-08, 1.319117e-08, 1.174979e-08, 
    1.039137e-08, 8.984961e-09, 7.719321e-09, 6.602429e-09, 5.60848e-09, 
    4.757383e-09, 4.0211e-09, 3.394431e-09, 2.900738e-09, 2.489959e-09,
  1.611962e-08, 1.55147e-08, 1.478447e-08, 1.385154e-08, 1.249944e-08, 
    1.129975e-08, 9.977325e-09, 8.749478e-09, 7.590658e-09, 6.577769e-09, 
    5.712053e-09, 4.926723e-09, 4.171027e-09, 3.538585e-09, 3.064397e-09,
  1.491231e-08, 1.223291e-08, 9.823267e-09, 7.702982e-09, 5.749539e-09, 
    4.101822e-09, 2.996365e-09, 2.347664e-09, 1.846078e-09, 1.524942e-09, 
    1.23165e-09, 1.012628e-09, 8.333558e-10, 6.677969e-10, 5.619149e-10,
  1.566898e-08, 1.344429e-08, 1.090755e-08, 8.637829e-09, 6.738379e-09, 
    4.910448e-09, 3.518252e-09, 2.611948e-09, 2.074187e-09, 1.684472e-09, 
    1.37708e-09, 1.116067e-09, 9.409891e-10, 7.717822e-10, 6.309235e-10,
  1.642822e-08, 1.443965e-08, 1.209188e-08, 9.634047e-09, 7.633905e-09, 
    5.839927e-09, 4.250347e-09, 3.054005e-09, 2.301941e-09, 1.83605e-09, 
    1.524617e-09, 1.254724e-09, 1.041353e-09, 8.72607e-10, 7.314801e-10,
  1.700544e-08, 1.530704e-08, 1.314089e-08, 1.073484e-08, 8.571272e-09, 
    6.731998e-09, 5.111081e-09, 3.700815e-09, 2.670596e-09, 2.02437e-09, 
    1.667084e-09, 1.404043e-09, 1.163715e-09, 9.860519e-10, 8.327586e-10,
  1.746767e-08, 1.592811e-08, 1.404941e-08, 1.177593e-08, 9.587372e-09, 
    7.591867e-09, 5.953083e-09, 4.442803e-09, 3.177745e-09, 2.317441e-09, 
    1.832927e-09, 1.541939e-09, 1.300336e-09, 1.091636e-09, 9.344787e-10,
  1.779637e-08, 1.638436e-08, 1.472308e-08, 1.269271e-08, 1.058737e-08, 
    8.472399e-09, 6.702747e-09, 5.197047e-09, 3.782669e-09, 2.703132e-09, 
    2.06098e-09, 1.710058e-09, 1.433765e-09, 1.214099e-09, 1.032455e-09,
  1.810244e-08, 1.68364e-08, 1.532295e-08, 1.347412e-08, 1.140234e-08, 
    9.337698e-09, 7.413842e-09, 5.908047e-09, 4.426355e-09, 3.181143e-09, 
    2.352323e-09, 1.903106e-09, 1.595001e-09, 1.357926e-09, 1.153014e-09,
  1.828621e-08, 1.721368e-08, 1.58552e-08, 1.413326e-08, 1.20819e-08, 
    1.008445e-08, 8.169693e-09, 6.672424e-09, 5.152605e-09, 3.790516e-09, 
    2.746131e-09, 2.150324e-09, 1.763231e-09, 1.505987e-09, 1.301561e-09,
  1.840949e-08, 1.746153e-08, 1.624367e-08, 1.456787e-08, 1.273039e-08, 
    1.074632e-08, 8.886175e-09, 7.380338e-09, 5.971216e-09, 4.498115e-09, 
    3.28596e-09, 2.472019e-09, 1.984746e-09, 1.657671e-09, 1.44513e-09,
  1.830978e-08, 1.760394e-08, 1.651189e-08, 1.50624e-08, 1.333472e-08, 
    1.142187e-08, 9.524543e-09, 8.097461e-09, 6.729844e-09, 5.267961e-09, 
    3.977803e-09, 2.944375e-09, 2.260164e-09, 1.846489e-09, 1.579131e-09,
  1.725959e-08, 1.550127e-08, 1.338287e-08, 1.137633e-08, 9.194616e-09, 
    6.864409e-09, 4.753399e-09, 3.339489e-09, 2.433658e-09, 1.702779e-09, 
    1.340294e-09, 1.245752e-09, 1.190644e-09, 1.096986e-09, 1.020146e-09,
  1.785424e-08, 1.653394e-08, 1.466395e-08, 1.275983e-08, 1.064442e-08, 
    8.363701e-09, 6.212405e-09, 4.397228e-09, 3.094982e-09, 2.178144e-09, 
    1.566353e-09, 1.318075e-09, 1.226657e-09, 1.168312e-09, 1.070682e-09,
  1.846072e-08, 1.737038e-08, 1.572839e-08, 1.391237e-08, 1.194249e-08, 
    9.79798e-09, 7.502849e-09, 5.617473e-09, 3.959816e-09, 2.771889e-09, 
    1.927421e-09, 1.47208e-09, 1.25266e-09, 1.183011e-09, 1.134983e-09,
  1.914845e-08, 1.80174e-08, 1.670615e-08, 1.510516e-08, 1.314841e-08, 
    1.112944e-08, 8.94277e-09, 6.830622e-09, 5.043362e-09, 3.574741e-09, 
    2.482224e-09, 1.764806e-09, 1.413152e-09, 1.192337e-09, 1.174701e-09,
  1.961437e-08, 1.853707e-08, 1.73896e-08, 1.602354e-08, 1.436203e-08, 
    1.246913e-08, 1.031593e-08, 8.226468e-09, 6.269196e-09, 4.585608e-09, 
    3.243527e-09, 2.259176e-09, 1.680256e-09, 1.350267e-09, 1.179771e-09,
  2.001123e-08, 1.91154e-08, 1.811177e-08, 1.691484e-08, 1.537945e-08, 
    1.369288e-08, 1.1682e-08, 9.547309e-09, 7.554822e-09, 5.746881e-09, 
    4.159578e-09, 2.902202e-09, 2.098121e-09, 1.60189e-09, 1.318907e-09,
  2.023078e-08, 1.949096e-08, 1.859738e-08, 1.761493e-08, 1.62756e-08, 
    1.478453e-08, 1.30344e-08, 1.093624e-08, 8.861745e-09, 6.984688e-09, 
    5.2714e-09, 3.749939e-09, 2.664953e-09, 2.002878e-09, 1.562564e-09,
  2.051475e-08, 1.996104e-08, 1.921687e-08, 1.833519e-08, 1.709254e-08, 
    1.573236e-08, 1.407375e-08, 1.224796e-08, 1.016797e-08, 8.160989e-09, 
    6.433105e-09, 4.799746e-09, 3.442969e-09, 2.531466e-09, 1.89662e-09,
  2.048328e-08, 1.997379e-08, 1.933084e-08, 1.8617e-08, 1.765747e-08, 
    1.650313e-08, 1.507672e-08, 1.331248e-08, 1.143053e-08, 9.394784e-09, 
    7.512481e-09, 5.912268e-09, 4.384697e-09, 3.2334e-09, 2.359024e-09,
  2.053459e-08, 2.011373e-08, 1.962228e-08, 1.904239e-08, 1.81254e-08, 
    1.710436e-08, 1.587798e-08, 1.433029e-08, 1.255738e-08, 1.061686e-08, 
    8.717767e-09, 6.97038e-09, 5.427758e-09, 3.994283e-09, 2.95758e-09,
  1.292933e-08, 9.899442e-09, 6.998155e-09, 4.293318e-09, 2.962125e-09, 
    2.252025e-09, 1.697559e-09, 1.216872e-09, 8.894818e-10, 7.181731e-10, 
    6.214675e-10, 5.791539e-10, 6.042061e-10, 6.770646e-10, 7.622529e-10,
  1.338167e-08, 1.095079e-08, 8.15358e-09, 5.185254e-09, 3.360942e-09, 
    2.477939e-09, 1.88593e-09, 1.368226e-09, 9.578234e-10, 7.686463e-10, 
    6.544381e-10, 5.851128e-10, 5.835833e-10, 6.394586e-10, 7.247416e-10,
  1.392088e-08, 1.183185e-08, 9.145277e-09, 6.2176e-09, 3.990776e-09, 
    2.777763e-09, 2.10201e-09, 1.535427e-09, 1.056401e-09, 8.192005e-10, 
    6.933533e-10, 6.104834e-10, 5.718681e-10, 6.052543e-10, 6.846888e-10,
  1.453667e-08, 1.253519e-08, 1.009797e-08, 7.303212e-09, 4.837259e-09, 
    3.25901e-09, 2.368787e-09, 1.706485e-09, 1.197709e-09, 8.889897e-10, 
    7.483817e-10, 6.519606e-10, 5.906645e-10, 5.875835e-10, 6.460203e-10,
  1.519339e-08, 1.315436e-08, 1.094977e-08, 8.369783e-09, 5.875594e-09, 
    3.942787e-09, 2.743368e-09, 1.949656e-09, 1.362045e-09, 9.920101e-10, 
    8.174116e-10, 7.048916e-10, 6.28293e-10, 5.886193e-10, 6.142318e-10,
  1.578792e-08, 1.381225e-08, 1.169389e-08, 9.388921e-09, 6.893777e-09, 
    4.809933e-09, 3.291849e-09, 2.265078e-09, 1.560362e-09, 1.12173e-09, 
    9.043815e-10, 7.771166e-10, 6.781267e-10, 6.099906e-10, 6.016488e-10,
  1.630289e-08, 1.436383e-08, 1.237763e-08, 1.030459e-08, 7.926165e-09, 
    5.775206e-09, 4.033551e-09, 2.723694e-09, 1.833188e-09, 1.281603e-09, 
    9.99922e-10, 8.623498e-10, 7.49318e-10, 6.562432e-10, 6.140378e-10,
  1.677513e-08, 1.493257e-08, 1.298919e-08, 1.107689e-08, 8.894715e-09, 
    6.832419e-09, 4.967922e-09, 3.346468e-09, 2.21634e-09, 1.525573e-09, 
    1.132564e-09, 9.467321e-10, 8.239918e-10, 7.221208e-10, 6.451886e-10,
  1.710755e-08, 1.547821e-08, 1.361951e-08, 1.175685e-08, 9.779572e-09, 
    7.867031e-09, 6.016306e-09, 4.1951e-09, 2.783738e-09, 1.874994e-09, 
    1.338976e-09, 1.054062e-09, 8.973933e-10, 7.909198e-10, 6.925031e-10,
  1.736077e-08, 1.604835e-08, 1.424625e-08, 1.240713e-08, 1.064454e-08, 
    8.941945e-09, 7.131962e-09, 5.198708e-09, 3.585132e-09, 2.428352e-09, 
    1.639761e-09, 1.212518e-09, 9.948387e-10, 8.595791e-10, 7.591879e-10,
  2.176251e-08, 2.107122e-08, 2.066751e-08, 2.005988e-08, 1.962374e-08, 
    1.803457e-08, 1.637056e-08, 1.446161e-08, 1.231491e-08, 9.907261e-09, 
    7.935767e-09, 6.723432e-09, 5.637386e-09, 4.456516e-09, 3.51723e-09,
  2.171778e-08, 2.091052e-08, 2.030044e-08, 1.951784e-08, 1.897507e-08, 
    1.740115e-08, 1.578575e-08, 1.396926e-08, 1.193958e-08, 9.687258e-09, 
    7.743381e-09, 6.486343e-09, 5.363241e-09, 4.229861e-09, 3.341578e-09,
  2.166491e-08, 2.069816e-08, 1.980801e-08, 1.900023e-08, 1.832488e-08, 
    1.681247e-08, 1.52365e-08, 1.342152e-08, 1.144129e-08, 9.341711e-09, 
    7.402529e-09, 6.122296e-09, 5.029202e-09, 3.966824e-09, 3.164347e-09,
  2.158088e-08, 2.053455e-08, 1.950179e-08, 1.865549e-08, 1.790644e-08, 
    1.634188e-08, 1.475757e-08, 1.294623e-08, 1.093717e-08, 8.917332e-09, 
    7.06651e-09, 5.763624e-09, 4.685935e-09, 3.696107e-09, 2.992181e-09,
  2.157504e-08, 2.039319e-08, 1.917724e-08, 1.833639e-08, 1.739574e-08, 
    1.583354e-08, 1.423351e-08, 1.230352e-08, 1.027833e-08, 8.421838e-09, 
    6.666356e-09, 5.347107e-09, 4.297496e-09, 3.431844e-09, 2.807929e-09,
  2.147299e-08, 2.012706e-08, 1.881313e-08, 1.786965e-08, 1.681927e-08, 
    1.524872e-08, 1.360616e-08, 1.150532e-08, 9.563204e-09, 7.869115e-09, 
    6.208823e-09, 4.872172e-09, 3.951947e-09, 3.181918e-09, 2.623429e-09,
  2.128284e-08, 1.982272e-08, 1.845388e-08, 1.738066e-08, 1.619796e-08, 
    1.451353e-08, 1.284198e-08, 1.057634e-08, 8.884435e-09, 7.359261e-09, 
    5.761412e-09, 4.465317e-09, 3.658482e-09, 2.973066e-09, 2.441935e-09,
  2.099651e-08, 1.946478e-08, 1.810185e-08, 1.692027e-08, 1.553464e-08, 
    1.372326e-08, 1.193623e-08, 9.720206e-09, 8.258444e-09, 6.858617e-09, 
    5.339415e-09, 4.130714e-09, 3.432779e-09, 2.781566e-09, 2.268288e-09,
  2.06599e-08, 1.918726e-08, 1.772228e-08, 1.648544e-08, 1.494733e-08, 
    1.275971e-08, 1.096857e-08, 8.928815e-09, 7.661598e-09, 6.408962e-09, 
    4.999478e-09, 3.924032e-09, 3.250769e-09, 2.583917e-09, 2.090612e-09,
  2.018405e-08, 1.875776e-08, 1.721885e-08, 1.599319e-08, 1.430379e-08, 
    1.172908e-08, 1.01305e-08, 8.264965e-09, 7.205532e-09, 6.096643e-09, 
    4.794793e-09, 3.760027e-09, 3.064452e-09, 2.392847e-09, 1.888801e-09,
  2.133732e-08, 2.121949e-08, 2.162931e-08, 2.194411e-08, 2.169631e-08, 
    2.070034e-08, 2.004865e-08, 1.93235e-08, 1.896771e-08, 1.819396e-08, 
    1.76191e-08, 1.706408e-08, 1.617271e-08, 1.516081e-08, 1.388693e-08,
  2.138751e-08, 2.162069e-08, 2.188692e-08, 2.267431e-08, 2.309185e-08, 
    2.265822e-08, 2.126947e-08, 2.003312e-08, 1.908646e-08, 1.826022e-08, 
    1.755642e-08, 1.743938e-08, 1.653941e-08, 1.552972e-08, 1.444652e-08,
  2.151191e-08, 2.173445e-08, 2.186673e-08, 2.241418e-08, 2.363866e-08, 
    2.388926e-08, 2.275316e-08, 2.112228e-08, 1.970158e-08, 1.886302e-08, 
    1.802433e-08, 1.74944e-08, 1.695391e-08, 1.585492e-08, 1.484942e-08,
  2.178551e-08, 2.199185e-08, 2.20986e-08, 2.228476e-08, 2.354377e-08, 
    2.452468e-08, 2.395922e-08, 2.241263e-08, 2.092678e-08, 1.974365e-08, 
    1.916862e-08, 1.819008e-08, 1.726852e-08, 1.622365e-08, 1.507991e-08,
  2.212733e-08, 2.227422e-08, 2.276117e-08, 2.270827e-08, 2.316048e-08, 
    2.441509e-08, 2.474505e-08, 2.404623e-08, 2.259857e-08, 2.058202e-08, 
    1.985625e-08, 1.926978e-08, 1.777899e-08, 1.636362e-08, 1.518923e-08,
  2.248796e-08, 2.257705e-08, 2.321856e-08, 2.349366e-08, 2.356391e-08, 
    2.412941e-08, 2.493246e-08, 2.522493e-08, 2.468297e-08, 2.233862e-08, 
    2.0656e-08, 1.966188e-08, 1.828813e-08, 1.647776e-08, 1.51692e-08,
  2.273222e-08, 2.299826e-08, 2.343585e-08, 2.404162e-08, 2.415207e-08, 
    2.433948e-08, 2.485431e-08, 2.571874e-08, 2.630741e-08, 2.401295e-08, 
    2.200638e-08, 2.045098e-08, 1.844636e-08, 1.658725e-08, 1.500776e-08,
  2.297437e-08, 2.33844e-08, 2.36627e-08, 2.424368e-08, 2.468445e-08, 
    2.489245e-08, 2.501414e-08, 2.53056e-08, 2.644995e-08, 2.462652e-08, 
    2.252283e-08, 2.112816e-08, 1.880507e-08, 1.656324e-08, 1.474223e-08,
  2.276149e-08, 2.369434e-08, 2.410319e-08, 2.427295e-08, 2.479379e-08, 
    2.505478e-08, 2.534451e-08, 2.49185e-08, 2.575888e-08, 2.457726e-08, 
    2.175556e-08, 2.0975e-08, 1.907866e-08, 1.645074e-08, 1.443568e-08,
  2.252836e-08, 2.356992e-08, 2.422546e-08, 2.444971e-08, 2.498834e-08, 
    2.516254e-08, 2.543523e-08, 2.449994e-08, 2.425909e-08, 2.346719e-08, 
    2.080563e-08, 1.953442e-08, 1.854927e-08, 1.60684e-08, 1.396428e-08,
  1.18502e-08, 1.090973e-08, 1.029592e-08, 9.621093e-09, 8.959014e-09, 
    8.490471e-09, 9.063577e-09, 9.924897e-09, 1.016368e-08, 9.495083e-09, 
    8.928475e-09, 8.714474e-09, 8.495063e-09, 8.212965e-09, 7.859604e-09,
  1.287769e-08, 1.184724e-08, 1.115385e-08, 1.047006e-08, 9.865097e-09, 
    8.999299e-09, 9.031695e-09, 9.903709e-09, 1.008333e-08, 1.015561e-08, 
    9.900445e-09, 9.617456e-09, 9.305123e-09, 9.047533e-09, 8.821316e-09,
  1.352962e-08, 1.303383e-08, 1.22989e-08, 1.161829e-08, 1.094573e-08, 
    1.004555e-08, 9.446231e-09, 9.880782e-09, 9.849249e-09, 9.982156e-09, 
    1.029623e-08, 1.05368e-08, 1.025482e-08, 9.825092e-09, 9.560834e-09,
  1.405592e-08, 1.391254e-08, 1.343596e-08, 1.282648e-08, 1.218762e-08, 
    1.155841e-08, 1.053704e-08, 1.033387e-08, 9.93998e-09, 1.017737e-08, 
    1.06966e-08, 1.128465e-08, 1.120868e-08, 1.086647e-08, 1.068773e-08,
  1.461328e-08, 1.444212e-08, 1.41742e-08, 1.381531e-08, 1.329908e-08, 
    1.295967e-08, 1.217609e-08, 1.146886e-08, 1.104829e-08, 1.05492e-08, 
    1.14037e-08, 1.197235e-08, 1.190471e-08, 1.195855e-08, 1.219096e-08,
  1.509821e-08, 1.479737e-08, 1.458774e-08, 1.445762e-08, 1.412395e-08, 
    1.387536e-08, 1.35364e-08, 1.300173e-08, 1.239858e-08, 1.156077e-08, 
    1.201225e-08, 1.265876e-08, 1.23871e-08, 1.28171e-08, 1.320961e-08,
  1.593266e-08, 1.54674e-08, 1.509544e-08, 1.487238e-08, 1.473039e-08, 
    1.44521e-08, 1.428391e-08, 1.391396e-08, 1.358571e-08, 1.281421e-08, 
    1.284917e-08, 1.346429e-08, 1.291832e-08, 1.358651e-08, 1.469509e-08,
  1.650789e-08, 1.610813e-08, 1.580862e-08, 1.566521e-08, 1.551686e-08, 
    1.532004e-08, 1.513502e-08, 1.497154e-08, 1.483263e-08, 1.443948e-08, 
    1.432093e-08, 1.47024e-08, 1.369525e-08, 1.441527e-08, 1.630266e-08,
  1.732639e-08, 1.669467e-08, 1.634583e-08, 1.629018e-08, 1.64086e-08, 
    1.633351e-08, 1.616194e-08, 1.622034e-08, 1.608454e-08, 1.594995e-08, 
    1.610074e-08, 1.659317e-08, 1.526549e-08, 1.590212e-08, 1.86391e-08,
  1.828725e-08, 1.78064e-08, 1.730364e-08, 1.690181e-08, 1.697198e-08, 
    1.717234e-08, 1.717639e-08, 1.722121e-08, 1.754291e-08, 1.735542e-08, 
    1.757884e-08, 1.825465e-08, 1.759299e-08, 1.815568e-08, 2.00239e-08,
  7.295664e-09, 6.501144e-09, 5.997294e-09, 5.460444e-09, 4.971884e-09, 
    4.50394e-09, 4.125399e-09, 3.891571e-09, 3.68605e-09, 3.523947e-09, 
    3.407866e-09, 3.313654e-09, 3.180151e-09, 2.988616e-09, 2.777425e-09,
  8.239607e-09, 7.263984e-09, 6.557764e-09, 6.092627e-09, 5.607937e-09, 
    5.152329e-09, 4.717984e-09, 4.358582e-09, 4.111155e-09, 3.979174e-09, 
    3.89141e-09, 3.79355e-09, 3.631097e-09, 3.457513e-09, 3.255216e-09,
  8.98123e-09, 8.182663e-09, 7.31765e-09, 6.770285e-09, 6.321236e-09, 
    5.822678e-09, 5.354273e-09, 4.966669e-09, 4.637419e-09, 4.427951e-09, 
    4.31318e-09, 4.193655e-09, 4.057298e-09, 3.913883e-09, 3.725968e-09,
  9.63423e-09, 8.941457e-09, 8.112065e-09, 7.457224e-09, 7.05435e-09, 
    6.607859e-09, 6.103551e-09, 5.652706e-09, 5.280838e-09, 5.002682e-09, 
    4.807117e-09, 4.673728e-09, 4.501568e-09, 4.324237e-09, 4.194342e-09,
  1.043335e-08, 9.660667e-09, 8.86759e-09, 8.116785e-09, 7.704865e-09, 
    7.330227e-09, 6.903755e-09, 6.513842e-09, 6.130094e-09, 5.825235e-09, 
    5.608502e-09, 5.395707e-09, 5.168588e-09, 4.961154e-09, 4.851466e-09,
  1.128496e-08, 1.042713e-08, 9.641504e-09, 8.828533e-09, 8.243701e-09, 
    7.838713e-09, 7.561811e-09, 7.270549e-09, 7.012189e-09, 6.694313e-09, 
    6.395579e-09, 6.134547e-09, 5.865759e-09, 5.695802e-09, 5.557285e-09,
  1.210656e-08, 1.122358e-08, 1.043488e-08, 9.595744e-09, 8.962812e-09, 
    8.305146e-09, 7.982038e-09, 7.82116e-09, 7.584998e-09, 7.357974e-09, 
    6.953183e-09, 6.686486e-09, 6.438572e-09, 6.279689e-09, 6.247497e-09,
  1.264831e-08, 1.201537e-08, 1.12189e-08, 1.044183e-08, 9.809161e-09, 
    9.167541e-09, 8.56735e-09, 8.257103e-09, 7.992818e-09, 7.679975e-09, 
    7.421008e-09, 7.131943e-09, 6.902015e-09, 6.777471e-09, 6.846369e-09,
  1.326004e-08, 1.25415e-08, 1.19218e-08, 1.120417e-08, 1.071431e-08, 
    1.013102e-08, 9.505908e-09, 8.9788e-09, 8.604538e-09, 8.259904e-09, 
    8.006681e-09, 7.741377e-09, 7.441006e-09, 7.253369e-09, 7.31504e-09,
  1.372565e-08, 1.311101e-08, 1.240568e-08, 1.177407e-08, 1.134378e-08, 
    1.089833e-08, 1.037228e-08, 9.81313e-09, 9.367064e-09, 9.048978e-09, 
    8.920916e-09, 8.668705e-09, 8.279172e-09, 7.903308e-09, 7.752512e-09,
  1.030325e-08, 9.479586e-09, 8.738438e-09, 8.119221e-09, 7.529135e-09, 
    7.005768e-09, 6.509927e-09, 5.862152e-09, 5.280753e-09, 4.766453e-09, 
    4.305027e-09, 3.896831e-09, 3.508481e-09, 3.178478e-09, 2.849471e-09,
  1.073758e-08, 9.902059e-09, 9.031655e-09, 8.350365e-09, 7.726438e-09, 
    7.243468e-09, 6.82815e-09, 6.301316e-09, 5.73278e-09, 5.230962e-09, 
    4.708251e-09, 4.246921e-09, 3.816529e-09, 3.472642e-09, 3.158226e-09,
  1.094329e-08, 1.042159e-08, 9.419821e-09, 8.628553e-09, 8.009719e-09, 
    7.457585e-09, 7.068266e-09, 6.668776e-09, 6.162091e-09, 5.648383e-09, 
    5.175913e-09, 4.695702e-09, 4.246142e-09, 3.808575e-09, 3.461362e-09,
  1.108531e-08, 1.076312e-08, 9.973713e-09, 9.096802e-09, 8.424851e-09, 
    7.812877e-09, 7.333637e-09, 6.966108e-09, 6.542086e-09, 6.060907e-09, 
    5.585966e-09, 5.132358e-09, 4.697996e-09, 4.252506e-09, 3.824392e-09,
  1.126791e-08, 1.104616e-08, 1.044001e-08, 9.628533e-09, 8.986692e-09, 
    8.297818e-09, 7.720783e-09, 7.306011e-09, 6.87972e-09, 6.45094e-09, 
    6.022408e-09, 5.573256e-09, 5.146636e-09, 4.715408e-09, 4.282773e-09,
  1.140733e-08, 1.122479e-08, 1.085585e-08, 9.998884e-09, 9.421805e-09, 
    8.89908e-09, 8.27059e-09, 7.718725e-09, 7.243109e-09, 6.817224e-09, 
    6.400441e-09, 6.007342e-09, 5.600671e-09, 5.198461e-09, 4.79746e-09,
  1.158894e-08, 1.120551e-08, 1.111854e-08, 1.036562e-08, 9.6838e-09, 
    9.230147e-09, 8.767274e-09, 8.282423e-09, 7.780724e-09, 7.294906e-09, 
    6.893623e-09, 6.480963e-09, 6.070031e-09, 5.674798e-09, 5.310352e-09,
  1.195063e-08, 1.127502e-08, 1.120325e-08, 1.070291e-08, 9.915061e-09, 
    9.51322e-09, 9.108883e-09, 8.701426e-09, 8.289266e-09, 7.888843e-09, 
    7.475328e-09, 7.06487e-09, 6.619973e-09, 6.186093e-09, 5.816559e-09,
  1.238713e-08, 1.153515e-08, 1.123381e-08, 1.093741e-08, 1.021298e-08, 
    9.73584e-09, 9.394329e-09, 9.060022e-09, 8.724657e-09, 8.367634e-09, 
    8.000497e-09, 7.617111e-09, 7.216018e-09, 6.776315e-09, 6.388319e-09,
  1.286168e-08, 1.189413e-08, 1.134945e-08, 1.109349e-08, 1.043796e-08, 
    9.988516e-09, 9.627911e-09, 9.352643e-09, 9.108911e-09, 8.795397e-09, 
    8.490856e-09, 8.176474e-09, 7.78163e-09, 7.381609e-09, 6.957321e-09,
  1.61189e-08, 1.495774e-08, 1.387513e-08, 1.29164e-08, 1.212006e-08, 
    1.129836e-08, 1.045117e-08, 9.423557e-09, 8.528567e-09, 7.831173e-09, 
    7.219828e-09, 6.667622e-09, 6.152671e-09, 5.561535e-09, 5.053609e-09,
  1.603105e-08, 1.511716e-08, 1.407656e-08, 1.304277e-08, 1.229281e-08, 
    1.15591e-08, 1.076161e-08, 9.872433e-09, 8.945644e-09, 8.1042e-09, 
    7.463955e-09, 6.888826e-09, 6.416967e-09, 5.902285e-09, 5.344027e-09,
  1.607081e-08, 1.526272e-08, 1.435184e-08, 1.322292e-08, 1.238791e-08, 
    1.171319e-08, 1.101089e-08, 1.021262e-08, 9.373298e-09, 8.449092e-09, 
    7.740445e-09, 7.124586e-09, 6.630587e-09, 6.203211e-09, 5.69972e-09,
  1.600535e-08, 1.528936e-08, 1.447379e-08, 1.345791e-08, 1.254207e-08, 
    1.179192e-08, 1.110035e-08, 1.045432e-08, 9.716497e-09, 8.867509e-09, 
    8.082833e-09, 7.410372e-09, 6.853323e-09, 6.420826e-09, 5.991482e-09,
  1.601222e-08, 1.527723e-08, 1.45053e-08, 1.357532e-08, 1.268311e-08, 
    1.191062e-08, 1.119466e-08, 1.056462e-08, 9.952149e-09, 9.26927e-09, 
    8.47754e-09, 7.782401e-09, 7.125511e-09, 6.650803e-09, 6.240784e-09,
  1.597377e-08, 1.525349e-08, 1.449781e-08, 1.366103e-08, 1.280078e-08, 
    1.203306e-08, 1.131489e-08, 1.071202e-08, 1.016389e-08, 9.568483e-09, 
    8.913613e-09, 8.190147e-09, 7.499115e-09, 6.908426e-09, 6.463643e-09,
  1.610342e-08, 1.529144e-08, 1.447229e-08, 1.367014e-08, 1.2847e-08, 
    1.212066e-08, 1.141106e-08, 1.080501e-08, 1.028196e-08, 9.775799e-09, 
    9.229005e-09, 8.583334e-09, 7.946357e-09, 7.333425e-09, 6.776828e-09,
  1.630574e-08, 1.53763e-08, 1.452985e-08, 1.364215e-08, 1.284898e-08, 
    1.213424e-08, 1.152692e-08, 1.093544e-08, 1.039423e-08, 9.938189e-09, 
    9.459934e-09, 8.916031e-09, 8.278154e-09, 7.733473e-09, 7.186045e-09,
  1.661476e-08, 1.548659e-08, 1.452315e-08, 1.363256e-08, 1.277968e-08, 
    1.210018e-08, 1.154625e-08, 1.104169e-08, 1.05096e-08, 1.004601e-08, 
    9.594249e-09, 9.132088e-09, 8.579006e-09, 8.038016e-09, 7.527467e-09,
  1.690071e-08, 1.569566e-08, 1.461641e-08, 1.364325e-08, 1.279112e-08, 
    1.209808e-08, 1.158313e-08, 1.10864e-08, 1.058938e-08, 1.016306e-08, 
    9.742539e-09, 9.359461e-09, 8.850694e-09, 8.301879e-09, 7.825603e-09,
  1.370037e-08, 1.282006e-08, 1.209674e-08, 1.13925e-08, 1.07837e-08, 
    1.016778e-08, 9.591518e-09, 8.922886e-09, 8.50968e-09, 7.926532e-09, 
    7.266774e-09, 6.749991e-09, 6.300414e-09, 5.716741e-09, 5.155704e-09,
  1.416457e-08, 1.336315e-08, 1.266756e-08, 1.194945e-08, 1.129817e-08, 
    1.068084e-08, 1.017836e-08, 9.530251e-09, 9.016868e-09, 8.564207e-09, 
    7.995845e-09, 7.420377e-09, 6.917545e-09, 6.429559e-09, 5.960207e-09,
  1.462516e-08, 1.388434e-08, 1.319514e-08, 1.259762e-08, 1.196206e-08, 
    1.128338e-08, 1.07425e-08, 1.016654e-08, 9.598514e-09, 9.136155e-09, 
    8.62062e-09, 8.052933e-09, 7.517762e-09, 7.002089e-09, 6.528168e-09,
  1.501656e-08, 1.435654e-08, 1.365463e-08, 1.305818e-08, 1.251788e-08, 
    1.19041e-08, 1.132726e-08, 1.072234e-08, 1.015522e-08, 9.615589e-09, 
    9.145132e-09, 8.584499e-09, 8.041442e-09, 7.52809e-09, 7.082565e-09,
  1.531806e-08, 1.470893e-08, 1.408272e-08, 1.347946e-08, 1.295151e-08, 
    1.239164e-08, 1.188376e-08, 1.135548e-08, 1.076806e-08, 1.023226e-08, 
    9.683687e-09, 9.159414e-09, 8.6557e-09, 8.147842e-09, 7.679095e-09,
  1.552073e-08, 1.50279e-08, 1.446086e-08, 1.383046e-08, 1.333079e-08, 
    1.278619e-08, 1.230035e-08, 1.183105e-08, 1.133632e-08, 1.077514e-08, 
    1.026082e-08, 9.718738e-09, 9.20863e-09, 8.735962e-09, 8.284643e-09,
  1.578626e-08, 1.522994e-08, 1.479131e-08, 1.421343e-08, 1.366327e-08, 
    1.315568e-08, 1.269192e-08, 1.224353e-08, 1.179113e-08, 1.13081e-08, 
    1.077769e-08, 1.026225e-08, 9.744955e-09, 9.239624e-09, 8.772966e-09,
  1.595556e-08, 1.546273e-08, 1.493182e-08, 1.44158e-08, 1.391876e-08, 
    1.345069e-08, 1.298873e-08, 1.258906e-08, 1.218519e-08, 1.174385e-08, 
    1.126664e-08, 1.078776e-08, 1.027663e-08, 9.765356e-09, 9.28237e-09,
  1.614624e-08, 1.559913e-08, 1.516289e-08, 1.459842e-08, 1.405549e-08, 
    1.359446e-08, 1.316653e-08, 1.27606e-08, 1.24087e-08, 1.201869e-08, 
    1.158626e-08, 1.113112e-08, 1.070976e-08, 1.022225e-08, 9.763862e-09,
  1.62829e-08, 1.579365e-08, 1.52004e-08, 1.478812e-08, 1.421234e-08, 
    1.368835e-08, 1.325525e-08, 1.286595e-08, 1.247688e-08, 1.213369e-08, 
    1.177533e-08, 1.136269e-08, 1.097942e-08, 1.057983e-08, 1.014075e-08,
  6.095002e-09, 4.972759e-09, 4.19625e-09, 3.441462e-09, 2.837511e-09, 
    2.369859e-09, 1.948114e-09, 1.638279e-09, 1.469808e-09, 1.393246e-09, 
    1.359545e-09, 1.329976e-09, 1.288075e-09, 1.224292e-09, 1.16191e-09,
  7.14071e-09, 5.908061e-09, 4.971272e-09, 4.209823e-09, 3.50818e-09, 
    2.978874e-09, 2.514045e-09, 2.089189e-09, 1.773382e-09, 1.562167e-09, 
    1.451335e-09, 1.394117e-09, 1.375094e-09, 1.359056e-09, 1.331528e-09,
  8.415896e-09, 6.975433e-09, 5.865224e-09, 4.970728e-09, 4.237306e-09, 
    3.64986e-09, 3.133221e-09, 2.665828e-09, 2.257997e-09, 1.920484e-09, 
    1.699398e-09, 1.556865e-09, 1.481464e-09, 1.440499e-09, 1.422183e-09,
  9.675848e-09, 8.229883e-09, 6.920108e-09, 5.855784e-09, 5.017034e-09, 
    4.360456e-09, 3.815276e-09, 3.315055e-09, 2.876445e-09, 2.474056e-09, 
    2.140107e-09, 1.891674e-09, 1.731505e-09, 1.63285e-09, 1.574277e-09,
  1.074051e-08, 9.422982e-09, 8.139361e-09, 6.903152e-09, 5.922498e-09, 
    5.182919e-09, 4.574627e-09, 4.032779e-09, 3.548759e-09, 3.111509e-09, 
    2.728334e-09, 2.392804e-09, 2.114812e-09, 1.931574e-09, 1.811981e-09,
  1.159571e-08, 1.038008e-08, 9.163799e-09, 7.960555e-09, 6.858666e-09, 
    6.026075e-09, 5.382408e-09, 4.84347e-09, 4.37013e-09, 3.919421e-09, 
    3.500264e-09, 3.119103e-09, 2.762485e-09, 2.464907e-09, 2.242916e-09,
  1.229921e-08, 1.120157e-08, 1.006887e-08, 8.923606e-09, 7.8676e-09, 
    6.923973e-09, 6.166707e-09, 5.581879e-09, 5.105184e-09, 4.697017e-09, 
    4.308033e-09, 3.947457e-09, 3.604501e-09, 3.281915e-09, 2.997502e-09,
  1.291281e-08, 1.194936e-08, 1.097582e-08, 9.915499e-09, 8.92036e-09, 
    7.997261e-09, 7.146831e-09, 6.438056e-09, 5.879615e-09, 5.43205e-09, 
    5.061916e-09, 4.730671e-09, 4.441105e-09, 4.158139e-09, 3.882932e-09,
  1.347057e-08, 1.262196e-08, 1.180633e-08, 1.090686e-08, 9.976445e-09, 
    9.093908e-09, 8.259287e-09, 7.515212e-09, 6.878585e-09, 6.361486e-09, 
    5.947708e-09, 5.609551e-09, 5.306903e-09, 5.035069e-09, 4.792336e-09,
  1.389696e-08, 1.318927e-08, 1.245769e-08, 1.171116e-08, 1.091383e-08, 
    1.012497e-08, 9.356802e-09, 8.626278e-09, 7.982273e-09, 7.428617e-09, 
    6.974541e-09, 6.600075e-09, 6.290854e-09, 6.016965e-09, 5.764205e-09,
  2.371746e-09, 2.083952e-09, 1.907391e-09, 1.784377e-09, 1.686111e-09, 
    1.560146e-09, 1.401786e-09, 1.246332e-09, 1.064911e-09, 8.808566e-10, 
    7.400891e-10, 6.369703e-10, 5.823503e-10, 5.463089e-10, 5.183402e-10,
  2.660441e-09, 2.336119e-09, 2.072797e-09, 1.878353e-09, 1.753934e-09, 
    1.67856e-09, 1.573757e-09, 1.407263e-09, 1.211683e-09, 1.037233e-09, 
    8.898671e-10, 7.619754e-10, 6.686121e-10, 6.067578e-10, 5.621038e-10,
  3.12435e-09, 2.598519e-09, 2.253874e-09, 2.017989e-09, 1.846086e-09, 
    1.744643e-09, 1.691776e-09, 1.549088e-09, 1.356966e-09, 1.204073e-09, 
    1.054971e-09, 9.108667e-10, 7.877513e-10, 6.872089e-10, 6.176019e-10,
  3.939985e-09, 3.060599e-09, 2.547209e-09, 2.195098e-09, 1.995066e-09, 
    1.857387e-09, 1.788771e-09, 1.683692e-09, 1.499325e-09, 1.355472e-09, 
    1.222307e-09, 1.072946e-09, 9.287374e-10, 8.007159e-10, 7.02666e-10,
  5.03407e-09, 3.828446e-09, 3.003803e-09, 2.492079e-09, 2.188245e-09, 
    1.998927e-09, 1.911241e-09, 1.807874e-09, 1.661678e-09, 1.51994e-09, 
    1.388402e-09, 1.245949e-09, 1.093784e-09, 9.556583e-10, 8.339422e-10,
  6.229841e-09, 4.834641e-09, 3.770008e-09, 2.99377e-09, 2.518733e-09, 
    2.210381e-09, 2.068278e-09, 1.917336e-09, 1.780769e-09, 1.671407e-09, 
    1.556225e-09, 1.437027e-09, 1.296705e-09, 1.155349e-09, 1.013575e-09,
  7.639761e-09, 6.008702e-09, 4.700943e-09, 3.75822e-09, 3.012906e-09, 
    2.566263e-09, 2.315016e-09, 2.109473e-09, 1.90182e-09, 1.79692e-09, 
    1.691606e-09, 1.584748e-09, 1.464573e-09, 1.337774e-09, 1.204112e-09,
  9.090425e-09, 7.370395e-09, 5.878274e-09, 4.691429e-09, 3.748469e-09, 
    3.039893e-09, 2.632788e-09, 2.373875e-09, 2.098347e-09, 1.947784e-09, 
    1.860706e-09, 1.770087e-09, 1.671262e-09, 1.558256e-09, 1.433084e-09,
  1.078505e-08, 8.740518e-09, 7.184102e-09, 5.815251e-09, 4.653217e-09, 
    3.725134e-09, 3.096877e-09, 2.691609e-09, 2.326897e-09, 2.089615e-09, 
    1.955575e-09, 1.865982e-09, 1.793776e-09, 1.730164e-09, 1.653017e-09,
  1.259951e-08, 1.036668e-08, 8.609698e-09, 7.117098e-09, 5.79285e-09, 
    4.583773e-09, 3.734894e-09, 3.191244e-09, 2.740353e-09, 2.391325e-09, 
    2.150499e-09, 1.996238e-09, 1.8841e-09, 1.818153e-09, 1.769775e-09,
  3.732414e-09, 2.90976e-09, 2.578159e-09, 2.277545e-09, 1.987815e-09, 
    1.777141e-09, 1.602472e-09, 1.423437e-09, 1.278172e-09, 1.159161e-09, 
    1.088002e-09, 1.030205e-09, 9.806645e-10, 9.653555e-10, 9.627675e-10,
  4.317857e-09, 3.201416e-09, 2.691836e-09, 2.366789e-09, 2.014422e-09, 
    1.837986e-09, 1.686834e-09, 1.506601e-09, 1.352588e-09, 1.226863e-09, 
    1.158552e-09, 1.101071e-09, 1.045119e-09, 1.006725e-09, 9.964111e-10,
  5.081979e-09, 3.728801e-09, 2.977696e-09, 2.511728e-09, 2.05418e-09, 
    1.876983e-09, 1.768914e-09, 1.609231e-09, 1.46025e-09, 1.317531e-09, 
    1.224603e-09, 1.175562e-09, 1.126908e-09, 1.078453e-09, 1.039946e-09,
  5.715919e-09, 4.36042e-09, 3.362948e-09, 2.751825e-09, 2.211211e-09, 
    1.949803e-09, 1.840562e-09, 1.699429e-09, 1.544364e-09, 1.430488e-09, 
    1.307937e-09, 1.22973e-09, 1.206297e-09, 1.174871e-09, 1.131934e-09,
  6.130626e-09, 4.897512e-09, 3.857042e-09, 3.08132e-09, 2.433989e-09, 
    2.061441e-09, 1.919239e-09, 1.771172e-09, 1.62412e-09, 1.515139e-09, 
    1.431359e-09, 1.321172e-09, 1.26074e-09, 1.24633e-09, 1.226982e-09,
  6.400679e-09, 5.36473e-09, 4.367986e-09, 3.58403e-09, 2.756574e-09, 
    2.240678e-09, 2.035277e-09, 1.871941e-09, 1.716854e-09, 1.605567e-09, 
    1.525724e-09, 1.46777e-09, 1.386325e-09, 1.332394e-09, 1.308111e-09,
  6.75755e-09, 5.781021e-09, 4.905229e-09, 4.113191e-09, 3.263537e-09, 
    2.522508e-09, 2.244263e-09, 2.043935e-09, 1.867008e-09, 1.730431e-09, 
    1.626396e-09, 1.553631e-09, 1.499167e-09, 1.444289e-09, 1.400222e-09,
  7.221807e-09, 6.29846e-09, 5.435574e-09, 4.653669e-09, 3.800463e-09, 
    2.993985e-09, 2.500385e-09, 2.232541e-09, 2.029899e-09, 1.871732e-09, 
    1.740411e-09, 1.653728e-09, 1.580676e-09, 1.530207e-09, 1.493327e-09,
  7.779036e-09, 6.852979e-09, 6.012306e-09, 5.18785e-09, 4.328804e-09, 
    3.453971e-09, 2.857196e-09, 2.439188e-09, 2.176387e-09, 1.991491e-09, 
    1.841007e-09, 1.725221e-09, 1.641262e-09, 1.582495e-09, 1.546008e-09,
  8.446649e-09, 7.455961e-09, 6.571839e-09, 5.783213e-09, 4.882918e-09, 
    3.964949e-09, 3.235419e-09, 2.730402e-09, 2.369477e-09, 2.127864e-09, 
    1.94626e-09, 1.806058e-09, 1.711369e-09, 1.64866e-09, 1.623329e-09,
  1.386882e-08, 1.226127e-08, 1.080304e-08, 9.172409e-09, 7.488386e-09, 
    5.788152e-09, 4.531019e-09, 3.475453e-09, 2.723489e-09, 2.234944e-09, 
    1.88548e-09, 1.69797e-09, 1.455257e-09, 1.204865e-09, 1.006995e-09,
  1.38923e-08, 1.262094e-08, 1.127755e-08, 9.78291e-09, 8.151735e-09, 
    6.449168e-09, 5.068642e-09, 3.920257e-09, 3.044305e-09, 2.448614e-09, 
    2.010828e-09, 1.756451e-09, 1.549733e-09, 1.338474e-09, 1.111506e-09,
  1.387486e-08, 1.281911e-08, 1.159204e-08, 1.01538e-08, 8.697269e-09, 
    7.075597e-09, 5.582855e-09, 4.352147e-09, 3.388771e-09, 2.70301e-09, 
    2.215709e-09, 1.883611e-09, 1.65195e-09, 1.452429e-09, 1.239206e-09,
  1.386999e-08, 1.295488e-08, 1.184403e-08, 1.043984e-08, 9.118638e-09, 
    7.638431e-09, 6.1328e-09, 4.762451e-09, 3.783204e-09, 2.988787e-09, 
    2.457134e-09, 2.054844e-09, 1.783949e-09, 1.561079e-09, 1.361252e-09,
  1.390308e-08, 1.304107e-08, 1.201431e-08, 1.064379e-08, 9.431813e-09, 
    8.102204e-09, 6.663307e-09, 5.163874e-09, 4.140314e-09, 3.310005e-09, 
    2.696183e-09, 2.258091e-09, 1.921818e-09, 1.685346e-09, 1.477991e-09,
  1.391711e-08, 1.306879e-08, 1.210539e-08, 1.082598e-08, 9.618375e-09, 
    8.438002e-09, 7.097678e-09, 5.622754e-09, 4.489419e-09, 3.636797e-09, 
    2.933066e-09, 2.469078e-09, 2.098586e-09, 1.812131e-09, 1.600879e-09,
  1.378958e-08, 1.298965e-08, 1.209741e-08, 1.093379e-08, 9.720262e-09, 
    8.615709e-09, 7.404434e-09, 6.057727e-09, 4.837005e-09, 3.974711e-09, 
    3.205041e-09, 2.66205e-09, 2.280309e-09, 1.953657e-09, 1.719123e-09,
  1.358383e-08, 1.280033e-08, 1.196825e-08, 1.092061e-08, 9.734733e-09, 
    8.68723e-09, 7.591043e-09, 6.373774e-09, 5.165855e-09, 4.255481e-09, 
    3.479742e-09, 2.866989e-09, 2.44986e-09, 2.118209e-09, 1.84173e-09,
  1.326947e-08, 1.250263e-08, 1.173217e-08, 1.082496e-08, 9.713943e-09, 
    8.694432e-09, 7.680705e-09, 6.584144e-09, 5.434942e-09, 4.509761e-09, 
    3.73096e-09, 3.082794e-09, 2.628095e-09, 2.289243e-09, 1.99098e-09,
  1.301526e-08, 1.221011e-08, 1.149124e-08, 1.064245e-08, 9.684286e-09, 
    8.695619e-09, 7.69991e-09, 6.710944e-09, 5.645681e-09, 4.714106e-09, 
    3.975897e-09, 3.299562e-09, 2.813178e-09, 2.444408e-09, 2.125758e-09,
  9.227585e-09, 7.591005e-09, 6.081587e-09, 4.803276e-09, 3.748959e-09, 
    2.811291e-09, 2.10254e-09, 1.687431e-09, 1.414737e-09, 1.223531e-09, 
    1.064287e-09, 9.166686e-10, 7.62778e-10, 6.197787e-10, 5.206359e-10,
  1.032643e-08, 8.66597e-09, 7.235526e-09, 5.883073e-09, 4.609213e-09, 
    3.477784e-09, 2.543444e-09, 1.950083e-09, 1.585699e-09, 1.32889e-09, 
    1.174223e-09, 1.033408e-09, 8.910001e-10, 7.50154e-10, 6.189987e-10,
  1.194245e-08, 9.92139e-09, 8.258252e-09, 6.872067e-09, 5.579199e-09, 
    4.327898e-09, 3.174761e-09, 2.312504e-09, 1.824107e-09, 1.470307e-09, 
    1.281416e-09, 1.141407e-09, 1.017289e-09, 8.833663e-10, 7.513117e-10,
  1.342562e-08, 1.144482e-08, 9.476396e-09, 7.904024e-09, 6.594021e-09, 
    5.257277e-09, 3.979233e-09, 2.848011e-09, 2.14944e-09, 1.691707e-09, 
    1.416702e-09, 1.255519e-09, 1.143305e-09, 1.01088e-09, 8.929271e-10,
  1.46262e-08, 1.284988e-08, 1.088368e-08, 9.05735e-09, 7.640645e-09, 
    6.302843e-09, 4.922602e-09, 3.598524e-09, 2.59326e-09, 1.982958e-09, 
    1.611128e-09, 1.378464e-09, 1.236347e-09, 1.112762e-09, 1.000784e-09,
  1.559198e-08, 1.419135e-08, 1.225278e-08, 1.036173e-08, 8.698834e-09, 
    7.320742e-09, 5.935733e-09, 4.487235e-09, 3.234202e-09, 2.373519e-09, 
    1.869316e-09, 1.555259e-09, 1.354003e-09, 1.203548e-09, 1.099648e-09,
  1.614882e-08, 1.522596e-08, 1.357008e-08, 1.164899e-08, 9.926453e-09, 
    8.371563e-09, 6.975282e-09, 5.51281e-09, 4.041879e-09, 2.904096e-09, 
    2.190255e-09, 1.778541e-09, 1.513803e-09, 1.329717e-09, 1.193105e-09,
  1.681037e-08, 1.600947e-08, 1.472343e-08, 1.296018e-08, 1.115095e-08, 
    9.512941e-09, 8.048565e-09, 6.555722e-09, 4.994092e-09, 3.627767e-09, 
    2.626885e-09, 2.066408e-09, 1.725986e-09, 1.493888e-09, 1.329241e-09,
  1.745545e-08, 1.680239e-08, 1.574395e-08, 1.4157e-08, 1.244921e-08, 
    1.071782e-08, 9.153802e-09, 7.652341e-09, 5.998417e-09, 4.486707e-09, 
    3.24104e-09, 2.44635e-09, 1.991882e-09, 1.693552e-09, 1.469722e-09,
  1.802232e-08, 1.748606e-08, 1.666691e-08, 1.52726e-08, 1.366502e-08, 
    1.195671e-08, 1.030071e-08, 8.763045e-09, 7.089731e-09, 5.419685e-09, 
    4.03476e-09, 2.954021e-09, 2.311758e-09, 1.923218e-09, 1.648635e-09,
  1.46488e-08, 1.20839e-08, 1.009124e-08, 7.876231e-09, 5.793638e-09, 
    4.166159e-09, 2.957889e-09, 1.972072e-09, 1.303689e-09, 9.715427e-10, 
    7.357965e-10, 5.767586e-10, 5.207442e-10, 4.823438e-10, 4.51611e-10,
  1.438687e-08, 1.163778e-08, 9.711592e-09, 7.583052e-09, 5.558936e-09, 
    3.964906e-09, 2.783641e-09, 1.80548e-09, 1.190652e-09, 8.949599e-10, 
    6.711347e-10, 5.324088e-10, 4.91527e-10, 4.653072e-10, 4.377845e-10,
  1.395235e-08, 1.109199e-08, 9.235389e-09, 7.139751e-09, 5.223192e-09, 
    3.718845e-09, 2.569155e-09, 1.638887e-09, 1.092739e-09, 8.25217e-10, 
    6.167236e-10, 5.028101e-10, 4.757236e-10, 4.55977e-10, 4.338312e-10,
  1.368902e-08, 1.077734e-08, 8.932844e-09, 6.861358e-09, 5.0612e-09, 
    3.60031e-09, 2.46722e-09, 1.56286e-09, 1.041465e-09, 7.690814e-10, 
    5.657612e-10, 4.773762e-10, 4.672228e-10, 4.547374e-10, 4.352904e-10,
  1.354296e-08, 1.057863e-08, 8.649592e-09, 6.561692e-09, 4.874623e-09, 
    3.512134e-09, 2.403727e-09, 1.510192e-09, 9.921808e-10, 7.095181e-10, 
    5.18278e-10, 4.484064e-10, 4.561868e-10, 4.526994e-10, 4.357151e-10,
  1.34284e-08, 1.042472e-08, 8.343049e-09, 6.206157e-09, 4.652509e-09, 
    3.431937e-09, 2.350527e-09, 1.460405e-09, 9.440554e-10, 6.625329e-10, 
    4.852272e-10, 4.272276e-10, 4.43881e-10, 4.455772e-10, 4.292397e-10,
  1.344238e-08, 1.031501e-08, 8.09099e-09, 5.867103e-09, 4.425122e-09, 
    3.356773e-09, 2.326276e-09, 1.430025e-09, 9.144007e-10, 6.379272e-10, 
    4.71472e-10, 4.220721e-10, 4.315005e-10, 4.295565e-10, 4.142806e-10,
  1.347992e-08, 1.035181e-08, 7.955284e-09, 5.593173e-09, 4.212035e-09, 
    3.289188e-09, 2.312386e-09, 1.417811e-09, 9.013256e-10, 6.37102e-10, 
    4.743749e-10, 4.243382e-10, 4.197387e-10, 4.109593e-10, 3.969686e-10,
  1.349606e-08, 1.048197e-08, 7.978533e-09, 5.447049e-09, 4.040361e-09, 
    3.225472e-09, 2.325272e-09, 1.449838e-09, 9.251467e-10, 6.486304e-10, 
    4.836698e-10, 4.322706e-10, 4.132782e-10, 3.958619e-10, 3.840404e-10,
  1.349489e-08, 1.067235e-08, 8.126376e-09, 5.443939e-09, 3.943253e-09, 
    3.194513e-09, 2.376426e-09, 1.520787e-09, 9.731017e-10, 6.727692e-10, 
    4.994809e-10, 4.417905e-10, 4.149012e-10, 3.938896e-10, 3.807553e-10,
  2.326914e-08, 2.338646e-08, 2.30362e-08, 2.226488e-08, 2.105798e-08, 
    1.980375e-08, 1.847134e-08, 1.734044e-08, 1.588194e-08, 1.42798e-08, 
    1.279685e-08, 1.151492e-08, 1.024987e-08, 9.084875e-09, 7.992342e-09,
  2.354735e-08, 2.345722e-08, 2.315488e-08, 2.242506e-08, 2.13239e-08, 
    1.982215e-08, 1.83927e-08, 1.734048e-08, 1.585855e-08, 1.431035e-08, 
    1.282331e-08, 1.148183e-08, 1.021196e-08, 9.043397e-09, 7.933113e-09,
  2.374968e-08, 2.344473e-08, 2.31724e-08, 2.251178e-08, 2.149785e-08, 
    1.986504e-08, 1.831724e-08, 1.722852e-08, 1.565911e-08, 1.408232e-08, 
    1.26771e-08, 1.133619e-08, 1.006991e-08, 8.930702e-09, 7.808138e-09,
  2.381111e-08, 2.363813e-08, 2.318355e-08, 2.255108e-08, 2.166323e-08, 
    1.989204e-08, 1.813686e-08, 1.703253e-08, 1.540831e-08, 1.381839e-08, 
    1.244782e-08, 1.108345e-08, 9.822918e-09, 8.698304e-09, 7.584064e-09,
  2.39694e-08, 2.382447e-08, 2.329991e-08, 2.256636e-08, 2.17269e-08, 
    1.986318e-08, 1.789764e-08, 1.670663e-08, 1.512237e-08, 1.349825e-08, 
    1.218982e-08, 1.083672e-08, 9.57006e-09, 8.412435e-09, 7.284696e-09,
  2.413025e-08, 2.390078e-08, 2.338048e-08, 2.265138e-08, 2.177415e-08, 
    1.985163e-08, 1.77207e-08, 1.643074e-08, 1.484901e-08, 1.31364e-08, 
    1.189084e-08, 1.059963e-08, 9.290458e-09, 8.08396e-09, 6.922978e-09,
  2.414405e-08, 2.393563e-08, 2.33539e-08, 2.264807e-08, 2.175054e-08, 
    1.981345e-08, 1.754193e-08, 1.615561e-08, 1.456984e-08, 1.27908e-08, 
    1.160483e-08, 1.034848e-08, 8.998198e-09, 7.707389e-09, 6.512571e-09,
  2.405772e-08, 2.377593e-08, 2.322108e-08, 2.255276e-08, 2.159357e-08, 
    1.966759e-08, 1.726585e-08, 1.586097e-08, 1.428028e-08, 1.246974e-08, 
    1.123159e-08, 1.002983e-08, 8.626428e-09, 7.293669e-09, 6.086077e-09,
  2.394156e-08, 2.354871e-08, 2.294509e-08, 2.229709e-08, 2.136225e-08, 
    1.94496e-08, 1.701965e-08, 1.550975e-08, 1.401209e-08, 1.219347e-08, 
    1.083068e-08, 9.635567e-09, 8.21265e-09, 6.857638e-09, 5.657323e-09,
  2.378814e-08, 2.330799e-08, 2.263491e-08, 2.191591e-08, 2.098436e-08, 
    1.911202e-08, 1.673585e-08, 1.521275e-08, 1.368729e-08, 1.190133e-08, 
    1.036697e-08, 9.183533e-09, 7.772625e-09, 6.432143e-09, 5.228177e-09,
  1.712162e-08, 1.541291e-08, 1.364595e-08, 1.143423e-08, 1.016461e-08, 
    8.924314e-09, 7.453454e-09, 6.391951e-09, 5.689095e-09, 4.906139e-09, 
    4.41776e-09, 4.171477e-09, 3.964794e-09, 3.632949e-09, 3.136504e-09,
  1.808175e-08, 1.676448e-08, 1.53486e-08, 1.348278e-08, 1.146928e-08, 
    1.006944e-08, 8.906642e-09, 7.713624e-09, 6.683281e-09, 6.006545e-09, 
    5.390377e-09, 4.841922e-09, 4.513844e-09, 4.261018e-09, 3.889415e-09,
  1.928545e-08, 1.784385e-08, 1.653044e-08, 1.504445e-08, 1.326076e-08, 
    1.140593e-08, 9.99027e-09, 8.94033e-09, 7.973795e-09, 7.047592e-09, 
    6.447567e-09, 5.877806e-09, 5.341061e-09, 4.930767e-09, 4.543717e-09,
  2.011455e-08, 1.888141e-08, 1.755415e-08, 1.632157e-08, 1.47936e-08, 
    1.324806e-08, 1.150006e-08, 1.012602e-08, 9.210775e-09, 8.393696e-09, 
    7.537638e-09, 6.93391e-09, 6.400862e-09, 5.856577e-09, 5.32572e-09,
  2.047422e-08, 1.952773e-08, 1.838843e-08, 1.724801e-08, 1.599829e-08, 
    1.460363e-08, 1.319346e-08, 1.16103e-08, 1.03583e-08, 9.550462e-09, 
    8.821957e-09, 8.013687e-09, 7.384152e-09, 6.850823e-09, 6.246175e-09,
  2.06343e-08, 1.989646e-08, 1.895935e-08, 1.797443e-08, 1.692767e-08, 
    1.573185e-08, 1.453402e-08, 1.316669e-08, 1.172111e-08, 1.063228e-08, 
    9.882752e-09, 9.253729e-09, 8.421812e-09, 7.775447e-09, 7.200685e-09,
  2.088137e-08, 2.014591e-08, 1.94523e-08, 1.859031e-08, 1.762106e-08, 
    1.662623e-08, 1.558939e-08, 1.452632e-08, 1.321194e-08, 1.188763e-08, 
    1.091763e-08, 1.026885e-08, 9.587834e-09, 8.824712e-09, 8.100964e-09,
  2.116287e-08, 2.052251e-08, 1.985528e-08, 1.909369e-08, 1.828721e-08, 
    1.736333e-08, 1.644965e-08, 1.550797e-08, 1.45322e-08, 1.330231e-08, 
    1.209415e-08, 1.121022e-08, 1.049746e-08, 9.879819e-09, 9.198081e-09,
  2.133365e-08, 2.078546e-08, 2.016529e-08, 1.951409e-08, 1.875231e-08, 
    1.798795e-08, 1.721751e-08, 1.635411e-08, 1.550519e-08, 1.45833e-08, 
    1.343856e-08, 1.231904e-08, 1.140657e-08, 1.071496e-08, 1.009272e-08,
  2.156157e-08, 2.103632e-08, 2.042833e-08, 1.984162e-08, 1.915745e-08, 
    1.841163e-08, 1.779042e-08, 1.704453e-08, 1.631341e-08, 1.552129e-08, 
    1.465279e-08, 1.34983e-08, 1.24115e-08, 1.15533e-08, 1.086609e-08,
  8.654376e-09, 5.631123e-09, 4.255833e-09, 3.544148e-09, 2.949968e-09, 
    2.37434e-09, 1.983629e-09, 1.627962e-09, 1.422317e-09, 1.248018e-09, 
    1.094324e-09, 1.007615e-09, 9.329963e-10, 7.789395e-10, 6.158309e-10,
  9.939779e-09, 7.174702e-09, 5.292508e-09, 4.018143e-09, 3.473851e-09, 
    2.790745e-09, 2.147433e-09, 1.798974e-09, 1.526373e-09, 1.375305e-09, 
    1.228681e-09, 1.082597e-09, 9.832217e-10, 9.157714e-10, 7.429579e-10,
  1.141549e-08, 8.639593e-09, 6.597606e-09, 4.886366e-09, 3.860626e-09, 
    3.296375e-09, 2.606054e-09, 2.043079e-09, 1.718821e-09, 1.506865e-09, 
    1.36733e-09, 1.225887e-09, 1.078533e-09, 9.712564e-10, 8.797963e-10,
  1.275904e-08, 1.021115e-08, 7.830798e-09, 6.011596e-09, 4.61153e-09, 
    3.721623e-09, 3.17576e-09, 2.540429e-09, 1.952122e-09, 1.687272e-09, 
    1.507572e-09, 1.367594e-09, 1.222648e-09, 1.091712e-09, 9.767878e-10,
  1.395855e-08, 1.164919e-08, 9.12795e-09, 7.14405e-09, 5.6439e-09, 
    4.412084e-09, 3.644947e-09, 3.084657e-09, 2.408879e-09, 1.932299e-09, 
    1.690462e-09, 1.51569e-09, 1.366114e-09, 1.250739e-09, 1.119781e-09,
  1.508638e-08, 1.29551e-08, 1.049287e-08, 8.23821e-09, 6.707898e-09, 
    5.389253e-09, 4.341456e-09, 3.548266e-09, 2.943768e-09, 2.366558e-09, 
    1.972185e-09, 1.7101e-09, 1.531492e-09, 1.392258e-09, 1.291132e-09,
  1.60679e-08, 1.40989e-08, 1.187624e-08, 9.527494e-09, 7.704365e-09, 
    6.395621e-09, 5.240666e-09, 4.236361e-09, 3.48432e-09, 2.892451e-09, 
    2.410045e-09, 2.011775e-09, 1.737036e-09, 1.566378e-09, 1.439567e-09,
  1.693395e-08, 1.508722e-08, 1.320203e-08, 1.085728e-08, 8.832395e-09, 
    7.411973e-09, 6.166125e-09, 5.151698e-09, 4.195887e-09, 3.464889e-09, 
    2.915584e-09, 2.447646e-09, 2.037984e-09, 1.773656e-09, 1.61408e-09,
  1.77107e-08, 1.599884e-08, 1.434332e-08, 1.22386e-08, 1.010747e-08, 
    8.46072e-09, 7.144245e-09, 6.053682e-09, 5.114256e-09, 4.183337e-09, 
    3.469176e-09, 2.934508e-09, 2.487011e-09, 2.081161e-09, 1.831057e-09,
  1.833404e-08, 1.677892e-08, 1.531385e-08, 1.353744e-08, 1.144087e-08, 
    9.566774e-09, 8.166838e-09, 6.95401e-09, 6.015262e-09, 5.095554e-09, 
    4.18553e-09, 3.462689e-09, 2.973456e-09, 2.556474e-09, 2.162525e-09,
  1.555565e-08, 1.108875e-08, 8.164373e-09, 5.461257e-09, 3.988956e-09, 
    2.899019e-09, 2.380457e-09, 1.962515e-09, 1.626564e-09, 1.352159e-09, 
    1.08526e-09, 8.866929e-10, 8.113855e-10, 7.825582e-10, 7.225953e-10,
  1.530379e-08, 1.145064e-08, 8.342352e-09, 5.656216e-09, 4.114221e-09, 
    3.067519e-09, 2.443884e-09, 1.965595e-09, 1.638796e-09, 1.39334e-09, 
    1.144058e-09, 9.418382e-10, 8.513864e-10, 8.174716e-10, 7.714331e-10,
  1.51695e-08, 1.167925e-08, 8.433068e-09, 5.773369e-09, 4.238661e-09, 
    3.210213e-09, 2.462976e-09, 1.980396e-09, 1.683937e-09, 1.428477e-09, 
    1.214204e-09, 1.014345e-09, 9.084117e-10, 8.598278e-10, 8.139805e-10,
  1.523039e-08, 1.194039e-08, 8.691472e-09, 5.987913e-09, 4.43784e-09, 
    3.334684e-09, 2.509524e-09, 2.054609e-09, 1.768426e-09, 1.482969e-09, 
    1.282834e-09, 1.091202e-09, 9.655589e-10, 8.984709e-10, 8.539192e-10,
  1.531707e-08, 1.221984e-08, 9.018255e-09, 6.244114e-09, 4.614275e-09, 
    3.454132e-09, 2.593e-09, 2.166299e-09, 1.865152e-09, 1.549807e-09, 
    1.344494e-09, 1.16753e-09, 1.027253e-09, 9.381774e-10, 8.858184e-10,
  1.539986e-08, 1.238582e-08, 9.288136e-09, 6.488194e-09, 4.796027e-09, 
    3.586474e-09, 2.692757e-09, 2.29787e-09, 1.955152e-09, 1.617111e-09, 
    1.399114e-09, 1.236142e-09, 1.087338e-09, 9.748277e-10, 9.098094e-10,
  1.540813e-08, 1.240846e-08, 9.495521e-09, 6.802632e-09, 5.014662e-09, 
    3.670877e-09, 2.808016e-09, 2.437496e-09, 2.029749e-09, 1.68278e-09, 
    1.446989e-09, 1.290446e-09, 1.140602e-09, 1.017817e-09, 9.387096e-10,
  1.528532e-08, 1.226236e-08, 9.710808e-09, 7.185218e-09, 5.249158e-09, 
    3.726945e-09, 2.928523e-09, 2.53796e-09, 2.080919e-09, 1.746603e-09, 
    1.503703e-09, 1.339166e-09, 1.199013e-09, 1.060183e-09, 9.781549e-10,
  1.493096e-08, 1.214726e-08, 1.005568e-08, 7.638907e-09, 5.481226e-09, 
    3.796223e-09, 3.052885e-09, 2.605427e-09, 2.130001e-09, 1.821075e-09, 
    1.557224e-09, 1.390829e-09, 1.257977e-09, 1.11483e-09, 1.017164e-09,
  1.454612e-08, 1.216951e-08, 1.046107e-08, 8.057828e-09, 5.654921e-09, 
    3.923262e-09, 3.192562e-09, 2.648859e-09, 2.183324e-09, 1.882408e-09, 
    1.61752e-09, 1.451568e-09, 1.299558e-09, 1.170241e-09, 1.058327e-09,
  2.365539e-08, 2.323198e-08, 2.158736e-08, 1.839521e-08, 1.378984e-08, 
    9.323362e-09, 5.761352e-09, 3.697408e-09, 2.783158e-09, 2.092467e-09, 
    1.574418e-09, 1.252893e-09, 1.016207e-09, 8.618097e-10, 6.282593e-10,
  2.333516e-08, 2.330264e-08, 2.213462e-08, 1.940463e-08, 1.505205e-08, 
    1.047578e-08, 6.678684e-09, 4.222956e-09, 3.003302e-09, 2.330171e-09, 
    1.719105e-09, 1.367393e-09, 1.101483e-09, 9.227651e-10, 7.194574e-10,
  2.297424e-08, 2.30001e-08, 2.223586e-08, 1.998013e-08, 1.60649e-08, 
    1.147657e-08, 7.559609e-09, 4.77097e-09, 3.248413e-09, 2.506084e-09, 
    1.866294e-09, 1.465344e-09, 1.178716e-09, 9.783454e-10, 7.862108e-10,
  2.273022e-08, 2.274441e-08, 2.208175e-08, 2.016622e-08, 1.674326e-08, 
    1.231022e-08, 8.382676e-09, 5.370813e-09, 3.55028e-09, 2.666048e-09, 
    2.002311e-09, 1.554872e-09, 1.248986e-09, 1.026654e-09, 8.487934e-10,
  2.242734e-08, 2.245871e-08, 2.195525e-08, 2.011313e-08, 1.704789e-08, 
    1.282301e-08, 9.008031e-09, 5.957961e-09, 3.880322e-09, 2.84484e-09, 
    2.133603e-09, 1.645655e-09, 1.317294e-09, 1.070753e-09, 8.928132e-10,
  2.22194e-08, 2.214828e-08, 2.170525e-08, 1.994698e-08, 1.706004e-08, 
    1.309306e-08, 9.410141e-09, 6.442397e-09, 4.184346e-09, 3.016962e-09, 
    2.25252e-09, 1.729518e-09, 1.385668e-09, 1.111839e-09, 9.316372e-10,
  2.205011e-08, 2.186782e-08, 2.139733e-08, 1.963022e-08, 1.682544e-08, 
    1.308397e-08, 9.577041e-09, 6.78643e-09, 4.44212e-09, 3.171978e-09, 
    2.344717e-09, 1.806295e-09, 1.447833e-09, 1.154127e-09, 9.562223e-10,
  2.194928e-08, 2.160224e-08, 2.09629e-08, 1.915881e-08, 1.6384e-08, 
    1.285635e-08, 9.522388e-09, 6.9396e-09, 4.66766e-09, 3.286751e-09, 
    2.443704e-09, 1.887218e-09, 1.509429e-09, 1.203389e-09, 9.904784e-10,
  2.182346e-08, 2.134316e-08, 2.037506e-08, 1.846342e-08, 1.571455e-08, 
    1.241535e-08, 9.302116e-09, 6.956098e-09, 4.805316e-09, 3.38169e-09, 
    2.542616e-09, 1.963068e-09, 1.563956e-09, 1.247008e-09, 1.030164e-09,
  2.173961e-08, 2.087904e-08, 1.961349e-08, 1.761831e-08, 1.491042e-08, 
    1.187253e-08, 9.020106e-09, 6.870008e-09, 4.859692e-09, 3.462565e-09, 
    2.617617e-09, 2.024373e-09, 1.61049e-09, 1.291092e-09, 1.075308e-09,
  1.46788e-08, 1.109461e-08, 8.610591e-09, 6.406697e-09, 4.611385e-09, 
    3.416573e-09, 2.696065e-09, 2.300119e-09, 1.897e-09, 1.539878e-09, 
    1.215242e-09, 1.039397e-09, 8.615272e-10, 7.227743e-10, 6.378814e-10,
  1.662921e-08, 1.332287e-08, 1.026036e-08, 7.737578e-09, 5.685941e-09, 
    4.095706e-09, 3.099371e-09, 2.517286e-09, 2.113054e-09, 1.729656e-09, 
    1.37235e-09, 1.127026e-09, 9.570197e-10, 8.036579e-10, 6.946776e-10,
  1.839961e-08, 1.52873e-08, 1.22392e-08, 9.332622e-09, 6.927885e-09, 
    5.008248e-09, 3.620701e-09, 2.819772e-09, 2.32776e-09, 1.918301e-09, 
    1.554165e-09, 1.236602e-09, 1.050844e-09, 8.863403e-10, 7.459752e-10,
  2.008865e-08, 1.702794e-08, 1.420595e-08, 1.120406e-08, 8.351194e-09, 
    6.100783e-09, 4.382681e-09, 3.231329e-09, 2.574016e-09, 2.132581e-09, 
    1.734709e-09, 1.383237e-09, 1.143586e-09, 9.795991e-10, 8.110211e-10,
  2.151285e-08, 1.877058e-08, 1.602713e-08, 1.319185e-08, 1.00925e-08, 
    7.450085e-09, 5.344252e-09, 3.803559e-09, 2.878878e-09, 2.359359e-09, 
    1.924038e-09, 1.567272e-09, 1.252007e-09, 1.071922e-09, 8.895847e-10,
  2.250892e-08, 2.03435e-08, 1.771157e-08, 1.506091e-08, 1.202523e-08, 
    8.938194e-09, 6.56276e-09, 4.579684e-09, 3.265664e-09, 2.593168e-09, 
    2.126965e-09, 1.748095e-09, 1.386431e-09, 1.160119e-09, 9.670824e-10,
  2.31215e-08, 2.159273e-08, 1.938708e-08, 1.684409e-08, 1.399733e-08, 
    1.073621e-08, 7.881019e-09, 5.650223e-09, 3.843651e-09, 2.870236e-09, 
    2.338457e-09, 1.9294e-09, 1.559866e-09, 1.257097e-09, 1.047249e-09,
  2.344965e-08, 2.248275e-08, 2.075641e-08, 1.857072e-08, 1.590265e-08, 
    1.268431e-08, 9.368754e-09, 6.792823e-09, 4.645409e-09, 3.224453e-09, 
    2.546455e-09, 2.115176e-09, 1.742248e-09, 1.366598e-09, 1.126855e-09,
  2.369831e-08, 2.323348e-08, 2.190486e-08, 2.005889e-08, 1.766946e-08, 
    1.471135e-08, 1.115258e-08, 8.04521e-09, 5.625385e-09, 3.728712e-09, 
    2.77874e-09, 2.296896e-09, 1.92478e-09, 1.494182e-09, 1.208592e-09,
  2.371601e-08, 2.364842e-08, 2.292382e-08, 2.135396e-08, 1.926561e-08, 
    1.659751e-08, 1.305397e-08, 9.493106e-09, 6.639228e-09, 4.437992e-09, 
    3.05583e-09, 2.477964e-09, 2.109856e-09, 1.639766e-09, 1.29148e-09,
  1.597307e-08, 1.354701e-08, 1.114743e-08, 8.806724e-09, 6.769946e-09, 
    5.187306e-09, 3.871445e-09, 2.853629e-09, 2.052853e-09, 1.555883e-09, 
    1.292124e-09, 1.035064e-09, 7.830848e-10, 5.647823e-10, 3.895237e-10,
  1.610638e-08, 1.38009e-08, 1.139589e-08, 9.004418e-09, 6.909381e-09, 
    5.315886e-09, 4.008495e-09, 2.971656e-09, 2.148736e-09, 1.607539e-09, 
    1.328875e-09, 1.092295e-09, 8.544427e-10, 6.314607e-10, 4.367451e-10,
  1.647105e-08, 1.407659e-08, 1.161907e-08, 9.132851e-09, 7.000533e-09, 
    5.348561e-09, 4.076184e-09, 3.037689e-09, 2.218566e-09, 1.648605e-09, 
    1.35423e-09, 1.138742e-09, 9.276338e-10, 7.091795e-10, 4.929296e-10,
  1.695611e-08, 1.445273e-08, 1.192912e-08, 9.328519e-09, 7.110978e-09, 
    5.406594e-09, 4.127353e-09, 3.097332e-09, 2.270573e-09, 1.685609e-09, 
    1.380984e-09, 1.178394e-09, 9.842754e-10, 7.799839e-10, 5.548316e-10,
  1.75777e-08, 1.491386e-08, 1.231834e-08, 9.612917e-09, 7.253562e-09, 
    5.472468e-09, 4.174265e-09, 3.159333e-09, 2.330113e-09, 1.721774e-09, 
    1.404858e-09, 1.209717e-09, 1.026464e-09, 8.339395e-10, 6.180007e-10,
  1.831678e-08, 1.543222e-08, 1.276614e-08, 9.942594e-09, 7.43114e-09, 
    5.518316e-09, 4.209725e-09, 3.216311e-09, 2.381175e-09, 1.75865e-09, 
    1.418349e-09, 1.23125e-09, 1.055595e-09, 8.730801e-10, 6.809477e-10,
  1.891847e-08, 1.601421e-08, 1.322777e-08, 1.02668e-08, 7.611145e-09, 
    5.596884e-09, 4.271677e-09, 3.264642e-09, 2.436242e-09, 1.807418e-09, 
    1.435852e-09, 1.235309e-09, 1.066822e-09, 9.055002e-10, 7.386109e-10,
  1.95416e-08, 1.661268e-08, 1.374543e-08, 1.073089e-08, 7.896344e-09, 
    5.691555e-09, 4.32039e-09, 3.322245e-09, 2.507014e-09, 1.865632e-09, 
    1.458572e-09, 1.238814e-09, 1.075683e-09, 9.347774e-10, 7.881764e-10,
  1.995722e-08, 1.725331e-08, 1.432721e-08, 1.129183e-08, 8.326364e-09, 
    5.841535e-09, 4.401663e-09, 3.396891e-09, 2.579804e-09, 1.940243e-09, 
    1.487565e-09, 1.24313e-09, 1.082873e-09, 9.60009e-10, 8.314934e-10,
  2.02855e-08, 1.788068e-08, 1.498708e-08, 1.193886e-08, 8.887517e-09, 
    6.126767e-09, 4.482126e-09, 3.457787e-09, 2.641013e-09, 2.016483e-09, 
    1.530738e-09, 1.255178e-09, 1.093489e-09, 9.803974e-10, 8.718134e-10,
  1.699492e-08, 1.668408e-08, 1.624496e-08, 1.492886e-08, 1.347598e-08, 
    1.225649e-08, 1.098718e-08, 9.29075e-09, 7.258402e-09, 5.729623e-09, 
    4.05892e-09, 2.536196e-09, 1.823733e-09, 1.474306e-09, 1.287995e-09,
  1.769958e-08, 1.744017e-08, 1.720011e-08, 1.600821e-08, 1.459114e-08, 
    1.325444e-08, 1.187002e-08, 1.04665e-08, 8.492933e-09, 6.665817e-09, 
    5.039334e-09, 3.449139e-09, 2.261742e-09, 1.676737e-09, 1.409879e-09,
  1.833561e-08, 1.777177e-08, 1.768503e-08, 1.703783e-08, 1.565167e-08, 
    1.427616e-08, 1.282132e-08, 1.144069e-08, 9.676896e-09, 7.814235e-09, 
    6.014665e-09, 4.383067e-09, 2.905072e-09, 1.971576e-09, 1.550965e-09,
  1.874245e-08, 1.823767e-08, 1.792564e-08, 1.765103e-08, 1.664538e-08, 
    1.530346e-08, 1.382238e-08, 1.233792e-08, 1.069693e-08, 8.919725e-09, 
    7.04284e-09, 5.264898e-09, 3.718049e-09, 2.410983e-09, 1.749803e-09,
  1.930724e-08, 1.870309e-08, 1.82954e-08, 1.804737e-08, 1.733618e-08, 
    1.622042e-08, 1.476346e-08, 1.323501e-08, 1.164795e-08, 9.948965e-09, 
    8.141385e-09, 6.219169e-09, 4.564613e-09, 3.0909e-09, 2.068679e-09,
  1.976237e-08, 1.918722e-08, 1.861962e-08, 1.83261e-08, 1.776194e-08, 
    1.696959e-08, 1.564114e-08, 1.413368e-08, 1.249996e-08, 1.086468e-08, 
    9.15857e-09, 7.259678e-09, 5.453793e-09, 3.870035e-09, 2.57366e-09,
  2.023988e-08, 1.97998e-08, 1.919148e-08, 1.877089e-08, 1.818087e-08, 
    1.749417e-08, 1.633255e-08, 1.494426e-08, 1.337609e-08, 1.176626e-08, 
    1.007081e-08, 8.267806e-09, 6.366988e-09, 4.732785e-09, 3.249319e-09,
  2.043147e-08, 2.015039e-08, 1.948673e-08, 1.91418e-08, 1.857976e-08, 
    1.802849e-08, 1.699238e-08, 1.566522e-08, 1.413854e-08, 1.260143e-08, 
    1.097071e-08, 9.194792e-09, 7.263563e-09, 5.53257e-09, 4.044341e-09,
  2.052099e-08, 2.044693e-08, 1.984858e-08, 1.928586e-08, 1.878921e-08, 
    1.823168e-08, 1.745209e-08, 1.626949e-08, 1.484894e-08, 1.330647e-08, 
    1.182401e-08, 1.019614e-08, 8.28109e-09, 6.314866e-09, 4.801374e-09,
  2.087985e-08, 2.066152e-08, 2.017052e-08, 1.955986e-08, 1.894401e-08, 
    1.844473e-08, 1.774277e-08, 1.668691e-08, 1.530833e-08, 1.382655e-08, 
    1.239315e-08, 1.102061e-08, 9.273045e-09, 7.254144e-09, 5.576557e-09,
  1.308565e-08, 1.097903e-08, 9.263085e-09, 7.524872e-09, 5.898925e-09, 
    4.398202e-09, 3.04866e-09, 2.15215e-09, 1.748725e-09, 1.533161e-09, 
    1.390887e-09, 1.264452e-09, 1.118922e-09, 8.236217e-10, 7.368829e-10,
  1.385231e-08, 1.206951e-08, 1.039287e-08, 8.563498e-09, 7.00729e-09, 
    5.451103e-09, 3.997225e-09, 2.792198e-09, 2.066773e-09, 1.703689e-09, 
    1.493084e-09, 1.355713e-09, 1.232928e-09, 9.988299e-10, 7.918083e-10,
  1.462577e-08, 1.309653e-08, 1.146059e-08, 9.707226e-09, 7.999863e-09, 
    6.541769e-09, 5.014776e-09, 3.622526e-09, 2.511671e-09, 1.919148e-09, 
    1.589945e-09, 1.395223e-09, 1.303867e-09, 1.122489e-09, 9.043948e-10,
  1.53128e-08, 1.401738e-08, 1.253459e-08, 1.08903e-08, 9.145153e-09, 
    7.60235e-09, 6.135931e-09, 4.667607e-09, 3.321866e-09, 2.336442e-09, 
    1.85414e-09, 1.551255e-09, 1.407862e-09, 1.286813e-09, 1.060302e-09,
  1.60654e-08, 1.478615e-08, 1.344949e-08, 1.204266e-08, 1.0403e-08, 
    8.739459e-09, 7.258686e-09, 5.782358e-09, 4.349782e-09, 3.061632e-09, 
    2.236092e-09, 1.797618e-09, 1.533511e-09, 1.389767e-09, 1.228881e-09,
  1.665228e-08, 1.5509e-08, 1.422619e-08, 1.294306e-08, 1.151924e-08, 
    9.995544e-09, 8.448771e-09, 6.965897e-09, 5.511833e-09, 4.065788e-09, 
    2.886239e-09, 2.166457e-09, 1.767495e-09, 1.515551e-09, 1.351337e-09,
  1.718203e-08, 1.619443e-08, 1.503127e-08, 1.379286e-08, 1.249674e-08, 
    1.107653e-08, 9.645857e-09, 8.217613e-09, 6.722599e-09, 5.284882e-09, 
    3.86682e-09, 2.788585e-09, 2.135749e-09, 1.745305e-09, 1.493743e-09,
  1.764117e-08, 1.673253e-08, 1.574863e-08, 1.460858e-08, 1.340593e-08, 
    1.213136e-08, 1.07871e-08, 9.439765e-09, 8.098168e-09, 6.555024e-09, 
    5.103282e-09, 3.699848e-09, 2.738304e-09, 2.123672e-09, 1.716925e-09,
  1.810214e-08, 1.730705e-08, 1.643059e-08, 1.537956e-08, 1.425145e-08, 
    1.304262e-08, 1.180979e-08, 1.05249e-08, 9.251304e-09, 7.975163e-09, 
    6.432064e-09, 4.981175e-09, 3.58397e-09, 2.70026e-09, 2.104292e-09,
  1.854136e-08, 1.777052e-08, 1.705969e-08, 1.617602e-08, 1.514596e-08, 
    1.401517e-08, 1.282354e-08, 1.163916e-08, 1.038457e-08, 9.155844e-09, 
    7.853458e-09, 6.33803e-09, 4.882451e-09, 3.526082e-09, 2.657929e-09,
  1.951699e-08, 1.750669e-08, 1.554947e-08, 1.328065e-08, 1.09109e-08, 
    8.271805e-09, 5.745007e-09, 3.807934e-09, 2.509853e-09, 1.854784e-09, 
    1.432315e-09, 1.112568e-09, 9.368716e-10, 7.976697e-10, 6.282611e-10,
  1.940006e-08, 1.827837e-08, 1.625876e-08, 1.413433e-08, 1.188898e-08, 
    9.433008e-09, 6.888903e-09, 4.706846e-09, 3.120643e-09, 2.143621e-09, 
    1.633007e-09, 1.280491e-09, 1.043587e-09, 8.848199e-10, 7.060296e-10,
  1.952863e-08, 1.866126e-08, 1.701019e-08, 1.486932e-08, 1.2788e-08, 
    1.046785e-08, 7.99067e-09, 5.65968e-09, 3.808797e-09, 2.55243e-09, 
    1.833909e-09, 1.454891e-09, 1.173628e-09, 9.698173e-10, 7.957829e-10,
  1.992327e-08, 1.905002e-08, 1.75424e-08, 1.561857e-08, 1.354041e-08, 
    1.135209e-08, 9.039534e-09, 6.684386e-09, 4.623932e-09, 3.083997e-09, 
    2.128395e-09, 1.624196e-09, 1.317254e-09, 1.075037e-09, 8.919153e-10,
  2.05678e-08, 1.942586e-08, 1.792285e-08, 1.629673e-08, 1.432829e-08, 
    1.220424e-08, 9.983224e-09, 7.709018e-09, 5.525084e-09, 3.748864e-09, 
    2.527269e-09, 1.8172e-09, 1.457183e-09, 1.196017e-09, 9.859082e-10,
  2.091048e-08, 1.986129e-08, 1.837192e-08, 1.682892e-08, 1.506997e-08, 
    1.299069e-08, 1.083879e-08, 8.688431e-09, 6.467919e-09, 4.560037e-09, 
    3.059849e-09, 2.093465e-09, 1.595397e-09, 1.304555e-09, 1.090324e-09,
  2.105793e-08, 2.012937e-08, 1.872339e-08, 1.726801e-08, 1.567239e-08, 
    1.37558e-08, 1.167211e-08, 9.633518e-09, 7.448314e-09, 5.419033e-09, 
    3.781977e-09, 2.554141e-09, 1.79799e-09, 1.428742e-09, 1.194639e-09,
  2.103456e-08, 2.020089e-08, 1.895978e-08, 1.766754e-08, 1.62045e-08, 
    1.443367e-08, 1.245818e-08, 1.052033e-08, 8.482613e-09, 6.360865e-09, 
    4.579938e-09, 3.19705e-09, 2.161752e-09, 1.589219e-09, 1.308783e-09,
  2.099607e-08, 2.014381e-08, 1.905019e-08, 1.791763e-08, 1.660909e-08, 
    1.501745e-08, 1.326196e-08, 1.136632e-08, 9.457397e-09, 7.434016e-09, 
    5.463328e-09, 3.939206e-09, 2.706058e-09, 1.865821e-09, 1.445329e-09,
  2.095619e-08, 1.993605e-08, 1.92344e-08, 1.82281e-08, 1.695359e-08, 
    1.55102e-08, 1.39491e-08, 1.220099e-08, 1.040953e-08, 8.522422e-09, 
    6.533775e-09, 4.804878e-09, 3.413406e-09, 2.328435e-09, 1.656826e-09,
  2.213566e-08, 2.163814e-08, 2.112897e-08, 1.99811e-08, 1.796756e-08, 
    1.531187e-08, 1.22143e-08, 8.754738e-09, 5.853658e-09, 3.840452e-09, 
    2.730124e-09, 2.057135e-09, 1.544085e-09, 1.381689e-09, 1.109137e-09,
  2.222395e-08, 2.202111e-08, 2.165233e-08, 2.086665e-08, 1.937887e-08, 
    1.734204e-08, 1.435996e-08, 1.104131e-08, 7.82982e-09, 5.140299e-09, 
    3.365967e-09, 2.504631e-09, 1.837968e-09, 1.474725e-09, 1.279207e-09,
  2.209591e-08, 2.224451e-08, 2.195656e-08, 2.145093e-08, 2.033046e-08, 
    1.887721e-08, 1.641218e-08, 1.314518e-08, 1.001546e-08, 6.854218e-09, 
    4.361716e-09, 3.078296e-09, 2.166944e-09, 1.656672e-09, 1.383946e-09,
  2.227251e-08, 2.232295e-08, 2.22907e-08, 2.193195e-08, 2.106981e-08, 
    1.988536e-08, 1.817351e-08, 1.526644e-08, 1.203914e-08, 8.899896e-09, 
    5.845441e-09, 3.813366e-09, 2.712055e-09, 1.931648e-09, 1.509142e-09,
  2.234926e-08, 2.246388e-08, 2.241995e-08, 2.23926e-08, 2.167986e-08, 
    2.06205e-08, 1.943334e-08, 1.715412e-08, 1.412648e-08, 1.096247e-08, 
    7.738965e-09, 4.952283e-09, 3.389622e-09, 2.34652e-09, 1.756936e-09,
  2.263888e-08, 2.260783e-08, 2.24976e-08, 2.256407e-08, 2.217528e-08, 
    2.122509e-08, 2.024787e-08, 1.868489e-08, 1.599725e-08, 1.293753e-08, 
    9.748116e-09, 6.627676e-09, 4.291823e-09, 2.943091e-09, 2.0599e-09,
  2.283995e-08, 2.299527e-08, 2.272605e-08, 2.282759e-08, 2.249846e-08, 
    2.170777e-08, 2.076867e-08, 1.970171e-08, 1.764914e-08, 1.480133e-08, 
    1.163503e-08, 8.471603e-09, 5.659257e-09, 3.74102e-09, 2.501703e-09,
  2.341251e-08, 2.333399e-08, 2.31422e-08, 2.309117e-08, 2.292916e-08, 
    2.219246e-08, 2.123441e-08, 2.031492e-08, 1.88475e-08, 1.644663e-08, 
    1.35031e-08, 1.028956e-08, 7.286318e-09, 4.78855e-09, 3.144071e-09,
  2.372587e-08, 2.36337e-08, 2.355685e-08, 2.350692e-08, 2.334663e-08, 
    2.269141e-08, 2.170161e-08, 2.08246e-08, 1.964781e-08, 1.77214e-08, 
    1.512681e-08, 1.205537e-08, 8.986417e-09, 6.236269e-09, 4.036929e-09,
  2.440572e-08, 2.43369e-08, 2.404952e-08, 2.393551e-08, 2.382616e-08, 
    2.338127e-08, 2.234656e-08, 2.125735e-08, 2.022644e-08, 1.869184e-08, 
    1.646473e-08, 1.372908e-08, 1.062983e-08, 7.734307e-09, 5.211727e-09,
  1.988928e-08, 1.897127e-08, 1.778763e-08, 1.624106e-08, 1.411886e-08, 
    1.199389e-08, 9.392441e-09, 6.786764e-09, 5.275693e-09, 4.175892e-09, 
    3.085469e-09, 2.212581e-09, 1.565579e-09, 1.069138e-09, 7.86775e-10,
  1.991745e-08, 1.919502e-08, 1.821381e-08, 1.685653e-08, 1.503465e-08, 
    1.314676e-08, 1.070644e-08, 8.062671e-09, 5.849551e-09, 4.628053e-09, 
    3.538446e-09, 2.542072e-09, 1.807838e-09, 1.249261e-09, 9.109833e-10,
  1.999201e-08, 1.933924e-08, 1.851632e-08, 1.750559e-08, 1.593486e-08, 
    1.419153e-08, 1.201379e-08, 9.41238e-09, 6.810571e-09, 5.102736e-09, 
    3.990532e-09, 2.945019e-09, 2.076282e-09, 1.448259e-09, 1.036179e-09,
  2.005303e-08, 1.955963e-08, 1.878936e-08, 1.800031e-08, 1.673418e-08, 
    1.509355e-08, 1.316844e-08, 1.068962e-08, 8.078757e-09, 5.865906e-09, 
    4.430631e-09, 3.404242e-09, 2.412526e-09, 1.677528e-09, 1.183098e-09,
  2.021848e-08, 1.98574e-08, 1.909285e-08, 1.841951e-08, 1.737713e-08, 
    1.584687e-08, 1.415252e-08, 1.19933e-08, 9.376427e-09, 7.012103e-09, 
    5.059113e-09, 3.890883e-09, 2.818819e-09, 1.956739e-09, 1.362498e-09,
  2.042836e-08, 2.011258e-08, 1.943213e-08, 1.878172e-08, 1.795723e-08, 
    1.656393e-08, 1.492013e-08, 1.322528e-08, 1.079735e-08, 8.349841e-09, 
    6.030918e-09, 4.458841e-09, 3.304908e-09, 2.293697e-09, 1.578931e-09,
  2.064038e-08, 2.031544e-08, 1.973812e-08, 1.910077e-08, 1.84176e-08, 
    1.728802e-08, 1.57364e-08, 1.4228e-08, 1.21966e-08, 9.769453e-09, 
    7.355502e-09, 5.269633e-09, 3.886484e-09, 2.708737e-09, 1.852683e-09,
  2.076978e-08, 2.05583e-08, 2.006488e-08, 1.941496e-08, 1.878863e-08, 
    1.792451e-08, 1.656018e-08, 1.511227e-08, 1.349095e-08, 1.117414e-08, 
    8.762535e-09, 6.407495e-09, 4.603133e-09, 3.252684e-09, 2.181761e-09,
  2.102727e-08, 2.079318e-08, 2.042451e-08, 1.983443e-08, 1.919797e-08, 
    1.852248e-08, 1.735556e-08, 1.595663e-08, 1.448012e-08, 1.262905e-08, 
    1.017263e-08, 7.774381e-09, 5.645353e-09, 3.956256e-09, 2.638582e-09,
  2.148191e-08, 2.130128e-08, 2.089839e-08, 2.029974e-08, 1.961349e-08, 
    1.901597e-08, 1.813969e-08, 1.687373e-08, 1.542471e-08, 1.377835e-08, 
    1.1697e-08, 9.178187e-09, 6.897463e-09, 4.925645e-09, 3.292054e-09,
  1.99188e-08, 1.984151e-08, 1.924321e-08, 1.754429e-08, 1.573247e-08, 
    1.438553e-08, 1.320482e-08, 1.168133e-08, 9.723508e-09, 7.830156e-09, 
    5.698412e-09, 4.141519e-09, 3.070839e-09, 2.149904e-09, 1.608454e-09,
  1.978674e-08, 1.989967e-08, 1.971438e-08, 1.844821e-08, 1.641827e-08, 
    1.491343e-08, 1.375987e-08, 1.240788e-08, 1.058901e-08, 8.828851e-09, 
    6.772667e-09, 4.937937e-09, 3.644675e-09, 2.553771e-09, 1.82045e-09,
  1.983566e-08, 1.988611e-08, 1.988173e-08, 1.903402e-08, 1.717917e-08, 
    1.546984e-08, 1.423967e-08, 1.298227e-08, 1.135536e-08, 9.672243e-09, 
    7.804876e-09, 5.808111e-09, 4.283642e-09, 3.037281e-09, 2.085608e-09,
  2.000864e-08, 1.995376e-08, 1.980877e-08, 1.938899e-08, 1.784032e-08, 
    1.605958e-08, 1.471331e-08, 1.354985e-08, 1.207165e-08, 1.044161e-08, 
    8.742282e-09, 6.711887e-09, 5.029527e-09, 3.606226e-09, 2.447923e-09,
  2.01806e-08, 1.995141e-08, 1.973763e-08, 1.938659e-08, 1.838193e-08, 
    1.668294e-08, 1.52468e-08, 1.404517e-08, 1.258898e-08, 1.11367e-08, 
    9.515682e-09, 7.609499e-09, 5.810492e-09, 4.270809e-09, 2.93313e-09,
  2.04653e-08, 2.009607e-08, 1.970161e-08, 1.941327e-08, 1.874108e-08, 
    1.72899e-08, 1.579661e-08, 1.45389e-08, 1.307128e-08, 1.163838e-08, 
    1.020637e-08, 8.514903e-09, 6.652745e-09, 4.965276e-09, 3.497321e-09,
  2.063996e-08, 2.028061e-08, 1.991192e-08, 1.951638e-08, 1.89415e-08, 
    1.774121e-08, 1.629371e-08, 1.506954e-08, 1.359368e-08, 1.212571e-08, 
    1.078419e-08, 9.257572e-09, 7.537751e-09, 5.681437e-09, 4.128016e-09,
  2.0864e-08, 2.044406e-08, 2.000357e-08, 1.967741e-08, 1.904944e-08, 
    1.802912e-08, 1.669365e-08, 1.560185e-08, 1.417419e-08, 1.270935e-08, 
    1.135719e-08, 9.88276e-09, 8.319445e-09, 6.455765e-09, 4.760836e-09,
  2.087606e-08, 2.071049e-08, 2.048782e-08, 1.98016e-08, 1.910596e-08, 
    1.828905e-08, 1.706447e-08, 1.60687e-08, 1.47394e-08, 1.329441e-08, 
    1.191858e-08, 1.049576e-08, 8.957302e-09, 7.222566e-09, 5.412304e-09,
  2.082259e-08, 2.093802e-08, 2.062462e-08, 2.014383e-08, 1.940045e-08, 
    1.851855e-08, 1.743864e-08, 1.650782e-08, 1.529835e-08, 1.384896e-08, 
    1.249249e-08, 1.107575e-08, 9.571077e-09, 7.899147e-09, 6.07311e-09,
  1.475145e-08, 1.349609e-08, 1.23208e-08, 1.056107e-08, 8.88532e-09, 
    7.180812e-09, 5.53309e-09, 4.214668e-09, 3.305992e-09, 2.659305e-09, 
    2.159251e-09, 1.706735e-09, 1.337038e-09, 1.079634e-09, 9.649594e-10,
  1.422933e-08, 1.29717e-08, 1.191957e-08, 1.036451e-08, 8.816979e-09, 
    7.226951e-09, 5.677057e-09, 4.359041e-09, 3.399518e-09, 2.700232e-09, 
    2.193372e-09, 1.768421e-09, 1.4274e-09, 1.176762e-09, 1.003694e-09,
  1.396896e-08, 1.274431e-08, 1.164397e-08, 1.023335e-08, 8.761031e-09, 
    7.217427e-09, 5.660734e-09, 4.337682e-09, 3.427927e-09, 2.73035e-09, 
    2.221664e-09, 1.799936e-09, 1.490024e-09, 1.258819e-09, 1.058391e-09,
  1.382305e-08, 1.268549e-08, 1.154485e-08, 1.014469e-08, 8.742489e-09, 
    7.223568e-09, 5.731805e-09, 4.4315e-09, 3.519872e-09, 2.831264e-09, 
    2.309877e-09, 1.896391e-09, 1.560869e-09, 1.33641e-09, 1.146452e-09,
  1.367648e-08, 1.270431e-08, 1.149372e-08, 1.016377e-08, 8.676063e-09, 
    7.21595e-09, 5.85009e-09, 4.608936e-09, 3.722248e-09, 3.017666e-09, 
    2.437852e-09, 2.007027e-09, 1.657753e-09, 1.437231e-09, 1.242116e-09,
  1.35792e-08, 1.277366e-08, 1.14834e-08, 1.015421e-08, 8.70165e-09, 
    7.231199e-09, 6.019642e-09, 4.916059e-09, 4.020642e-09, 3.295432e-09, 
    2.605581e-09, 2.161548e-09, 1.817026e-09, 1.57018e-09, 1.364664e-09,
  1.354021e-08, 1.275725e-08, 1.146253e-08, 1.013324e-08, 8.831041e-09, 
    7.570765e-09, 6.422337e-09, 5.288189e-09, 4.296826e-09, 3.564866e-09, 
    2.910396e-09, 2.372165e-09, 2.018598e-09, 1.734788e-09, 1.53256e-09,
  1.358723e-08, 1.278566e-08, 1.150056e-08, 1.033069e-08, 9.258928e-09, 
    8.094757e-09, 6.960484e-09, 5.694153e-09, 4.579737e-09, 3.869574e-09, 
    3.267799e-09, 2.678648e-09, 2.264112e-09, 1.950069e-09, 1.722953e-09,
  1.380908e-08, 1.297035e-08, 1.176717e-08, 1.0685e-08, 9.739035e-09, 
    8.621853e-09, 7.409576e-09, 6.098086e-09, 4.974203e-09, 4.259346e-09, 
    3.64779e-09, 3.058917e-09, 2.580119e-09, 2.226203e-09, 1.914843e-09,
  1.415815e-08, 1.329487e-08, 1.221888e-08, 1.11747e-08, 1.020705e-08, 
    8.987445e-09, 7.658752e-09, 6.488183e-09, 5.463764e-09, 4.704725e-09, 
    4.064924e-09, 3.467681e-09, 2.97422e-09, 2.558373e-09, 2.194657e-09,
  2.284175e-08, 2.211716e-08, 2.177404e-08, 2.137067e-08, 2.046492e-08, 
    1.899901e-08, 1.685292e-08, 1.407063e-08, 1.123153e-08, 8.650282e-09, 
    6.333293e-09, 4.635584e-09, 3.512108e-09, 2.762709e-09, 2.337793e-09,
  2.255829e-08, 2.205991e-08, 2.177896e-08, 2.145016e-08, 2.060403e-08, 
    1.916508e-08, 1.70601e-08, 1.437936e-08, 1.1662e-08, 9.095038e-09, 
    6.840365e-09, 5.047818e-09, 3.783801e-09, 2.930095e-09, 2.439054e-09,
  2.252096e-08, 2.200092e-08, 2.171459e-08, 2.140306e-08, 2.054456e-08, 
    1.906496e-08, 1.694404e-08, 1.444735e-08, 1.194381e-08, 9.440037e-09, 
    7.224689e-09, 5.441545e-09, 4.050033e-09, 3.098553e-09, 2.540424e-09,
  2.252779e-08, 2.190956e-08, 2.162271e-08, 2.131239e-08, 2.049335e-08, 
    1.907222e-08, 1.690334e-08, 1.457651e-08, 1.219145e-08, 9.771337e-09, 
    7.551101e-09, 5.781194e-09, 4.349724e-09, 3.269157e-09, 2.628658e-09,
  2.236265e-08, 2.180343e-08, 2.139712e-08, 2.117446e-08, 2.041132e-08, 
    1.904327e-08, 1.685786e-08, 1.460028e-08, 1.233946e-08, 9.939642e-09, 
    7.766117e-09, 6.051858e-09, 4.619898e-09, 3.428387e-09, 2.697019e-09,
  2.233201e-08, 2.177523e-08, 2.115401e-08, 2.1028e-08, 2.027183e-08, 
    1.881504e-08, 1.664432e-08, 1.449142e-08, 1.227137e-08, 9.933228e-09, 
    7.866102e-09, 6.243331e-09, 4.83761e-09, 3.566564e-09, 2.763328e-09,
  2.211985e-08, 2.146835e-08, 2.073669e-08, 2.062914e-08, 1.978014e-08, 
    1.825647e-08, 1.6249e-08, 1.417871e-08, 1.21309e-08, 9.865284e-09, 
    7.889085e-09, 6.354738e-09, 4.977585e-09, 3.710712e-09, 2.86159e-09,
  2.156928e-08, 2.102098e-08, 2.022483e-08, 2.001875e-08, 1.889964e-08, 
    1.737678e-08, 1.556357e-08, 1.37992e-08, 1.194715e-08, 9.763595e-09, 
    7.888421e-09, 6.384753e-09, 5.038208e-09, 3.804827e-09, 2.95582e-09,
  2.06089e-08, 2.0213e-08, 1.947873e-08, 1.90629e-08, 1.764658e-08, 
    1.63643e-08, 1.493481e-08, 1.338012e-08, 1.167734e-08, 9.616645e-09, 
    7.844367e-09, 6.335918e-09, 5.009466e-09, 3.853198e-09, 3.032909e-09,
  1.963662e-08, 1.931856e-08, 1.84717e-08, 1.764558e-08, 1.650677e-08, 
    1.564352e-08, 1.42719e-08, 1.28489e-08, 1.128995e-08, 9.307391e-09, 
    7.669418e-09, 6.195692e-09, 4.927707e-09, 3.846266e-09, 3.060588e-09,
  2.161814e-08, 2.04241e-08, 1.877489e-08, 1.668881e-08, 1.389837e-08, 
    1.14228e-08, 9.204197e-09, 7.172644e-09, 5.303877e-09, 3.508165e-09, 
    2.699675e-09, 2.217277e-09, 1.826673e-09, 1.535802e-09, 1.324431e-09,
  2.171842e-08, 2.098322e-08, 1.948327e-08, 1.769376e-08, 1.518907e-08, 
    1.263395e-08, 1.033071e-08, 8.18354e-09, 6.321927e-09, 4.428362e-09, 
    3.089344e-09, 2.475493e-09, 2.050711e-09, 1.702881e-09, 1.464349e-09,
  2.193947e-08, 2.137796e-08, 2.014835e-08, 1.856509e-08, 1.637376e-08, 
    1.379854e-08, 1.135048e-08, 9.245039e-09, 7.272267e-09, 5.386775e-09, 
    3.72318e-09, 2.730926e-09, 2.295056e-09, 1.896139e-09, 1.604645e-09,
  2.213704e-08, 2.170062e-08, 2.068363e-08, 1.930652e-08, 1.735377e-08, 
    1.495711e-08, 1.246578e-08, 1.023121e-08, 8.279833e-09, 6.353371e-09, 
    4.590761e-09, 3.168445e-09, 2.56089e-09, 2.142836e-09, 1.803778e-09,
  2.229609e-08, 2.190867e-08, 2.115599e-08, 1.985844e-08, 1.819626e-08, 
    1.589315e-08, 1.352814e-08, 1.124406e-08, 9.292354e-09, 7.287325e-09, 
    5.48142e-09, 3.837686e-09, 2.841717e-09, 2.399744e-09, 2.018707e-09,
  2.236199e-08, 2.199777e-08, 2.137332e-08, 2.02976e-08, 1.879858e-08, 
    1.672358e-08, 1.444249e-08, 1.219143e-08, 1.022025e-08, 8.252439e-09, 
    6.386764e-09, 4.665066e-09, 3.299182e-09, 2.633209e-09, 2.225639e-09,
  2.232418e-08, 2.205151e-08, 2.157612e-08, 2.048614e-08, 1.908994e-08, 
    1.731073e-08, 1.529485e-08, 1.310862e-08, 1.109668e-08, 9.183304e-09, 
    7.235197e-09, 5.477705e-09, 3.927522e-09, 2.9633e-09, 2.460957e-09,
  2.218822e-08, 2.19426e-08, 2.148486e-08, 2.06397e-08, 1.941337e-08, 
    1.773954e-08, 1.592523e-08, 1.387273e-08, 1.190642e-08, 1.003208e-08, 
    8.071211e-09, 6.255547e-09, 4.628392e-09, 3.402282e-09, 2.707419e-09,
  2.22046e-08, 2.189629e-08, 2.151585e-08, 2.073896e-08, 1.954103e-08, 
    1.805541e-08, 1.640116e-08, 1.44996e-08, 1.262291e-08, 1.083153e-08, 
    8.870193e-09, 7.025942e-09, 5.350092e-09, 3.99439e-09, 3.07444e-09,
  2.222614e-08, 2.204364e-08, 2.166044e-08, 2.086046e-08, 1.977151e-08, 
    1.834617e-08, 1.67682e-08, 1.504658e-08, 1.322476e-08, 1.152639e-08, 
    9.623867e-09, 7.769188e-09, 6.06392e-09, 4.596837e-09, 3.543071e-09,
  1.899213e-08, 1.76775e-08, 1.630702e-08, 1.436134e-08, 1.216341e-08, 
    9.970116e-09, 8.469522e-09, 6.7265e-09, 5.066582e-09, 3.903111e-09, 
    2.840473e-09, 2.049365e-09, 1.521892e-09, 1.256748e-09, 1.063894e-09,
  2.036216e-08, 1.905225e-08, 1.778302e-08, 1.619901e-08, 1.411863e-08, 
    1.179545e-08, 9.786912e-09, 8.228769e-09, 6.53068e-09, 5.009523e-09, 
    3.631316e-09, 2.59283e-09, 1.802548e-09, 1.408255e-09, 1.187438e-09,
  2.140439e-08, 2.030892e-08, 1.912962e-08, 1.768556e-08, 1.590396e-08, 
    1.386909e-08, 1.136429e-08, 9.462072e-09, 7.759493e-09, 6.25131e-09, 
    4.758689e-09, 3.452796e-09, 2.399172e-09, 1.716251e-09, 1.403028e-09,
  2.233454e-08, 2.134769e-08, 2.018546e-08, 1.909226e-08, 1.746673e-08, 
    1.57414e-08, 1.362687e-08, 1.114406e-08, 9.107705e-09, 7.420435e-09, 
    5.94624e-09, 4.596414e-09, 3.372383e-09, 2.350202e-09, 1.75658e-09,
  2.31533e-08, 2.233351e-08, 2.116509e-08, 2.013428e-08, 1.87523e-08, 
    1.729242e-08, 1.541775e-08, 1.32317e-08, 1.07238e-08, 8.649058e-09, 
    7.016093e-09, 5.648226e-09, 4.43907e-09, 3.240054e-09, 2.320923e-09,
  2.37463e-08, 2.310212e-08, 2.20805e-08, 2.118771e-08, 1.993896e-08, 
    1.865826e-08, 1.699827e-08, 1.497509e-08, 1.265735e-08, 1.015002e-08, 
    8.133424e-09, 6.615631e-09, 5.471626e-09, 4.25042e-09, 3.093917e-09,
  2.41872e-08, 2.36466e-08, 2.27921e-08, 2.203148e-08, 2.09822e-08, 
    1.962711e-08, 1.82725e-08, 1.647662e-08, 1.436939e-08, 1.201104e-08, 
    9.543914e-09, 7.609207e-09, 6.339626e-09, 5.251248e-09, 3.984565e-09,
  2.434622e-08, 2.407699e-08, 2.334702e-08, 2.273802e-08, 2.184039e-08, 
    2.066677e-08, 1.917436e-08, 1.765203e-08, 1.578161e-08, 1.355661e-08, 
    1.130041e-08, 8.930471e-09, 7.159884e-09, 6.01119e-09, 4.919373e-09,
  2.442258e-08, 2.420421e-08, 2.365487e-08, 2.328093e-08, 2.252698e-08, 
    2.153219e-08, 2.02133e-08, 1.860749e-08, 1.68733e-08, 1.483478e-08, 
    1.270307e-08, 1.052724e-08, 8.330695e-09, 6.73487e-09, 5.611818e-09,
  2.446969e-08, 2.423127e-08, 2.383411e-08, 2.360821e-08, 2.304832e-08, 
    2.212709e-08, 2.09172e-08, 1.944925e-08, 1.780184e-08, 1.596658e-08, 
    1.393941e-08, 1.181633e-08, 9.720043e-09, 7.773526e-09, 6.255401e-09,
  2.723227e-09, 2.074772e-09, 1.772695e-09, 1.464477e-09, 1.110032e-09, 
    7.835349e-10, 5.88101e-10, 5.300004e-10, 5.114758e-10, 4.736925e-10, 
    4.286289e-10, 3.769536e-10, 3.401469e-10, 3.090376e-10, 2.649339e-10,
  3.429032e-09, 2.652721e-09, 2.074874e-09, 1.758669e-09, 1.464464e-09, 
    1.134958e-09, 8.213082e-10, 6.079275e-10, 5.040811e-10, 4.520801e-10, 
    4.223002e-10, 3.862052e-10, 3.485206e-10, 3.13134e-10, 2.811224e-10,
  4.468557e-09, 3.455466e-09, 2.614625e-09, 2.053207e-09, 1.728587e-09, 
    1.44018e-09, 1.14938e-09, 8.634827e-10, 6.426055e-10, 5.1725e-10, 
    4.533963e-10, 4.306194e-10, 4.133983e-10, 3.80453e-10, 3.372333e-10,
  5.93494e-09, 4.523023e-09, 3.529941e-09, 2.677903e-09, 2.115262e-09, 
    1.773758e-09, 1.496692e-09, 1.219743e-09, 9.334776e-10, 6.972591e-10, 
    5.630209e-10, 4.796638e-10, 4.473347e-10, 4.21538e-10, 3.866432e-10,
  7.478905e-09, 5.926682e-09, 4.634932e-09, 3.591032e-09, 2.768518e-09, 
    2.202474e-09, 1.842491e-09, 1.556477e-09, 1.270992e-09, 9.858516e-10, 
    7.73802e-10, 6.296649e-10, 5.200271e-10, 4.596412e-10, 4.284566e-10,
  9.216784e-09, 7.478365e-09, 6.005318e-09, 4.743083e-09, 3.722411e-09, 
    2.91112e-09, 2.332026e-09, 1.933971e-09, 1.623689e-09, 1.34808e-09, 
    1.096105e-09, 8.977302e-10, 7.32926e-10, 5.945481e-10, 5.10291e-10,
  1.117329e-08, 9.189998e-09, 7.544498e-09, 6.110674e-09, 4.912475e-09, 
    3.918042e-09, 3.125627e-09, 2.527198e-09, 2.079366e-09, 1.737033e-09, 
    1.465185e-09, 1.221485e-09, 1.019799e-09, 8.270435e-10, 6.724333e-10,
  1.324183e-08, 1.109331e-08, 9.220343e-09, 7.626357e-09, 6.266244e-09, 
    5.124255e-09, 4.160361e-09, 3.388382e-09, 2.768784e-09, 2.273133e-09, 
    1.896667e-09, 1.603608e-09, 1.338144e-09, 1.096803e-09, 8.839178e-10,
  1.531396e-08, 1.318926e-08, 1.116456e-08, 9.36602e-09, 7.781711e-09, 
    6.450676e-09, 5.344496e-09, 4.406502e-09, 3.625414e-09, 2.999461e-09, 
    2.479404e-09, 2.072313e-09, 1.734494e-09, 1.426904e-09, 1.145044e-09,
  1.748424e-08, 1.524328e-08, 1.321382e-08, 1.133042e-08, 9.664286e-09, 
    8.086706e-09, 6.763758e-09, 5.665703e-09, 4.716344e-09, 3.890626e-09, 
    3.230706e-09, 2.69752e-09, 2.271119e-09, 1.894217e-09, 1.554397e-09,
  4.920299e-09, 3.44288e-09, 2.504241e-09, 1.931852e-09, 1.603374e-09, 
    1.39817e-09, 1.232894e-09, 9.935403e-10, 7.264128e-10, 5.977353e-10, 
    5.128277e-10, 4.21309e-10, 3.38316e-10, 2.187635e-10, 9.656921e-11,
  5.36531e-09, 3.819757e-09, 2.786356e-09, 2.087331e-09, 1.700102e-09, 
    1.453168e-09, 1.295386e-09, 1.113328e-09, 8.699745e-10, 6.616624e-10, 
    5.552929e-10, 4.590767e-10, 3.687431e-10, 2.900716e-10, 1.895327e-10,
  5.959428e-09, 4.295613e-09, 3.06447e-09, 2.288391e-09, 1.819187e-09, 
    1.535379e-09, 1.353356e-09, 1.191014e-09, 9.891536e-10, 7.648333e-10, 
    6.050548e-10, 5.060425e-10, 4.159296e-10, 3.213995e-10, 2.596914e-10,
  6.634211e-09, 4.819362e-09, 3.448523e-09, 2.500117e-09, 1.951153e-09, 
    1.609222e-09, 1.402896e-09, 1.250273e-09, 1.078543e-09, 8.787759e-10, 
    6.879644e-10, 5.574092e-10, 4.634225e-10, 3.732271e-10, 2.861705e-10,
  7.314481e-09, 5.346632e-09, 3.853278e-09, 2.77735e-09, 2.117175e-09, 
    1.704534e-09, 1.459805e-09, 1.298479e-09, 1.147862e-09, 9.656044e-10, 
    7.73214e-10, 6.294749e-10, 5.123609e-10, 4.154082e-10, 3.237992e-10,
  8.049414e-09, 5.888313e-09, 4.256203e-09, 3.072629e-09, 2.316717e-09, 
    1.847915e-09, 1.537881e-09, 1.367382e-09, 1.220803e-09, 1.042395e-09, 
    8.497394e-10, 6.988087e-10, 5.716255e-10, 4.614847e-10, 3.663704e-10,
  8.738709e-09, 6.524955e-09, 4.727051e-09, 3.394242e-09, 2.527375e-09, 
    2.004301e-09, 1.647091e-09, 1.44007e-09, 1.297577e-09, 1.126788e-09, 
    9.314469e-10, 7.678885e-10, 6.323755e-10, 5.158e-10, 4.108021e-10,
  9.478251e-09, 7.125444e-09, 5.223586e-09, 3.746966e-09, 2.757536e-09, 
    2.168036e-09, 1.784023e-09, 1.528999e-09, 1.378894e-09, 1.213545e-09, 
    1.024377e-09, 8.55838e-10, 7.137404e-10, 5.813037e-10, 4.646612e-10,
  1.042313e-08, 7.850684e-09, 5.71663e-09, 4.149963e-09, 3.009649e-09, 
    2.323572e-09, 1.919116e-09, 1.635284e-09, 1.475378e-09, 1.314083e-09, 
    1.130677e-09, 9.531925e-10, 7.99158e-10, 6.578715e-10, 5.237896e-10,
  1.138974e-08, 8.691553e-09, 6.315676e-09, 4.559195e-09, 3.334238e-09, 
    2.500253e-09, 2.046103e-09, 1.733137e-09, 1.558952e-09, 1.421857e-09, 
    1.250105e-09, 1.073939e-09, 9.014204e-10, 7.351474e-10, 5.835581e-10,
  2.011136e-08, 1.698308e-08, 1.39324e-08, 1.08946e-08, 8.000525e-09, 
    5.562053e-09, 3.759782e-09, 2.625468e-09, 1.82119e-09, 1.398494e-09, 
    1.176928e-09, 1.050733e-09, 8.524424e-10, 6.890469e-10, 5.073605e-10,
  2.09078e-08, 1.79476e-08, 1.490424e-08, 1.184684e-08, 9.185871e-09, 
    6.53363e-09, 4.469817e-09, 3.095422e-09, 2.121124e-09, 1.603262e-09, 
    1.283389e-09, 1.082581e-09, 9.089902e-10, 7.329308e-10, 5.892085e-10,
  2.152563e-08, 1.878229e-08, 1.580092e-08, 1.274679e-08, 9.963871e-09, 
    7.462371e-09, 5.175549e-09, 3.577066e-09, 2.474484e-09, 1.823789e-09, 
    1.417021e-09, 1.146326e-09, 9.60383e-10, 7.855863e-10, 6.38596e-10,
  2.211499e-08, 1.954916e-08, 1.668271e-08, 1.350797e-08, 1.067608e-08, 
    8.221043e-09, 5.838563e-09, 4.099967e-09, 2.855293e-09, 2.059853e-09, 
    1.547767e-09, 1.250818e-09, 1.025166e-09, 8.505437e-10, 6.978005e-10,
  2.266031e-08, 2.020481e-08, 1.743282e-08, 1.429648e-08, 1.134566e-08, 
    8.818362e-09, 6.493366e-09, 4.59814e-09, 3.205896e-09, 2.311614e-09, 
    1.717301e-09, 1.352648e-09, 1.103626e-09, 9.100377e-10, 7.582081e-10,
  2.305074e-08, 2.082057e-08, 1.81233e-08, 1.505326e-08, 1.186418e-08, 
    9.322135e-09, 6.983534e-09, 4.995527e-09, 3.527983e-09, 2.540756e-09, 
    1.896152e-09, 1.456157e-09, 1.178865e-09, 9.721512e-10, 8.177952e-10,
  2.339084e-08, 2.12871e-08, 1.874935e-08, 1.569925e-08, 1.246852e-08, 
    9.735045e-09, 7.381101e-09, 5.34163e-09, 3.798031e-09, 2.731296e-09, 
    2.059837e-09, 1.57346e-09, 1.260379e-09, 1.037357e-09, 8.731733e-10,
  2.365528e-08, 2.172715e-08, 1.930975e-08, 1.628852e-08, 1.302579e-08, 
    1.016041e-08, 7.692003e-09, 5.616716e-09, 4.018321e-09, 2.873659e-09, 
    2.200997e-09, 1.691753e-09, 1.351581e-09, 1.112216e-09, 9.322562e-10,
  2.383763e-08, 2.20842e-08, 1.98303e-08, 1.682433e-08, 1.353419e-08, 
    1.050581e-08, 7.997276e-09, 5.816961e-09, 4.197343e-09, 2.998602e-09, 
    2.323557e-09, 1.811622e-09, 1.437367e-09, 1.192705e-09, 9.869781e-10,
  2.39385e-08, 2.240962e-08, 2.024278e-08, 1.737123e-08, 1.400294e-08, 
    1.086591e-08, 8.250327e-09, 5.994626e-09, 4.337234e-09, 3.116759e-09, 
    2.408785e-09, 1.918969e-09, 1.521068e-09, 1.274973e-09, 1.064491e-09,
  1.476427e-08, 1.220027e-08, 9.50392e-09, 6.906632e-09, 5.042119e-09, 
    3.563909e-09, 2.281559e-09, 1.578746e-09, 1.507392e-09, 1.304276e-09, 
    1.143513e-09, 9.615323e-10, 8.618864e-10, 7.844242e-10, 6.651679e-10,
  1.620214e-08, 1.413364e-08, 1.15136e-08, 8.794772e-09, 6.517141e-09, 
    4.694935e-09, 3.284992e-09, 2.169828e-09, 1.62961e-09, 1.447842e-09, 
    1.277665e-09, 1.04238e-09, 9.180929e-10, 7.892744e-10, 6.685821e-10,
  1.763981e-08, 1.554221e-08, 1.345661e-08, 1.06819e-08, 8.199454e-09, 
    6.066354e-09, 4.246889e-09, 2.983195e-09, 2.072609e-09, 1.588671e-09, 
    1.429177e-09, 1.176811e-09, 1.006131e-09, 9.007316e-10, 7.386347e-10,
  1.891039e-08, 1.706966e-08, 1.50561e-08, 1.263403e-08, 9.967448e-09, 
    7.638321e-09, 5.576252e-09, 3.883241e-09, 2.777395e-09, 1.95773e-09, 
    1.582852e-09, 1.373433e-09, 1.116841e-09, 9.961066e-10, 8.656909e-10,
  1.991768e-08, 1.835131e-08, 1.653438e-08, 1.434315e-08, 1.181582e-08, 
    9.323156e-09, 7.058191e-09, 5.045805e-09, 3.57568e-09, 2.587665e-09, 
    1.876947e-09, 1.534762e-09, 1.27563e-09, 1.051954e-09, 9.447932e-10,
  2.067914e-08, 1.934172e-08, 1.794917e-08, 1.588549e-08, 1.352547e-08, 
    1.110597e-08, 8.628755e-09, 6.404435e-09, 4.496584e-09, 3.270269e-09, 
    2.371642e-09, 1.755445e-09, 1.438333e-09, 1.160947e-09, 9.983491e-10,
  2.126913e-08, 2.014398e-08, 1.900414e-08, 1.737197e-08, 1.514437e-08, 
    1.273758e-08, 1.036279e-08, 7.880317e-09, 5.630739e-09, 4.00683e-09, 
    2.980404e-09, 2.148582e-09, 1.634101e-09, 1.30114e-09, 1.076219e-09,
  2.191155e-08, 2.085863e-08, 1.982231e-08, 1.85085e-08, 1.670034e-08, 
    1.431932e-08, 1.194615e-08, 9.49048e-09, 6.966591e-09, 4.876346e-09, 
    3.59794e-09, 2.687179e-09, 1.944315e-09, 1.482663e-09, 1.173729e-09,
  2.238496e-08, 2.147474e-08, 2.056326e-08, 1.942621e-08, 1.792237e-08, 
    1.587591e-08, 1.34478e-08, 1.10079e-08, 8.373728e-09, 5.947369e-09, 
    4.252292e-09, 3.237013e-09, 2.383243e-09, 1.74474e-09, 1.30741e-09,
  2.288937e-08, 2.204866e-08, 2.12484e-08, 2.021468e-08, 1.896915e-08, 
    1.715921e-08, 1.490633e-08, 1.242803e-08, 9.798652e-09, 7.132052e-09, 
    5.06161e-09, 3.743629e-09, 2.852347e-09, 2.078816e-09, 1.517541e-09,
  1.158657e-08, 7.909382e-09, 4.658848e-09, 2.767504e-09, 2.121478e-09, 
    1.584435e-09, 1.040982e-09, 8.699546e-10, 7.265097e-10, 6.199314e-10, 
    5.177136e-10, 4.486303e-10, 4.262871e-10, 4.204698e-10, 3.731297e-10,
  1.304566e-08, 9.670525e-09, 6.346554e-09, 3.589101e-09, 2.43728e-09, 
    1.933242e-09, 1.396276e-09, 9.898331e-10, 8.455613e-10, 7.000946e-10, 
    5.798053e-10, 4.920216e-10, 4.581832e-10, 4.35347e-10, 3.979928e-10,
  1.452839e-08, 1.124528e-08, 7.874944e-09, 4.848537e-09, 2.967784e-09, 
    2.211154e-09, 1.773543e-09, 1.249795e-09, 9.412695e-10, 8.146694e-10, 
    6.545999e-10, 5.347833e-10, 4.848705e-10, 4.589476e-10, 4.338627e-10,
  1.601093e-08, 1.27245e-08, 9.422929e-09, 6.237678e-09, 3.798328e-09, 
    2.602119e-09, 2.035678e-09, 1.607267e-09, 1.091275e-09, 8.798458e-10, 
    7.535463e-10, 5.903747e-10, 5.125779e-10, 4.970421e-10, 4.787524e-10,
  1.72841e-08, 1.41067e-08, 1.101178e-08, 7.627736e-09, 4.884912e-09, 
    3.181081e-09, 2.338214e-09, 1.907907e-09, 1.425138e-09, 9.885573e-10, 
    8.420821e-10, 6.800926e-10, 5.370617e-10, 5.100643e-10, 5.260097e-10,
  1.860447e-08, 1.526956e-08, 1.241136e-08, 9.087738e-09, 6.031099e-09, 
    3.971274e-09, 2.779395e-09, 2.131384e-09, 1.777244e-09, 1.24449e-09, 
    9.404749e-10, 7.708525e-10, 5.965189e-10, 5.205232e-10, 5.373241e-10,
  1.981785e-08, 1.640655e-08, 1.37197e-08, 1.046143e-08, 7.255487e-09, 
    4.802962e-09, 3.33749e-09, 2.41013e-09, 2.004652e-09, 1.576354e-09, 
    1.115258e-09, 8.67846e-10, 6.727679e-10, 5.495399e-10, 5.338433e-10,
  2.070504e-08, 1.760592e-08, 1.482489e-08, 1.184298e-08, 8.488782e-09, 
    5.742443e-09, 3.949476e-09, 2.79943e-09, 2.185093e-09, 1.86555e-09, 
    1.393869e-09, 1.008225e-09, 7.689549e-10, 6.034052e-10, 5.452237e-10,
  2.122411e-08, 1.872006e-08, 1.593647e-08, 1.31146e-08, 9.733265e-09, 
    6.765579e-09, 4.645971e-09, 3.29133e-09, 2.456253e-09, 2.059357e-09, 
    1.658844e-09, 1.22026e-09, 8.923089e-10, 6.864661e-10, 5.790738e-10,
  2.156308e-08, 1.962546e-08, 1.692422e-08, 1.426675e-08, 1.108476e-08, 
    7.788218e-09, 5.432713e-09, 3.822295e-09, 2.830441e-09, 2.268685e-09, 
    1.876725e-09, 1.467161e-09, 1.069323e-09, 8.044008e-10, 6.476303e-10,
  8.42256e-09, 5.400014e-09, 2.62225e-09, 1.471623e-09, 1.159315e-09, 
    1.007197e-09, 8.753765e-10, 6.960514e-10, 5.418506e-10, 4.299034e-10, 
    2.951465e-10, 2.448736e-10, 2.919195e-10, 3.41432e-10, 3.405987e-10,
  1.048179e-08, 7.35708e-09, 4.205343e-09, 2.021333e-09, 1.31864e-09, 
    1.102687e-09, 9.625483e-10, 8.065391e-10, 6.473007e-10, 5.100889e-10, 
    3.582269e-10, 2.607789e-10, 2.646307e-10, 3.28417e-10, 3.571713e-10,
  1.298391e-08, 9.229203e-09, 6.126232e-09, 3.093035e-09, 1.587321e-09, 
    1.227889e-09, 1.047269e-09, 9.098181e-10, 7.414431e-10, 6.010653e-10, 
    4.371817e-10, 3.099999e-10, 2.668225e-10, 3.236226e-10, 3.859994e-10,
  1.545914e-08, 1.152769e-08, 8.121146e-09, 4.752953e-09, 2.29204e-09, 
    1.399761e-09, 1.139897e-09, 9.992032e-10, 8.409786e-10, 6.992131e-10, 
    5.207592e-10, 3.697625e-10, 2.935852e-10, 3.15518e-10, 3.982812e-10,
  1.767313e-08, 1.403613e-08, 1.01451e-08, 6.765165e-09, 3.455215e-09, 
    1.771648e-09, 1.265433e-09, 1.079294e-09, 9.384669e-10, 7.946482e-10, 
    6.237727e-10, 4.299004e-10, 3.37371e-10, 3.162427e-10, 3.857248e-10,
  1.956704e-08, 1.635766e-08, 1.247035e-08, 8.812094e-09, 5.115385e-09, 
    2.527303e-09, 1.477532e-09, 1.14684e-09, 1.032325e-09, 8.890558e-10, 
    7.39581e-10, 5.126557e-10, 3.917107e-10, 3.337144e-10, 3.617471e-10,
  2.112472e-08, 1.832801e-08, 1.482141e-08, 1.076637e-08, 7.097115e-09, 
    3.647324e-09, 1.895251e-09, 1.263055e-09, 1.090208e-09, 9.710458e-10, 
    8.498161e-10, 6.249013e-10, 4.599175e-10, 3.681984e-10, 3.529916e-10,
  2.242578e-08, 1.999734e-08, 1.703446e-08, 1.304057e-08, 9.119177e-09, 
    5.200598e-09, 2.600866e-09, 1.492664e-09, 1.131008e-09, 1.048173e-09, 
    9.460694e-10, 7.53183e-10, 5.479048e-10, 4.228564e-10, 3.651727e-10,
  2.348244e-08, 2.144215e-08, 1.886557e-08, 1.525229e-08, 1.110779e-08, 
    7.06778e-09, 3.605618e-09, 1.911314e-09, 1.247029e-09, 1.088595e-09, 
    1.021195e-09, 8.833285e-10, 6.535549e-10, 4.948391e-10, 3.973924e-10,
  2.433839e-08, 2.260558e-08, 2.052566e-08, 1.740326e-08, 1.32157e-08, 
    9.085158e-09, 5.015845e-09, 2.542793e-09, 1.4738e-09, 1.129445e-09, 
    1.067072e-09, 9.908907e-10, 7.803809e-10, 5.809739e-10, 4.472307e-10,
  7.209653e-09, 4.393482e-09, 2.77089e-09, 1.864439e-09, 1.471505e-09, 
    1.219378e-09, 1.014915e-09, 8.134912e-10, 6.819274e-10, 6.485086e-10, 
    6.56066e-10, 7.346918e-10, 7.957006e-10, 8.433944e-10, 8.607765e-10,
  7.779091e-09, 4.979261e-09, 3.076188e-09, 2.013399e-09, 1.545574e-09, 
    1.276949e-09, 1.06488e-09, 8.512575e-10, 6.966716e-10, 6.389038e-10, 
    6.346372e-10, 7.075117e-10, 7.963685e-10, 8.451191e-10, 8.649749e-10,
  9.115362e-09, 5.659261e-09, 3.406508e-09, 2.157391e-09, 1.60075e-09, 
    1.317071e-09, 1.099996e-09, 8.963816e-10, 7.149649e-10, 6.25759e-10, 
    6.138701e-10, 6.734253e-10, 7.770413e-10, 8.285243e-10, 8.623569e-10,
  1.089458e-08, 6.666415e-09, 3.871953e-09, 2.358014e-09, 1.674584e-09, 
    1.36e-09, 1.149586e-09, 9.704202e-10, 7.500255e-10, 6.451314e-10, 
    6.067629e-10, 6.452602e-10, 7.391395e-10, 8.11835e-10, 8.589262e-10,
  1.292303e-08, 7.905213e-09, 4.528307e-09, 2.641564e-09, 1.789494e-09, 
    1.414804e-09, 1.20285e-09, 1.063523e-09, 8.146732e-10, 6.774905e-10, 
    6.1621e-10, 6.281692e-10, 7.020483e-10, 7.89339e-10, 8.423593e-10,
  1.507822e-08, 9.433998e-09, 5.393542e-09, 3.023032e-09, 1.956539e-09, 
    1.488662e-09, 1.244619e-09, 1.113457e-09, 8.847265e-10, 6.918509e-10, 
    6.377779e-10, 6.162932e-10, 6.698676e-10, 7.486656e-10, 8.209327e-10,
  1.708631e-08, 1.126525e-08, 6.52609e-09, 3.566496e-09, 2.195917e-09, 
    1.584517e-09, 1.292747e-09, 1.14519e-09, 9.666322e-10, 7.446374e-10, 
    6.633101e-10, 6.173282e-10, 6.415959e-10, 7.079652e-10, 7.927898e-10,
  1.865014e-08, 1.325558e-08, 7.944288e-09, 4.302879e-09, 2.516875e-09, 
    1.72319e-09, 1.357243e-09, 1.168706e-09, 1.024325e-09, 7.882009e-10, 
    6.64284e-10, 6.229058e-10, 6.230876e-10, 6.752457e-10, 7.55293e-10,
  1.97272e-08, 1.53802e-08, 9.65002e-09, 5.279718e-09, 2.965542e-09, 
    1.923089e-09, 1.447089e-09, 1.216553e-09, 1.065792e-09, 8.569194e-10, 
    6.942777e-10, 6.39868e-10, 6.166264e-10, 6.449631e-10, 7.195346e-10,
  2.043136e-08, 1.717706e-08, 1.174787e-08, 6.505216e-09, 3.562112e-09, 
    2.179513e-09, 1.573401e-09, 1.292332e-09, 1.114745e-09, 9.195168e-10, 
    7.373297e-10, 6.42353e-10, 6.14082e-10, 6.252404e-10, 6.846047e-10,
  2.343167e-08, 2.221043e-08, 2.014257e-08, 1.751778e-08, 1.502195e-08, 
    1.263208e-08, 1.034364e-08, 8.293734e-09, 6.466188e-09, 5.010091e-09, 
    3.899932e-09, 2.938697e-09, 2.155676e-09, 1.672799e-09, 1.341888e-09,
  2.366834e-08, 2.265446e-08, 2.070052e-08, 1.808097e-08, 1.54657e-08, 
    1.296088e-08, 1.062027e-08, 8.488898e-09, 6.606806e-09, 5.069934e-09, 
    3.900248e-09, 2.89894e-09, 2.086482e-09, 1.586899e-09, 1.270789e-09,
  2.38359e-08, 2.291814e-08, 2.111335e-08, 1.855466e-08, 1.602991e-08, 
    1.336984e-08, 1.089746e-08, 8.682081e-09, 6.717286e-09, 5.077423e-09, 
    3.845544e-09, 2.832813e-09, 2.012784e-09, 1.513923e-09, 1.218736e-09,
  2.402225e-08, 2.310848e-08, 2.160075e-08, 1.903391e-08, 1.654751e-08, 
    1.381569e-08, 1.123429e-08, 8.914109e-09, 6.878458e-09, 5.122171e-09, 
    3.808137e-09, 2.776946e-09, 1.951902e-09, 1.468867e-09, 1.19307e-09,
  2.426554e-08, 2.342972e-08, 2.189652e-08, 1.959666e-08, 1.701028e-08, 
    1.439831e-08, 1.161963e-08, 9.215626e-09, 7.080083e-09, 5.239851e-09, 
    3.843049e-09, 2.76549e-09, 1.923785e-09, 1.434212e-09, 1.173091e-09,
  2.468534e-08, 2.358798e-08, 2.22623e-08, 2.005772e-08, 1.751617e-08, 
    1.499707e-08, 1.209797e-08, 9.539005e-09, 7.321891e-09, 5.415973e-09, 
    3.919845e-09, 2.76889e-09, 1.887027e-09, 1.392066e-09, 1.156333e-09,
  2.532387e-08, 2.391633e-08, 2.261906e-08, 2.046286e-08, 1.794956e-08, 
    1.555127e-08, 1.266564e-08, 9.915129e-09, 7.585334e-09, 5.588296e-09, 
    4.02351e-09, 2.791039e-09, 1.868001e-09, 1.359669e-09, 1.149192e-09,
  2.612759e-08, 2.466563e-08, 2.301453e-08, 2.10558e-08, 1.831344e-08, 
    1.598493e-08, 1.329862e-08, 1.034244e-08, 7.88316e-09, 5.781634e-09, 
    4.148176e-09, 2.854572e-09, 1.875502e-09, 1.340827e-09, 1.137247e-09,
  2.674348e-08, 2.523007e-08, 2.372998e-08, 2.174583e-08, 1.896647e-08, 
    1.636694e-08, 1.385406e-08, 1.086874e-08, 8.216318e-09, 5.997802e-09, 
    4.284272e-09, 2.95499e-09, 1.909613e-09, 1.334978e-09, 1.129189e-09,
  2.684758e-08, 2.588424e-08, 2.463602e-08, 2.245024e-08, 1.975222e-08, 
    1.690756e-08, 1.434129e-08, 1.150369e-08, 8.606961e-09, 6.257212e-09, 
    4.450729e-09, 3.083392e-09, 1.966478e-09, 1.338736e-09, 1.115128e-09,
  1.57862e-08, 1.512837e-08, 1.462246e-08, 1.387686e-08, 1.321057e-08, 
    1.270287e-08, 1.226451e-08, 1.157551e-08, 1.080035e-08, 1.011503e-08, 
    9.374041e-09, 8.56854e-09, 7.575468e-09, 6.713842e-09, 6.060554e-09,
  1.612156e-08, 1.574704e-08, 1.533265e-08, 1.451465e-08, 1.36896e-08, 
    1.308458e-08, 1.271058e-08, 1.21493e-08, 1.13687e-08, 1.068517e-08, 
    9.926998e-09, 9.206327e-09, 8.237598e-09, 7.171023e-09, 6.370562e-09,
  1.652598e-08, 1.616519e-08, 1.593886e-08, 1.52424e-08, 1.421027e-08, 
    1.348712e-08, 1.314697e-08, 1.271553e-08, 1.197984e-08, 1.125986e-08, 
    1.051738e-08, 9.740354e-09, 8.825123e-09, 7.690504e-09, 6.695009e-09,
  1.68411e-08, 1.655965e-08, 1.637847e-08, 1.603391e-08, 1.489277e-08, 
    1.391726e-08, 1.351369e-08, 1.324918e-08, 1.259077e-08, 1.182316e-08, 
    1.104648e-08, 1.025896e-08, 9.368176e-09, 8.21893e-09, 7.081833e-09,
  1.722337e-08, 1.692053e-08, 1.675358e-08, 1.657106e-08, 1.564632e-08, 
    1.4484e-08, 1.384996e-08, 1.368546e-08, 1.319327e-08, 1.241234e-08, 
    1.157409e-08, 1.077216e-08, 9.843764e-09, 8.714194e-09, 7.482898e-09,
  1.79445e-08, 1.751375e-08, 1.726096e-08, 1.706963e-08, 1.644197e-08, 
    1.512383e-08, 1.424012e-08, 1.402591e-08, 1.368913e-08, 1.29983e-08, 
    1.207979e-08, 1.12471e-08, 1.024967e-08, 9.112268e-09, 7.84594e-09,
  1.867394e-08, 1.824335e-08, 1.797145e-08, 1.745796e-08, 1.716185e-08, 
    1.589924e-08, 1.464505e-08, 1.429476e-08, 1.41789e-08, 1.357415e-08, 
    1.262155e-08, 1.167988e-08, 1.06552e-08, 9.448271e-09, 8.174596e-09,
  1.943704e-08, 1.886703e-08, 1.871621e-08, 1.81306e-08, 1.769934e-08, 
    1.668651e-08, 1.524672e-08, 1.442457e-08, 1.437559e-08, 1.404049e-08, 
    1.309753e-08, 1.211075e-08, 1.101492e-08, 9.752575e-09, 8.470288e-09,
  1.994918e-08, 1.933443e-08, 1.918089e-08, 1.875332e-08, 1.810924e-08, 
    1.730651e-08, 1.594657e-08, 1.471178e-08, 1.44926e-08, 1.433999e-08, 
    1.356399e-08, 1.254705e-08, 1.136133e-08, 1.001443e-08, 8.704539e-09,
  2.060426e-08, 1.99574e-08, 1.947929e-08, 1.923961e-08, 1.868192e-08, 
    1.790344e-08, 1.662794e-08, 1.510105e-08, 1.453013e-08, 1.45058e-08, 
    1.395094e-08, 1.292535e-08, 1.171564e-08, 1.025994e-08, 8.909568e-09,
  2.266997e-08, 2.075111e-08, 1.926318e-08, 1.743253e-08, 1.590007e-08, 
    1.403507e-08, 1.232608e-08, 1.049299e-08, 8.543827e-09, 6.722481e-09, 
    5.323753e-09, 4.277674e-09, 3.475567e-09, 2.861517e-09, 2.410468e-09,
  2.2259e-08, 2.102846e-08, 1.973533e-08, 1.750987e-08, 1.575834e-08, 
    1.398531e-08, 1.228608e-08, 1.060974e-08, 8.739424e-09, 6.922563e-09, 
    5.480149e-09, 4.438457e-09, 3.649794e-09, 3.019019e-09, 2.548411e-09,
  2.209554e-08, 2.099382e-08, 1.948779e-08, 1.728604e-08, 1.555153e-08, 
    1.390272e-08, 1.221599e-08, 1.070365e-08, 9.032219e-09, 7.241298e-09, 
    5.762727e-09, 4.668677e-09, 3.835177e-09, 3.203324e-09, 2.740072e-09,
  2.17947e-08, 2.040077e-08, 1.882868e-08, 1.678491e-08, 1.517984e-08, 
    1.359023e-08, 1.215932e-08, 1.085984e-08, 9.332939e-09, 7.628046e-09, 
    6.112226e-09, 4.959996e-09, 4.05787e-09, 3.399688e-09, 2.896354e-09,
  2.149262e-08, 1.9695e-08, 1.835089e-08, 1.632894e-08, 1.469766e-08, 
    1.342936e-08, 1.219209e-08, 1.092816e-08, 9.558545e-09, 7.972287e-09, 
    6.519698e-09, 5.281908e-09, 4.271735e-09, 3.54107e-09, 3.011543e-09,
  2.116037e-08, 1.915032e-08, 1.801408e-08, 1.609769e-08, 1.463644e-08, 
    1.361848e-08, 1.231018e-08, 1.096621e-08, 9.729194e-09, 8.331591e-09, 
    6.930471e-09, 5.630394e-09, 4.510653e-09, 3.686627e-09, 3.091198e-09,
  2.071457e-08, 1.881929e-08, 1.774501e-08, 1.62531e-08, 1.500297e-08, 
    1.385592e-08, 1.241897e-08, 1.104513e-08, 9.89184e-09, 8.654848e-09, 
    7.336522e-09, 6.070942e-09, 4.869869e-09, 3.90725e-09, 3.235497e-09,
  2.065308e-08, 1.888268e-08, 1.771842e-08, 1.668226e-08, 1.547498e-08, 
    1.401604e-08, 1.256008e-08, 1.12703e-08, 1.014271e-08, 8.994082e-09, 
    7.76317e-09, 6.57985e-09, 5.366665e-09, 4.288364e-09, 3.474981e-09,
  2.0966e-08, 1.916871e-08, 1.804432e-08, 1.701615e-08, 1.567987e-08, 
    1.414783e-08, 1.277323e-08, 1.160168e-08, 1.04571e-08, 9.353434e-09, 
    8.196765e-09, 7.103439e-09, 5.962208e-09, 4.802851e-09, 3.827155e-09,
  2.176909e-08, 1.975776e-08, 1.837419e-08, 1.722455e-08, 1.581703e-08, 
    1.440313e-08, 1.305945e-08, 1.194189e-08, 1.084586e-08, 9.756395e-09, 
    8.609805e-09, 7.585106e-09, 6.513297e-09, 5.411096e-09, 4.289626e-09,
  2.36699e-08, 2.3391e-08, 2.325418e-08, 2.329829e-08, 2.357014e-08, 
    2.3786e-08, 2.365225e-08, 2.244585e-08, 2.083932e-08, 1.916086e-08, 
    1.747403e-08, 1.568018e-08, 1.395751e-08, 1.281391e-08, 1.135132e-08,
  2.380407e-08, 2.409175e-08, 2.378987e-08, 2.326241e-08, 2.314727e-08, 
    2.333657e-08, 2.353254e-08, 2.293737e-08, 2.182628e-08, 2.016895e-08, 
    1.839446e-08, 1.663724e-08, 1.466899e-08, 1.323332e-08, 1.186435e-08,
  2.453866e-08, 2.448131e-08, 2.450246e-08, 2.396915e-08, 2.331051e-08, 
    2.334904e-08, 2.346429e-08, 2.330819e-08, 2.254047e-08, 2.129738e-08, 
    1.935357e-08, 1.740125e-08, 1.546152e-08, 1.378852e-08, 1.236602e-08,
  2.637841e-08, 2.558085e-08, 2.552522e-08, 2.492817e-08, 2.395341e-08, 
    2.349055e-08, 2.349596e-08, 2.332493e-08, 2.290196e-08, 2.20037e-08, 
    2.036247e-08, 1.827902e-08, 1.609551e-08, 1.428261e-08, 1.274105e-08,
  2.736834e-08, 2.663676e-08, 2.613428e-08, 2.554087e-08, 2.458511e-08, 
    2.370915e-08, 2.340193e-08, 2.327412e-08, 2.301318e-08, 2.243106e-08, 
    2.117387e-08, 1.923715e-08, 1.693086e-08, 1.485508e-08, 1.304417e-08,
  2.738702e-08, 2.679324e-08, 2.647711e-08, 2.573099e-08, 2.488595e-08, 
    2.392411e-08, 2.333228e-08, 2.318629e-08, 2.295547e-08, 2.264366e-08, 
    2.182394e-08, 2.014837e-08, 1.769713e-08, 1.547485e-08, 1.344971e-08,
  2.67897e-08, 2.665385e-08, 2.671789e-08, 2.598062e-08, 2.540367e-08, 
    2.437088e-08, 2.347094e-08, 2.308335e-08, 2.279727e-08, 2.251174e-08, 
    2.204464e-08, 2.077074e-08, 1.844706e-08, 1.605797e-08, 1.38142e-08,
  2.607584e-08, 2.62114e-08, 2.663273e-08, 2.645969e-08, 2.585265e-08, 
    2.47702e-08, 2.380603e-08, 2.315031e-08, 2.26539e-08, 2.232212e-08, 
    2.19973e-08, 2.100657e-08, 1.901143e-08, 1.663419e-08, 1.424061e-08,
  2.637648e-08, 2.608796e-08, 2.639303e-08, 2.668472e-08, 2.614093e-08, 
    2.494246e-08, 2.401277e-08, 2.342108e-08, 2.280282e-08, 2.216515e-08, 
    2.161999e-08, 2.073437e-08, 1.906355e-08, 1.704737e-08, 1.467915e-08,
  2.620822e-08, 2.608889e-08, 2.604035e-08, 2.610412e-08, 2.544373e-08, 
    2.45561e-08, 2.396223e-08, 2.344935e-08, 2.30278e-08, 2.239084e-08, 
    2.158068e-08, 2.055861e-08, 1.900213e-08, 1.721113e-08, 1.5003e-08,
  2.528158e-08, 2.506346e-08, 2.443454e-08, 2.371603e-08, 2.273816e-08, 
    2.193984e-08, 2.105231e-08, 2.015819e-08, 1.870952e-08, 1.764329e-08, 
    1.717448e-08, 1.699957e-08, 1.649091e-08, 1.51054e-08, 1.337817e-08,
  2.477113e-08, 2.476846e-08, 2.430299e-08, 2.369514e-08, 2.257643e-08, 
    2.180557e-08, 2.104276e-08, 2.020675e-08, 1.900745e-08, 1.791639e-08, 
    1.72684e-08, 1.702103e-08, 1.680932e-08, 1.586979e-08, 1.40349e-08,
  2.475357e-08, 2.474303e-08, 2.426879e-08, 2.358851e-08, 2.250841e-08, 
    2.165107e-08, 2.097298e-08, 2.035056e-08, 1.927612e-08, 1.82296e-08, 
    1.747766e-08, 1.701226e-08, 1.691808e-08, 1.631243e-08, 1.477719e-08,
  2.469359e-08, 2.473246e-08, 2.423439e-08, 2.34937e-08, 2.234212e-08, 
    2.153983e-08, 2.080091e-08, 2.033095e-08, 1.954618e-08, 1.84925e-08, 
    1.766789e-08, 1.708129e-08, 1.688179e-08, 1.647771e-08, 1.534705e-08,
  2.469259e-08, 2.458243e-08, 2.403647e-08, 2.335515e-08, 2.232916e-08, 
    2.160125e-08, 2.080376e-08, 2.035708e-08, 1.974004e-08, 1.883629e-08, 
    1.794906e-08, 1.719911e-08, 1.684408e-08, 1.653918e-08, 1.565547e-08,
  2.440086e-08, 2.418893e-08, 2.389444e-08, 2.336728e-08, 2.23919e-08, 
    2.169257e-08, 2.085306e-08, 2.035297e-08, 1.991365e-08, 1.900951e-08, 
    1.820228e-08, 1.738712e-08, 1.690394e-08, 1.65611e-08, 1.582208e-08,
  2.450678e-08, 2.416454e-08, 2.360632e-08, 2.338873e-08, 2.263952e-08, 
    2.184717e-08, 2.094032e-08, 2.029623e-08, 1.999012e-08, 1.925796e-08, 
    1.838943e-08, 1.756955e-08, 1.697276e-08, 1.663057e-08, 1.598729e-08,
  2.44507e-08, 2.435559e-08, 2.380312e-08, 2.328331e-08, 2.290921e-08, 
    2.211828e-08, 2.110606e-08, 2.028147e-08, 2.003735e-08, 1.946001e-08, 
    1.873349e-08, 1.781754e-08, 1.701501e-08, 1.655559e-08, 1.60616e-08,
  2.425021e-08, 2.444004e-08, 2.407865e-08, 2.366315e-08, 2.300815e-08, 
    2.239264e-08, 2.145699e-08, 2.03447e-08, 2.002657e-08, 1.962563e-08, 
    1.91135e-08, 1.821953e-08, 1.726276e-08, 1.649175e-08, 1.600003e-08,
  2.41078e-08, 2.418965e-08, 2.412766e-08, 2.405642e-08, 2.365058e-08, 
    2.276645e-08, 2.192298e-08, 2.062399e-08, 2.011766e-08, 1.979358e-08, 
    1.937053e-08, 1.859062e-08, 1.765475e-08, 1.665028e-08, 1.596986e-08,
  2.011125e-08, 1.926096e-08, 1.795977e-08, 1.685462e-08, 1.596929e-08, 
    1.506054e-08, 1.406633e-08, 1.309853e-08, 1.240311e-08, 1.153179e-08, 
    1.07538e-08, 9.787168e-09, 8.964268e-09, 8.605633e-09, 8.463512e-09,
  2.17297e-08, 2.080962e-08, 1.961798e-08, 1.836742e-08, 1.739009e-08, 
    1.651636e-08, 1.554751e-08, 1.445533e-08, 1.359849e-08, 1.283334e-08, 
    1.200684e-08, 1.124253e-08, 1.030896e-08, 9.63861e-09, 9.371005e-09,
  2.376429e-08, 2.233704e-08, 2.109337e-08, 1.999201e-08, 1.894269e-08, 
    1.795018e-08, 1.69541e-08, 1.595704e-08, 1.486441e-08, 1.402503e-08, 
    1.318902e-08, 1.247291e-08, 1.169264e-08, 1.093947e-08, 1.044201e-08,
  2.544029e-08, 2.389479e-08, 2.254801e-08, 2.149295e-08, 2.053519e-08, 
    1.941839e-08, 1.83192e-08, 1.736716e-08, 1.620103e-08, 1.526609e-08, 
    1.432807e-08, 1.3593e-08, 1.291213e-08, 1.218787e-08, 1.156484e-08,
  2.641282e-08, 2.524512e-08, 2.378665e-08, 2.288551e-08, 2.188669e-08, 
    2.071314e-08, 1.954103e-08, 1.860822e-08, 1.754238e-08, 1.65383e-08, 
    1.557171e-08, 1.466523e-08, 1.405848e-08, 1.346088e-08, 1.278445e-08,
  2.737091e-08, 2.634318e-08, 2.517115e-08, 2.411642e-08, 2.296308e-08, 
    2.153039e-08, 2.051668e-08, 1.962269e-08, 1.874334e-08, 1.778498e-08, 
    1.688301e-08, 1.584575e-08, 1.523277e-08, 1.467046e-08, 1.404527e-08,
  2.829533e-08, 2.686622e-08, 2.602635e-08, 2.51926e-08, 2.373735e-08, 
    2.234539e-08, 2.135112e-08, 2.048756e-08, 1.976649e-08, 1.89129e-08, 
    1.816693e-08, 1.717896e-08, 1.651045e-08, 1.591588e-08, 1.528322e-08,
  2.876976e-08, 2.724931e-08, 2.65358e-08, 2.563234e-08, 2.432435e-08, 
    2.30763e-08, 2.222478e-08, 2.127016e-08, 2.059995e-08, 1.986675e-08, 
    1.92423e-08, 1.840077e-08, 1.7687e-08, 1.70788e-08, 1.647802e-08,
  2.916772e-08, 2.732053e-08, 2.645448e-08, 2.590595e-08, 2.500065e-08, 
    2.395758e-08, 2.288972e-08, 2.190521e-08, 2.116993e-08, 2.063403e-08, 
    2.020843e-08, 1.953457e-08, 1.884404e-08, 1.817632e-08, 1.758967e-08,
  2.904045e-08, 2.765098e-08, 2.653781e-08, 2.606759e-08, 2.548611e-08, 
    2.459679e-08, 2.350017e-08, 2.237792e-08, 2.154246e-08, 2.104282e-08, 
    2.084698e-08, 2.030298e-08, 1.965573e-08, 1.910653e-08, 1.853428e-08,
  1.340145e-08, 1.102562e-08, 9.356998e-09, 7.160351e-09, 5.59541e-09, 
    4.468446e-09, 3.60587e-09, 2.94553e-09, 2.439168e-09, 2.035291e-09, 
    1.637633e-09, 1.2583e-09, 9.819726e-10, 7.907932e-10, 6.21427e-10,
  1.41993e-08, 1.213575e-08, 1.029016e-08, 8.398144e-09, 6.483597e-09, 
    5.132252e-09, 4.16242e-09, 3.387848e-09, 2.787419e-09, 2.347831e-09, 
    1.948282e-09, 1.563842e-09, 1.21092e-09, 9.605363e-10, 7.738304e-10,
  1.525687e-08, 1.339762e-08, 1.147549e-08, 9.551299e-09, 7.687381e-09, 
    5.973121e-09, 4.822096e-09, 3.997049e-09, 3.282838e-09, 2.734275e-09, 
    2.317226e-09, 1.933223e-09, 1.558945e-09, 1.218281e-09, 9.797873e-10,
  1.588289e-08, 1.457195e-08, 1.273812e-08, 1.081587e-08, 8.865936e-09, 
    7.064402e-09, 5.567474e-09, 4.59458e-09, 3.84478e-09, 3.196451e-09, 
    2.677024e-09, 2.257935e-09, 1.894226e-09, 1.52162e-09, 1.199471e-09,
  1.637399e-08, 1.537031e-08, 1.382554e-08, 1.200547e-08, 1.016747e-08, 
    8.32472e-09, 6.600305e-09, 5.30166e-09, 4.453688e-09, 3.764782e-09, 
    3.165926e-09, 2.650855e-09, 2.238211e-09, 1.874039e-09, 1.516158e-09,
  1.682772e-08, 1.613795e-08, 1.477829e-08, 1.319093e-08, 1.141795e-08, 
    9.671965e-09, 7.922694e-09, 6.331987e-09, 5.183637e-09, 4.400952e-09, 
    3.770264e-09, 3.193737e-09, 2.68714e-09, 2.272679e-09, 1.912618e-09,
  1.750159e-08, 1.688817e-08, 1.580727e-08, 1.436267e-08, 1.274689e-08, 
    1.101313e-08, 9.327992e-09, 7.66109e-09, 6.212426e-09, 5.149507e-09, 
    4.417648e-09, 3.816288e-09, 3.251554e-09, 2.764847e-09, 2.354429e-09,
  1.827975e-08, 1.761506e-08, 1.674221e-08, 1.54608e-08, 1.404884e-08, 
    1.243405e-08, 1.07608e-08, 9.113377e-09, 7.565326e-09, 6.205856e-09, 
    5.167428e-09, 4.453631e-09, 3.874788e-09, 3.332976e-09, 2.878729e-09,
  1.934403e-08, 1.848629e-08, 1.765352e-08, 1.652218e-08, 1.521535e-08, 
    1.38109e-08, 1.224305e-08, 1.063864e-08, 9.039391e-09, 7.613683e-09, 
    6.32007e-09, 5.284171e-09, 4.556218e-09, 4.005142e-09, 3.503404e-09,
  1.999469e-08, 1.913225e-08, 1.836268e-08, 1.747034e-08, 1.633752e-08, 
    1.504673e-08, 1.365309e-08, 1.217889e-08, 1.060499e-08, 9.063542e-09, 
    7.726919e-09, 6.545803e-09, 5.574881e-09, 4.850657e-09, 4.295545e-09,
  2.122994e-08, 2.078519e-08, 1.925145e-08, 1.587656e-08, 1.456786e-08, 
    1.330176e-08, 1.196376e-08, 1.025493e-08, 8.63334e-09, 7.246589e-09, 
    6.090447e-09, 5.384164e-09, 4.31862e-09, 3.318799e-09, 2.574035e-09,
  2.234961e-08, 2.134644e-08, 1.985031e-08, 1.736304e-08, 1.516692e-08, 
    1.389695e-08, 1.263587e-08, 1.102358e-08, 9.418818e-09, 7.876434e-09, 
    6.617848e-09, 5.701457e-09, 4.867433e-09, 3.849248e-09, 2.987857e-09,
  2.353164e-08, 2.205831e-08, 2.056705e-08, 1.851161e-08, 1.599952e-08, 
    1.44581e-08, 1.329398e-08, 1.188335e-08, 1.027367e-08, 8.651623e-09, 
    7.264655e-09, 6.194671e-09, 5.360079e-09, 4.431809e-09, 3.476795e-09,
  2.379836e-08, 2.349253e-08, 2.087562e-08, 1.93476e-08, 1.710371e-08, 
    1.510164e-08, 1.37994e-08, 1.260602e-08, 1.11139e-08, 9.547467e-09, 
    7.950035e-09, 6.748421e-09, 5.790251e-09, 4.989914e-09, 4.047001e-09,
  2.347354e-08, 2.436389e-08, 2.198528e-08, 1.980012e-08, 1.820287e-08, 
    1.599156e-08, 1.44272e-08, 1.31602e-08, 1.185868e-08, 1.040818e-08, 
    8.829375e-09, 7.353608e-09, 6.297779e-09, 5.377786e-09, 4.582614e-09,
  2.325763e-08, 2.460114e-08, 2.351139e-08, 2.013999e-08, 1.891253e-08, 
    1.710559e-08, 1.51767e-08, 1.373576e-08, 1.242761e-08, 1.114299e-08, 
    9.718479e-09, 8.148078e-09, 6.854742e-09, 5.863343e-09, 4.998519e-09,
  2.287318e-08, 2.400252e-08, 2.4359e-08, 2.102572e-08, 1.924338e-08, 
    1.788491e-08, 1.614214e-08, 1.437431e-08, 1.297189e-08, 1.166787e-08, 
    1.043466e-08, 9.027574e-09, 7.541788e-09, 6.37625e-09, 5.455066e-09,
  2.237602e-08, 2.319574e-08, 2.432179e-08, 2.227904e-08, 1.943221e-08, 
    1.839653e-08, 1.693103e-08, 1.517729e-08, 1.355572e-08, 1.218685e-08, 
    1.098093e-08, 9.738444e-09, 8.372689e-09, 6.979965e-09, 5.952138e-09,
  2.163569e-08, 2.244046e-08, 2.354092e-08, 2.328269e-08, 1.99378e-08, 
    1.852989e-08, 1.757734e-08, 1.602028e-08, 1.417474e-08, 1.265951e-08, 
    1.147717e-08, 1.032002e-08, 9.124824e-09, 7.741041e-09, 6.496673e-09,
  2.091064e-08, 2.166054e-08, 2.275317e-08, 2.318587e-08, 2.0915e-08, 
    1.860389e-08, 1.794188e-08, 1.685862e-08, 1.49345e-08, 1.330969e-08, 
    1.193808e-08, 1.082194e-08, 9.691933e-09, 8.477882e-09, 7.193478e-09,
  1.849957e-08, 1.767336e-08, 1.697929e-08, 1.620297e-08, 1.533873e-08, 
    1.455548e-08, 1.351343e-08, 1.266412e-08, 1.173636e-08, 1.059384e-08, 
    9.293225e-09, 8.232368e-09, 6.94573e-09, 5.837785e-09, 4.761389e-09,
  1.911791e-08, 1.812212e-08, 1.734024e-08, 1.66834e-08, 1.5724e-08, 
    1.487034e-08, 1.396046e-08, 1.305647e-08, 1.234899e-08, 1.145909e-08, 
    1.024674e-08, 8.955697e-09, 7.868333e-09, 6.707053e-09, 5.705494e-09,
  1.972962e-08, 1.889094e-08, 1.778081e-08, 1.708899e-08, 1.633896e-08, 
    1.53149e-08, 1.446412e-08, 1.355223e-08, 1.283265e-08, 1.223752e-08, 
    1.124388e-08, 9.99934e-09, 8.637469e-09, 7.604913e-09, 6.536342e-09,
  2.042465e-08, 1.948626e-08, 1.845178e-08, 1.742962e-08, 1.671383e-08, 
    1.592798e-08, 1.489386e-08, 1.411579e-08, 1.323651e-08, 1.27011e-08, 
    1.201834e-08, 1.096831e-08, 9.580063e-09, 8.376898e-09, 7.412609e-09,
  2.156338e-08, 2.025222e-08, 1.910749e-08, 1.796355e-08, 1.69771e-08, 
    1.632647e-08, 1.547158e-08, 1.45691e-08, 1.376529e-08, 1.304375e-08, 
    1.250666e-08, 1.180398e-08, 1.064387e-08, 9.243913e-09, 8.163926e-09,
  2.225517e-08, 2.12706e-08, 1.990402e-08, 1.868191e-08, 1.74275e-08, 
    1.659526e-08, 1.59391e-08, 1.512767e-08, 1.426938e-08, 1.356091e-08, 
    1.28567e-08, 1.237017e-08, 1.150015e-08, 1.033326e-08, 8.999064e-09,
  2.295053e-08, 2.202979e-08, 2.07304e-08, 1.945284e-08, 1.810621e-08, 
    1.694923e-08, 1.62038e-08, 1.561961e-08, 1.476587e-08, 1.409047e-08, 
    1.330123e-08, 1.280003e-08, 1.21624e-08, 1.123954e-08, 1.003948e-08,
  2.37808e-08, 2.286767e-08, 2.156109e-08, 2.024703e-08, 1.900666e-08, 
    1.750277e-08, 1.650136e-08, 1.592428e-08, 1.524811e-08, 1.452355e-08, 
    1.38316e-08, 1.313104e-08, 1.260541e-08, 1.192099e-08, 1.10161e-08,
  2.438581e-08, 2.356635e-08, 2.25107e-08, 2.104241e-08, 1.982216e-08, 
    1.843202e-08, 1.688201e-08, 1.618944e-08, 1.560736e-08, 1.494591e-08, 
    1.426118e-08, 1.363874e-08, 1.289112e-08, 1.235669e-08, 1.171655e-08,
  2.465028e-08, 2.418771e-08, 2.331864e-08, 2.207201e-08, 2.056925e-08, 
    1.942647e-08, 1.768086e-08, 1.645741e-08, 1.582476e-08, 1.525942e-08, 
    1.459343e-08, 1.407474e-08, 1.340181e-08, 1.274904e-08, 1.217491e-08,
  2.098211e-08, 1.996162e-08, 1.944506e-08, 1.875781e-08, 1.881591e-08, 
    1.844981e-08, 1.757052e-08, 1.657319e-08, 1.566871e-08, 1.484351e-08, 
    1.368465e-08, 1.215181e-08, 1.087444e-08, 9.747427e-09, 8.175831e-09,
  2.095812e-08, 2.027582e-08, 1.945691e-08, 1.882146e-08, 1.870312e-08, 
    1.865658e-08, 1.813979e-08, 1.725804e-08, 1.636947e-08, 1.53897e-08, 
    1.447001e-08, 1.323539e-08, 1.171819e-08, 1.049069e-08, 9.169402e-09,
  2.079604e-08, 2.036835e-08, 1.955054e-08, 1.881011e-08, 1.856082e-08, 
    1.85704e-08, 1.843747e-08, 1.789121e-08, 1.70719e-08, 1.621476e-08, 
    1.525865e-08, 1.428071e-08, 1.291264e-08, 1.134872e-08, 1.014316e-08,
  2.041445e-08, 2.033194e-08, 1.970891e-08, 1.881551e-08, 1.841321e-08, 
    1.836193e-08, 1.841648e-08, 1.825116e-08, 1.768751e-08, 1.696572e-08, 
    1.604554e-08, 1.510056e-08, 1.405942e-08, 1.242876e-08, 1.096395e-08,
  2.013628e-08, 2.022333e-08, 1.98139e-08, 1.890181e-08, 1.826688e-08, 
    1.812999e-08, 1.828892e-08, 1.838766e-08, 1.810695e-08, 1.762158e-08, 
    1.684244e-08, 1.590042e-08, 1.496705e-08, 1.366612e-08, 1.189588e-08,
  2.007365e-08, 2.020944e-08, 1.978053e-08, 1.903865e-08, 1.824613e-08, 
    1.788675e-08, 1.791454e-08, 1.822781e-08, 1.819309e-08, 1.80188e-08, 
    1.754864e-08, 1.672037e-08, 1.576652e-08, 1.473161e-08, 1.309908e-08,
  2.040918e-08, 2.027148e-08, 1.975893e-08, 1.912337e-08, 1.830254e-08, 
    1.778619e-08, 1.761861e-08, 1.792136e-08, 1.811522e-08, 1.81264e-08, 
    1.796604e-08, 1.738803e-08, 1.653331e-08, 1.558248e-08, 1.425707e-08,
  2.089828e-08, 2.055989e-08, 1.983727e-08, 1.921509e-08, 1.840841e-08, 
    1.778751e-08, 1.741654e-08, 1.753854e-08, 1.790324e-08, 1.805421e-08, 
    1.809388e-08, 1.785156e-08, 1.710821e-08, 1.638617e-08, 1.511024e-08,
  2.143351e-08, 2.095895e-08, 2.00783e-08, 1.934623e-08, 1.861927e-08, 
    1.789805e-08, 1.739556e-08, 1.728588e-08, 1.76742e-08, 1.795664e-08, 
    1.807425e-08, 1.80236e-08, 1.759137e-08, 1.693476e-08, 1.592893e-08,
  2.198887e-08, 2.151354e-08, 2.03436e-08, 1.954312e-08, 1.883877e-08, 
    1.813699e-08, 1.739955e-08, 1.719824e-08, 1.745582e-08, 1.786174e-08, 
    1.80789e-08, 1.816289e-08, 1.787155e-08, 1.741206e-08, 1.666368e-08,
  2.360514e-08, 2.224435e-08, 2.142441e-08, 2.061263e-08, 2.030612e-08, 
    1.991977e-08, 1.985971e-08, 1.915396e-08, 1.852161e-08, 1.824659e-08, 
    1.767016e-08, 1.716359e-08, 1.688062e-08, 1.618709e-08, 1.558305e-08,
  2.44828e-08, 2.296809e-08, 2.191407e-08, 2.096093e-08, 2.054992e-08, 
    2.017584e-08, 2.000195e-08, 1.990708e-08, 1.931164e-08, 1.845081e-08, 
    1.788412e-08, 1.728298e-08, 1.710393e-08, 1.659469e-08, 1.605545e-08,
  2.540103e-08, 2.359892e-08, 2.245536e-08, 2.155254e-08, 2.078873e-08, 
    2.071241e-08, 2.031218e-08, 2.064833e-08, 2.032119e-08, 1.887971e-08, 
    1.812297e-08, 1.747861e-08, 1.725157e-08, 1.694299e-08, 1.642448e-08,
  2.663837e-08, 2.448406e-08, 2.290094e-08, 2.214449e-08, 2.13292e-08, 
    2.129471e-08, 2.096671e-08, 2.134656e-08, 2.125021e-08, 1.94475e-08, 
    1.841487e-08, 1.764761e-08, 1.71942e-08, 1.720535e-08, 1.661532e-08,
  2.753829e-08, 2.567135e-08, 2.366603e-08, 2.265361e-08, 2.188052e-08, 
    2.188521e-08, 2.164256e-08, 2.20105e-08, 2.220066e-08, 1.992094e-08, 
    1.860677e-08, 1.785905e-08, 1.715766e-08, 1.719354e-08, 1.679775e-08,
  2.759782e-08, 2.647523e-08, 2.47085e-08, 2.320209e-08, 2.236882e-08, 
    2.242605e-08, 2.237877e-08, 2.271839e-08, 2.274722e-08, 2.031372e-08, 
    1.867273e-08, 1.790453e-08, 1.709465e-08, 1.70079e-08, 1.682099e-08,
  2.747115e-08, 2.688028e-08, 2.545432e-08, 2.394478e-08, 2.275413e-08, 
    2.280645e-08, 2.290046e-08, 2.37497e-08, 2.31099e-08, 2.032316e-08, 
    1.8689e-08, 1.789188e-08, 1.704127e-08, 1.673377e-08, 1.673789e-08,
  2.789168e-08, 2.690263e-08, 2.590783e-08, 2.456619e-08, 2.322175e-08, 
    2.305744e-08, 2.331806e-08, 2.446409e-08, 2.342759e-08, 1.999884e-08, 
    1.851317e-08, 1.775774e-08, 1.688075e-08, 1.644651e-08, 1.648811e-08,
  2.871527e-08, 2.716688e-08, 2.631731e-08, 2.513192e-08, 2.363639e-08, 
    2.316805e-08, 2.34901e-08, 2.489699e-08, 2.357557e-08, 1.952373e-08, 
    1.820386e-08, 1.764073e-08, 1.679482e-08, 1.624731e-08, 1.617179e-08,
  2.93973e-08, 2.755809e-08, 2.65253e-08, 2.566545e-08, 2.408834e-08, 
    2.334319e-08, 2.349595e-08, 2.521964e-08, 2.362985e-08, 1.914603e-08, 
    1.786468e-08, 1.743546e-08, 1.673452e-08, 1.61537e-08, 1.592919e-08,
  1.519873e-08, 1.43176e-08, 1.359786e-08, 1.323305e-08, 1.311358e-08, 
    1.311772e-08, 1.317325e-08, 1.324844e-08, 1.32757e-08, 1.272673e-08, 
    1.198773e-08, 1.140457e-08, 1.097203e-08, 1.04968e-08, 1.016049e-08,
  1.524587e-08, 1.445757e-08, 1.386067e-08, 1.354041e-08, 1.340574e-08, 
    1.335659e-08, 1.353908e-08, 1.359377e-08, 1.371867e-08, 1.339014e-08, 
    1.271347e-08, 1.20703e-08, 1.162638e-08, 1.102373e-08, 1.06627e-08,
  1.538647e-08, 1.47117e-08, 1.421811e-08, 1.389036e-08, 1.375736e-08, 
    1.366741e-08, 1.379029e-08, 1.407027e-08, 1.413988e-08, 1.401636e-08, 
    1.341066e-08, 1.275306e-08, 1.227832e-08, 1.1739e-08, 1.119054e-08,
  1.573409e-08, 1.496704e-08, 1.443073e-08, 1.406019e-08, 1.387312e-08, 
    1.38025e-08, 1.384909e-08, 1.432979e-08, 1.451149e-08, 1.454801e-08, 
    1.403256e-08, 1.347656e-08, 1.296658e-08, 1.246122e-08, 1.179616e-08,
  1.625806e-08, 1.535681e-08, 1.464251e-08, 1.412002e-08, 1.387609e-08, 
    1.389881e-08, 1.396749e-08, 1.45454e-08, 1.491558e-08, 1.497853e-08, 
    1.46397e-08, 1.405563e-08, 1.366624e-08, 1.327533e-08, 1.259963e-08,
  1.692421e-08, 1.584365e-08, 1.492707e-08, 1.420247e-08, 1.387633e-08, 
    1.396633e-08, 1.413638e-08, 1.474227e-08, 1.54636e-08, 1.541841e-08, 
    1.51875e-08, 1.46535e-08, 1.42427e-08, 1.395847e-08, 1.349743e-08,
  1.764111e-08, 1.644319e-08, 1.535378e-08, 1.438909e-08, 1.400844e-08, 
    1.408807e-08, 1.441218e-08, 1.495365e-08, 1.597336e-08, 1.611434e-08, 
    1.576452e-08, 1.524753e-08, 1.482209e-08, 1.455408e-08, 1.41837e-08,
  1.816459e-08, 1.707237e-08, 1.586315e-08, 1.46586e-08, 1.422063e-08, 
    1.423921e-08, 1.470665e-08, 1.538126e-08, 1.650299e-08, 1.690217e-08, 
    1.64789e-08, 1.590066e-08, 1.547073e-08, 1.516246e-08, 1.474039e-08,
  1.851948e-08, 1.766349e-08, 1.646596e-08, 1.504226e-08, 1.449325e-08, 
    1.449583e-08, 1.497791e-08, 1.580361e-08, 1.714455e-08, 1.765205e-08, 
    1.728168e-08, 1.670189e-08, 1.611152e-08, 1.588265e-08, 1.533678e-08,
  1.881458e-08, 1.812199e-08, 1.701915e-08, 1.562772e-08, 1.483583e-08, 
    1.481067e-08, 1.527577e-08, 1.628966e-08, 1.796652e-08, 1.832029e-08, 
    1.811003e-08, 1.760597e-08, 1.684929e-08, 1.640292e-08, 1.59371e-08,
  2.169985e-08, 2.110752e-08, 2.073832e-08, 2.057706e-08, 1.985264e-08, 
    1.852285e-08, 1.732483e-08, 1.566889e-08, 1.374136e-08, 1.176136e-08, 
    1.016056e-08, 8.883958e-09, 7.917853e-09, 6.751664e-09, 5.533999e-09,
  2.196516e-08, 2.111042e-08, 2.053075e-08, 2.031574e-08, 1.957553e-08, 
    1.830726e-08, 1.719589e-08, 1.561635e-08, 1.356924e-08, 1.15825e-08, 
    1.009141e-08, 8.915112e-09, 7.926761e-09, 6.799554e-09, 5.594177e-09,
  2.208121e-08, 2.112103e-08, 2.039173e-08, 2.004825e-08, 1.921363e-08, 
    1.800121e-08, 1.702734e-08, 1.553531e-08, 1.345721e-08, 1.150479e-08, 
    1.009464e-08, 8.980471e-09, 7.987365e-09, 6.902088e-09, 5.71646e-09,
  2.213025e-08, 2.109359e-08, 2.024214e-08, 1.978097e-08, 1.885594e-08, 
    1.760717e-08, 1.672306e-08, 1.534533e-08, 1.337059e-08, 1.145857e-08, 
    1.011855e-08, 9.065886e-09, 8.072775e-09, 6.999266e-09, 5.849976e-09,
  2.206691e-08, 2.100565e-08, 2.007464e-08, 1.949995e-08, 1.8601e-08, 
    1.726477e-08, 1.633085e-08, 1.509033e-08, 1.3254e-08, 1.14423e-08, 
    1.019545e-08, 9.163988e-09, 8.156165e-09, 7.122153e-09, 6.01283e-09,
  2.189463e-08, 2.087428e-08, 1.990567e-08, 1.926942e-08, 1.834858e-08, 
    1.695739e-08, 1.593576e-08, 1.48003e-08, 1.318327e-08, 1.145895e-08, 
    1.02365e-08, 9.223905e-09, 8.226727e-09, 7.257651e-09, 6.185092e-09,
  2.171932e-08, 2.07019e-08, 1.973542e-08, 1.899691e-08, 1.809931e-08, 
    1.667177e-08, 1.559409e-08, 1.450765e-08, 1.307317e-08, 1.151088e-08, 
    1.031226e-08, 9.274145e-09, 8.314378e-09, 7.407757e-09, 6.400271e-09,
  2.154696e-08, 2.055694e-08, 1.955384e-08, 1.875483e-08, 1.783103e-08, 
    1.641591e-08, 1.521625e-08, 1.425454e-08, 1.29494e-08, 1.154132e-08, 
    1.036249e-08, 9.368009e-09, 8.42319e-09, 7.590294e-09, 6.653718e-09,
  2.145137e-08, 2.044071e-08, 1.941206e-08, 1.850557e-08, 1.757157e-08, 
    1.61561e-08, 1.492255e-08, 1.398052e-08, 1.281626e-08, 1.154519e-08, 
    1.04362e-08, 9.46207e-09, 8.576652e-09, 7.781531e-09, 6.947586e-09,
  2.142416e-08, 2.039225e-08, 1.929287e-08, 1.825546e-08, 1.726239e-08, 
    1.587921e-08, 1.463378e-08, 1.36779e-08, 1.263265e-08, 1.149774e-08, 
    1.047461e-08, 9.558474e-09, 8.729406e-09, 7.984721e-09, 7.256465e-09,
  1.822964e-08, 1.75469e-08, 1.71195e-08, 1.681833e-08, 1.631446e-08, 
    1.595396e-08, 1.596569e-08, 1.612052e-08, 1.647891e-08, 1.661487e-08, 
    1.65823e-08, 1.601422e-08, 1.483993e-08, 1.340682e-08, 1.188675e-08,
  1.83662e-08, 1.769915e-08, 1.711174e-08, 1.703929e-08, 1.67083e-08, 
    1.638802e-08, 1.642826e-08, 1.663722e-08, 1.694793e-08, 1.696452e-08, 
    1.680793e-08, 1.615641e-08, 1.487077e-08, 1.330826e-08, 1.16778e-08,
  1.846579e-08, 1.789346e-08, 1.721192e-08, 1.722861e-08, 1.708086e-08, 
    1.681664e-08, 1.68756e-08, 1.720496e-08, 1.753511e-08, 1.739721e-08, 
    1.705186e-08, 1.628874e-08, 1.48867e-08, 1.324116e-08, 1.149244e-08,
  1.859954e-08, 1.812739e-08, 1.740837e-08, 1.739925e-08, 1.742759e-08, 
    1.718588e-08, 1.728109e-08, 1.777629e-08, 1.810013e-08, 1.781303e-08, 
    1.727581e-08, 1.632779e-08, 1.489545e-08, 1.317516e-08, 1.132378e-08,
  1.883602e-08, 1.835604e-08, 1.766157e-08, 1.763358e-08, 1.772789e-08, 
    1.755491e-08, 1.77373e-08, 1.831762e-08, 1.863619e-08, 1.822719e-08, 
    1.755516e-08, 1.643157e-08, 1.486343e-08, 1.312951e-08, 1.117822e-08,
  1.919123e-08, 1.864635e-08, 1.791286e-08, 1.789265e-08, 1.813441e-08, 
    1.796069e-08, 1.819552e-08, 1.881416e-08, 1.912336e-08, 1.857914e-08, 
    1.77343e-08, 1.65192e-08, 1.48912e-08, 1.308843e-08, 1.104435e-08,
  1.951474e-08, 1.895236e-08, 1.813424e-08, 1.812499e-08, 1.861025e-08, 
    1.850466e-08, 1.868856e-08, 1.933461e-08, 1.961771e-08, 1.883103e-08, 
    1.793673e-08, 1.664352e-08, 1.497242e-08, 1.306707e-08, 1.093167e-08,
  1.986973e-08, 1.918519e-08, 1.832617e-08, 1.826476e-08, 1.905299e-08, 
    1.904988e-08, 1.917941e-08, 1.978823e-08, 2.014635e-08, 1.904888e-08, 
    1.801135e-08, 1.675523e-08, 1.50784e-08, 1.308847e-08, 1.085145e-08,
  2.00249e-08, 1.936877e-08, 1.852098e-08, 1.829734e-08, 1.93218e-08, 
    1.960972e-08, 1.969351e-08, 2.022056e-08, 2.056898e-08, 1.929606e-08, 
    1.80227e-08, 1.683086e-08, 1.518934e-08, 1.31736e-08, 1.08323e-08,
  2.009938e-08, 1.944255e-08, 1.86942e-08, 1.840062e-08, 1.936211e-08, 
    1.99574e-08, 2.010961e-08, 2.057305e-08, 2.092253e-08, 1.955138e-08, 
    1.800062e-08, 1.676819e-08, 1.525875e-08, 1.329459e-08, 1.086854e-08,
  1.681168e-08, 1.784068e-08, 1.839645e-08, 1.864873e-08, 1.894678e-08, 
    1.893686e-08, 1.863599e-08, 1.812716e-08, 1.812221e-08, 1.76238e-08, 
    1.641089e-08, 1.546899e-08, 1.444227e-08, 1.424241e-08, 1.401051e-08,
  1.709271e-08, 1.812189e-08, 1.881756e-08, 1.897753e-08, 1.934548e-08, 
    1.91856e-08, 1.877804e-08, 1.803872e-08, 1.774339e-08, 1.746676e-08, 
    1.628226e-08, 1.540266e-08, 1.430958e-08, 1.386355e-08, 1.373511e-08,
  1.71536e-08, 1.844817e-08, 1.934515e-08, 1.932441e-08, 1.966253e-08, 
    1.938846e-08, 1.889476e-08, 1.80399e-08, 1.754049e-08, 1.714867e-08, 
    1.610415e-08, 1.526206e-08, 1.416288e-08, 1.350778e-08, 1.338579e-08,
  1.721178e-08, 1.870887e-08, 1.982261e-08, 1.970253e-08, 1.986486e-08, 
    1.960933e-08, 1.90133e-08, 1.794011e-08, 1.730394e-08, 1.69131e-08, 
    1.586703e-08, 1.505314e-08, 1.398931e-08, 1.315184e-08, 1.295229e-08,
  1.733684e-08, 1.896044e-08, 2.043379e-08, 2.018431e-08, 2.005851e-08, 
    1.968138e-08, 1.908341e-08, 1.792872e-08, 1.712633e-08, 1.663237e-08, 
    1.569499e-08, 1.477701e-08, 1.376102e-08, 1.282983e-08, 1.24772e-08,
  1.760809e-08, 1.909807e-08, 2.094433e-08, 2.080358e-08, 2.034655e-08, 
    1.975993e-08, 1.910065e-08, 1.785307e-08, 1.687851e-08, 1.638561e-08, 
    1.55406e-08, 1.461482e-08, 1.357316e-08, 1.255651e-08, 1.204865e-08,
  1.783966e-08, 1.931661e-08, 2.135942e-08, 2.135729e-08, 2.069018e-08, 
    1.978501e-08, 1.904146e-08, 1.7695e-08, 1.65407e-08, 1.609199e-08, 
    1.537058e-08, 1.45087e-08, 1.343164e-08, 1.234183e-08, 1.164953e-08,
  1.812147e-08, 1.94834e-08, 2.158623e-08, 2.184111e-08, 2.10251e-08, 
    1.988e-08, 1.888e-08, 1.75675e-08, 1.61828e-08, 1.568928e-08, 
    1.523377e-08, 1.448574e-08, 1.335322e-08, 1.225017e-08, 1.136669e-08,
  1.841541e-08, 1.960174e-08, 2.169291e-08, 2.209541e-08, 2.120786e-08, 
    2.005216e-08, 1.881243e-08, 1.74358e-08, 1.591241e-08, 1.527425e-08, 
    1.505033e-08, 1.443387e-08, 1.341689e-08, 1.217927e-08, 1.115717e-08,
  1.866133e-08, 1.978201e-08, 2.168594e-08, 2.222519e-08, 2.120022e-08, 
    2.0053e-08, 1.883798e-08, 1.739131e-08, 1.582288e-08, 1.493861e-08, 
    1.486437e-08, 1.447474e-08, 1.352041e-08, 1.229815e-08, 1.108779e-08,
  1.922452e-08, 1.898968e-08, 1.870964e-08, 1.836667e-08, 1.824284e-08, 
    1.820317e-08, 1.825167e-08, 1.836117e-08, 1.864306e-08, 1.825292e-08, 
    1.770323e-08, 1.733338e-08, 1.744724e-08, 1.753143e-08, 1.651301e-08,
  1.916344e-08, 1.893414e-08, 1.871824e-08, 1.839831e-08, 1.81611e-08, 
    1.786937e-08, 1.791168e-08, 1.797435e-08, 1.839189e-08, 1.825795e-08, 
    1.766035e-08, 1.714814e-08, 1.723688e-08, 1.739814e-08, 1.670743e-08,
  1.901448e-08, 1.869233e-08, 1.842708e-08, 1.81251e-08, 1.78587e-08, 
    1.760732e-08, 1.769262e-08, 1.768642e-08, 1.807484e-08, 1.826792e-08, 
    1.788517e-08, 1.724683e-08, 1.716946e-08, 1.727862e-08, 1.686215e-08,
  1.860551e-08, 1.815278e-08, 1.777743e-08, 1.761165e-08, 1.751669e-08, 
    1.736583e-08, 1.748211e-08, 1.752946e-08, 1.787305e-08, 1.823367e-08, 
    1.79926e-08, 1.744884e-08, 1.720916e-08, 1.712093e-08, 1.700485e-08,
  1.779635e-08, 1.736638e-08, 1.704978e-08, 1.696876e-08, 1.709053e-08, 
    1.717522e-08, 1.739114e-08, 1.755217e-08, 1.773736e-08, 1.810724e-08, 
    1.811199e-08, 1.766784e-08, 1.731159e-08, 1.700643e-08, 1.686849e-08,
  1.68852e-08, 1.643205e-08, 1.622735e-08, 1.63813e-08, 1.673071e-08, 
    1.707979e-08, 1.743832e-08, 1.762979e-08, 1.767821e-08, 1.783743e-08, 
    1.798986e-08, 1.780168e-08, 1.739195e-08, 1.697675e-08, 1.674594e-08,
  1.583405e-08, 1.557834e-08, 1.564166e-08, 1.600762e-08, 1.650211e-08, 
    1.713656e-08, 1.770242e-08, 1.788934e-08, 1.76818e-08, 1.767337e-08, 
    1.772966e-08, 1.775183e-08, 1.744939e-08, 1.684601e-08, 1.65021e-08,
  1.515656e-08, 1.505614e-08, 1.532499e-08, 1.600552e-08, 1.663562e-08, 
    1.715934e-08, 1.781198e-08, 1.834375e-08, 1.812671e-08, 1.771877e-08, 
    1.743206e-08, 1.759285e-08, 1.738181e-08, 1.687787e-08, 1.636168e-08,
  1.476925e-08, 1.47921e-08, 1.517055e-08, 1.618525e-08, 1.702036e-08, 
    1.765069e-08, 1.824018e-08, 1.883457e-08, 1.883955e-08, 1.826327e-08, 
    1.762831e-08, 1.740369e-08, 1.737154e-08, 1.681567e-08, 1.62088e-08,
  1.467922e-08, 1.453731e-08, 1.49748e-08, 1.643212e-08, 1.774968e-08, 
    1.836172e-08, 1.901667e-08, 1.945828e-08, 1.962703e-08, 1.882324e-08, 
    1.779486e-08, 1.754236e-08, 1.727821e-08, 1.689748e-08, 1.617383e-08,
  2.544691e-08, 2.514843e-08, 2.394611e-08, 2.285967e-08, 2.17002e-08, 
    2.065595e-08, 2.021924e-08, 2.054143e-08, 2.099688e-08, 2.140904e-08, 
    2.145802e-08, 2.02033e-08, 1.942049e-08, 1.982994e-08, 2.092484e-08,
  2.623772e-08, 2.502475e-08, 2.426879e-08, 2.350709e-08, 2.247657e-08, 
    2.139063e-08, 2.072186e-08, 2.037388e-08, 2.056465e-08, 2.079913e-08, 
    2.094566e-08, 1.997795e-08, 1.920175e-08, 1.93813e-08, 2.053847e-08,
  2.762015e-08, 2.562403e-08, 2.452733e-08, 2.352195e-08, 2.297271e-08, 
    2.222199e-08, 2.133677e-08, 2.057105e-08, 2.052344e-08, 2.055582e-08, 
    2.055706e-08, 1.985692e-08, 1.91758e-08, 1.910199e-08, 2.00164e-08,
  2.719577e-08, 2.660608e-08, 2.542852e-08, 2.36524e-08, 2.265394e-08, 
    2.224629e-08, 2.168462e-08, 2.096519e-08, 2.059309e-08, 2.041677e-08, 
    2.006714e-08, 1.964899e-08, 1.918825e-08, 1.905274e-08, 1.961902e-08,
  2.646557e-08, 2.621579e-08, 2.602574e-08, 2.419368e-08, 2.242586e-08, 
    2.179551e-08, 2.152658e-08, 2.094196e-08, 2.037558e-08, 2.012175e-08, 
    1.969024e-08, 1.948557e-08, 1.919378e-08, 1.904153e-08, 1.938425e-08,
  2.612786e-08, 2.547487e-08, 2.566062e-08, 2.450787e-08, 2.25739e-08, 
    2.140511e-08, 2.087943e-08, 2.055463e-08, 2.016253e-08, 1.988642e-08, 
    1.945301e-08, 1.93893e-08, 1.922245e-08, 1.913092e-08, 1.937319e-08,
  2.571192e-08, 2.491356e-08, 2.475544e-08, 2.406142e-08, 2.262267e-08, 
    2.137267e-08, 2.055756e-08, 2.036998e-08, 1.994678e-08, 1.970153e-08, 
    1.953761e-08, 1.942654e-08, 1.927891e-08, 1.920373e-08, 1.947499e-08,
  2.499784e-08, 2.435972e-08, 2.344312e-08, 2.317532e-08, 2.217869e-08, 
    2.144788e-08, 2.069626e-08, 2.021455e-08, 1.973529e-08, 1.955753e-08, 
    2.000573e-08, 1.993562e-08, 1.944594e-08, 1.925586e-08, 1.951268e-08,
  2.44015e-08, 2.366747e-08, 2.261227e-08, 2.215799e-08, 2.159799e-08, 
    2.112396e-08, 2.068635e-08, 2.025873e-08, 1.978635e-08, 1.944578e-08, 
    2.002537e-08, 2.013062e-08, 1.96312e-08, 1.934405e-08, 1.938831e-08,
  2.422432e-08, 2.314935e-08, 2.210892e-08, 2.151797e-08, 2.09262e-08, 
    2.046174e-08, 2.009632e-08, 1.984639e-08, 1.960133e-08, 1.927793e-08, 
    1.942507e-08, 2.003455e-08, 1.963457e-08, 1.950881e-08, 1.937523e-08,
  2.248211e-08, 2.072554e-08, 1.91139e-08, 1.742793e-08, 1.572701e-08, 
    1.430228e-08, 1.302434e-08, 1.233087e-08, 1.256085e-08, 1.310992e-08, 
    1.494377e-08, 1.688935e-08, 1.64768e-08, 1.483623e-08, 1.433406e-08,
  2.283199e-08, 2.16041e-08, 2.000411e-08, 1.847151e-08, 1.694225e-08, 
    1.548399e-08, 1.432183e-08, 1.321133e-08, 1.305016e-08, 1.31287e-08, 
    1.453331e-08, 1.66729e-08, 1.684126e-08, 1.558656e-08, 1.485167e-08,
  2.383637e-08, 2.211212e-08, 2.06515e-08, 1.934275e-08, 1.805469e-08, 
    1.664919e-08, 1.554243e-08, 1.449534e-08, 1.405384e-08, 1.40108e-08, 
    1.470319e-08, 1.683694e-08, 1.702711e-08, 1.62472e-08, 1.532654e-08,
  2.459844e-08, 2.340508e-08, 2.156831e-08, 1.986231e-08, 1.882638e-08, 
    1.772604e-08, 1.680647e-08, 1.594633e-08, 1.557265e-08, 1.543413e-08, 
    1.574163e-08, 1.715477e-08, 1.751889e-08, 1.677851e-08, 1.578757e-08,
  2.440471e-08, 2.415358e-08, 2.294399e-08, 2.10306e-08, 1.936911e-08, 
    1.838138e-08, 1.764915e-08, 1.708099e-08, 1.687354e-08, 1.67662e-08, 
    1.673649e-08, 1.740656e-08, 1.78225e-08, 1.728228e-08, 1.623754e-08,
  2.315428e-08, 2.440091e-08, 2.375447e-08, 2.244075e-08, 2.052331e-08, 
    1.90939e-08, 1.832953e-08, 1.796083e-08, 1.776542e-08, 1.800877e-08, 
    1.795297e-08, 1.780368e-08, 1.816987e-08, 1.768144e-08, 1.651766e-08,
  2.247874e-08, 2.343305e-08, 2.390121e-08, 2.31795e-08, 2.174679e-08, 
    1.999175e-08, 1.891804e-08, 1.845393e-08, 1.834979e-08, 1.85161e-08, 
    1.860268e-08, 1.822287e-08, 1.836184e-08, 1.824854e-08, 1.704814e-08,
  2.245986e-08, 2.287469e-08, 2.343346e-08, 2.351598e-08, 2.259592e-08, 
    2.111814e-08, 1.974935e-08, 1.901812e-08, 1.875911e-08, 1.872326e-08, 
    1.852767e-08, 1.851464e-08, 1.846856e-08, 1.868439e-08, 1.776326e-08,
  2.255423e-08, 2.253622e-08, 2.296787e-08, 2.326899e-08, 2.279435e-08, 
    2.184011e-08, 2.061936e-08, 1.958432e-08, 1.90199e-08, 1.887376e-08, 
    1.859257e-08, 1.873358e-08, 1.856838e-08, 1.88865e-08, 1.866653e-08,
  2.291185e-08, 2.239346e-08, 2.254903e-08, 2.28544e-08, 2.268077e-08, 
    2.219815e-08, 2.155519e-08, 2.06767e-08, 1.996942e-08, 1.963152e-08, 
    1.943785e-08, 1.92365e-08, 1.905051e-08, 1.896743e-08, 1.930358e-08,
  2.397799e-08, 2.3942e-08, 2.393953e-08, 2.34565e-08, 2.238156e-08, 
    2.098488e-08, 1.999533e-08, 1.899262e-08, 1.770817e-08, 1.772388e-08, 
    1.836303e-08, 1.893905e-08, 1.835008e-08, 1.670499e-08, 1.565531e-08,
  2.61325e-08, 2.413654e-08, 2.390526e-08, 2.374691e-08, 2.269396e-08, 
    2.126392e-08, 2.0082e-08, 1.947765e-08, 1.8395e-08, 1.768585e-08, 
    1.801711e-08, 1.878033e-08, 1.863436e-08, 1.733947e-08, 1.589992e-08,
  2.680712e-08, 2.54828e-08, 2.381172e-08, 2.360364e-08, 2.304583e-08, 
    2.184567e-08, 2.019372e-08, 1.925681e-08, 1.892525e-08, 1.824251e-08, 
    1.767749e-08, 1.870818e-08, 1.849241e-08, 1.79292e-08, 1.616554e-08,
  2.624183e-08, 2.587036e-08, 2.468844e-08, 2.366982e-08, 2.307509e-08, 
    2.25023e-08, 2.108961e-08, 1.926017e-08, 1.827362e-08, 1.834203e-08, 
    1.7889e-08, 1.850744e-08, 1.868464e-08, 1.812229e-08, 1.652302e-08,
  2.557287e-08, 2.599589e-08, 2.510986e-08, 2.429823e-08, 2.325654e-08, 
    2.231092e-08, 2.183904e-08, 2.010254e-08, 1.818723e-08, 1.760227e-08, 
    1.778026e-08, 1.799008e-08, 1.886111e-08, 1.843717e-08, 1.692294e-08,
  2.511039e-08, 2.565649e-08, 2.53966e-08, 2.455169e-08, 2.362961e-08, 
    2.259143e-08, 2.160553e-08, 2.088343e-08, 1.891671e-08, 1.754241e-08, 
    1.72281e-08, 1.76899e-08, 1.861106e-08, 1.878045e-08, 1.734288e-08,
  2.492983e-08, 2.537135e-08, 2.534889e-08, 2.464145e-08, 2.367582e-08, 
    2.278961e-08, 2.1626e-08, 2.089632e-08, 1.963658e-08, 1.808911e-08, 
    1.72367e-08, 1.72923e-08, 1.792292e-08, 1.892897e-08, 1.7659e-08,
  2.48152e-08, 2.504705e-08, 2.515953e-08, 2.454192e-08, 2.359271e-08, 
    2.279957e-08, 2.175979e-08, 2.070819e-08, 1.990225e-08, 1.854958e-08, 
    1.749529e-08, 1.708574e-08, 1.748028e-08, 1.844492e-08, 1.777437e-08,
  2.450134e-08, 2.472625e-08, 2.484434e-08, 2.432907e-08, 2.337103e-08, 
    2.257042e-08, 2.156336e-08, 2.052978e-08, 1.968996e-08, 1.862664e-08, 
    1.766502e-08, 1.705107e-08, 1.705624e-08, 1.782994e-08, 1.768103e-08,
  2.428001e-08, 2.444682e-08, 2.456805e-08, 2.41114e-08, 2.318953e-08, 
    2.23544e-08, 2.142293e-08, 2.03146e-08, 1.949617e-08, 1.861451e-08, 
    1.760461e-08, 1.707261e-08, 1.670263e-08, 1.705535e-08, 1.720437e-08,
  1.755446e-08, 1.509694e-08, 1.589814e-08, 1.668573e-08, 1.584891e-08, 
    1.407288e-08, 1.316189e-08, 1.241945e-08, 1.164178e-08, 1.120455e-08, 
    1.028729e-08, 1.025073e-08, 1.069957e-08, 1.282204e-08, 1.453147e-08,
  1.978866e-08, 1.97992e-08, 1.630937e-08, 1.573368e-08, 1.65846e-08, 
    1.673416e-08, 1.518859e-08, 1.400064e-08, 1.24879e-08, 1.188363e-08, 
    1.100281e-08, 1.073161e-08, 1.11951e-08, 1.139907e-08, 1.405987e-08,
  2.040401e-08, 2.018736e-08, 2.080301e-08, 1.770841e-08, 1.606373e-08, 
    1.68442e-08, 1.761239e-08, 1.69997e-08, 1.465611e-08, 1.273959e-08, 
    1.22164e-08, 1.115764e-08, 1.13559e-08, 1.215672e-08, 1.269933e-08,
  2.387605e-08, 2.204929e-08, 2.101774e-08, 2.130405e-08, 1.903705e-08, 
    1.660566e-08, 1.696254e-08, 1.793611e-08, 1.832305e-08, 1.597932e-08, 
    1.368234e-08, 1.262297e-08, 1.166204e-08, 1.23906e-08, 1.283321e-08,
  2.531772e-08, 2.449413e-08, 2.304494e-08, 2.209803e-08, 2.207718e-08, 
    2.025052e-08, 1.725971e-08, 1.676299e-08, 1.777179e-08, 1.862853e-08, 
    1.742102e-08, 1.499364e-08, 1.32971e-08, 1.264513e-08, 1.326744e-08,
  2.554353e-08, 2.520164e-08, 2.458125e-08, 2.383719e-08, 2.282645e-08, 
    2.259889e-08, 2.130654e-08, 1.810638e-08, 1.654865e-08, 1.752488e-08, 
    1.861851e-08, 1.842772e-08, 1.617386e-08, 1.401504e-08, 1.368811e-08,
  2.564816e-08, 2.539656e-08, 2.515169e-08, 2.487044e-08, 2.432273e-08, 
    2.319392e-08, 2.309311e-08, 2.201626e-08, 1.878225e-08, 1.650377e-08, 
    1.744719e-08, 1.855775e-08, 1.872379e-08, 1.711443e-08, 1.47623e-08,
  2.592366e-08, 2.558629e-08, 2.525972e-08, 2.524536e-08, 2.521861e-08, 
    2.449978e-08, 2.341222e-08, 2.323539e-08, 2.236536e-08, 1.944961e-08, 
    1.680278e-08, 1.738475e-08, 1.829968e-08, 1.871063e-08, 1.716169e-08,
  2.560235e-08, 2.565081e-08, 2.558157e-08, 2.539704e-08, 2.531739e-08, 
    2.531788e-08, 2.443518e-08, 2.322498e-08, 2.304853e-08, 2.232023e-08, 
    1.999054e-08, 1.762727e-08, 1.721729e-08, 1.821666e-08, 1.860172e-08,
  2.443982e-08, 2.496734e-08, 2.554411e-08, 2.587036e-08, 2.570712e-08, 
    2.561287e-08, 2.513679e-08, 2.419299e-08, 2.290481e-08, 2.280888e-08, 
    2.20269e-08, 2.00315e-08, 1.809733e-08, 1.709897e-08, 1.829499e-08,
  1.249278e-08, 1.156133e-08, 1.052087e-08, 9.69661e-09, 9.35226e-09, 
    9.003218e-09, 8.751733e-09, 8.242576e-09, 7.900541e-09, 7.304804e-09, 
    6.86723e-09, 6.500547e-09, 6.319445e-09, 6.348629e-09, 6.471834e-09,
  1.315488e-08, 1.22345e-08, 1.142244e-08, 1.033753e-08, 9.546713e-09, 
    9.209715e-09, 9.031393e-09, 8.639572e-09, 8.266563e-09, 7.752162e-09, 
    7.222576e-09, 6.819115e-09, 6.503964e-09, 6.393523e-09, 6.281123e-09,
  1.372173e-08, 1.301722e-08, 1.198671e-08, 1.113185e-08, 1.023099e-08, 
    9.406399e-09, 9.123418e-09, 8.932889e-09, 8.530794e-09, 8.147937e-09, 
    7.59078e-09, 7.196528e-09, 6.775106e-09, 6.613521e-09, 6.416509e-09,
  1.397876e-08, 1.373743e-08, 1.259699e-08, 1.159643e-08, 1.087314e-08, 
    1.009928e-08, 9.394968e-09, 9.094154e-09, 8.864401e-09, 8.422213e-09, 
    7.891483e-09, 7.437331e-09, 7.048592e-09, 6.82704e-09, 6.680991e-09,
  1.41175e-08, 1.397887e-08, 1.349699e-08, 1.223615e-08, 1.128271e-08, 
    1.058889e-08, 9.913535e-09, 9.435208e-09, 9.079606e-09, 8.828875e-09, 
    8.303888e-09, 7.739987e-09, 7.258788e-09, 7.010879e-09, 6.893607e-09,
  1.449219e-08, 1.403814e-08, 1.378783e-08, 1.30865e-08, 1.201955e-08, 
    1.106161e-08, 1.037184e-08, 9.817093e-09, 9.542624e-09, 9.143415e-09, 
    8.787076e-09, 8.236734e-09, 7.671595e-09, 7.319235e-09, 7.126715e-09,
  1.525844e-08, 1.457758e-08, 1.38703e-08, 1.349696e-08, 1.275898e-08, 
    1.181006e-08, 1.085622e-08, 1.011928e-08, 9.780922e-09, 9.59603e-09, 
    9.169535e-09, 8.859313e-09, 8.225955e-09, 7.829037e-09, 7.684213e-09,
  1.579964e-08, 1.524017e-08, 1.462447e-08, 1.391118e-08, 1.318896e-08, 
    1.235835e-08, 1.151966e-08, 1.064687e-08, 9.960784e-09, 9.742757e-09, 
    9.452447e-09, 9.150565e-09, 9.006726e-09, 8.45506e-09, 8.33595e-09,
  1.653515e-08, 1.577639e-08, 1.518875e-08, 1.466876e-08, 1.402133e-08, 
    1.303183e-08, 1.21015e-08, 1.136385e-08, 1.053007e-08, 9.856525e-09, 
    9.668424e-09, 9.307148e-09, 9.383866e-09, 9.228435e-09, 8.93862e-09,
  1.826412e-08, 1.684457e-08, 1.587712e-08, 1.52554e-08, 1.480669e-08, 
    1.408071e-08, 1.287233e-08, 1.195447e-08, 1.129205e-08, 1.04104e-08, 
    9.875071e-09, 9.623908e-09, 9.389177e-09, 9.592084e-09, 9.512181e-09,
  2.088506e-08, 1.714195e-08, 1.498117e-08, 1.329481e-08, 1.214793e-08, 
    1.147795e-08, 1.082036e-08, 1.016662e-08, 9.571931e-09, 9.190232e-09, 
    8.906497e-09, 8.604333e-09, 8.198076e-09, 7.777215e-09, 7.334335e-09,
  2.083336e-08, 1.657189e-08, 1.453213e-08, 1.285738e-08, 1.178598e-08, 
    1.109382e-08, 1.048065e-08, 9.848407e-09, 9.282556e-09, 8.913844e-09, 
    8.667786e-09, 8.446975e-09, 8.164547e-09, 7.847565e-09, 7.497419e-09,
  2.088284e-08, 1.630216e-08, 1.420914e-08, 1.24141e-08, 1.134361e-08, 
    1.07196e-08, 1.011022e-08, 9.501921e-09, 8.987702e-09, 8.708811e-09, 
    8.466909e-09, 8.270931e-09, 8.088197e-09, 7.854415e-09, 7.582979e-09,
  2.06711e-08, 1.615411e-08, 1.396468e-08, 1.199918e-08, 1.090878e-08, 
    1.03159e-08, 9.756293e-09, 9.255655e-09, 8.807354e-09, 8.52538e-09, 
    8.323196e-09, 8.133597e-09, 8.039564e-09, 7.880935e-09, 7.652078e-09,
  2.030104e-08, 1.59808e-08, 1.36448e-08, 1.157571e-08, 1.051779e-08, 
    1.000319e-08, 9.456504e-09, 9.012529e-09, 8.636301e-09, 8.417341e-09, 
    8.272104e-09, 8.090914e-09, 7.975249e-09, 7.918685e-09, 7.734971e-09,
  1.96787e-08, 1.562596e-08, 1.335547e-08, 1.129998e-08, 1.026122e-08, 
    9.70013e-09, 9.188873e-09, 8.788835e-09, 8.490365e-09, 8.330434e-09, 
    8.294593e-09, 8.23238e-09, 8.0775e-09, 8.017255e-09, 7.875744e-09,
  1.888989e-08, 1.521447e-08, 1.310004e-08, 1.122494e-08, 1.013985e-08, 
    9.540696e-09, 9.032078e-09, 8.642906e-09, 8.38763e-09, 8.310707e-09, 
    8.306382e-09, 8.416299e-09, 8.304232e-09, 8.227043e-09, 8.103759e-09,
  1.813784e-08, 1.479106e-08, 1.291976e-08, 1.120879e-08, 1.010471e-08, 
    9.417931e-09, 8.943521e-09, 8.59856e-09, 8.39552e-09, 8.394792e-09, 
    8.418388e-09, 8.602576e-09, 8.62449e-09, 8.491877e-09, 8.434756e-09,
  1.759568e-08, 1.445458e-08, 1.27823e-08, 1.121043e-08, 1.014617e-08, 
    9.42368e-09, 9.000763e-09, 8.664923e-09, 8.488406e-09, 8.518589e-09, 
    8.527923e-09, 8.772961e-09, 9.047639e-09, 8.907268e-09, 8.764934e-09,
  1.716751e-08, 1.424347e-08, 1.266384e-08, 1.119771e-08, 1.024237e-08, 
    9.507303e-09, 9.131528e-09, 8.858868e-09, 8.712175e-09, 8.758158e-09, 
    8.788223e-09, 8.924594e-09, 9.250742e-09, 9.373673e-09, 9.208706e-09,
  2.057524e-08, 1.859138e-08, 1.777051e-08, 1.792539e-08, 1.675071e-08, 
    1.560869e-08, 1.613937e-08, 1.619386e-08, 1.675617e-08, 1.725294e-08, 
    1.815753e-08, 1.856871e-08, 1.795e-08, 1.631243e-08, 1.46029e-08,
  2.117177e-08, 1.990369e-08, 1.834943e-08, 1.825794e-08, 1.775183e-08, 
    1.644575e-08, 1.607553e-08, 1.606749e-08, 1.710711e-08, 1.830268e-08, 
    1.865948e-08, 1.82631e-08, 1.739979e-08, 1.604631e-08, 1.46708e-08,
  2.105746e-08, 2.085254e-08, 2.004364e-08, 1.913548e-08, 1.852133e-08, 
    1.729024e-08, 1.624266e-08, 1.583318e-08, 1.695777e-08, 1.858821e-08, 
    1.908937e-08, 1.827906e-08, 1.690418e-08, 1.566436e-08, 1.446278e-08,
  2.124673e-08, 2.16331e-08, 2.130355e-08, 1.998315e-08, 1.9666e-08, 
    1.855501e-08, 1.724326e-08, 1.634635e-08, 1.688388e-08, 1.84043e-08, 
    1.897267e-08, 1.807089e-08, 1.658771e-08, 1.531681e-08, 1.419263e-08,
  2.171437e-08, 2.215984e-08, 2.187221e-08, 2.076885e-08, 2.011984e-08, 
    1.94205e-08, 1.853667e-08, 1.746426e-08, 1.731254e-08, 1.836399e-08, 
    1.843251e-08, 1.763212e-08, 1.625337e-08, 1.49482e-08, 1.389809e-08,
  2.278725e-08, 2.26548e-08, 2.215649e-08, 2.108295e-08, 2.015727e-08, 
    1.948243e-08, 1.921481e-08, 1.846717e-08, 1.786311e-08, 1.855909e-08, 
    1.784611e-08, 1.713179e-08, 1.584496e-08, 1.457187e-08, 1.350622e-08,
  2.43182e-08, 2.354304e-08, 2.202717e-08, 2.106466e-08, 2.000332e-08, 
    1.923959e-08, 1.928119e-08, 1.917217e-08, 1.819132e-08, 1.8323e-08, 
    1.7349e-08, 1.646122e-08, 1.534108e-08, 1.410438e-08, 1.299805e-08,
  2.576521e-08, 2.475058e-08, 2.215515e-08, 2.071284e-08, 1.974201e-08, 
    1.907064e-08, 1.923851e-08, 1.926433e-08, 1.818909e-08, 1.779747e-08, 
    1.665116e-08, 1.586903e-08, 1.484627e-08, 1.353072e-08, 1.242664e-08,
  2.705822e-08, 2.557766e-08, 2.327173e-08, 2.080104e-08, 1.943726e-08, 
    1.884482e-08, 1.903387e-08, 1.88298e-08, 1.78345e-08, 1.697933e-08, 
    1.594984e-08, 1.530092e-08, 1.424661e-08, 1.289615e-08, 1.188607e-08,
  2.759968e-08, 2.585305e-08, 2.390662e-08, 2.172703e-08, 1.92866e-08, 
    1.859291e-08, 1.883046e-08, 1.824436e-08, 1.725599e-08, 1.63402e-08, 
    1.542314e-08, 1.469626e-08, 1.359575e-08, 1.229619e-08, 1.138466e-08,
  9.561727e-09, 9.129518e-09, 9.046667e-09, 8.873963e-09, 8.655899e-09, 
    8.359506e-09, 8.214898e-09, 8.006809e-09, 8.139136e-09, 8.049132e-09, 
    8.415185e-09, 8.893628e-09, 9.217301e-09, 9.724922e-09, 1.01192e-08,
  9.993265e-09, 9.60027e-09, 9.292052e-09, 9.142553e-09, 9.012188e-09, 
    8.839132e-09, 8.760024e-09, 8.428265e-09, 8.505647e-09, 8.601089e-09, 
    9.162573e-09, 9.579383e-09, 9.750583e-09, 1.001994e-08, 1.048583e-08,
  1.032256e-08, 9.968545e-09, 9.553503e-09, 9.322129e-09, 9.16194e-09, 
    9.116288e-09, 9.104787e-09, 8.832711e-09, 9.009155e-09, 9.292706e-09, 
    1.018084e-08, 1.077237e-08, 1.101536e-08, 1.100972e-08, 1.144571e-08,
  1.084709e-08, 1.0416e-08, 9.885176e-09, 9.529053e-09, 9.260561e-09, 
    9.170734e-09, 9.159183e-09, 9.107874e-09, 9.495069e-09, 9.785341e-09, 
    1.069933e-08, 1.168469e-08, 1.219632e-08, 1.228817e-08, 1.26652e-08,
  1.116205e-08, 1.081305e-08, 1.037057e-08, 9.930248e-09, 9.597223e-09, 
    9.477374e-09, 9.430636e-09, 9.522001e-09, 9.961088e-09, 1.027723e-08, 
    1.072133e-08, 1.220742e-08, 1.304311e-08, 1.32618e-08, 1.34621e-08,
  1.146833e-08, 1.0989e-08, 1.082998e-08, 1.057982e-08, 1.020033e-08, 
    9.978508e-09, 9.834742e-09, 9.884844e-09, 1.027966e-08, 1.066655e-08, 
    1.106406e-08, 1.253256e-08, 1.357826e-08, 1.381973e-08, 1.41572e-08,
  1.172797e-08, 1.122738e-08, 1.117603e-08, 1.127777e-08, 1.129466e-08, 
    1.113361e-08, 1.089015e-08, 1.06962e-08, 1.073511e-08, 1.09789e-08, 
    1.124676e-08, 1.266968e-08, 1.378913e-08, 1.404988e-08, 1.460831e-08,
  1.190256e-08, 1.140124e-08, 1.131217e-08, 1.167158e-08, 1.20322e-08, 
    1.206527e-08, 1.201342e-08, 1.199279e-08, 1.186511e-08, 1.183463e-08, 
    1.211145e-08, 1.334623e-08, 1.432475e-08, 1.462876e-08, 1.526629e-08,
  1.229076e-08, 1.204819e-08, 1.165661e-08, 1.179802e-08, 1.229119e-08, 
    1.242104e-08, 1.237887e-08, 1.258301e-08, 1.235017e-08, 1.235622e-08, 
    1.288366e-08, 1.415639e-08, 1.492019e-08, 1.512662e-08, 1.581325e-08,
  1.28181e-08, 1.225841e-08, 1.210199e-08, 1.229201e-08, 1.264355e-08, 
    1.287792e-08, 1.276892e-08, 1.291375e-08, 1.277095e-08, 1.263331e-08, 
    1.336066e-08, 1.481599e-08, 1.548501e-08, 1.556966e-08, 1.618083e-08,
  7.050491e-09, 6.367919e-09, 5.973362e-09, 5.438425e-09, 5.104738e-09, 
    4.701311e-09, 4.527263e-09, 4.235969e-09, 3.987002e-09, 3.848564e-09, 
    3.787047e-09, 3.798368e-09, 3.783412e-09, 3.761838e-09, 3.734979e-09,
  7.017817e-09, 6.41234e-09, 6.011431e-09, 5.482337e-09, 5.20097e-09, 
    4.784387e-09, 4.596926e-09, 4.443867e-09, 4.394785e-09, 4.34344e-09, 
    4.295327e-09, 4.343644e-09, 4.356384e-09, 4.286399e-09, 4.120538e-09,
  7.010826e-09, 6.404873e-09, 6.02071e-09, 5.54925e-09, 5.302466e-09, 
    4.977642e-09, 4.811799e-09, 4.708375e-09, 4.732398e-09, 4.843551e-09, 
    4.805443e-09, 4.655332e-09, 4.505017e-09, 4.536311e-09, 4.575672e-09,
  7.024784e-09, 6.421762e-09, 6.09406e-09, 5.620532e-09, 5.377434e-09, 
    5.070292e-09, 5.005053e-09, 5.069578e-09, 5.164051e-09, 5.185212e-09, 
    5.14068e-09, 4.980773e-09, 4.91185e-09, 4.952919e-09, 5.040658e-09,
  7.142069e-09, 6.579673e-09, 6.292533e-09, 5.912622e-09, 5.69865e-09, 
    5.546968e-09, 5.404874e-09, 5.333637e-09, 5.429557e-09, 5.491141e-09, 
    5.391835e-09, 5.366273e-09, 5.361908e-09, 5.394711e-09, 5.637478e-09,
  7.320548e-09, 6.90485e-09, 6.677888e-09, 6.298122e-09, 6.157305e-09, 
    5.972043e-09, 6.094051e-09, 6.029708e-09, 5.917807e-09, 5.770711e-09, 
    5.702676e-09, 5.773102e-09, 5.906315e-09, 6.020551e-09, 6.191303e-09,
  7.552484e-09, 7.158591e-09, 6.932253e-09, 6.701992e-09, 6.621146e-09, 
    6.45251e-09, 6.289838e-09, 6.329911e-09, 6.225334e-09, 6.161184e-09, 
    5.985977e-09, 6.125123e-09, 6.218883e-09, 6.39268e-09, 6.516907e-09,
  7.702966e-09, 7.34264e-09, 7.095722e-09, 6.88346e-09, 6.627111e-09, 
    6.609074e-09, 6.567914e-09, 6.585362e-09, 6.585363e-09, 6.737969e-09, 
    6.735389e-09, 6.765387e-09, 6.761503e-09, 6.955823e-09, 7.017401e-09,
  7.840737e-09, 7.393948e-09, 7.019771e-09, 6.864408e-09, 6.83613e-09, 
    6.8383e-09, 6.941116e-09, 7.120732e-09, 7.06225e-09, 6.984947e-09, 
    7.094057e-09, 7.171749e-09, 7.341403e-09, 7.527093e-09, 7.858648e-09,
  8.231875e-09, 7.805909e-09, 7.517608e-09, 7.554593e-09, 7.407726e-09, 
    7.508421e-09, 7.587156e-09, 7.708773e-09, 7.73533e-09, 7.57251e-09, 
    7.514255e-09, 7.706791e-09, 7.843252e-09, 8.186905e-09, 8.594855e-09,
  1.344609e-08, 1.330914e-08, 1.294771e-08, 1.245103e-08, 1.209029e-08, 
    1.180308e-08, 1.122988e-08, 1.092318e-08, 1.061579e-08, 1.036839e-08, 
    1.024736e-08, 9.837672e-09, 9.423625e-09, 9.047267e-09, 8.71009e-09,
  1.238812e-08, 1.2538e-08, 1.219756e-08, 1.188187e-08, 1.160265e-08, 
    1.120479e-08, 1.074856e-08, 1.027202e-08, 9.807835e-09, 9.467067e-09, 
    9.218287e-09, 8.841673e-09, 8.504205e-09, 8.137413e-09, 7.928851e-09,
  1.150154e-08, 1.117461e-08, 1.087449e-08, 1.061911e-08, 1.029507e-08, 
    9.933804e-09, 9.528564e-09, 9.137709e-09, 8.785046e-09, 8.455696e-09, 
    8.20912e-09, 7.958355e-09, 7.674639e-09, 7.395419e-09, 7.166131e-09,
  1.004627e-08, 9.853227e-09, 9.745888e-09, 9.257077e-09, 8.805394e-09, 
    8.416179e-09, 8.251279e-09, 8.038689e-09, 7.785495e-09, 7.539878e-09, 
    7.32137e-09, 7.093683e-09, 6.923229e-09, 6.743288e-09, 6.559258e-09,
  8.338414e-09, 8.270773e-09, 8.148177e-09, 7.843154e-09, 7.538331e-09, 
    7.247015e-09, 7.130784e-09, 6.77518e-09, 6.602273e-09, 6.4117e-09, 
    6.331478e-09, 6.142756e-09, 6.067305e-09, 5.988142e-09, 5.814447e-09,
  7.127959e-09, 6.92522e-09, 6.703525e-09, 6.630252e-09, 6.56511e-09, 
    6.474055e-09, 6.309424e-09, 6.132058e-09, 5.897955e-09, 5.616859e-09, 
    5.592363e-09, 5.469482e-09, 5.456767e-09, 5.475639e-09, 5.352335e-09,
  6.02532e-09, 5.740019e-09, 5.639521e-09, 5.713078e-09, 5.786983e-09, 
    5.744881e-09, 5.668062e-09, 5.629509e-09, 5.561721e-09, 5.267786e-09, 
    5.205228e-09, 5.078581e-09, 5.141724e-09, 5.151329e-09, 5.107326e-09,
  5.312507e-09, 5.220889e-09, 5.116513e-09, 5.20775e-09, 5.259098e-09, 
    5.293677e-09, 5.42507e-09, 5.279017e-09, 5.196892e-09, 5.200907e-09, 
    5.203491e-09, 5.063011e-09, 5.031653e-09, 5.009387e-09, 4.912221e-09,
  4.994334e-09, 4.976355e-09, 5.048987e-09, 5.084113e-09, 5.058963e-09, 
    5.054435e-09, 5.232458e-09, 5.481069e-09, 5.265277e-09, 5.144904e-09, 
    5.223199e-09, 5.178235e-09, 5.113386e-09, 5.122946e-09, 5.0404e-09,
  5.239863e-09, 5.420638e-09, 5.267887e-09, 5.301128e-09, 5.301717e-09, 
    5.556542e-09, 5.51115e-09, 5.616565e-09, 5.618871e-09, 5.522574e-09, 
    5.462664e-09, 5.440233e-09, 5.478709e-09, 5.486303e-09, 5.571344e-09,
  2.534746e-08, 2.502467e-08, 2.485959e-08, 2.414463e-08, 2.330308e-08, 
    2.240262e-08, 2.206748e-08, 2.142347e-08, 2.09189e-08, 2.040421e-08, 
    1.987309e-08, 1.921248e-08, 1.862518e-08, 1.785255e-08, 1.725895e-08,
  2.516656e-08, 2.50537e-08, 2.482629e-08, 2.391024e-08, 2.333419e-08, 
    2.270012e-08, 2.252399e-08, 2.17941e-08, 2.123399e-08, 2.031331e-08, 
    1.954876e-08, 1.884241e-08, 1.824675e-08, 1.748086e-08, 1.68154e-08,
  2.455525e-08, 2.449989e-08, 2.422826e-08, 2.360221e-08, 2.300176e-08, 
    2.231762e-08, 2.220338e-08, 2.159227e-08, 2.087423e-08, 1.976625e-08, 
    1.891974e-08, 1.834626e-08, 1.784423e-08, 1.713192e-08, 1.651371e-08,
  2.294827e-08, 2.274087e-08, 2.249239e-08, 2.20385e-08, 2.154124e-08, 
    2.124667e-08, 2.107986e-08, 2.022363e-08, 1.942685e-08, 1.839062e-08, 
    1.790037e-08, 1.761346e-08, 1.727028e-08, 1.674978e-08, 1.630814e-08,
  2.101438e-08, 2.114387e-08, 2.076648e-08, 2.036726e-08, 2.006789e-08, 
    1.96662e-08, 1.917312e-08, 1.843394e-08, 1.793563e-08, 1.739593e-08, 
    1.714046e-08, 1.694684e-08, 1.657186e-08, 1.612641e-08, 1.568756e-08,
  1.906841e-08, 1.941318e-08, 1.928916e-08, 1.932851e-08, 1.901608e-08, 
    1.863269e-08, 1.797393e-08, 1.738023e-08, 1.687295e-08, 1.649838e-08, 
    1.647136e-08, 1.62703e-08, 1.597263e-08, 1.559593e-08, 1.521597e-08,
  1.730744e-08, 1.780109e-08, 1.772845e-08, 1.782165e-08, 1.754771e-08, 
    1.719802e-08, 1.682529e-08, 1.653261e-08, 1.61222e-08, 1.578599e-08, 
    1.557162e-08, 1.527581e-08, 1.513545e-08, 1.481481e-08, 1.443228e-08,
  1.467961e-08, 1.569875e-08, 1.576994e-08, 1.582746e-08, 1.569708e-08, 
    1.558685e-08, 1.546291e-08, 1.519797e-08, 1.498752e-08, 1.489667e-08, 
    1.467098e-08, 1.444721e-08, 1.423461e-08, 1.39694e-08, 1.382267e-08,
  1.081598e-08, 1.223063e-08, 1.284216e-08, 1.328643e-08, 1.345251e-08, 
    1.360439e-08, 1.363425e-08, 1.373602e-08, 1.376065e-08, 1.374527e-08, 
    1.367166e-08, 1.354254e-08, 1.346014e-08, 1.329901e-08, 1.313216e-08,
  8.118691e-09, 9.462024e-09, 1.023499e-08, 1.078991e-08, 1.122915e-08, 
    1.153883e-08, 1.188828e-08, 1.206824e-08, 1.223806e-08, 1.238462e-08, 
    1.244042e-08, 1.251362e-08, 1.238962e-08, 1.236713e-08, 1.24975e-08,
  2.222664e-08, 2.21705e-08, 2.17137e-08, 2.128787e-08, 2.079062e-08, 
    2.008565e-08, 1.95775e-08, 1.919058e-08, 1.890654e-08, 1.863455e-08, 
    1.838252e-08, 1.796448e-08, 1.738662e-08, 1.679673e-08, 1.55917e-08,
  2.242892e-08, 2.223896e-08, 2.211596e-08, 2.135347e-08, 2.072621e-08, 
    2.005494e-08, 1.955949e-08, 1.921234e-08, 1.910328e-08, 1.907811e-08, 
    1.894357e-08, 1.864696e-08, 1.820476e-08, 1.763276e-08, 1.693739e-08,
  2.187697e-08, 2.138334e-08, 2.157639e-08, 2.128392e-08, 2.102361e-08, 
    2.049044e-08, 2.021746e-08, 1.991363e-08, 1.954462e-08, 1.94361e-08, 
    1.93392e-08, 1.909759e-08, 1.862131e-08, 1.801441e-08, 1.757212e-08,
  2.21457e-08, 2.189181e-08, 2.206157e-08, 2.183752e-08, 2.189133e-08, 
    2.155192e-08, 2.112293e-08, 2.085036e-08, 2.053988e-08, 2.01875e-08, 
    1.989191e-08, 1.957815e-08, 1.919036e-08, 1.865994e-08, 1.812982e-08,
  2.227437e-08, 2.237285e-08, 2.289786e-08, 2.293053e-08, 2.288902e-08, 
    2.265922e-08, 2.218786e-08, 2.16762e-08, 2.101972e-08, 2.048052e-08, 
    2.006328e-08, 1.980074e-08, 1.941642e-08, 1.898109e-08, 1.848202e-08,
  2.387881e-08, 2.408058e-08, 2.448583e-08, 2.422352e-08, 2.386561e-08, 
    2.348831e-08, 2.282675e-08, 2.228618e-08, 2.174759e-08, 2.119804e-08, 
    2.081917e-08, 2.042301e-08, 1.996482e-08, 1.949268e-08, 1.882642e-08,
  2.527844e-08, 2.544528e-08, 2.529574e-08, 2.443279e-08, 2.384464e-08, 
    2.357977e-08, 2.31538e-08, 2.275596e-08, 2.234163e-08, 2.185863e-08, 
    2.127843e-08, 2.080763e-08, 2.036219e-08, 1.991674e-08, 1.936244e-08,
  2.50518e-08, 2.392842e-08, 2.355913e-08, 2.272461e-08, 2.247713e-08, 
    2.26863e-08, 2.283283e-08, 2.30373e-08, 2.298609e-08, 2.256588e-08, 
    2.20333e-08, 2.141557e-08, 2.071811e-08, 2.009694e-08, 1.940364e-08,
  2.208044e-08, 2.201099e-08, 2.199478e-08, 2.183983e-08, 2.196796e-08, 
    2.230554e-08, 2.254727e-08, 2.283756e-08, 2.289858e-08, 2.284895e-08, 
    2.244753e-08, 2.183935e-08, 2.114075e-08, 2.068353e-08, 1.985758e-08,
  2.036099e-08, 2.092155e-08, 2.10511e-08, 2.147531e-08, 2.178015e-08, 
    2.208553e-08, 2.221011e-08, 2.229397e-08, 2.23637e-08, 2.241068e-08, 
    2.254494e-08, 2.234216e-08, 2.1698e-08, 2.099284e-08, 2.046518e-08,
  2.175666e-08, 2.160121e-08, 2.051382e-08, 1.91893e-08, 1.803465e-08, 
    1.700173e-08, 1.630537e-08, 1.572362e-08, 1.523829e-08, 1.507028e-08, 
    1.493386e-08, 1.472517e-08, 1.38283e-08, 1.200713e-08, 1.058093e-08,
  2.117855e-08, 2.081922e-08, 1.95941e-08, 1.849007e-08, 1.739737e-08, 
    1.654187e-08, 1.568133e-08, 1.507072e-08, 1.481845e-08, 1.476117e-08, 
    1.453253e-08, 1.448934e-08, 1.35661e-08, 1.194727e-08, 1.044154e-08,
  2.028462e-08, 1.989661e-08, 1.892604e-08, 1.799202e-08, 1.710599e-08, 
    1.619457e-08, 1.531451e-08, 1.476848e-08, 1.438692e-08, 1.423966e-08, 
    1.421819e-08, 1.417069e-08, 1.35025e-08, 1.187285e-08, 1.036419e-08,
  1.911439e-08, 1.86388e-08, 1.77651e-08, 1.719818e-08, 1.668354e-08, 
    1.610392e-08, 1.53116e-08, 1.474631e-08, 1.421074e-08, 1.382662e-08, 
    1.412603e-08, 1.397457e-08, 1.322883e-08, 1.197784e-08, 1.044865e-08,
  1.906585e-08, 1.831103e-08, 1.743864e-08, 1.680992e-08, 1.631739e-08, 
    1.575237e-08, 1.524976e-08, 1.485764e-08, 1.441378e-08, 1.379096e-08, 
    1.385049e-08, 1.399058e-08, 1.328045e-08, 1.196221e-08, 1.052747e-08,
  1.868805e-08, 1.779473e-08, 1.721236e-08, 1.674915e-08, 1.62507e-08, 
    1.569762e-08, 1.505443e-08, 1.461601e-08, 1.421908e-08, 1.372513e-08, 
    1.377687e-08, 1.380196e-08, 1.330712e-08, 1.238667e-08, 1.082814e-08,
  1.924426e-08, 1.839399e-08, 1.770795e-08, 1.711545e-08, 1.660413e-08, 
    1.595294e-08, 1.531957e-08, 1.478718e-08, 1.425346e-08, 1.379042e-08, 
    1.345519e-08, 1.360171e-08, 1.360146e-08, 1.257291e-08, 1.130556e-08,
  2.105621e-08, 1.981642e-08, 1.90095e-08, 1.830468e-08, 1.761059e-08, 
    1.687366e-08, 1.604584e-08, 1.517331e-08, 1.449365e-08, 1.398387e-08, 
    1.360462e-08, 1.329062e-08, 1.329438e-08, 1.305003e-08, 1.174824e-08,
  2.305999e-08, 2.168339e-08, 2.070364e-08, 2.006246e-08, 1.926227e-08, 
    1.838219e-08, 1.740704e-08, 1.648174e-08, 1.554577e-08, 1.456138e-08, 
    1.386338e-08, 1.330739e-08, 1.332708e-08, 1.292836e-08, 1.222927e-08,
  2.330262e-08, 2.258949e-08, 2.201727e-08, 2.146388e-08, 2.06918e-08, 
    1.994925e-08, 1.91351e-08, 1.789109e-08, 1.672107e-08, 1.578529e-08, 
    1.487988e-08, 1.380644e-08, 1.320817e-08, 1.317535e-08, 1.249939e-08,
  2.445386e-08, 2.436164e-08, 2.36457e-08, 2.283856e-08, 2.254059e-08, 
    2.24058e-08, 2.217732e-08, 2.167194e-08, 2.140611e-08, 2.093409e-08, 
    2.049246e-08, 1.989813e-08, 1.914958e-08, 1.827486e-08, 1.767689e-08,
  2.452103e-08, 2.418212e-08, 2.362995e-08, 2.30769e-08, 2.27878e-08, 
    2.243939e-08, 2.211921e-08, 2.17361e-08, 2.15161e-08, 2.126238e-08, 
    2.08656e-08, 1.994148e-08, 1.899234e-08, 1.812045e-08, 1.750931e-08,
  2.461572e-08, 2.381522e-08, 2.328394e-08, 2.284555e-08, 2.2424e-08, 
    2.196828e-08, 2.183229e-08, 2.172979e-08, 2.173676e-08, 2.128615e-08, 
    2.059788e-08, 1.955947e-08, 1.868318e-08, 1.779751e-08, 1.713581e-08,
  2.456483e-08, 2.348315e-08, 2.282315e-08, 2.234101e-08, 2.190278e-08, 
    2.164383e-08, 2.168341e-08, 2.165756e-08, 2.147483e-08, 2.084021e-08, 
    2.009574e-08, 1.900881e-08, 1.815391e-08, 1.731078e-08, 1.677744e-08,
  2.425777e-08, 2.325212e-08, 2.262535e-08, 2.211221e-08, 2.174503e-08, 
    2.14928e-08, 2.153326e-08, 2.143661e-08, 2.094105e-08, 2.00549e-08, 
    1.9397e-08, 1.841288e-08, 1.757132e-08, 1.685009e-08, 1.639989e-08,
  2.380308e-08, 2.316544e-08, 2.256703e-08, 2.196263e-08, 2.160204e-08, 
    2.120168e-08, 2.118673e-08, 2.085917e-08, 2.012441e-08, 1.91435e-08, 
    1.87513e-08, 1.780981e-08, 1.700369e-08, 1.635857e-08, 1.594976e-08,
  2.369177e-08, 2.311451e-08, 2.23849e-08, 2.185916e-08, 2.13312e-08, 
    2.086248e-08, 2.059129e-08, 1.991291e-08, 1.913235e-08, 1.830689e-08, 
    1.80428e-08, 1.727862e-08, 1.650838e-08, 1.584884e-08, 1.542243e-08,
  2.322805e-08, 2.274372e-08, 2.198204e-08, 2.127135e-08, 2.06288e-08, 
    2.000636e-08, 1.965986e-08, 1.891499e-08, 1.817919e-08, 1.748107e-08, 
    1.731389e-08, 1.684713e-08, 1.609491e-08, 1.537631e-08, 1.487486e-08,
  2.30657e-08, 2.22803e-08, 2.126416e-08, 2.058515e-08, 1.979828e-08, 
    1.917287e-08, 1.851111e-08, 1.776021e-08, 1.711252e-08, 1.665086e-08, 
    1.667589e-08, 1.637881e-08, 1.573554e-08, 1.492797e-08, 1.436977e-08,
  2.222691e-08, 2.136957e-08, 2.050563e-08, 1.953754e-08, 1.871699e-08, 
    1.794506e-08, 1.749805e-08, 1.690609e-08, 1.639116e-08, 1.576739e-08, 
    1.584326e-08, 1.583992e-08, 1.529061e-08, 1.453575e-08, 1.39523e-08,
  2.284837e-08, 2.231254e-08, 2.194763e-08, 2.048597e-08, 1.975084e-08, 
    1.936635e-08, 1.875912e-08, 1.839657e-08, 1.842743e-08, 1.858734e-08, 
    1.860292e-08, 1.872057e-08, 1.938762e-08, 2.000367e-08, 1.990908e-08,
  2.317687e-08, 2.239229e-08, 2.18001e-08, 2.080412e-08, 2.021436e-08, 
    1.960984e-08, 1.899007e-08, 1.877259e-08, 1.870058e-08, 1.86997e-08, 
    1.867953e-08, 1.881379e-08, 1.934679e-08, 1.987632e-08, 1.981518e-08,
  2.286505e-08, 2.224803e-08, 2.169285e-08, 2.084226e-08, 2.068617e-08, 
    2.047398e-08, 1.952339e-08, 1.893848e-08, 1.86444e-08, 1.852156e-08, 
    1.851053e-08, 1.873603e-08, 1.928231e-08, 1.976019e-08, 1.980031e-08,
  2.22413e-08, 2.183328e-08, 2.127884e-08, 2.069439e-08, 2.042947e-08, 
    1.981866e-08, 1.902023e-08, 1.866762e-08, 1.83419e-08, 1.831711e-08, 
    1.842604e-08, 1.875396e-08, 1.926944e-08, 1.966452e-08, 1.974805e-08,
  2.172636e-08, 2.123987e-08, 2.050775e-08, 1.983453e-08, 1.958825e-08, 
    1.895619e-08, 1.847032e-08, 1.832003e-08, 1.818229e-08, 1.826191e-08, 
    1.837289e-08, 1.871134e-08, 1.929527e-08, 1.9659e-08, 1.976879e-08,
  2.119177e-08, 2.048235e-08, 1.964194e-08, 1.886993e-08, 1.859568e-08, 
    1.826396e-08, 1.820823e-08, 1.83432e-08, 1.832537e-08, 1.846714e-08, 
    1.859102e-08, 1.885703e-08, 1.931381e-08, 1.965221e-08, 1.975066e-08,
  2.077005e-08, 2.00013e-08, 1.908892e-08, 1.855565e-08, 1.840631e-08, 
    1.831553e-08, 1.847341e-08, 1.859271e-08, 1.866051e-08, 1.874599e-08, 
    1.878786e-08, 1.889626e-08, 1.932055e-08, 1.960731e-08, 1.970833e-08,
  2.07599e-08, 1.997052e-08, 1.91664e-08, 1.878163e-08, 1.872214e-08, 
    1.87839e-08, 1.900609e-08, 1.910444e-08, 1.903129e-08, 1.90969e-08, 
    1.908147e-08, 1.909769e-08, 1.932676e-08, 1.94826e-08, 1.960431e-08,
  2.105503e-08, 2.035798e-08, 1.98106e-08, 1.942487e-08, 1.933591e-08, 
    1.937896e-08, 1.960688e-08, 1.958951e-08, 1.953626e-08, 1.951623e-08, 
    1.933138e-08, 1.91451e-08, 1.924019e-08, 1.934059e-08, 1.950686e-08,
  2.137286e-08, 2.069236e-08, 2.047295e-08, 2.013697e-08, 2.000861e-08, 
    1.996252e-08, 1.990295e-08, 1.975934e-08, 1.973515e-08, 1.964894e-08, 
    1.938996e-08, 1.922635e-08, 1.918263e-08, 1.925064e-08, 1.931442e-08,
  2.628126e-08, 2.641185e-08, 2.513727e-08, 2.375811e-08, 2.261876e-08, 
    2.168867e-08, 2.084689e-08, 2.038463e-08, 1.993448e-08, 1.95555e-08, 
    1.94258e-08, 1.93479e-08, 1.955298e-08, 1.940216e-08, 1.864138e-08,
  2.594702e-08, 2.595539e-08, 2.503652e-08, 2.372933e-08, 2.244322e-08, 
    2.142191e-08, 2.05773e-08, 2.027505e-08, 1.986204e-08, 1.945143e-08, 
    1.935753e-08, 1.948427e-08, 1.972621e-08, 1.997896e-08, 1.93343e-08,
  2.539224e-08, 2.499208e-08, 2.401719e-08, 2.286063e-08, 2.195738e-08, 
    2.113837e-08, 2.050826e-08, 2.014748e-08, 1.969512e-08, 1.933009e-08, 
    1.927787e-08, 1.940698e-08, 1.966872e-08, 2.014345e-08, 1.984326e-08,
  2.423542e-08, 2.401375e-08, 2.285008e-08, 2.187685e-08, 2.111811e-08, 
    2.057648e-08, 2.020734e-08, 2.00588e-08, 1.962437e-08, 1.931017e-08, 
    1.922505e-08, 1.936805e-08, 1.951073e-08, 2.028262e-08, 2.016415e-08,
  2.283739e-08, 2.248489e-08, 2.154215e-08, 2.096821e-08, 2.038804e-08, 
    2.001086e-08, 1.979895e-08, 1.969208e-08, 1.939621e-08, 1.922178e-08, 
    1.919751e-08, 1.926052e-08, 1.941812e-08, 2.021997e-08, 2.048094e-08,
  2.144053e-08, 2.113026e-08, 2.034553e-08, 2.00043e-08, 1.968224e-08, 
    1.943055e-08, 1.928076e-08, 1.916232e-08, 1.898278e-08, 1.907724e-08, 
    1.908404e-08, 1.920063e-08, 1.933302e-08, 2.010173e-08, 2.067318e-08,
  2.071326e-08, 2.029716e-08, 1.955855e-08, 1.943317e-08, 1.919382e-08, 
    1.905545e-08, 1.871099e-08, 1.870658e-08, 1.875185e-08, 1.879398e-08, 
    1.890318e-08, 1.914655e-08, 1.928851e-08, 2.000909e-08, 2.0772e-08,
  2.049364e-08, 2.0158e-08, 1.953565e-08, 1.931715e-08, 1.895379e-08, 
    1.87483e-08, 1.865968e-08, 1.864828e-08, 1.856671e-08, 1.864107e-08, 
    1.878096e-08, 1.905268e-08, 1.931725e-08, 1.994386e-08, 2.078459e-08,
  2.024012e-08, 1.993912e-08, 1.955543e-08, 1.952429e-08, 1.921343e-08, 
    1.897995e-08, 1.871341e-08, 1.863903e-08, 1.866887e-08, 1.86715e-08, 
    1.872843e-08, 1.899632e-08, 1.930967e-08, 2.004975e-08, 2.086317e-08,
  1.997923e-08, 1.978719e-08, 1.964027e-08, 1.971131e-08, 1.949586e-08, 
    1.932179e-08, 1.928351e-08, 1.92223e-08, 1.91413e-08, 1.903574e-08, 
    1.890237e-08, 1.911096e-08, 1.946075e-08, 2.010776e-08, 2.097276e-08,
  2.61391e-08, 2.59834e-08, 2.598386e-08, 2.61911e-08, 2.615273e-08, 
    2.621145e-08, 2.566594e-08, 2.489537e-08, 2.497722e-08, 2.404962e-08, 
    2.138159e-08, 1.793264e-08, 1.573578e-08, 1.401036e-08, 1.243645e-08,
  2.661048e-08, 2.660326e-08, 2.662214e-08, 2.652643e-08, 2.615057e-08, 
    2.59053e-08, 2.555692e-08, 2.501217e-08, 2.500702e-08, 2.439645e-08, 
    2.19747e-08, 1.881402e-08, 1.619607e-08, 1.442006e-08, 1.291407e-08,
  2.777715e-08, 2.738425e-08, 2.729725e-08, 2.680769e-08, 2.661811e-08, 
    2.613088e-08, 2.554136e-08, 2.484465e-08, 2.477132e-08, 2.422977e-08, 
    2.238105e-08, 1.955641e-08, 1.687668e-08, 1.486503e-08, 1.330996e-08,
  2.886931e-08, 2.82625e-08, 2.761662e-08, 2.711509e-08, 2.663271e-08, 
    2.597941e-08, 2.530774e-08, 2.472187e-08, 2.45142e-08, 2.402062e-08, 
    2.260579e-08, 2.024662e-08, 1.760103e-08, 1.533633e-08, 1.363889e-08,
  2.994974e-08, 2.919151e-08, 2.84514e-08, 2.775719e-08, 2.707523e-08, 
    2.590652e-08, 2.509743e-08, 2.466546e-08, 2.451882e-08, 2.374101e-08, 
    2.236518e-08, 2.046814e-08, 1.814257e-08, 1.584075e-08, 1.394561e-08,
  2.869603e-08, 2.857347e-08, 2.804168e-08, 2.77709e-08, 2.669543e-08, 
    2.559379e-08, 2.518878e-08, 2.473892e-08, 2.439481e-08, 2.32243e-08, 
    2.195198e-08, 2.029709e-08, 1.854753e-08, 1.64682e-08, 1.428892e-08,
  2.586002e-08, 2.645953e-08, 2.66906e-08, 2.70327e-08, 2.595058e-08, 
    2.526084e-08, 2.496943e-08, 2.453032e-08, 2.402159e-08, 2.267002e-08, 
    2.152731e-08, 2.008892e-08, 1.86757e-08, 1.705039e-08, 1.479557e-08,
  2.421901e-08, 2.475823e-08, 2.545217e-08, 2.57812e-08, 2.495725e-08, 
    2.452219e-08, 2.429502e-08, 2.389635e-08, 2.309772e-08, 2.18106e-08, 
    2.100351e-08, 1.98623e-08, 1.876747e-08, 1.761761e-08, 1.546174e-08,
  2.378646e-08, 2.403793e-08, 2.45635e-08, 2.46412e-08, 2.386417e-08, 
    2.346448e-08, 2.292986e-08, 2.25982e-08, 2.209069e-08, 2.094912e-08, 
    2.048842e-08, 1.969803e-08, 1.878975e-08, 1.815435e-08, 1.629068e-08,
  2.299947e-08, 2.314846e-08, 2.360479e-08, 2.353333e-08, 2.281912e-08, 
    2.237196e-08, 2.187624e-08, 2.170619e-08, 2.130126e-08, 2.04026e-08, 
    2.009187e-08, 1.950597e-08, 1.875009e-08, 1.850566e-08, 1.719208e-08,
  2.580333e-08, 2.447507e-08, 2.513813e-08, 2.626265e-08, 2.721868e-08, 
    2.785353e-08, 2.64494e-08, 2.371121e-08, 2.148559e-08, 1.878864e-08, 
    1.687802e-08, 1.620161e-08, 1.593888e-08, 1.521421e-08, 1.471522e-08,
  2.628502e-08, 2.516532e-08, 2.47094e-08, 2.561492e-08, 2.668963e-08, 
    2.790489e-08, 2.764022e-08, 2.50157e-08, 2.255018e-08, 2.017042e-08, 
    1.743618e-08, 1.657596e-08, 1.626351e-08, 1.547822e-08, 1.497629e-08,
  2.617443e-08, 2.543698e-08, 2.468271e-08, 2.507856e-08, 2.588006e-08, 
    2.790098e-08, 2.815131e-08, 2.629404e-08, 2.373619e-08, 2.148002e-08, 
    1.853389e-08, 1.701632e-08, 1.659765e-08, 1.586631e-08, 1.528506e-08,
  2.635175e-08, 2.569563e-08, 2.500438e-08, 2.501979e-08, 2.546651e-08, 
    2.756244e-08, 2.850956e-08, 2.758886e-08, 2.495543e-08, 2.256735e-08, 
    1.968204e-08, 1.756466e-08, 1.697347e-08, 1.624158e-08, 1.55662e-08,
  2.661642e-08, 2.581729e-08, 2.515834e-08, 2.516904e-08, 2.524047e-08, 
    2.712879e-08, 2.887594e-08, 2.878203e-08, 2.657408e-08, 2.377225e-08, 
    2.094633e-08, 1.817924e-08, 1.733558e-08, 1.661447e-08, 1.577543e-08,
  2.744263e-08, 2.639013e-08, 2.60705e-08, 2.596083e-08, 2.532532e-08, 
    2.702422e-08, 2.880773e-08, 2.934228e-08, 2.780612e-08, 2.467849e-08, 
    2.198897e-08, 1.88785e-08, 1.766528e-08, 1.696526e-08, 1.603043e-08,
  2.821509e-08, 2.717153e-08, 2.692319e-08, 2.630221e-08, 2.585649e-08, 
    2.737474e-08, 2.868686e-08, 2.923464e-08, 2.886497e-08, 2.581082e-08, 
    2.293944e-08, 1.9629e-08, 1.798301e-08, 1.722109e-08, 1.625197e-08,
  2.845238e-08, 2.741368e-08, 2.714755e-08, 2.659358e-08, 2.651455e-08, 
    2.757088e-08, 2.843757e-08, 2.926657e-08, 2.931775e-08, 2.638581e-08, 
    2.335986e-08, 2.021939e-08, 1.82633e-08, 1.744484e-08, 1.651633e-08,
  2.870662e-08, 2.768511e-08, 2.772754e-08, 2.733423e-08, 2.725166e-08, 
    2.804334e-08, 2.823606e-08, 2.922054e-08, 2.915604e-08, 2.678716e-08, 
    2.341639e-08, 2.055449e-08, 1.848533e-08, 1.760296e-08, 1.676138e-08,
  2.907062e-08, 2.802315e-08, 2.804575e-08, 2.760702e-08, 2.764011e-08, 
    2.761972e-08, 2.777961e-08, 2.875726e-08, 2.873251e-08, 2.675855e-08, 
    2.313317e-08, 2.069703e-08, 1.869608e-08, 1.77216e-08, 1.691327e-08,
  2.535845e-08, 2.538887e-08, 2.389501e-08, 2.157317e-08, 2.025771e-08, 
    1.909977e-08, 1.844912e-08, 1.800783e-08, 1.700953e-08, 1.534416e-08, 
    1.373075e-08, 1.209445e-08, 1.115168e-08, 1.013381e-08, 9.292346e-09,
  2.641394e-08, 2.587502e-08, 2.542839e-08, 2.364584e-08, 2.158083e-08, 
    1.997035e-08, 1.912973e-08, 1.836403e-08, 1.756727e-08, 1.577042e-08, 
    1.39812e-08, 1.226273e-08, 1.125257e-08, 1.032895e-08, 9.460154e-09,
  2.690388e-08, 2.656786e-08, 2.625591e-08, 2.535747e-08, 2.358011e-08, 
    2.116807e-08, 1.9637e-08, 1.883793e-08, 1.807664e-08, 1.631416e-08, 
    1.430071e-08, 1.251473e-08, 1.13523e-08, 1.051081e-08, 9.658888e-09,
  2.67743e-08, 2.677672e-08, 2.685212e-08, 2.629303e-08, 2.525451e-08, 
    2.30039e-08, 2.050579e-08, 1.949751e-08, 1.863845e-08, 1.694579e-08, 
    1.478215e-08, 1.276676e-08, 1.15028e-08, 1.063717e-08, 9.809531e-09,
  2.712377e-08, 2.670106e-08, 2.692368e-08, 2.675071e-08, 2.619869e-08, 
    2.466236e-08, 2.195096e-08, 2.020113e-08, 1.920162e-08, 1.75233e-08, 
    1.544841e-08, 1.31063e-08, 1.165178e-08, 1.073526e-08, 9.921218e-09,
  2.702737e-08, 2.705267e-08, 2.689617e-08, 2.705143e-08, 2.661379e-08, 
    2.590941e-08, 2.346895e-08, 2.095949e-08, 1.972905e-08, 1.806411e-08, 
    1.604486e-08, 1.357266e-08, 1.183016e-08, 1.080605e-08, 9.998309e-09,
  2.626197e-08, 2.690013e-08, 2.69445e-08, 2.696675e-08, 2.688983e-08, 
    2.632549e-08, 2.465341e-08, 2.222864e-08, 2.012967e-08, 1.854092e-08, 
    1.658308e-08, 1.411683e-08, 1.209752e-08, 1.094858e-08, 1.007001e-08,
  2.578923e-08, 2.639001e-08, 2.685621e-08, 2.695037e-08, 2.69789e-08, 
    2.672975e-08, 2.558725e-08, 2.329674e-08, 2.09367e-08, 1.892818e-08, 
    1.704971e-08, 1.470679e-08, 1.245659e-08, 1.113493e-08, 1.014855e-08,
  2.550657e-08, 2.572018e-08, 2.649053e-08, 2.670209e-08, 2.695324e-08, 
    2.704465e-08, 2.643205e-08, 2.43669e-08, 2.166736e-08, 1.955822e-08, 
    1.739786e-08, 1.528405e-08, 1.289056e-08, 1.136148e-08, 1.028523e-08,
  2.515822e-08, 2.5144e-08, 2.613008e-08, 2.645915e-08, 2.689319e-08, 
    2.741419e-08, 2.70543e-08, 2.53066e-08, 2.248441e-08, 2.014849e-08, 
    1.789734e-08, 1.587331e-08, 1.3373e-08, 1.16646e-08, 1.048689e-08,
  2.059665e-08, 2.00953e-08, 2.008546e-08, 1.916998e-08, 1.81138e-08, 
    1.699524e-08, 1.603833e-08, 1.49936e-08, 1.374269e-08, 1.262723e-08, 
    1.156104e-08, 1.043279e-08, 9.445153e-09, 8.533144e-09, 7.600447e-09,
  1.997908e-08, 1.974253e-08, 2.006052e-08, 1.902401e-08, 1.785009e-08, 
    1.691054e-08, 1.597807e-08, 1.515123e-08, 1.405787e-08, 1.30202e-08, 
    1.199151e-08, 1.083904e-08, 9.798418e-09, 8.780967e-09, 7.757983e-09,
  2.024353e-08, 1.948354e-08, 1.985247e-08, 1.901166e-08, 1.778763e-08, 
    1.686103e-08, 1.592326e-08, 1.508931e-08, 1.418078e-08, 1.327868e-08, 
    1.228508e-08, 1.115558e-08, 1.009838e-08, 9.026635e-09, 7.907917e-09,
  2.081426e-08, 1.96331e-08, 1.96827e-08, 1.915294e-08, 1.792138e-08, 
    1.697154e-08, 1.591051e-08, 1.50203e-08, 1.416474e-08, 1.337056e-08, 
    1.250008e-08, 1.143538e-08, 1.037607e-08, 9.257685e-09, 8.037826e-09,
  2.094591e-08, 1.984293e-08, 1.94445e-08, 1.928062e-08, 1.810317e-08, 
    1.707539e-08, 1.592924e-08, 1.498696e-08, 1.414701e-08, 1.340244e-08, 
    1.258632e-08, 1.159612e-08, 1.061683e-08, 9.459686e-09, 8.181627e-09,
  2.105291e-08, 2.021232e-08, 1.945564e-08, 1.940362e-08, 1.859757e-08, 
    1.740774e-08, 1.618735e-08, 1.504341e-08, 1.413664e-08, 1.346149e-08, 
    1.27138e-08, 1.177464e-08, 1.084754e-08, 9.651553e-09, 8.319669e-09,
  2.121853e-08, 2.047281e-08, 1.983409e-08, 1.946918e-08, 1.904274e-08, 
    1.793001e-08, 1.671982e-08, 1.53759e-08, 1.420414e-08, 1.350874e-08, 
    1.279402e-08, 1.189523e-08, 1.102949e-08, 9.837682e-09, 8.463775e-09,
  2.131167e-08, 2.074744e-08, 2.021962e-08, 1.986579e-08, 1.926253e-08, 
    1.827903e-08, 1.716595e-08, 1.582616e-08, 1.437718e-08, 1.352322e-08, 
    1.290022e-08, 1.201613e-08, 1.120015e-08, 1.005785e-08, 8.63536e-09,
  2.187758e-08, 2.129426e-08, 2.059394e-08, 2.032351e-08, 1.965775e-08, 
    1.868379e-08, 1.760069e-08, 1.624805e-08, 1.465949e-08, 1.369671e-08, 
    1.305185e-08, 1.220377e-08, 1.138891e-08, 1.03065e-08, 8.848749e-09,
  2.245384e-08, 2.186862e-08, 2.114669e-08, 2.066368e-08, 2.013602e-08, 
    1.908303e-08, 1.810264e-08, 1.667556e-08, 1.496895e-08, 1.382215e-08, 
    1.322548e-08, 1.243688e-08, 1.165531e-08, 1.055875e-08, 9.129898e-09,
  2.531348e-08, 2.479984e-08, 2.425463e-08, 2.301278e-08, 2.168248e-08, 
    2.060752e-08, 1.952261e-08, 1.826208e-08, 1.674158e-08, 1.555179e-08, 
    1.445096e-08, 1.306607e-08, 1.194261e-08, 1.100668e-08, 1.004228e-08,
  2.526903e-08, 2.468883e-08, 2.387635e-08, 2.258059e-08, 2.141565e-08, 
    2.031139e-08, 1.911653e-08, 1.777432e-08, 1.639448e-08, 1.529351e-08, 
    1.43394e-08, 1.30772e-08, 1.193227e-08, 1.10551e-08, 1.012449e-08,
  2.504992e-08, 2.433057e-08, 2.345855e-08, 2.212401e-08, 2.098655e-08, 
    1.990928e-08, 1.868123e-08, 1.744683e-08, 1.617914e-08, 1.517658e-08, 
    1.423903e-08, 1.302793e-08, 1.179309e-08, 1.08974e-08, 1.007461e-08,
  2.446468e-08, 2.378314e-08, 2.272406e-08, 2.151449e-08, 2.057888e-08, 
    1.950113e-08, 1.836285e-08, 1.714273e-08, 1.593629e-08, 1.488215e-08, 
    1.38194e-08, 1.238629e-08, 1.128712e-08, 1.058967e-08, 9.911719e-09,
  2.384075e-08, 2.324166e-08, 2.225893e-08, 2.120285e-08, 2.024061e-08, 
    1.911224e-08, 1.792271e-08, 1.68189e-08, 1.564112e-08, 1.438013e-08, 
    1.305322e-08, 1.181438e-08, 1.082945e-08, 1.009224e-08, 9.805462e-09,
  2.328062e-08, 2.252121e-08, 2.161693e-08, 2.075933e-08, 1.973163e-08, 
    1.859114e-08, 1.755462e-08, 1.639252e-08, 1.502939e-08, 1.371107e-08, 
    1.259767e-08, 1.153391e-08, 1.054847e-08, 9.919199e-09, 9.695871e-09,
  2.25753e-08, 2.16738e-08, 2.090235e-08, 2.015312e-08, 1.916265e-08, 
    1.81145e-08, 1.700459e-08, 1.574697e-08, 1.441551e-08, 1.309914e-08, 
    1.20583e-08, 1.08055e-08, 1.00121e-08, 9.869975e-09, 9.721712e-09,
  2.217589e-08, 2.101901e-08, 2.018705e-08, 1.93669e-08, 1.845581e-08, 
    1.741553e-08, 1.624701e-08, 1.506986e-08, 1.384478e-08, 1.241983e-08, 
    1.126312e-08, 1.026816e-08, 9.768927e-09, 9.71337e-09, 9.730016e-09,
  2.153382e-08, 2.049827e-08, 1.94922e-08, 1.85634e-08, 1.774948e-08, 
    1.684422e-08, 1.565384e-08, 1.46081e-08, 1.338068e-08, 1.185555e-08, 
    1.083418e-08, 1.004507e-08, 9.627782e-09, 9.758038e-09, 9.797163e-09,
  2.069779e-08, 1.965566e-08, 1.886508e-08, 1.806337e-08, 1.713517e-08, 
    1.633855e-08, 1.534752e-08, 1.430492e-08, 1.306654e-08, 1.163856e-08, 
    1.060512e-08, 9.987263e-09, 9.784897e-09, 9.940544e-09, 1.006965e-08,
  2.415058e-08, 2.341407e-08, 2.237616e-08, 2.121057e-08, 2.007814e-08, 
    1.88753e-08, 1.764171e-08, 1.632408e-08, 1.489016e-08, 1.330467e-08, 
    1.210847e-08, 1.098309e-08, 1.012035e-08, 8.980764e-09, 7.813918e-09,
  2.45728e-08, 2.42522e-08, 2.340364e-08, 2.221301e-08, 2.121597e-08, 
    2.009553e-08, 1.897503e-08, 1.782677e-08, 1.669423e-08, 1.502838e-08, 
    1.360429e-08, 1.232676e-08, 1.130714e-08, 1.027655e-08, 9.08057e-09,
  2.540118e-08, 2.495919e-08, 2.436173e-08, 2.343068e-08, 2.232814e-08, 
    2.12382e-08, 2.017212e-08, 1.896282e-08, 1.802827e-08, 1.670976e-08, 
    1.521811e-08, 1.379747e-08, 1.259918e-08, 1.154784e-08, 1.037387e-08,
  2.610496e-08, 2.57044e-08, 2.498247e-08, 2.410495e-08, 2.319893e-08, 
    2.238278e-08, 2.153599e-08, 2.029564e-08, 1.919428e-08, 1.7961e-08, 
    1.665339e-08, 1.519404e-08, 1.376357e-08, 1.26282e-08, 1.152764e-08,
  2.676752e-08, 2.642158e-08, 2.596745e-08, 2.517721e-08, 2.403505e-08, 
    2.305168e-08, 2.234198e-08, 2.137557e-08, 2.026964e-08, 1.902412e-08, 
    1.767871e-08, 1.642057e-08, 1.507283e-08, 1.384478e-08, 1.267599e-08,
  2.784971e-08, 2.738337e-08, 2.69302e-08, 2.614675e-08, 2.511224e-08, 
    2.409889e-08, 2.320965e-08, 2.228625e-08, 2.117032e-08, 1.990155e-08, 
    1.851162e-08, 1.738866e-08, 1.609424e-08, 1.483172e-08, 1.369239e-08,
  2.881081e-08, 2.810891e-08, 2.721836e-08, 2.642177e-08, 2.555423e-08, 
    2.462903e-08, 2.381675e-08, 2.306181e-08, 2.209367e-08, 2.085533e-08, 
    1.939479e-08, 1.809183e-08, 1.699838e-08, 1.590533e-08, 1.466958e-08,
  2.860555e-08, 2.804561e-08, 2.719276e-08, 2.660299e-08, 2.585459e-08, 
    2.513214e-08, 2.43858e-08, 2.357529e-08, 2.255284e-08, 2.132543e-08, 
    1.996134e-08, 1.876115e-08, 1.757941e-08, 1.649053e-08, 1.548843e-08,
  2.817696e-08, 2.771286e-08, 2.689781e-08, 2.631673e-08, 2.547507e-08, 
    2.460436e-08, 2.36505e-08, 2.279934e-08, 2.200615e-08, 2.116388e-08, 
    2.011009e-08, 1.897949e-08, 1.804748e-08, 1.705661e-08, 1.593253e-08,
  2.71748e-08, 2.657495e-08, 2.548066e-08, 2.473996e-08, 2.36802e-08, 
    2.299061e-08, 2.250022e-08, 2.202488e-08, 2.135688e-08, 2.060647e-08, 
    1.969178e-08, 1.897458e-08, 1.828041e-08, 1.730161e-08, 1.618006e-08,
  1.84242e-08, 1.7944e-08, 1.723744e-08, 1.617511e-08, 1.564917e-08, 
    1.483893e-08, 1.346324e-08, 1.202814e-08, 1.102937e-08, 9.882934e-09, 
    8.544378e-09, 7.29447e-09, 5.969505e-09, 4.973634e-09, 4.263301e-09,
  1.898698e-08, 1.84787e-08, 1.78042e-08, 1.670114e-08, 1.589784e-08, 
    1.536415e-08, 1.426918e-08, 1.276261e-08, 1.145233e-08, 1.031111e-08, 
    9.111336e-09, 7.835128e-09, 6.564514e-09, 5.377426e-09, 4.544208e-09,
  1.951847e-08, 1.901823e-08, 1.833298e-08, 1.7265e-08, 1.637402e-08, 
    1.568802e-08, 1.501452e-08, 1.367714e-08, 1.216654e-08, 1.0921e-08, 
    9.773566e-09, 8.515187e-09, 7.224725e-09, 5.883761e-09, 4.885034e-09,
  2.032775e-08, 1.968531e-08, 1.913941e-08, 1.815395e-08, 1.703784e-08, 
    1.619529e-08, 1.557042e-08, 1.459898e-08, 1.316529e-08, 1.173084e-08, 
    1.054669e-08, 9.285177e-09, 7.965058e-09, 6.556445e-09, 5.332296e-09,
  2.142571e-08, 2.040077e-08, 1.988088e-08, 1.914787e-08, 1.802611e-08, 
    1.700575e-08, 1.615679e-08, 1.538504e-08, 1.428174e-08, 1.278034e-08, 
    1.142873e-08, 1.016699e-08, 8.781226e-09, 7.352903e-09, 5.949787e-09,
  2.261768e-08, 2.130638e-08, 2.066261e-08, 2.01215e-08, 1.923784e-08, 
    1.791351e-08, 1.697298e-08, 1.611218e-08, 1.516212e-08, 1.38931e-08, 
    1.242487e-08, 1.105269e-08, 9.671686e-09, 8.191549e-09, 6.68361e-09,
  2.382081e-08, 2.222279e-08, 2.148361e-08, 2.098229e-08, 2.043132e-08, 
    1.930405e-08, 1.79306e-08, 1.687649e-08, 1.591819e-08, 1.486673e-08, 
    1.350045e-08, 1.202769e-08, 1.061293e-08, 9.108805e-09, 7.558617e-09,
  2.455296e-08, 2.332903e-08, 2.222741e-08, 2.168051e-08, 2.121751e-08, 
    2.044946e-08, 1.926898e-08, 1.776939e-08, 1.65581e-08, 1.554855e-08, 
    1.448383e-08, 1.299429e-08, 1.154241e-08, 1.004555e-08, 8.478848e-09,
  2.48816e-08, 2.403551e-08, 2.30854e-08, 2.242108e-08, 2.193787e-08, 
    2.143278e-08, 2.052218e-08, 1.914315e-08, 1.756458e-08, 1.621584e-08, 
    1.522984e-08, 1.410456e-08, 1.25494e-08, 1.09652e-08, 9.347352e-09,
  2.510145e-08, 2.440762e-08, 2.350819e-08, 2.280316e-08, 2.232097e-08, 
    2.194053e-08, 2.142347e-08, 2.049988e-08, 1.898296e-08, 1.728426e-08, 
    1.585975e-08, 1.485835e-08, 1.355523e-08, 1.206359e-08, 1.034308e-08,
  1.505181e-08, 1.413322e-08, 1.358091e-08, 1.307517e-08, 1.293528e-08, 
    1.277108e-08, 1.244778e-08, 1.192947e-08, 1.126926e-08, 1.065241e-08, 
    9.851948e-09, 9.029955e-09, 8.139871e-09, 7.450554e-09, 6.628613e-09,
  1.47413e-08, 1.407501e-08, 1.356757e-08, 1.313419e-08, 1.295708e-08, 
    1.283332e-08, 1.255866e-08, 1.218414e-08, 1.166193e-08, 1.107692e-08, 
    1.044567e-08, 9.651739e-09, 8.638513e-09, 7.796367e-09, 7.112198e-09,
  1.463612e-08, 1.397907e-08, 1.349491e-08, 1.309181e-08, 1.288496e-08, 
    1.282616e-08, 1.265306e-08, 1.234711e-08, 1.193112e-08, 1.133861e-08, 
    1.081382e-08, 1.027193e-08, 9.360084e-09, 8.297771e-09, 7.491262e-09,
  1.444822e-08, 1.390854e-08, 1.338896e-08, 1.298953e-08, 1.273292e-08, 
    1.269353e-08, 1.266928e-08, 1.249352e-08, 1.217582e-08, 1.166395e-08, 
    1.107263e-08, 1.070137e-08, 1.004465e-08, 8.954751e-09, 7.949267e-09,
  1.431262e-08, 1.390571e-08, 1.340467e-08, 1.294225e-08, 1.259387e-08, 
    1.252555e-08, 1.254013e-08, 1.239847e-08, 1.22083e-08, 1.188211e-08, 
    1.139778e-08, 1.098759e-08, 1.060386e-08, 9.692473e-09, 8.582783e-09,
  1.432032e-08, 1.398102e-08, 1.34925e-08, 1.299358e-08, 1.261184e-08, 
    1.248804e-08, 1.245331e-08, 1.238125e-08, 1.215691e-08, 1.195604e-08, 
    1.159562e-08, 1.125485e-08, 1.096856e-08, 1.036394e-08, 9.298954e-09,
  1.456372e-08, 1.40863e-08, 1.365187e-08, 1.326514e-08, 1.279886e-08, 
    1.256598e-08, 1.240771e-08, 1.232739e-08, 1.216761e-08, 1.2027e-08, 
    1.177937e-08, 1.148018e-08, 1.118958e-08, 1.086009e-08, 1.00026e-08,
  1.546183e-08, 1.443637e-08, 1.383456e-08, 1.356413e-08, 1.328666e-08, 
    1.296715e-08, 1.270193e-08, 1.249335e-08, 1.236494e-08, 1.216223e-08, 
    1.201591e-08, 1.173961e-08, 1.145121e-08, 1.120702e-08, 1.064254e-08,
  1.64905e-08, 1.54602e-08, 1.440775e-08, 1.396314e-08, 1.370979e-08, 
    1.342886e-08, 1.322397e-08, 1.301199e-08, 1.285568e-08, 1.275549e-08, 
    1.244256e-08, 1.221488e-08, 1.185214e-08, 1.153259e-08, 1.111418e-08,
  1.773191e-08, 1.657954e-08, 1.555292e-08, 1.471812e-08, 1.429141e-08, 
    1.391171e-08, 1.369915e-08, 1.355482e-08, 1.335853e-08, 1.324117e-08, 
    1.306827e-08, 1.278793e-08, 1.240987e-08, 1.197475e-08, 1.156451e-08,
  2.709094e-08, 2.406304e-08, 2.26021e-08, 2.181515e-08, 2.172623e-08, 
    2.150773e-08, 2.107546e-08, 2.000493e-08, 1.901574e-08, 1.785108e-08, 
    1.608973e-08, 1.46625e-08, 1.35949e-08, 1.197835e-08, 9.959783e-09,
  2.794155e-08, 2.475624e-08, 2.263114e-08, 2.133607e-08, 2.07305e-08, 
    2.049451e-08, 2.033398e-08, 1.954549e-08, 1.895925e-08, 1.793125e-08, 
    1.665561e-08, 1.493485e-08, 1.373473e-08, 1.233751e-08, 1.049895e-08,
  2.859604e-08, 2.538062e-08, 2.265618e-08, 2.084179e-08, 1.990146e-08, 
    1.945074e-08, 1.963439e-08, 1.886407e-08, 1.838754e-08, 1.754636e-08, 
    1.644697e-08, 1.504301e-08, 1.3771e-08, 1.249572e-08, 1.091373e-08,
  2.891817e-08, 2.593386e-08, 2.280186e-08, 2.051854e-08, 1.928677e-08, 
    1.872221e-08, 1.876266e-08, 1.832254e-08, 1.760275e-08, 1.698339e-08, 
    1.594658e-08, 1.481958e-08, 1.372951e-08, 1.255467e-08, 1.119232e-08,
  2.899947e-08, 2.597141e-08, 2.257896e-08, 2.018591e-08, 1.897202e-08, 
    1.832711e-08, 1.82524e-08, 1.776271e-08, 1.700979e-08, 1.628287e-08, 
    1.535453e-08, 1.437275e-08, 1.344265e-08, 1.238432e-08, 1.132086e-08,
  2.83906e-08, 2.537745e-08, 2.213379e-08, 1.996015e-08, 1.876021e-08, 
    1.804879e-08, 1.779389e-08, 1.727437e-08, 1.654294e-08, 1.585451e-08, 
    1.488044e-08, 1.392473e-08, 1.309306e-08, 1.219205e-08, 1.13042e-08,
  2.703112e-08, 2.449161e-08, 2.176322e-08, 1.988836e-08, 1.847619e-08, 
    1.764138e-08, 1.722452e-08, 1.664899e-08, 1.595988e-08, 1.541447e-08, 
    1.458551e-08, 1.358197e-08, 1.270529e-08, 1.192029e-08, 1.1207e-08,
  2.581082e-08, 2.382633e-08, 2.146663e-08, 1.966531e-08, 1.830829e-08, 
    1.731049e-08, 1.667256e-08, 1.600464e-08, 1.542433e-08, 1.491025e-08, 
    1.421632e-08, 1.335157e-08, 1.242992e-08, 1.166462e-08, 1.111047e-08,
  2.485747e-08, 2.341446e-08, 2.117917e-08, 1.95369e-08, 1.821328e-08, 
    1.707071e-08, 1.637629e-08, 1.573423e-08, 1.508377e-08, 1.447315e-08, 
    1.384266e-08, 1.319876e-08, 1.230546e-08, 1.150407e-08, 1.103938e-08,
  2.464614e-08, 2.321281e-08, 2.089807e-08, 1.922063e-08, 1.813254e-08, 
    1.721224e-08, 1.647632e-08, 1.57106e-08, 1.500613e-08, 1.433125e-08, 
    1.361562e-08, 1.296163e-08, 1.220763e-08, 1.146884e-08, 1.101714e-08,
  2.305009e-08, 2.165222e-08, 2.137061e-08, 2.046174e-08, 1.910494e-08, 
    1.678807e-08, 1.62067e-08, 1.555078e-08, 1.512579e-08, 1.493318e-08, 
    1.484651e-08, 1.498477e-08, 1.513877e-08, 1.521904e-08, 1.462124e-08,
  2.409295e-08, 2.257767e-08, 2.15968e-08, 2.0755e-08, 2.026401e-08, 
    1.834371e-08, 1.68703e-08, 1.613203e-08, 1.584639e-08, 1.552389e-08, 
    1.515378e-08, 1.513295e-08, 1.5316e-08, 1.55391e-08, 1.527771e-08,
  2.529658e-08, 2.346816e-08, 2.211328e-08, 2.102371e-08, 2.079826e-08, 
    1.924159e-08, 1.782918e-08, 1.688923e-08, 1.634667e-08, 1.631498e-08, 
    1.582816e-08, 1.554393e-08, 1.547126e-08, 1.572262e-08, 1.57722e-08,
  2.584645e-08, 2.434052e-08, 2.276778e-08, 2.15206e-08, 2.095692e-08, 
    2.01066e-08, 1.832929e-08, 1.728105e-08, 1.701894e-08, 1.681722e-08, 
    1.685671e-08, 1.601064e-08, 1.581686e-08, 1.595019e-08, 1.618396e-08,
  2.563587e-08, 2.533813e-08, 2.327935e-08, 2.187881e-08, 2.117764e-08, 
    2.059749e-08, 1.911522e-08, 1.753816e-08, 1.73359e-08, 1.736976e-08, 
    1.755184e-08, 1.702848e-08, 1.633544e-08, 1.634767e-08, 1.659901e-08,
  2.535465e-08, 2.561431e-08, 2.418436e-08, 2.218949e-08, 2.114091e-08, 
    2.071267e-08, 2.01261e-08, 1.812935e-08, 1.751121e-08, 1.773058e-08, 
    1.810813e-08, 1.78894e-08, 1.707975e-08, 1.668702e-08, 1.690455e-08,
  2.551556e-08, 2.548558e-08, 2.462882e-08, 2.291636e-08, 2.114873e-08, 
    2.040066e-08, 2.043829e-08, 1.934658e-08, 1.809112e-08, 1.797572e-08, 
    1.859457e-08, 1.863664e-08, 1.820183e-08, 1.732521e-08, 1.731297e-08,
  2.631182e-08, 2.574507e-08, 2.488289e-08, 2.34726e-08, 2.167418e-08, 
    2.018878e-08, 1.99945e-08, 1.987611e-08, 1.916397e-08, 1.845217e-08, 
    1.894204e-08, 1.927126e-08, 1.898353e-08, 1.807971e-08, 1.763786e-08,
  2.707674e-08, 2.620075e-08, 2.534711e-08, 2.384283e-08, 2.229598e-08, 
    2.043447e-08, 1.938361e-08, 1.918269e-08, 1.912161e-08, 1.903603e-08, 
    1.917108e-08, 1.952856e-08, 1.958244e-08, 1.894641e-08, 1.819095e-08,
  2.755135e-08, 2.668531e-08, 2.57853e-08, 2.395054e-08, 2.277883e-08, 
    2.087641e-08, 1.920694e-08, 1.845609e-08, 1.842816e-08, 1.895312e-08, 
    1.935075e-08, 1.971485e-08, 1.98813e-08, 1.961513e-08, 1.899344e-08,
  1.696427e-08, 1.608858e-08, 1.606626e-08, 1.666282e-08, 1.679457e-08, 
    1.596517e-08, 1.495362e-08, 1.387656e-08, 1.281781e-08, 1.19659e-08, 
    1.156192e-08, 1.161646e-08, 1.183921e-08, 1.180062e-08, 1.16843e-08,
  1.816336e-08, 1.712485e-08, 1.62439e-08, 1.611381e-08, 1.661861e-08, 
    1.651586e-08, 1.52763e-08, 1.432009e-08, 1.351347e-08, 1.238095e-08, 
    1.173691e-08, 1.16303e-08, 1.183513e-08, 1.191779e-08, 1.185045e-08,
  1.919323e-08, 1.822886e-08, 1.722979e-08, 1.665459e-08, 1.645947e-08, 
    1.681572e-08, 1.590275e-08, 1.4805e-08, 1.404407e-08, 1.294326e-08, 
    1.203512e-08, 1.16438e-08, 1.168922e-08, 1.198463e-08, 1.196942e-08,
  2.04237e-08, 1.969997e-08, 1.820562e-08, 1.73922e-08, 1.697711e-08, 
    1.703771e-08, 1.658421e-08, 1.536105e-08, 1.466088e-08, 1.35394e-08, 
    1.253229e-08, 1.177333e-08, 1.146102e-08, 1.178161e-08, 1.199155e-08,
  2.071557e-08, 2.085e-08, 2.017094e-08, 1.853313e-08, 1.76852e-08, 
    1.736855e-08, 1.711306e-08, 1.606629e-08, 1.519079e-08, 1.414584e-08, 
    1.308708e-08, 1.230636e-08, 1.144001e-08, 1.151377e-08, 1.195834e-08,
  2.130683e-08, 2.104523e-08, 2.107102e-08, 2.064871e-08, 1.921815e-08, 
    1.811891e-08, 1.76248e-08, 1.677295e-08, 1.576063e-08, 1.484461e-08, 
    1.368066e-08, 1.272323e-08, 1.190216e-08, 1.138911e-08, 1.180653e-08,
  2.351419e-08, 2.19133e-08, 2.136522e-08, 2.148114e-08, 2.136376e-08, 
    1.990532e-08, 1.846684e-08, 1.748856e-08, 1.638286e-08, 1.542823e-08, 
    1.441786e-08, 1.335024e-08, 1.250073e-08, 1.171886e-08, 1.173114e-08,
  2.433285e-08, 2.363743e-08, 2.212379e-08, 2.159524e-08, 2.189125e-08, 
    2.180092e-08, 2.043164e-08, 1.848389e-08, 1.719087e-08, 1.604062e-08, 
    1.508471e-08, 1.417604e-08, 1.323887e-08, 1.245054e-08, 1.186184e-08,
  2.514432e-08, 2.40979e-08, 2.35387e-08, 2.231014e-08, 2.188027e-08, 
    2.208559e-08, 2.203649e-08, 2.062303e-08, 1.840129e-08, 1.672847e-08, 
    1.564312e-08, 1.48224e-08, 1.402998e-08, 1.317623e-08, 1.245609e-08,
  2.555449e-08, 2.438478e-08, 2.350373e-08, 2.301041e-08, 2.226979e-08, 
    2.199395e-08, 2.22036e-08, 2.196674e-08, 2.061348e-08, 1.815356e-08, 
    1.633912e-08, 1.542736e-08, 1.468322e-08, 1.389284e-08, 1.322697e-08,
  2.056487e-08, 2.009232e-08, 1.928373e-08, 1.864959e-08, 1.731082e-08, 
    1.600575e-08, 1.480603e-08, 1.417214e-08, 1.378846e-08, 1.326991e-08, 
    1.271069e-08, 1.180206e-08, 1.121931e-08, 1.089872e-08, 1.029588e-08,
  2.010356e-08, 1.946396e-08, 1.892427e-08, 1.859981e-08, 1.763032e-08, 
    1.651641e-08, 1.487906e-08, 1.413963e-08, 1.377383e-08, 1.351461e-08, 
    1.321539e-08, 1.248464e-08, 1.15614e-08, 1.083087e-08, 1.049957e-08,
  2.03189e-08, 1.928128e-08, 1.868364e-08, 1.827579e-08, 1.750817e-08, 
    1.678834e-08, 1.539337e-08, 1.416908e-08, 1.359534e-08, 1.331844e-08, 
    1.31929e-08, 1.265623e-08, 1.180045e-08, 1.082063e-08, 1.050012e-08,
  2.122115e-08, 1.948731e-08, 1.871761e-08, 1.817112e-08, 1.725911e-08, 
    1.660982e-08, 1.575211e-08, 1.456075e-08, 1.367761e-08, 1.32004e-08, 
    1.299556e-08, 1.250132e-08, 1.187453e-08, 1.100287e-08, 1.064052e-08,
  2.132013e-08, 1.999534e-08, 1.894112e-08, 1.824818e-08, 1.71981e-08, 
    1.651284e-08, 1.578854e-08, 1.50512e-08, 1.402355e-08, 1.326734e-08, 
    1.294198e-08, 1.234394e-08, 1.178834e-08, 1.109084e-08, 1.073467e-08,
  2.126794e-08, 1.992143e-08, 1.896396e-08, 1.835368e-08, 1.727566e-08, 
    1.640087e-08, 1.567818e-08, 1.50104e-08, 1.419667e-08, 1.328676e-08, 
    1.280349e-08, 1.231755e-08, 1.175878e-08, 1.119318e-08, 1.077356e-08,
  2.113896e-08, 1.980972e-08, 1.875727e-08, 1.80497e-08, 1.712069e-08, 
    1.622405e-08, 1.53434e-08, 1.463221e-08, 1.400179e-08, 1.320261e-08, 
    1.271618e-08, 1.240843e-08, 1.187712e-08, 1.126012e-08, 1.0862e-08,
  2.099694e-08, 1.967604e-08, 1.86343e-08, 1.800927e-08, 1.711142e-08, 
    1.609862e-08, 1.511543e-08, 1.433355e-08, 1.374693e-08, 1.298215e-08, 
    1.25254e-08, 1.223284e-08, 1.18042e-08, 1.136016e-08, 1.09479e-08,
  2.093031e-08, 1.969239e-08, 1.861759e-08, 1.789765e-08, 1.693848e-08, 
    1.614763e-08, 1.520035e-08, 1.427398e-08, 1.357494e-08, 1.279549e-08, 
    1.211113e-08, 1.190213e-08, 1.160123e-08, 1.146928e-08, 1.128313e-08,
  2.060112e-08, 1.953999e-08, 1.870745e-08, 1.806109e-08, 1.698094e-08, 
    1.59325e-08, 1.512001e-08, 1.424172e-08, 1.345527e-08, 1.266462e-08, 
    1.186461e-08, 1.141298e-08, 1.122208e-08, 1.135019e-08, 1.161458e-08,
  1.797491e-08, 1.787496e-08, 1.751483e-08, 1.717037e-08, 1.680113e-08, 
    1.627313e-08, 1.597633e-08, 1.506259e-08, 1.38159e-08, 1.251367e-08, 
    1.189367e-08, 1.088976e-08, 1.05911e-08, 1.130196e-08, 1.370584e-08,
  1.796465e-08, 1.81068e-08, 1.802684e-08, 1.756706e-08, 1.711673e-08, 
    1.678658e-08, 1.648386e-08, 1.610837e-08, 1.546764e-08, 1.428184e-08, 
    1.318183e-08, 1.253694e-08, 1.21898e-08, 1.220972e-08, 1.405751e-08,
  1.815249e-08, 1.832417e-08, 1.840013e-08, 1.815191e-08, 1.767489e-08, 
    1.720582e-08, 1.689321e-08, 1.657044e-08, 1.636604e-08, 1.586651e-08, 
    1.503902e-08, 1.418184e-08, 1.41482e-08, 1.424378e-08, 1.493117e-08,
  1.842258e-08, 1.848926e-08, 1.879366e-08, 1.878963e-08, 1.843103e-08, 
    1.787624e-08, 1.744053e-08, 1.692973e-08, 1.650043e-08, 1.637306e-08, 
    1.614812e-08, 1.556733e-08, 1.563232e-08, 1.592534e-08, 1.583734e-08,
  1.983524e-08, 1.960277e-08, 1.881478e-08, 1.899397e-08, 1.902538e-08, 
    1.862299e-08, 1.802797e-08, 1.742442e-08, 1.686465e-08, 1.648355e-08, 
    1.671975e-08, 1.657012e-08, 1.639684e-08, 1.591449e-08, 1.610628e-08,
  2.067551e-08, 2.046429e-08, 2.018195e-08, 1.933162e-08, 1.900463e-08, 
    1.902793e-08, 1.889629e-08, 1.82575e-08, 1.779305e-08, 1.726516e-08, 
    1.706901e-08, 1.704419e-08, 1.683519e-08, 1.605258e-08, 1.58498e-08,
  2.130697e-08, 2.113839e-08, 2.089452e-08, 2.066025e-08, 2.003186e-08, 
    1.93237e-08, 1.922931e-08, 1.920479e-08, 1.903742e-08, 1.842256e-08, 
    1.783798e-08, 1.761096e-08, 1.749225e-08, 1.667229e-08, 1.532637e-08,
  2.168737e-08, 2.16452e-08, 2.154994e-08, 2.131912e-08, 2.066797e-08, 
    2.025924e-08, 1.992144e-08, 1.962347e-08, 1.957889e-08, 1.961982e-08, 
    1.896206e-08, 1.846363e-08, 1.801967e-08, 1.731285e-08, 1.529458e-08,
  2.196169e-08, 2.211829e-08, 2.205827e-08, 2.197605e-08, 2.149784e-08, 
    2.0757e-08, 2.024724e-08, 2.004337e-08, 1.981053e-08, 1.995546e-08, 
    1.988163e-08, 1.949534e-08, 1.869855e-08, 1.783033e-08, 1.58403e-08,
  2.259247e-08, 2.242227e-08, 2.245635e-08, 2.246584e-08, 2.200943e-08, 
    2.140467e-08, 2.054515e-08, 2.009836e-08, 1.969728e-08, 1.965964e-08, 
    1.986148e-08, 1.984711e-08, 1.921929e-08, 1.83245e-08, 1.654969e-08,
  1.208423e-08, 1.147213e-08, 1.100294e-08, 1.012915e-08, 9.807033e-09, 
    9.882434e-09, 1.008727e-08, 1.014964e-08, 1.018163e-08, 1.031207e-08, 
    1.037575e-08, 1.046335e-08, 1.054748e-08, 1.092069e-08, 1.109125e-08,
  1.223588e-08, 1.173483e-08, 1.131956e-08, 1.080935e-08, 1.030196e-08, 
    1.021934e-08, 1.036184e-08, 1.054182e-08, 1.062735e-08, 1.077326e-08, 
    1.090109e-08, 1.098572e-08, 1.104365e-08, 1.131104e-08, 1.172589e-08,
  1.217686e-08, 1.189909e-08, 1.14516e-08, 1.110393e-08, 1.062812e-08, 
    1.047086e-08, 1.060113e-08, 1.076655e-08, 1.105675e-08, 1.126012e-08, 
    1.156353e-08, 1.165979e-08, 1.182536e-08, 1.19715e-08, 1.233504e-08,
  1.215079e-08, 1.203944e-08, 1.174296e-08, 1.136825e-08, 1.092772e-08, 
    1.065976e-08, 1.071819e-08, 1.094539e-08, 1.131949e-08, 1.160266e-08, 
    1.209435e-08, 1.230967e-08, 1.25919e-08, 1.274366e-08, 1.300616e-08,
  1.263142e-08, 1.226327e-08, 1.20655e-08, 1.18469e-08, 1.146537e-08, 
    1.107356e-08, 1.09758e-08, 1.111982e-08, 1.14921e-08, 1.184547e-08, 
    1.239525e-08, 1.276283e-08, 1.314119e-08, 1.350569e-08, 1.365784e-08,
  1.312633e-08, 1.27235e-08, 1.235331e-08, 1.20995e-08, 1.18361e-08, 
    1.154838e-08, 1.133522e-08, 1.138445e-08, 1.168629e-08, 1.202627e-08, 
    1.248549e-08, 1.299847e-08, 1.356949e-08, 1.410685e-08, 1.438181e-08,
  1.372625e-08, 1.333146e-08, 1.302613e-08, 1.279069e-08, 1.233569e-08, 
    1.197889e-08, 1.168064e-08, 1.154115e-08, 1.163731e-08, 1.201439e-08, 
    1.257245e-08, 1.306207e-08, 1.398598e-08, 1.468515e-08, 1.512919e-08,
  1.462658e-08, 1.398339e-08, 1.360254e-08, 1.340483e-08, 1.316206e-08, 
    1.277171e-08, 1.240883e-08, 1.202909e-08, 1.189218e-08, 1.213859e-08, 
    1.251873e-08, 1.321576e-08, 1.425682e-08, 1.520259e-08, 1.575005e-08,
  1.572532e-08, 1.493503e-08, 1.443465e-08, 1.417693e-08, 1.383545e-08, 
    1.350475e-08, 1.322883e-08, 1.287612e-08, 1.260948e-08, 1.269206e-08, 
    1.290728e-08, 1.353996e-08, 1.466619e-08, 1.569975e-08, 1.627591e-08,
  1.726674e-08, 1.617249e-08, 1.534733e-08, 1.513832e-08, 1.507155e-08, 
    1.470939e-08, 1.427382e-08, 1.384029e-08, 1.349761e-08, 1.360558e-08, 
    1.386391e-08, 1.439054e-08, 1.515717e-08, 1.654472e-08, 1.68205e-08,
  1.046006e-08, 9.168367e-09, 8.201464e-09, 7.281364e-09, 6.688359e-09, 
    6.149168e-09, 5.963189e-09, 5.76836e-09, 5.676728e-09, 5.706324e-09, 
    5.69807e-09, 5.687752e-09, 5.699226e-09, 5.836586e-09, 5.91443e-09,
  1.134634e-08, 1.00098e-08, 9.074668e-09, 8.00291e-09, 7.15539e-09, 
    6.496192e-09, 6.120756e-09, 5.940524e-09, 5.922304e-09, 5.994703e-09, 
    5.992611e-09, 5.961142e-09, 5.866914e-09, 5.959814e-09, 5.96625e-09,
  1.19998e-08, 1.104935e-08, 1.001699e-08, 8.90023e-09, 7.929866e-09, 
    7.102137e-09, 6.569584e-09, 6.223604e-09, 6.289536e-09, 6.444498e-09, 
    6.439385e-09, 6.348913e-09, 6.229666e-09, 6.128678e-09, 6.115014e-09,
  1.246358e-08, 1.17465e-08, 1.099787e-08, 9.823574e-09, 8.64349e-09, 
    7.874582e-09, 7.243049e-09, 6.703367e-09, 6.709176e-09, 6.893883e-09, 
    6.872134e-09, 6.678387e-09, 6.596874e-09, 6.387474e-09, 6.464298e-09,
  1.283847e-08, 1.216484e-08, 1.137007e-08, 1.050479e-08, 9.367407e-09, 
    8.575093e-09, 8.020409e-09, 7.454398e-09, 7.113304e-09, 7.231096e-09, 
    7.21645e-09, 7.051548e-09, 6.929828e-09, 6.739684e-09, 6.931747e-09,
  1.327786e-08, 1.26326e-08, 1.180362e-08, 1.097268e-08, 1.004884e-08, 
    9.181709e-09, 8.701851e-09, 8.241549e-09, 7.714116e-09, 7.559544e-09, 
    7.600488e-09, 7.396455e-09, 7.199957e-09, 7.05377e-09, 7.449211e-09,
  1.357542e-08, 1.309468e-08, 1.23745e-08, 1.14379e-08, 1.058848e-08, 
    9.739338e-09, 9.229771e-09, 8.941552e-09, 8.529224e-09, 8.05496e-09, 
    8.024253e-09, 7.887152e-09, 7.516517e-09, 7.437749e-09, 7.994925e-09,
  1.395002e-08, 1.335084e-08, 1.281458e-08, 1.205014e-08, 1.113463e-08, 
    1.030192e-08, 9.707509e-09, 9.424894e-09, 9.240307e-09, 8.727903e-09, 
    8.495126e-09, 8.310146e-09, 7.910101e-09, 7.877281e-09, 8.451564e-09,
  1.446987e-08, 1.363629e-08, 1.314822e-08, 1.251334e-08, 1.175171e-08, 
    1.09654e-08, 1.026372e-08, 9.910507e-09, 9.682542e-09, 9.409945e-09, 
    9.064325e-09, 8.713804e-09, 8.400126e-09, 8.465062e-09, 9.18241e-09,
  1.532644e-08, 1.407698e-08, 1.340605e-08, 1.282894e-08, 1.215179e-08, 
    1.146782e-08, 1.07898e-08, 1.031466e-08, 9.953649e-09, 9.802024e-09, 
    9.647822e-09, 9.321043e-09, 8.992778e-09, 9.199697e-09, 9.809849e-09,
  1.464212e-08, 1.343625e-08, 1.226008e-08, 1.065555e-08, 9.193798e-09, 
    8.161177e-09, 7.463818e-09, 6.797961e-09, 6.123535e-09, 5.634249e-09, 
    5.140566e-09, 4.777606e-09, 4.584682e-09, 4.554324e-09, 4.549324e-09,
  1.418984e-08, 1.298747e-08, 1.157343e-08, 9.744389e-09, 8.540298e-09, 
    7.601637e-09, 6.872392e-09, 6.197367e-09, 5.620411e-09, 5.195099e-09, 
    4.775445e-09, 4.516703e-09, 4.46388e-09, 4.443056e-09, 4.465621e-09,
  1.392168e-08, 1.254601e-08, 1.089926e-08, 9.029301e-09, 7.947134e-09, 
    7.01681e-09, 6.266643e-09, 5.702072e-09, 5.206801e-09, 4.863442e-09, 
    4.553292e-09, 4.357957e-09, 4.324247e-09, 4.390281e-09, 4.394232e-09,
  1.35531e-08, 1.227048e-08, 1.047161e-08, 8.62016e-09, 7.545127e-09, 
    6.553736e-09, 5.832325e-09, 5.303811e-09, 4.874618e-09, 4.617253e-09, 
    4.372427e-09, 4.223566e-09, 4.239199e-09, 4.340234e-09, 4.352148e-09,
  1.316784e-08, 1.200135e-08, 1.020535e-08, 8.436446e-09, 7.215954e-09, 
    6.178871e-09, 5.407036e-09, 5.024985e-09, 4.723614e-09, 4.505132e-09, 
    4.248445e-09, 4.142153e-09, 4.193374e-09, 4.366857e-09, 4.338999e-09,
  1.292216e-08, 1.186087e-08, 1.014798e-08, 8.379088e-09, 7.172778e-09, 
    5.953381e-09, 5.257092e-09, 4.859265e-09, 4.630611e-09, 4.408257e-09, 
    4.172453e-09, 4.054861e-09, 4.187816e-09, 4.364507e-09, 4.388259e-09,
  1.294044e-08, 1.179904e-08, 1.021488e-08, 8.431974e-09, 7.151485e-09, 
    5.99773e-09, 5.322158e-09, 4.841219e-09, 4.574604e-09, 4.378582e-09, 
    4.134506e-09, 4.032475e-09, 4.219634e-09, 4.423564e-09, 4.509058e-09,
  1.308492e-08, 1.188653e-08, 1.040136e-08, 8.689089e-09, 7.290454e-09, 
    6.189974e-09, 5.538217e-09, 4.957843e-09, 4.563576e-09, 4.328469e-09, 
    4.11487e-09, 4.029903e-09, 4.27062e-09, 4.469003e-09, 4.681316e-09,
  1.337286e-08, 1.215997e-08, 1.060034e-08, 8.991853e-09, 7.68382e-09, 
    6.492999e-09, 5.820397e-09, 5.134721e-09, 4.694483e-09, 4.372151e-09, 
    4.115654e-09, 4.065355e-09, 4.317782e-09, 4.498857e-09, 4.832118e-09,
  1.371669e-08, 1.24631e-08, 1.095559e-08, 9.317514e-09, 8.111272e-09, 
    6.945916e-09, 6.165238e-09, 5.416375e-09, 4.848419e-09, 4.433138e-09, 
    4.217954e-09, 4.158051e-09, 4.344921e-09, 4.513194e-09, 4.957435e-09,
  2.371024e-08, 2.193186e-08, 2.026754e-08, 1.860007e-08, 1.665816e-08, 
    1.553403e-08, 1.54625e-08, 1.586847e-08, 1.665553e-08, 1.67811e-08, 
    1.641618e-08, 1.58761e-08, 1.504923e-08, 1.422414e-08, 1.344681e-08,
  2.399553e-08, 2.260384e-08, 2.081272e-08, 1.900207e-08, 1.686059e-08, 
    1.571691e-08, 1.569778e-08, 1.599828e-08, 1.65301e-08, 1.656754e-08, 
    1.596137e-08, 1.51315e-08, 1.415337e-08, 1.325072e-08, 1.236444e-08,
  2.426374e-08, 2.317128e-08, 2.132984e-08, 1.921563e-08, 1.700554e-08, 
    1.582063e-08, 1.576037e-08, 1.595196e-08, 1.6222e-08, 1.603627e-08, 
    1.541143e-08, 1.447478e-08, 1.33046e-08, 1.239685e-08, 1.142866e-08,
  2.430068e-08, 2.348389e-08, 2.15144e-08, 1.913231e-08, 1.700522e-08, 
    1.583605e-08, 1.567334e-08, 1.569736e-08, 1.581146e-08, 1.54552e-08, 
    1.488494e-08, 1.361989e-08, 1.244121e-08, 1.143167e-08, 1.062046e-08,
  2.415772e-08, 2.340116e-08, 2.132373e-08, 1.891074e-08, 1.695468e-08, 
    1.580115e-08, 1.544352e-08, 1.532027e-08, 1.521308e-08, 1.484236e-08, 
    1.420688e-08, 1.26649e-08, 1.147152e-08, 1.051112e-08, 1.000286e-08,
  2.396381e-08, 2.305792e-08, 2.089634e-08, 1.855876e-08, 1.678084e-08, 
    1.564191e-08, 1.5128e-08, 1.485842e-08, 1.458526e-08, 1.436335e-08, 
    1.325305e-08, 1.167743e-08, 1.053363e-08, 9.802954e-09, 9.498433e-09,
  2.369621e-08, 2.253399e-08, 2.031989e-08, 1.81343e-08, 1.655575e-08, 
    1.53925e-08, 1.473122e-08, 1.43813e-08, 1.404061e-08, 1.385563e-08, 
    1.222181e-08, 1.072795e-08, 9.712154e-09, 9.198798e-09, 8.871486e-09,
  2.333729e-08, 2.19814e-08, 1.977971e-08, 1.767265e-08, 1.62795e-08, 
    1.508722e-08, 1.436342e-08, 1.392949e-08, 1.35764e-08, 1.327563e-08, 
    1.126334e-08, 9.800315e-09, 9.040269e-09, 8.600788e-09, 8.24823e-09,
  2.287892e-08, 2.136932e-08, 1.92114e-08, 1.721869e-08, 1.589862e-08, 
    1.479572e-08, 1.408428e-08, 1.357019e-08, 1.319993e-08, 1.241961e-08, 
    1.025061e-08, 9.020027e-09, 8.396633e-09, 7.981694e-09, 7.680197e-09,
  2.231622e-08, 2.080424e-08, 1.8591e-08, 1.673757e-08, 1.558533e-08, 
    1.450492e-08, 1.389009e-08, 1.317471e-08, 1.280741e-08, 1.134109e-08, 
    9.326681e-09, 8.341924e-09, 7.830632e-09, 7.439722e-09, 7.253314e-09,
  2.311167e-08, 2.18544e-08, 2.090093e-08, 1.938023e-08, 1.812221e-08, 
    1.697793e-08, 1.594339e-08, 1.513063e-08, 1.444802e-08, 1.362396e-08, 
    1.281847e-08, 1.241066e-08, 1.204261e-08, 1.19723e-08, 1.217983e-08,
  2.390877e-08, 2.246728e-08, 2.122498e-08, 1.971341e-08, 1.826817e-08, 
    1.698754e-08, 1.57235e-08, 1.475766e-08, 1.413728e-08, 1.334539e-08, 
    1.274179e-08, 1.237525e-08, 1.216536e-08, 1.238411e-08, 1.267847e-08,
  2.452369e-08, 2.300485e-08, 2.153252e-08, 1.993627e-08, 1.843972e-08, 
    1.705345e-08, 1.56614e-08, 1.455062e-08, 1.389957e-08, 1.323609e-08, 
    1.277625e-08, 1.237362e-08, 1.234399e-08, 1.269054e-08, 1.315231e-08,
  2.486777e-08, 2.343363e-08, 2.166524e-08, 1.994956e-08, 1.847775e-08, 
    1.712176e-08, 1.54911e-08, 1.428942e-08, 1.359442e-08, 1.309148e-08, 
    1.266183e-08, 1.240283e-08, 1.250316e-08, 1.302833e-08, 1.354751e-08,
  2.492887e-08, 2.37945e-08, 2.174353e-08, 1.986901e-08, 1.836751e-08, 
    1.710341e-08, 1.54554e-08, 1.417091e-08, 1.349843e-08, 1.302031e-08, 
    1.251767e-08, 1.248713e-08, 1.284779e-08, 1.354707e-08, 1.397474e-08,
  2.478787e-08, 2.395482e-08, 2.181633e-08, 1.974458e-08, 1.813193e-08, 
    1.690035e-08, 1.536252e-08, 1.408783e-08, 1.339058e-08, 1.282979e-08, 
    1.257824e-08, 1.265325e-08, 1.320255e-08, 1.3804e-08, 1.414168e-08,
  2.447053e-08, 2.37412e-08, 2.17813e-08, 1.960407e-08, 1.782781e-08, 
    1.65981e-08, 1.52144e-08, 1.400384e-08, 1.326117e-08, 1.264006e-08, 
    1.270865e-08, 1.296151e-08, 1.360347e-08, 1.416125e-08, 1.397817e-08,
  2.388003e-08, 2.335754e-08, 2.161123e-08, 1.952144e-08, 1.755687e-08, 
    1.629095e-08, 1.506062e-08, 1.387458e-08, 1.310345e-08, 1.249844e-08, 
    1.282955e-08, 1.323415e-08, 1.379088e-08, 1.409535e-08, 1.365127e-08,
  2.338686e-08, 2.29645e-08, 2.141852e-08, 1.930877e-08, 1.724183e-08, 
    1.601394e-08, 1.48391e-08, 1.3738e-08, 1.295552e-08, 1.251439e-08, 
    1.306354e-08, 1.36071e-08, 1.407247e-08, 1.398517e-08, 1.322798e-08,
  2.318188e-08, 2.266607e-08, 2.123782e-08, 1.917684e-08, 1.698582e-08, 
    1.574746e-08, 1.46567e-08, 1.361275e-08, 1.278574e-08, 1.265097e-08, 
    1.338987e-08, 1.382286e-08, 1.404228e-08, 1.365711e-08, 1.296496e-08,
  1.69919e-08, 1.667226e-08, 1.647241e-08, 1.610437e-08, 1.575915e-08, 
    1.534196e-08, 1.494723e-08, 1.468192e-08, 1.445354e-08, 1.436551e-08, 
    1.424695e-08, 1.411673e-08, 1.373403e-08, 1.338323e-08, 1.302967e-08,
  1.712471e-08, 1.680144e-08, 1.659539e-08, 1.61632e-08, 1.572116e-08, 
    1.531196e-08, 1.499446e-08, 1.47701e-08, 1.460221e-08, 1.454873e-08, 
    1.447341e-08, 1.436216e-08, 1.392398e-08, 1.356426e-08, 1.320828e-08,
  1.731806e-08, 1.694477e-08, 1.664415e-08, 1.619801e-08, 1.579236e-08, 
    1.541328e-08, 1.509635e-08, 1.487304e-08, 1.478902e-08, 1.474229e-08, 
    1.464129e-08, 1.456222e-08, 1.415771e-08, 1.377019e-08, 1.339802e-08,
  1.761885e-08, 1.726106e-08, 1.683816e-08, 1.638329e-08, 1.598678e-08, 
    1.556209e-08, 1.522693e-08, 1.49873e-08, 1.497081e-08, 1.497293e-08, 
    1.487309e-08, 1.47766e-08, 1.438759e-08, 1.398889e-08, 1.361021e-08,
  1.797451e-08, 1.760605e-08, 1.710228e-08, 1.66139e-08, 1.623423e-08, 
    1.577544e-08, 1.537191e-08, 1.509792e-08, 1.509935e-08, 1.516191e-08, 
    1.509142e-08, 1.503534e-08, 1.459223e-08, 1.409256e-08, 1.375932e-08,
  1.825355e-08, 1.798772e-08, 1.7446e-08, 1.689785e-08, 1.66356e-08, 
    1.616321e-08, 1.568846e-08, 1.525178e-08, 1.52396e-08, 1.537719e-08, 
    1.531003e-08, 1.521587e-08, 1.471679e-08, 1.418102e-08, 1.382626e-08,
  1.858387e-08, 1.855931e-08, 1.7936e-08, 1.728373e-08, 1.70425e-08, 
    1.66988e-08, 1.609615e-08, 1.547212e-08, 1.529876e-08, 1.549919e-08, 
    1.541787e-08, 1.532996e-08, 1.487825e-08, 1.43094e-08, 1.394598e-08,
  1.907522e-08, 1.911048e-08, 1.858804e-08, 1.780544e-08, 1.747874e-08, 
    1.718087e-08, 1.658298e-08, 1.577417e-08, 1.54314e-08, 1.555845e-08, 
    1.551334e-08, 1.537149e-08, 1.498866e-08, 1.444131e-08, 1.401807e-08,
  1.956489e-08, 1.953298e-08, 1.919392e-08, 1.846015e-08, 1.796379e-08, 
    1.762819e-08, 1.712332e-08, 1.615852e-08, 1.559465e-08, 1.564177e-08, 
    1.553819e-08, 1.536645e-08, 1.504726e-08, 1.451471e-08, 1.405017e-08,
  2.000471e-08, 1.980589e-08, 1.974876e-08, 1.910028e-08, 1.844148e-08, 
    1.802256e-08, 1.754888e-08, 1.668766e-08, 1.584595e-08, 1.57016e-08, 
    1.554709e-08, 1.526754e-08, 1.499765e-08, 1.451276e-08, 1.399736e-08,
  1.552387e-08, 1.501142e-08, 1.459846e-08, 1.430145e-08, 1.444736e-08, 
    1.448373e-08, 1.477163e-08, 1.483768e-08, 1.541517e-08, 1.537192e-08, 
    1.489582e-08, 1.447375e-08, 1.42245e-08, 1.440945e-08, 1.433266e-08,
  1.562262e-08, 1.519254e-08, 1.494212e-08, 1.463125e-08, 1.468029e-08, 
    1.469412e-08, 1.48341e-08, 1.511191e-08, 1.57775e-08, 1.561715e-08, 
    1.465614e-08, 1.398805e-08, 1.394673e-08, 1.428995e-08, 1.416591e-08,
  1.562082e-08, 1.534383e-08, 1.519559e-08, 1.492443e-08, 1.491832e-08, 
    1.490865e-08, 1.507102e-08, 1.534439e-08, 1.608389e-08, 1.565254e-08, 
    1.444256e-08, 1.37053e-08, 1.395212e-08, 1.425564e-08, 1.405662e-08,
  1.576053e-08, 1.555847e-08, 1.553954e-08, 1.525284e-08, 1.520498e-08, 
    1.517661e-08, 1.537846e-08, 1.576201e-08, 1.607006e-08, 1.558794e-08, 
    1.444995e-08, 1.382148e-08, 1.407792e-08, 1.4243e-08, 1.399011e-08,
  1.600425e-08, 1.584645e-08, 1.585389e-08, 1.558057e-08, 1.542131e-08, 
    1.546758e-08, 1.559148e-08, 1.587832e-08, 1.607145e-08, 1.556683e-08, 
    1.470496e-08, 1.405049e-08, 1.422501e-08, 1.422769e-08, 1.388608e-08,
  1.62952e-08, 1.61027e-08, 1.615507e-08, 1.58568e-08, 1.56716e-08, 
    1.575974e-08, 1.584893e-08, 1.613915e-08, 1.610325e-08, 1.570139e-08, 
    1.510125e-08, 1.451418e-08, 1.435381e-08, 1.41865e-08, 1.378248e-08,
  1.663727e-08, 1.639989e-08, 1.628234e-08, 1.610744e-08, 1.59637e-08, 
    1.615511e-08, 1.616837e-08, 1.631582e-08, 1.629762e-08, 1.594118e-08, 
    1.553263e-08, 1.496288e-08, 1.454721e-08, 1.417074e-08, 1.372867e-08,
  1.691192e-08, 1.656937e-08, 1.639388e-08, 1.629949e-08, 1.62869e-08, 
    1.645985e-08, 1.652775e-08, 1.650384e-08, 1.652785e-08, 1.6173e-08, 
    1.590898e-08, 1.538852e-08, 1.478478e-08, 1.421993e-08, 1.367866e-08,
  1.726941e-08, 1.680989e-08, 1.6522e-08, 1.655491e-08, 1.655449e-08, 
    1.669817e-08, 1.669624e-08, 1.673469e-08, 1.675468e-08, 1.635425e-08, 
    1.603834e-08, 1.565677e-08, 1.504275e-08, 1.43205e-08, 1.3691e-08,
  1.765573e-08, 1.701709e-08, 1.66698e-08, 1.67078e-08, 1.681781e-08, 
    1.697505e-08, 1.689707e-08, 1.698482e-08, 1.696572e-08, 1.645498e-08, 
    1.610459e-08, 1.584196e-08, 1.524211e-08, 1.447418e-08, 1.366234e-08,
  1.34264e-08, 1.217523e-08, 1.128086e-08, 1.03641e-08, 9.877256e-09, 
    9.442013e-09, 9.259539e-09, 9.428446e-09, 9.494808e-09, 9.914713e-09, 
    1.007506e-08, 1.049575e-08, 1.124035e-08, 1.18215e-08, 1.272014e-08,
  1.270198e-08, 1.15992e-08, 1.085892e-08, 9.988433e-09, 9.556943e-09, 
    9.277732e-09, 9.334652e-09, 9.668431e-09, 9.772736e-09, 1.01204e-08, 
    1.038641e-08, 1.085011e-08, 1.17425e-08, 1.233901e-08, 1.332312e-08,
  1.213537e-08, 1.106334e-08, 1.034904e-08, 9.629176e-09, 9.350103e-09, 
    9.273479e-09, 9.484443e-09, 9.867626e-09, 1.006617e-08, 1.04801e-08, 
    1.083198e-08, 1.133418e-08, 1.234017e-08, 1.289664e-08, 1.394385e-08,
  1.16148e-08, 1.059377e-08, 1.000656e-08, 9.431784e-09, 9.272886e-09, 
    9.353212e-09, 9.570939e-09, 1.008564e-08, 1.044818e-08, 1.088407e-08, 
    1.148845e-08, 1.215566e-08, 1.31947e-08, 1.358935e-08, 1.459639e-08,
  1.129768e-08, 1.033755e-08, 9.818198e-09, 9.388611e-09, 9.344954e-09, 
    9.430384e-09, 9.73743e-09, 1.049816e-08, 1.094014e-08, 1.143344e-08, 
    1.23976e-08, 1.306748e-08, 1.423173e-08, 1.427508e-08, 1.460537e-08,
  1.107675e-08, 1.016801e-08, 9.852292e-09, 9.630202e-09, 9.547549e-09, 
    9.796786e-09, 1.020925e-08, 1.09594e-08, 1.155424e-08, 1.229659e-08, 
    1.348077e-08, 1.402828e-08, 1.491451e-08, 1.440894e-08, 1.444597e-08,
  1.085655e-08, 1.017664e-08, 1.010775e-08, 9.849439e-09, 1.005329e-08, 
    1.04002e-08, 1.083963e-08, 1.165865e-08, 1.245123e-08, 1.315204e-08, 
    1.462236e-08, 1.489144e-08, 1.517513e-08, 1.455665e-08, 1.434745e-08,
  1.089928e-08, 1.05657e-08, 1.057255e-08, 1.0515e-08, 1.071158e-08, 
    1.10622e-08, 1.149227e-08, 1.217985e-08, 1.30657e-08, 1.398273e-08, 
    1.499498e-08, 1.56875e-08, 1.529361e-08, 1.46195e-08, 1.434822e-08,
  1.124497e-08, 1.106117e-08, 1.110877e-08, 1.113493e-08, 1.120046e-08, 
    1.148877e-08, 1.193945e-08, 1.27065e-08, 1.344603e-08, 1.411586e-08, 
    1.539665e-08, 1.61799e-08, 1.568009e-08, 1.476413e-08, 1.424254e-08,
  1.152573e-08, 1.153574e-08, 1.161199e-08, 1.147919e-08, 1.165539e-08, 
    1.191005e-08, 1.250207e-08, 1.308403e-08, 1.350093e-08, 1.422072e-08, 
    1.600434e-08, 1.681669e-08, 1.614541e-08, 1.492539e-08, 1.41464e-08,
  2.506566e-08, 2.425951e-08, 2.180427e-08, 1.942771e-08, 1.703858e-08, 
    1.489489e-08, 1.290241e-08, 1.224533e-08, 1.135099e-08, 1.080441e-08, 
    1.022957e-08, 9.587319e-09, 8.938853e-09, 8.560141e-09, 8.396083e-09,
  2.416345e-08, 2.249847e-08, 2.054143e-08, 1.802247e-08, 1.562734e-08, 
    1.353623e-08, 1.217454e-08, 1.14755e-08, 1.047241e-08, 9.773262e-09, 
    9.324615e-09, 9.192717e-09, 8.923895e-09, 8.602797e-09, 8.390337e-09,
  2.393114e-08, 2.160004e-08, 1.957354e-08, 1.706359e-08, 1.465984e-08, 
    1.271917e-08, 1.158632e-08, 1.083233e-08, 9.860175e-09, 9.428958e-09, 
    9.271941e-09, 9.182514e-09, 8.939428e-09, 8.560931e-09, 8.192925e-09,
  2.247434e-08, 2.044009e-08, 1.831704e-08, 1.584366e-08, 1.355775e-08, 
    1.189248e-08, 1.101432e-08, 1.036016e-08, 9.778556e-09, 9.402153e-09, 
    9.21093e-09, 9.078807e-09, 8.822101e-09, 8.466919e-09, 8.312624e-09,
  2.026087e-08, 1.904272e-08, 1.636703e-08, 1.42526e-08, 1.262724e-08, 
    1.165778e-08, 1.095686e-08, 1.029756e-08, 9.718294e-09, 9.279544e-09, 
    9.083768e-09, 8.944046e-09, 8.679177e-09, 8.620213e-09, 8.821202e-09,
  1.837134e-08, 1.699294e-08, 1.44176e-08, 1.346471e-08, 1.225223e-08, 
    1.145507e-08, 1.069214e-08, 1.008175e-08, 9.559948e-09, 9.203857e-09, 
    9.046164e-09, 8.915553e-09, 8.943144e-09, 9.079731e-09, 9.417639e-09,
  1.663317e-08, 1.522579e-08, 1.336773e-08, 1.271949e-08, 1.150619e-08, 
    1.091181e-08, 1.023059e-08, 9.856383e-09, 9.471059e-09, 9.135305e-09, 
    9.156299e-09, 9.201734e-09, 9.330742e-09, 9.593575e-09, 1.003324e-08,
  1.550229e-08, 1.380959e-08, 1.25802e-08, 1.187054e-08, 1.074174e-08, 
    1.030928e-08, 9.814098e-09, 9.683203e-09, 9.295283e-09, 9.236365e-09, 
    9.582847e-09, 9.717469e-09, 9.804844e-09, 1.006252e-08, 1.054407e-08,
  1.420182e-08, 1.283441e-08, 1.192384e-08, 1.089398e-08, 1.015052e-08, 
    9.884866e-09, 9.670461e-09, 9.474053e-09, 9.455441e-09, 9.559589e-09, 
    1.003591e-08, 1.027623e-08, 1.021468e-08, 1.041788e-08, 1.100231e-08,
  1.294353e-08, 1.173108e-08, 1.096656e-08, 1.009896e-08, 9.699741e-09, 
    9.589638e-09, 9.260615e-09, 9.663445e-09, 9.897467e-09, 1.015743e-08, 
    1.058628e-08, 1.060805e-08, 1.053312e-08, 1.085322e-08, 1.145848e-08,
  2.926051e-08, 2.876636e-08, 2.805016e-08, 2.696052e-08, 2.516993e-08, 
    2.34518e-08, 2.161299e-08, 2.009496e-08, 1.865619e-08, 1.804662e-08, 
    1.709242e-08, 1.574219e-08, 1.460061e-08, 1.397542e-08, 1.304848e-08,
  2.952177e-08, 2.940232e-08, 2.828211e-08, 2.702099e-08, 2.484466e-08, 
    2.303402e-08, 2.120348e-08, 1.983037e-08, 1.865318e-08, 1.783045e-08, 
    1.692028e-08, 1.567044e-08, 1.452339e-08, 1.360357e-08, 1.275652e-08,
  2.99908e-08, 2.966445e-08, 2.858306e-08, 2.689793e-08, 2.448164e-08, 
    2.276936e-08, 2.089646e-08, 1.963427e-08, 1.833562e-08, 1.741986e-08, 
    1.664018e-08, 1.541583e-08, 1.40832e-08, 1.311368e-08, 1.234972e-08,
  3.03495e-08, 2.97002e-08, 2.83166e-08, 2.633941e-08, 2.435748e-08, 
    2.257213e-08, 2.065927e-08, 1.93408e-08, 1.793804e-08, 1.692888e-08, 
    1.602877e-08, 1.488903e-08, 1.362007e-08, 1.257766e-08, 1.181017e-08,
  3.016092e-08, 2.892965e-08, 2.713711e-08, 2.587587e-08, 2.368593e-08, 
    2.196312e-08, 2.005012e-08, 1.862646e-08, 1.707418e-08, 1.601339e-08, 
    1.493653e-08, 1.36303e-08, 1.235731e-08, 1.176173e-08, 1.139502e-08,
  2.87203e-08, 2.734816e-08, 2.575081e-08, 2.436572e-08, 2.244255e-08, 
    2.105595e-08, 1.939923e-08, 1.79945e-08, 1.637611e-08, 1.522714e-08, 
    1.41111e-08, 1.311762e-08, 1.230234e-08, 1.176542e-08, 1.134314e-08,
  2.653631e-08, 2.602713e-08, 2.385962e-08, 2.322689e-08, 2.136581e-08, 
    2.035041e-08, 1.87534e-08, 1.740812e-08, 1.591245e-08, 1.498431e-08, 
    1.395496e-08, 1.306713e-08, 1.230619e-08, 1.183428e-08, 1.144736e-08,
  2.477214e-08, 2.39171e-08, 2.243657e-08, 2.215892e-08, 2.027237e-08, 
    1.955149e-08, 1.786531e-08, 1.670172e-08, 1.541232e-08, 1.461995e-08, 
    1.369374e-08, 1.290616e-08, 1.229492e-08, 1.191056e-08, 1.159734e-08,
  2.212703e-08, 2.179411e-08, 2.055216e-08, 2.02426e-08, 1.875426e-08, 
    1.809331e-08, 1.652197e-08, 1.56838e-08, 1.459898e-08, 1.405242e-08, 
    1.32366e-08, 1.272488e-08, 1.232745e-08, 1.202401e-08, 1.170866e-08,
  1.934008e-08, 1.887899e-08, 1.789873e-08, 1.76668e-08, 1.676704e-08, 
    1.646057e-08, 1.530152e-08, 1.485186e-08, 1.408638e-08, 1.365686e-08, 
    1.299285e-08, 1.258929e-08, 1.217966e-08, 1.19388e-08, 1.182853e-08,
  3.446413e-08, 3.379773e-08, 3.259408e-08, 3.16971e-08, 3.087552e-08, 
    2.960526e-08, 2.806137e-08, 2.615471e-08, 2.35626e-08, 2.24751e-08, 
    2.237899e-08, 2.262602e-08, 2.243842e-08, 2.227067e-08, 2.126716e-08,
  3.491489e-08, 3.467339e-08, 3.328268e-08, 3.150311e-08, 3.138906e-08, 
    2.894016e-08, 2.692721e-08, 2.476585e-08, 2.247528e-08, 2.151371e-08, 
    2.152501e-08, 2.162962e-08, 2.19265e-08, 2.206824e-08, 2.121809e-08,
  3.45457e-08, 3.442964e-08, 3.352344e-08, 3.163273e-08, 3.088221e-08, 
    3.052126e-08, 2.721561e-08, 2.505123e-08, 2.275363e-08, 2.156113e-08, 
    2.11883e-08, 2.115676e-08, 2.116228e-08, 2.139967e-08, 2.048277e-08,
  3.440265e-08, 3.445209e-08, 3.362814e-08, 3.208508e-08, 3.080691e-08, 
    2.995277e-08, 2.74695e-08, 2.470687e-08, 2.234991e-08, 2.140499e-08, 
    2.102036e-08, 2.07123e-08, 2.067086e-08, 2.085461e-08, 1.955552e-08,
  3.434488e-08, 3.433175e-08, 3.315196e-08, 3.219175e-08, 3.08634e-08, 
    2.967042e-08, 2.716871e-08, 2.473146e-08, 2.263291e-08, 2.158551e-08, 
    2.120812e-08, 2.071098e-08, 2.036152e-08, 2.016006e-08, 1.912788e-08,
  3.447316e-08, 3.405892e-08, 3.312085e-08, 3.240634e-08, 3.100891e-08, 
    2.952897e-08, 2.710497e-08, 2.504628e-08, 2.293564e-08, 2.192434e-08, 
    2.126762e-08, 2.057215e-08, 1.998913e-08, 1.971159e-08, 1.860306e-08,
  3.404121e-08, 3.383565e-08, 3.28908e-08, 3.23055e-08, 3.12236e-08, 
    2.987917e-08, 2.733903e-08, 2.533828e-08, 2.344996e-08, 2.238593e-08, 
    2.145001e-08, 2.056019e-08, 1.983732e-08, 1.929659e-08, 1.793519e-08,
  3.272205e-08, 3.286307e-08, 3.227304e-08, 3.259061e-08, 3.152299e-08, 
    2.96343e-08, 2.741414e-08, 2.588545e-08, 2.402405e-08, 2.296697e-08, 
    2.177524e-08, 2.072885e-08, 1.967828e-08, 1.888565e-08, 1.746405e-08,
  3.142606e-08, 3.197978e-08, 3.178684e-08, 3.179378e-08, 2.992468e-08, 
    2.888167e-08, 2.710745e-08, 2.593038e-08, 2.399691e-08, 2.296235e-08, 
    2.171818e-08, 2.063553e-08, 1.950963e-08, 1.849351e-08, 1.709386e-08,
  2.934052e-08, 2.956655e-08, 2.92287e-08, 2.919353e-08, 2.812853e-08, 
    2.75462e-08, 2.601005e-08, 2.515782e-08, 2.340002e-08, 2.254172e-08, 
    2.130562e-08, 2.020277e-08, 1.898056e-08, 1.811565e-08, 1.685249e-08,
  3.171683e-08, 3.26702e-08, 3.24733e-08, 3.143067e-08, 2.978433e-08, 
    2.807121e-08, 2.676066e-08, 2.586733e-08, 2.52297e-08, 2.396983e-08, 
    2.246131e-08, 2.058911e-08, 1.824699e-08, 1.638595e-08, 1.486977e-08,
  3.197774e-08, 3.365333e-08, 3.349638e-08, 3.24259e-08, 3.071477e-08, 
    2.876065e-08, 2.654349e-08, 2.482302e-08, 2.313577e-08, 2.208529e-08, 
    2.122988e-08, 2.053426e-08, 1.97178e-08, 1.837889e-08, 1.662868e-08,
  3.133849e-08, 3.234954e-08, 3.219802e-08, 3.163142e-08, 3.043329e-08, 
    2.899564e-08, 2.732928e-08, 2.575409e-08, 2.432446e-08, 2.324797e-08, 
    2.1933e-08, 2.058079e-08, 1.988382e-08, 1.968451e-08, 1.87745e-08,
  3.296008e-08, 3.398633e-08, 3.469716e-08, 3.446951e-08, 3.322556e-08, 
    3.197737e-08, 3.008299e-08, 2.815931e-08, 2.629416e-08, 2.492662e-08, 
    2.348361e-08, 2.241853e-08, 2.106208e-08, 1.93427e-08, 1.880468e-08,
  3.426449e-08, 3.520691e-08, 3.563416e-08, 3.53402e-08, 3.397111e-08, 
    3.301471e-08, 3.188768e-08, 3.057322e-08, 2.873856e-08, 2.654907e-08, 
    2.516827e-08, 2.363105e-08, 2.213066e-08, 2.071521e-08, 1.954767e-08,
  3.341268e-08, 3.432838e-08, 3.546832e-08, 3.61811e-08, 3.612595e-08, 
    3.587033e-08, 3.527947e-08, 3.375466e-08, 3.182111e-08, 3.039739e-08, 
    2.846158e-08, 2.66941e-08, 2.487244e-08, 2.240644e-08, 2.052899e-08,
  3.247255e-08, 3.471292e-08, 3.632503e-08, 3.73632e-08, 3.827273e-08, 
    3.898331e-08, 3.850351e-08, 3.74338e-08, 3.521724e-08, 3.272752e-08, 
    3.138621e-08, 2.914577e-08, 2.643954e-08, 2.467371e-08, 2.291086e-08,
  3.227941e-08, 3.33377e-08, 3.362852e-08, 3.431639e-08, 3.540237e-08, 
    3.601606e-08, 3.720086e-08, 3.731187e-08, 3.657962e-08, 3.475373e-08, 
    3.261487e-08, 3.112472e-08, 2.910227e-08, 2.624647e-08, 2.411827e-08,
  3.06554e-08, 3.014369e-08, 3.10481e-08, 3.100924e-08, 3.192723e-08, 
    3.238361e-08, 3.357881e-08, 3.415145e-08, 3.464145e-08, 3.432716e-08, 
    3.350175e-08, 3.196774e-08, 2.985816e-08, 2.827794e-08, 2.529177e-08,
  2.835493e-08, 2.831696e-08, 2.908792e-08, 2.934712e-08, 3.026591e-08, 
    3.06445e-08, 3.148644e-08, 3.238736e-08, 3.319842e-08, 3.337618e-08, 
    3.262848e-08, 3.108149e-08, 2.952634e-08, 2.754571e-08, 2.622478e-08,
  1.244271e-08, 1.282215e-08, 1.325035e-08, 1.358223e-08, 1.374687e-08, 
    1.362475e-08, 1.356145e-08, 1.341874e-08, 1.329026e-08, 1.316773e-08, 
    1.331287e-08, 1.338282e-08, 1.380248e-08, 1.345178e-08, 1.332236e-08,
  1.464515e-08, 1.481238e-08, 1.51086e-08, 1.540686e-08, 1.598628e-08, 
    1.631059e-08, 1.618906e-08, 1.586156e-08, 1.525086e-08, 1.456303e-08, 
    1.396962e-08, 1.364247e-08, 1.353131e-08, 1.308888e-08, 1.249791e-08,
  1.68056e-08, 1.736666e-08, 1.780634e-08, 1.827535e-08, 1.86181e-08, 
    1.890356e-08, 1.856516e-08, 1.793749e-08, 1.660152e-08, 1.519191e-08, 
    1.413085e-08, 1.347953e-08, 1.322535e-08, 1.33102e-08, 1.264488e-08,
  1.761883e-08, 1.865305e-08, 1.935685e-08, 2.013734e-08, 2.039591e-08, 
    2.063413e-08, 2.045102e-08, 1.980582e-08, 1.858327e-08, 1.667565e-08, 
    1.544716e-08, 1.440744e-08, 1.379436e-08, 1.369176e-08, 1.372584e-08,
  1.826155e-08, 1.911024e-08, 1.996097e-08, 2.091956e-08, 2.158084e-08, 
    2.226154e-08, 2.213895e-08, 2.14825e-08, 2.059173e-08, 1.951057e-08, 
    1.768215e-08, 1.614391e-08, 1.512145e-08, 1.439348e-08, 1.425859e-08,
  2.142381e-08, 2.184166e-08, 2.207282e-08, 2.283717e-08, 2.319311e-08, 
    2.398492e-08, 2.459537e-08, 2.47826e-08, 2.432544e-08, 2.304907e-08, 
    2.143178e-08, 1.900325e-08, 1.716564e-08, 1.588747e-08, 1.543706e-08,
  2.285459e-08, 2.278647e-08, 2.258094e-08, 2.324583e-08, 2.435821e-08, 
    2.608705e-08, 2.788453e-08, 2.965544e-08, 3.009075e-08, 2.918147e-08, 
    2.683783e-08, 2.435825e-08, 2.166042e-08, 1.881205e-08, 1.698001e-08,
  2.152725e-08, 2.229096e-08, 2.397743e-08, 2.665124e-08, 2.987311e-08, 
    3.330996e-08, 3.567924e-08, 3.823921e-08, 3.890428e-08, 3.798826e-08, 
    3.605066e-08, 3.243766e-08, 2.767528e-08, 2.457886e-08, 2.130803e-08,
  2.281698e-08, 2.497475e-08, 2.814601e-08, 3.018167e-08, 3.321154e-08, 
    3.501034e-08, 3.819015e-08, 3.955203e-08, 4.250661e-08, 4.239705e-08, 
    4.142388e-08, 3.836036e-08, 3.466296e-08, 2.871221e-08, 2.490429e-08,
  2.388211e-08, 2.709689e-08, 2.878332e-08, 2.983467e-08, 3.087468e-08, 
    3.244693e-08, 3.485752e-08, 3.527369e-08, 3.716366e-08, 3.808588e-08, 
    3.844344e-08, 3.758234e-08, 3.681816e-08, 3.561928e-08, 2.935982e-08,
  1.209348e-08, 1.072382e-08, 9.604904e-09, 8.952254e-09, 8.473112e-09, 
    8.172462e-09, 8.142377e-09, 8.06163e-09, 8.266619e-09, 8.65139e-09, 
    9.610107e-09, 1.052219e-08, 1.114964e-08, 1.083072e-08, 1.055686e-08,
  1.195859e-08, 1.083289e-08, 9.760702e-09, 9.038739e-09, 8.639994e-09, 
    8.420441e-09, 8.394659e-09, 8.305878e-09, 8.415261e-09, 8.65266e-09, 
    9.326459e-09, 1.010684e-08, 1.096063e-08, 1.106266e-08, 1.054499e-08,
  1.210596e-08, 1.10998e-08, 1.001668e-08, 9.248287e-09, 8.899532e-09, 
    8.796871e-09, 8.730233e-09, 8.501401e-09, 8.381851e-09, 8.491002e-09, 
    8.990996e-09, 9.535653e-09, 1.035027e-08, 1.091247e-08, 1.06894e-08,
  1.226278e-08, 1.167213e-08, 1.070237e-08, 9.69083e-09, 8.934103e-09, 
    8.758117e-09, 8.857819e-09, 8.761601e-09, 8.582773e-09, 8.369105e-09, 
    8.535997e-09, 9.072362e-09, 9.626227e-09, 1.036037e-08, 1.059303e-08,
  1.249041e-08, 1.209466e-08, 1.154739e-08, 1.085675e-08, 1.020204e-08, 
    9.652823e-09, 9.445499e-09, 9.347779e-09, 9.059947e-09, 8.527795e-09, 
    8.319946e-09, 8.404363e-09, 8.875515e-09, 9.190756e-09, 9.936737e-09,
  1.268527e-08, 1.226778e-08, 1.177531e-08, 1.151515e-08, 1.13026e-08, 
    1.129372e-08, 1.112541e-08, 1.098401e-08, 1.083114e-08, 1.014412e-08, 
    9.416952e-09, 8.78259e-09, 8.631806e-09, 8.78069e-09, 8.885806e-09,
  1.265905e-08, 1.246444e-08, 1.244621e-08, 1.260946e-08, 1.275514e-08, 
    1.299271e-08, 1.307685e-08, 1.281861e-08, 1.226829e-08, 1.147497e-08, 
    1.045809e-08, 9.580309e-09, 8.938957e-09, 8.805986e-09, 8.719369e-09,
  1.347644e-08, 1.368334e-08, 1.445965e-08, 1.514253e-08, 1.593562e-08, 
    1.698599e-08, 1.730694e-08, 1.717138e-08, 1.604414e-08, 1.474416e-08, 
    1.291938e-08, 1.113216e-08, 9.835039e-09, 9.299783e-09, 8.829819e-09,
  1.472661e-08, 1.482731e-08, 1.593295e-08, 1.797832e-08, 1.995332e-08, 
    2.293991e-08, 2.298824e-08, 2.353019e-08, 2.298155e-08, 2.11911e-08, 
    1.884248e-08, 1.600589e-08, 1.332418e-08, 1.081848e-08, 9.920551e-09,
  1.36702e-08, 1.547025e-08, 1.798287e-08, 2.240051e-08, 2.659773e-08, 
    2.71947e-08, 2.855408e-08, 2.869155e-08, 2.83681e-08, 2.622616e-08, 
    2.413655e-08, 2.156109e-08, 1.854451e-08, 1.500902e-08, 1.161458e-08,
  2.383313e-08, 2.185447e-08, 1.987362e-08, 1.762681e-08, 1.624582e-08, 
    1.470767e-08, 1.331263e-08, 1.174276e-08, 1.021708e-08, 9.14318e-09, 
    8.688119e-09, 8.865594e-09, 9.479627e-09, 9.862665e-09, 9.752323e-09,
  2.454325e-08, 2.232755e-08, 2.053333e-08, 1.838377e-08, 1.647912e-08, 
    1.495549e-08, 1.346946e-08, 1.183292e-08, 1.023802e-08, 9.078345e-09, 
    8.489005e-09, 8.827061e-09, 9.65931e-09, 1.01648e-08, 1.003263e-08,
  2.498094e-08, 2.265155e-08, 2.103156e-08, 1.92185e-08, 1.692659e-08, 
    1.513018e-08, 1.362313e-08, 1.196285e-08, 1.026529e-08, 9.016262e-09, 
    8.311795e-09, 8.615999e-09, 9.729805e-09, 1.042248e-08, 1.033641e-08,
  2.47617e-08, 2.261171e-08, 2.109548e-08, 1.942582e-08, 1.723656e-08, 
    1.539198e-08, 1.375411e-08, 1.206183e-08, 1.035156e-08, 8.982107e-09, 
    8.179943e-09, 8.364125e-09, 9.609695e-09, 1.060823e-08, 1.062507e-08,
  2.403837e-08, 2.239328e-08, 2.098851e-08, 1.960973e-08, 1.759916e-08, 
    1.565449e-08, 1.399341e-08, 1.223735e-08, 1.049696e-08, 8.951893e-09, 
    8.05115e-09, 8.113619e-09, 9.433404e-09, 1.06655e-08, 1.086057e-08,
  2.260579e-08, 2.15171e-08, 2.021275e-08, 1.921219e-08, 1.758372e-08, 
    1.569032e-08, 1.400702e-08, 1.231344e-08, 1.064541e-08, 8.988359e-09, 
    7.962687e-09, 7.885317e-09, 9.223114e-09, 1.056001e-08, 1.09636e-08,
  2.109706e-08, 2.053383e-08, 1.956988e-08, 1.877697e-08, 1.745157e-08, 
    1.58928e-08, 1.432407e-08, 1.256398e-08, 1.091495e-08, 9.170659e-09, 
    8.004576e-09, 7.757604e-09, 9.034765e-09, 1.043501e-08, 1.097737e-08,
  1.976552e-08, 1.955624e-08, 1.881379e-08, 1.831855e-08, 1.715396e-08, 
    1.576659e-08, 1.438767e-08, 1.275836e-08, 1.11555e-08, 9.356036e-09, 
    8.155125e-09, 7.75058e-09, 8.907501e-09, 1.028659e-08, 1.089776e-08,
  1.92527e-08, 1.912082e-08, 1.854378e-08, 1.80912e-08, 1.729719e-08, 
    1.61913e-08, 1.502827e-08, 1.328474e-08, 1.152194e-08, 9.519887e-09, 
    8.227034e-09, 7.756504e-09, 8.737966e-09, 1.014159e-08, 1.081219e-08,
  1.850596e-08, 1.8248e-08, 1.783576e-08, 1.742843e-08, 1.681297e-08, 
    1.612578e-08, 1.542916e-08, 1.396141e-08, 1.206473e-08, 9.933228e-09, 
    8.524469e-09, 7.927677e-09, 8.67638e-09, 9.902873e-09, 1.071055e-08,
  3.23126e-08, 3.199415e-08, 3.036475e-08, 2.748085e-08, 2.413788e-08, 
    2.046664e-08, 1.783659e-08, 1.623537e-08, 1.502251e-08, 1.313332e-08, 
    1.150689e-08, 1.06368e-08, 1.001372e-08, 9.3053e-09, 8.647803e-09,
  3.367046e-08, 3.270357e-08, 3.134449e-08, 2.928578e-08, 2.571296e-08, 
    2.159403e-08, 1.842924e-08, 1.650948e-08, 1.528029e-08, 1.348999e-08, 
    1.177263e-08, 1.068088e-08, 9.945005e-09, 9.253582e-09, 8.668692e-09,
  3.447876e-08, 3.342574e-08, 3.223016e-08, 3.085681e-08, 2.754787e-08, 
    2.282121e-08, 1.911741e-08, 1.694685e-08, 1.553934e-08, 1.377982e-08, 
    1.198827e-08, 1.072096e-08, 9.865962e-09, 9.176479e-09, 8.655504e-09,
  3.445284e-08, 3.337803e-08, 3.25902e-08, 3.19597e-08, 2.940368e-08, 
    2.424079e-08, 1.999888e-08, 1.737458e-08, 1.571205e-08, 1.400897e-08, 
    1.220977e-08, 1.076933e-08, 9.783344e-09, 9.085094e-09, 8.636203e-09,
  3.401619e-08, 3.295657e-08, 3.262818e-08, 3.286219e-08, 3.100456e-08, 
    2.574616e-08, 2.100556e-08, 1.783168e-08, 1.588334e-08, 1.412058e-08, 
    1.234069e-08, 1.080128e-08, 9.712757e-09, 8.976802e-09, 8.602229e-09,
  3.337991e-08, 3.279034e-08, 3.218346e-08, 3.318435e-08, 3.175334e-08, 
    2.708544e-08, 2.211109e-08, 1.836209e-08, 1.601722e-08, 1.419392e-08, 
    1.243175e-08, 1.080499e-08, 9.612249e-09, 8.855594e-09, 8.553625e-09,
  3.283707e-08, 3.283793e-08, 3.178462e-08, 3.345139e-08, 3.216043e-08, 
    2.822919e-08, 2.310644e-08, 1.887209e-08, 1.609294e-08, 1.415745e-08, 
    1.240936e-08, 1.07699e-08, 9.514062e-09, 8.735356e-09, 8.489909e-09,
  3.20022e-08, 3.223253e-08, 3.113808e-08, 3.330319e-08, 3.274588e-08, 
    2.879371e-08, 2.371512e-08, 1.920417e-08, 1.612456e-08, 1.412429e-08, 
    1.234475e-08, 1.068145e-08, 9.383097e-09, 8.606948e-09, 8.424087e-09,
  3.114983e-08, 3.158037e-08, 3.04719e-08, 3.269382e-08, 3.226893e-08, 
    2.8605e-08, 2.385713e-08, 1.927899e-08, 1.603516e-08, 1.398353e-08, 
    1.219566e-08, 1.053343e-08, 9.250616e-09, 8.488784e-09, 8.354403e-09,
  2.998977e-08, 3.04511e-08, 2.967939e-08, 3.183264e-08, 3.145885e-08, 
    2.780201e-08, 2.347691e-08, 1.91934e-08, 1.594483e-08, 1.383486e-08, 
    1.195808e-08, 1.033323e-08, 9.096624e-09, 8.377305e-09, 8.297039e-09,
  2.431276e-08, 2.131886e-08, 1.825345e-08, 1.639248e-08, 1.549314e-08, 
    1.527145e-08, 1.614333e-08, 1.752633e-08, 1.837006e-08, 1.862935e-08, 
    1.692356e-08, 1.403906e-08, 1.219009e-08, 1.156643e-08, 1.137633e-08,
  2.760828e-08, 2.33405e-08, 1.966084e-08, 1.690237e-08, 1.578745e-08, 
    1.538612e-08, 1.592945e-08, 1.72241e-08, 1.818044e-08, 1.900275e-08, 
    1.752931e-08, 1.469481e-08, 1.246751e-08, 1.172529e-08, 1.15504e-08,
  3.034751e-08, 2.584962e-08, 2.181955e-08, 1.817984e-08, 1.610224e-08, 
    1.546316e-08, 1.579175e-08, 1.687271e-08, 1.766784e-08, 1.921961e-08, 
    1.8081e-08, 1.536591e-08, 1.276408e-08, 1.178768e-08, 1.164582e-08,
  3.190633e-08, 2.835966e-08, 2.396824e-08, 1.994013e-08, 1.690059e-08, 
    1.549625e-08, 1.571143e-08, 1.660881e-08, 1.733776e-08, 1.907229e-08, 
    1.865884e-08, 1.600242e-08, 1.31016e-08, 1.184408e-08, 1.162791e-08,
  3.292601e-08, 3.078627e-08, 2.598432e-08, 2.192252e-08, 1.821023e-08, 
    1.58162e-08, 1.556873e-08, 1.645725e-08, 1.700406e-08, 1.87841e-08, 
    1.907319e-08, 1.663348e-08, 1.347955e-08, 1.189861e-08, 1.155736e-08,
  3.339045e-08, 3.212014e-08, 2.795083e-08, 2.386678e-08, 1.98907e-08, 
    1.659992e-08, 1.543058e-08, 1.625492e-08, 1.675961e-08, 1.832784e-08, 
    1.938122e-08, 1.716257e-08, 1.389397e-08, 1.201004e-08, 1.149542e-08,
  3.381523e-08, 3.286466e-08, 2.968229e-08, 2.562749e-08, 2.160628e-08, 
    1.780042e-08, 1.55712e-08, 1.611668e-08, 1.657028e-08, 1.785511e-08, 
    1.965353e-08, 1.767866e-08, 1.427607e-08, 1.2156e-08, 1.145493e-08,
  3.408293e-08, 3.339355e-08, 3.131684e-08, 2.727457e-08, 2.331982e-08, 
    1.910886e-08, 1.597468e-08, 1.600818e-08, 1.647506e-08, 1.739309e-08, 
    1.981438e-08, 1.810991e-08, 1.465101e-08, 1.233282e-08, 1.145483e-08,
  3.449469e-08, 3.356581e-08, 3.262976e-08, 2.880465e-08, 2.495224e-08, 
    2.066523e-08, 1.666178e-08, 1.605485e-08, 1.646996e-08, 1.711391e-08, 
    1.978304e-08, 1.849245e-08, 1.498655e-08, 1.249578e-08, 1.146606e-08,
  3.497438e-08, 3.389066e-08, 3.340398e-08, 3.015384e-08, 2.613707e-08, 
    2.209971e-08, 1.75207e-08, 1.612607e-08, 1.649765e-08, 1.701497e-08, 
    1.965825e-08, 1.879714e-08, 1.52927e-08, 1.266335e-08, 1.149978e-08,
  2.708807e-08, 2.64264e-08, 2.543089e-08, 2.432257e-08, 2.339589e-08, 
    2.205218e-08, 2.030006e-08, 1.803389e-08, 1.577112e-08, 1.434889e-08, 
    1.345744e-08, 1.27851e-08, 1.225443e-08, 1.201537e-08, 1.163952e-08,
  2.682845e-08, 2.671653e-08, 2.575317e-08, 2.452701e-08, 2.340288e-08, 
    2.209885e-08, 2.034238e-08, 1.815795e-08, 1.586023e-08, 1.452087e-08, 
    1.367936e-08, 1.308586e-08, 1.247824e-08, 1.21008e-08, 1.168756e-08,
  2.667822e-08, 2.701682e-08, 2.62153e-08, 2.484228e-08, 2.353155e-08, 
    2.211386e-08, 2.030499e-08, 1.822898e-08, 1.597216e-08, 1.464513e-08, 
    1.386021e-08, 1.335928e-08, 1.277074e-08, 1.228444e-08, 1.175499e-08,
  2.668272e-08, 2.719546e-08, 2.670076e-08, 2.532457e-08, 2.382993e-08, 
    2.216007e-08, 2.025987e-08, 1.824832e-08, 1.604185e-08, 1.475882e-08, 
    1.39771e-08, 1.356733e-08, 1.306522e-08, 1.250377e-08, 1.194283e-08,
  2.656193e-08, 2.725539e-08, 2.727204e-08, 2.587324e-08, 2.415086e-08, 
    2.221e-08, 2.017774e-08, 1.817673e-08, 1.610308e-08, 1.486606e-08, 
    1.41064e-08, 1.372316e-08, 1.332556e-08, 1.277775e-08, 1.217654e-08,
  2.655339e-08, 2.724216e-08, 2.776926e-08, 2.647341e-08, 2.451689e-08, 
    2.230772e-08, 2.00843e-08, 1.807575e-08, 1.610659e-08, 1.496118e-08, 
    1.424983e-08, 1.385706e-08, 1.352848e-08, 1.301698e-08, 1.243478e-08,
  2.644859e-08, 2.739069e-08, 2.821777e-08, 2.704484e-08, 2.486307e-08, 
    2.23918e-08, 1.993596e-08, 1.789769e-08, 1.608736e-08, 1.504511e-08, 
    1.44011e-08, 1.40051e-08, 1.371865e-08, 1.322333e-08, 1.267522e-08,
  2.632186e-08, 2.75269e-08, 2.857439e-08, 2.764918e-08, 2.520575e-08, 
    2.241421e-08, 1.975082e-08, 1.768249e-08, 1.598624e-08, 1.508661e-08, 
    1.454587e-08, 1.413194e-08, 1.386692e-08, 1.338559e-08, 1.287285e-08,
  2.625528e-08, 2.782591e-08, 2.884669e-08, 2.818178e-08, 2.548012e-08, 
    2.235904e-08, 1.948075e-08, 1.739193e-08, 1.586621e-08, 1.508812e-08, 
    1.467066e-08, 1.427351e-08, 1.401234e-08, 1.353084e-08, 1.301663e-08,
  2.634519e-08, 2.816551e-08, 2.901767e-08, 2.871637e-08, 2.575573e-08, 
    2.221763e-08, 1.910216e-08, 1.703861e-08, 1.564237e-08, 1.503909e-08, 
    1.481251e-08, 1.442714e-08, 1.41476e-08, 1.368812e-08, 1.314256e-08,
  2.220008e-08, 2.265989e-08, 2.291332e-08, 2.284092e-08, 2.286319e-08, 
    2.310861e-08, 2.344347e-08, 2.402759e-08, 2.412155e-08, 2.404586e-08, 
    2.321176e-08, 2.253801e-08, 2.193186e-08, 2.145319e-08, 2.123102e-08,
  2.251739e-08, 2.263149e-08, 2.293381e-08, 2.299098e-08, 2.291715e-08, 
    2.319838e-08, 2.361925e-08, 2.422849e-08, 2.440659e-08, 2.419142e-08, 
    2.350014e-08, 2.276933e-08, 2.21215e-08, 2.172616e-08, 2.115909e-08,
  2.287749e-08, 2.289975e-08, 2.301974e-08, 2.305563e-08, 2.300433e-08, 
    2.323092e-08, 2.37516e-08, 2.442136e-08, 2.463224e-08, 2.428226e-08, 
    2.359719e-08, 2.293885e-08, 2.22812e-08, 2.174056e-08, 2.127137e-08,
  2.310753e-08, 2.314634e-08, 2.322901e-08, 2.317923e-08, 2.312178e-08, 
    2.331082e-08, 2.39354e-08, 2.463615e-08, 2.483621e-08, 2.433716e-08, 
    2.353665e-08, 2.283183e-08, 2.217848e-08, 2.171413e-08, 2.123418e-08,
  2.330137e-08, 2.324757e-08, 2.342623e-08, 2.341714e-08, 2.32447e-08, 
    2.338359e-08, 2.410977e-08, 2.486589e-08, 2.492293e-08, 2.429814e-08, 
    2.339872e-08, 2.267435e-08, 2.190018e-08, 2.162825e-08, 2.114342e-08,
  2.363089e-08, 2.35196e-08, 2.366779e-08, 2.362182e-08, 2.336371e-08, 
    2.350355e-08, 2.438279e-08, 2.513926e-08, 2.510349e-08, 2.427445e-08, 
    2.327263e-08, 2.242252e-08, 2.160282e-08, 2.111396e-08, 2.078529e-08,
  2.384431e-08, 2.369993e-08, 2.384819e-08, 2.378636e-08, 2.355864e-08, 
    2.366802e-08, 2.464497e-08, 2.548377e-08, 2.51686e-08, 2.40552e-08, 
    2.272344e-08, 2.18449e-08, 2.107765e-08, 2.050556e-08, 2.024683e-08,
  2.404865e-08, 2.392341e-08, 2.408171e-08, 2.404957e-08, 2.367523e-08, 
    2.371559e-08, 2.493236e-08, 2.562273e-08, 2.501252e-08, 2.360467e-08, 
    2.221143e-08, 2.099236e-08, 2.006744e-08, 1.956977e-08, 1.94504e-08,
  2.417881e-08, 2.401856e-08, 2.435431e-08, 2.431029e-08, 2.379665e-08, 
    2.385447e-08, 2.517958e-08, 2.570373e-08, 2.474543e-08, 2.30059e-08, 
    2.129329e-08, 1.994938e-08, 1.904391e-08, 1.868624e-08, 1.870357e-08,
  2.463441e-08, 2.428645e-08, 2.458298e-08, 2.442872e-08, 2.386304e-08, 
    2.400954e-08, 2.544112e-08, 2.57776e-08, 2.435804e-08, 2.215158e-08, 
    2.018369e-08, 1.873509e-08, 1.780663e-08, 1.760749e-08, 1.770724e-08,
  2.358149e-08, 2.290103e-08, 2.209736e-08, 2.141695e-08, 2.051533e-08, 
    2.016245e-08, 2.011037e-08, 1.928166e-08, 1.799869e-08, 1.722391e-08, 
    1.635936e-08, 1.547412e-08, 1.639609e-08, 1.906839e-08, 1.894729e-08,
  2.341465e-08, 2.310424e-08, 2.248416e-08, 2.188976e-08, 2.091011e-08, 
    2.019473e-08, 2.003968e-08, 1.980312e-08, 1.887213e-08, 1.775835e-08, 
    1.72014e-08, 1.626349e-08, 1.602681e-08, 1.723311e-08, 1.932303e-08,
  2.303899e-08, 2.305854e-08, 2.253296e-08, 2.20852e-08, 2.128118e-08, 
    2.023636e-08, 1.980762e-08, 1.989348e-08, 1.957975e-08, 1.8454e-08, 
    1.783961e-08, 1.722087e-08, 1.639923e-08, 1.690192e-08, 1.833313e-08,
  2.300128e-08, 2.292297e-08, 2.253322e-08, 2.205232e-08, 2.141813e-08, 
    2.043371e-08, 1.947106e-08, 1.931038e-08, 1.963476e-08, 1.921474e-08, 
    1.857075e-08, 1.818505e-08, 1.733547e-08, 1.69095e-08, 1.763348e-08,
  2.338935e-08, 2.295332e-08, 2.252724e-08, 2.199618e-08, 2.146263e-08, 
    2.072065e-08, 1.964474e-08, 1.909365e-08, 1.936414e-08, 1.958277e-08, 
    1.919103e-08, 1.903193e-08, 1.834412e-08, 1.775482e-08, 1.742909e-08,
  2.363273e-08, 2.309114e-08, 2.259097e-08, 2.198683e-08, 2.142161e-08, 
    2.092191e-08, 1.995814e-08, 1.917974e-08, 1.927139e-08, 1.958755e-08, 
    1.960136e-08, 1.954445e-08, 1.920674e-08, 1.886578e-08, 1.814647e-08,
  2.380768e-08, 2.315391e-08, 2.266087e-08, 2.205234e-08, 2.139731e-08, 
    2.106968e-08, 2.045009e-08, 1.958891e-08, 1.944355e-08, 1.979594e-08, 
    1.997059e-08, 2.018006e-08, 2.006644e-08, 1.995788e-08, 1.935043e-08,
  2.395624e-08, 2.332062e-08, 2.26875e-08, 2.199342e-08, 2.13474e-08, 
    2.112177e-08, 2.076834e-08, 2.012416e-08, 1.984906e-08, 2.010907e-08, 
    2.045977e-08, 2.087896e-08, 2.111514e-08, 2.093642e-08, 2.067419e-08,
  2.394812e-08, 2.327692e-08, 2.276399e-08, 2.21924e-08, 2.158024e-08, 
    2.125099e-08, 2.103913e-08, 2.079265e-08, 2.041149e-08, 2.052619e-08, 
    2.091216e-08, 2.133659e-08, 2.190045e-08, 2.171268e-08, 2.170036e-08,
  2.394295e-08, 2.326506e-08, 2.266122e-08, 2.216108e-08, 2.159167e-08, 
    2.13917e-08, 2.128139e-08, 2.113039e-08, 2.116926e-08, 2.132216e-08, 
    2.164508e-08, 2.182658e-08, 2.23859e-08, 2.239212e-08, 2.252591e-08,
  2.131287e-08, 2.070679e-08, 2.029275e-08, 1.964235e-08, 1.896603e-08, 
    1.847957e-08, 1.793117e-08, 1.736722e-08, 1.773232e-08, 1.796287e-08, 
    1.722985e-08, 1.696402e-08, 1.707262e-08, 1.646396e-08, 1.489142e-08,
  2.351582e-08, 2.330886e-08, 2.254065e-08, 2.189148e-08, 2.057323e-08, 
    1.996981e-08, 1.912179e-08, 1.84618e-08, 1.834148e-08, 1.884359e-08, 
    1.806153e-08, 1.716396e-08, 1.703469e-08, 1.692753e-08, 1.56006e-08,
  2.586419e-08, 2.556326e-08, 2.501342e-08, 2.414053e-08, 2.321378e-08, 
    2.199462e-08, 2.10951e-08, 2.003902e-08, 1.931143e-08, 1.939903e-08, 
    1.866057e-08, 1.756722e-08, 1.719276e-08, 1.712986e-08, 1.628618e-08,
  2.783446e-08, 2.776707e-08, 2.748296e-08, 2.612122e-08, 2.482851e-08, 
    2.389523e-08, 2.261514e-08, 2.185946e-08, 2.0994e-08, 2.047402e-08, 
    1.934486e-08, 1.830463e-08, 1.741378e-08, 1.721117e-08, 1.69068e-08,
  2.873395e-08, 2.891742e-08, 2.934692e-08, 2.897405e-08, 2.697163e-08, 
    2.525614e-08, 2.38627e-08, 2.249953e-08, 2.204406e-08, 2.155099e-08, 
    2.036029e-08, 1.881716e-08, 1.786871e-08, 1.7243e-08, 1.728173e-08,
  2.946654e-08, 2.907396e-08, 2.952173e-08, 3.07338e-08, 3.082907e-08, 
    2.857931e-08, 2.587015e-08, 2.360709e-08, 2.220732e-08, 2.181346e-08, 
    2.127781e-08, 1.98181e-08, 1.834493e-08, 1.750563e-08, 1.733513e-08,
  2.853164e-08, 2.820336e-08, 2.798803e-08, 2.819451e-08, 2.958656e-08, 
    3.065032e-08, 2.901045e-08, 2.590545e-08, 2.338253e-08, 2.18647e-08, 
    2.124234e-08, 2.054277e-08, 1.891257e-08, 1.778731e-08, 1.727199e-08,
  2.764437e-08, 2.774201e-08, 2.767765e-08, 2.774852e-08, 2.750474e-08, 
    2.884869e-08, 2.954497e-08, 2.807842e-08, 2.493195e-08, 2.28353e-08, 
    2.117871e-08, 2.056364e-08, 1.923546e-08, 1.81866e-08, 1.734905e-08,
  2.790064e-08, 2.750363e-08, 2.760525e-08, 2.771967e-08, 2.762252e-08, 
    2.71675e-08, 2.829915e-08, 2.853571e-08, 2.641421e-08, 2.417005e-08, 
    2.188744e-08, 2.055411e-08, 1.949784e-08, 1.860209e-08, 1.774827e-08,
  2.732072e-08, 2.725841e-08, 2.720268e-08, 2.731324e-08, 2.735238e-08, 
    2.742359e-08, 2.693e-08, 2.774347e-08, 2.683885e-08, 2.473696e-08, 
    2.280286e-08, 2.089694e-08, 1.969054e-08, 1.897572e-08, 1.816477e-08,
  7.280887e-09, 6.985624e-09, 6.86793e-09, 6.909472e-09, 7.005454e-09, 
    7.27554e-09, 7.414614e-09, 7.781792e-09, 8.114489e-09, 9.364452e-09, 
    1.020702e-08, 1.046333e-08, 1.111874e-08, 1.238158e-08, 1.42085e-08,
  7.77697e-09, 7.657374e-09, 7.498012e-09, 7.397568e-09, 7.401388e-09, 
    7.605004e-09, 7.77079e-09, 8.142341e-09, 8.494101e-09, 9.369737e-09, 
    1.04605e-08, 1.056675e-08, 1.109274e-08, 1.193444e-08, 1.357181e-08,
  8.566132e-09, 8.579101e-09, 8.609256e-09, 8.425105e-09, 8.375476e-09, 
    8.292579e-09, 8.492012e-09, 8.563808e-09, 9.110007e-09, 9.288612e-09, 
    1.066438e-08, 1.095606e-08, 1.116692e-08, 1.177817e-08, 1.321487e-08,
  1.048071e-08, 1.060572e-08, 1.084464e-08, 1.092544e-08, 1.083938e-08, 
    1.067167e-08, 1.049984e-08, 1.014305e-08, 1.032301e-08, 1.00079e-08, 
    1.057975e-08, 1.10377e-08, 1.104933e-08, 1.14987e-08, 1.261789e-08,
  1.305184e-08, 1.319695e-08, 1.35055e-08, 1.372607e-08, 1.384737e-08, 
    1.37158e-08, 1.363019e-08, 1.340598e-08, 1.298088e-08, 1.320385e-08, 
    1.255786e-08, 1.247857e-08, 1.139522e-08, 1.162294e-08, 1.244479e-08,
  1.574816e-08, 1.60739e-08, 1.627498e-08, 1.633246e-08, 1.602697e-08, 
    1.567889e-08, 1.499745e-08, 1.482247e-08, 1.425467e-08, 1.430597e-08, 
    1.386244e-08, 1.377255e-08, 1.226277e-08, 1.180644e-08, 1.220479e-08,
  1.896244e-08, 2.013553e-08, 2.06379e-08, 2.13497e-08, 2.141868e-08, 
    2.085625e-08, 1.990652e-08, 1.842396e-08, 1.737696e-08, 1.639119e-08, 
    1.560925e-08, 1.505039e-08, 1.382612e-08, 1.233792e-08, 1.248393e-08,
  2.208068e-08, 2.323158e-08, 2.397711e-08, 2.414248e-08, 2.467356e-08, 
    2.460659e-08, 2.454398e-08, 2.332523e-08, 2.130278e-08, 1.963638e-08, 
    1.759502e-08, 1.643248e-08, 1.519489e-08, 1.299693e-08, 1.297956e-08,
  2.410516e-08, 2.485008e-08, 2.52248e-08, 2.601916e-08, 2.618876e-08, 
    2.667129e-08, 2.667468e-08, 2.711221e-08, 2.629068e-08, 2.433507e-08, 
    2.140276e-08, 1.831902e-08, 1.664115e-08, 1.370695e-08, 1.345042e-08,
  2.476485e-08, 2.543949e-08, 2.618104e-08, 2.676142e-08, 2.739439e-08, 
    2.754217e-08, 2.810614e-08, 2.820549e-08, 2.860881e-08, 2.833969e-08, 
    2.661694e-08, 2.206458e-08, 1.893985e-08, 1.490353e-08, 1.386635e-08,
  1.67137e-08, 1.618437e-08, 1.564324e-08, 1.497571e-08, 1.417971e-08, 
    1.33568e-08, 1.261743e-08, 1.187322e-08, 1.097494e-08, 1.009678e-08, 
    9.479233e-09, 9.106215e-09, 9.034611e-09, 9.193748e-09, 9.683363e-09,
  1.695499e-08, 1.650663e-08, 1.584181e-08, 1.503591e-08, 1.410749e-08, 
    1.313064e-08, 1.234443e-08, 1.159172e-08, 1.074061e-08, 9.847592e-09, 
    9.072824e-09, 8.645956e-09, 8.532634e-09, 8.674024e-09, 9.059181e-09,
  1.732616e-08, 1.677e-08, 1.61134e-08, 1.52924e-08, 1.430427e-08, 
    1.318773e-08, 1.219425e-08, 1.137429e-08, 1.057097e-08, 9.666423e-09, 
    8.816601e-09, 8.320956e-09, 8.141193e-09, 8.324184e-09, 8.66152e-09,
  1.71526e-08, 1.6662e-08, 1.604e-08, 1.533999e-08, 1.458255e-08, 
    1.364251e-08, 1.254575e-08, 1.150829e-08, 1.058756e-08, 9.717316e-09, 
    8.75771e-09, 8.057039e-09, 7.826971e-09, 7.888691e-09, 8.212342e-09,
  1.672484e-08, 1.628569e-08, 1.579546e-08, 1.525094e-08, 1.458115e-08, 
    1.385621e-08, 1.295015e-08, 1.196601e-08, 1.096868e-08, 1.000773e-08, 
    9.041051e-09, 8.187619e-09, 7.728533e-09, 7.618001e-09, 7.745125e-09,
  1.63182e-08, 1.57938e-08, 1.535995e-08, 1.495459e-08, 1.448822e-08, 
    1.397499e-08, 1.331616e-08, 1.2484e-08, 1.14416e-08, 1.033472e-08, 
    9.262233e-09, 8.306771e-09, 7.662941e-09, 7.384152e-09, 7.415563e-09,
  1.617643e-08, 1.568105e-08, 1.517771e-08, 1.480092e-08, 1.435882e-08, 
    1.397173e-08, 1.363209e-08, 1.312361e-08, 1.246181e-08, 1.145194e-08, 
    1.029642e-08, 8.978366e-09, 7.94858e-09, 7.293556e-09, 7.141971e-09,
  1.635401e-08, 1.58771e-08, 1.550151e-08, 1.509983e-08, 1.479033e-08, 
    1.423796e-08, 1.384587e-08, 1.33114e-08, 1.280177e-08, 1.210186e-08, 
    1.104844e-08, 9.841512e-09, 8.575356e-09, 7.533801e-09, 7.086902e-09,
  1.687913e-08, 1.646796e-08, 1.614432e-08, 1.604093e-08, 1.584572e-08, 
    1.566682e-08, 1.521574e-08, 1.476526e-08, 1.428951e-08, 1.373295e-08, 
    1.287024e-08, 1.149545e-08, 9.693101e-09, 8.273583e-09, 7.350674e-09,
  1.780798e-08, 1.7294e-08, 1.698933e-08, 1.682692e-08, 1.691952e-08, 
    1.672442e-08, 1.681078e-08, 1.63552e-08, 1.609752e-08, 1.547129e-08, 
    1.471532e-08, 1.375564e-08, 1.188842e-08, 9.347765e-09, 7.952431e-09,
  1.912795e-08, 1.894527e-08, 1.889975e-08, 1.896348e-08, 1.875449e-08, 
    1.834775e-08, 1.789392e-08, 1.756258e-08, 1.718243e-08, 1.678579e-08, 
    1.641408e-08, 1.609236e-08, 1.581095e-08, 1.563899e-08, 1.570824e-08,
  1.892931e-08, 1.895301e-08, 1.872442e-08, 1.85476e-08, 1.847636e-08, 
    1.827103e-08, 1.792369e-08, 1.757374e-08, 1.724825e-08, 1.692199e-08, 
    1.667059e-08, 1.621154e-08, 1.575245e-08, 1.54085e-08, 1.542035e-08,
  1.871886e-08, 1.874827e-08, 1.856375e-08, 1.833549e-08, 1.822537e-08, 
    1.824841e-08, 1.817016e-08, 1.805354e-08, 1.778135e-08, 1.735049e-08, 
    1.684797e-08, 1.64026e-08, 1.596877e-08, 1.532964e-08, 1.507991e-08,
  1.878111e-08, 1.860668e-08, 1.840799e-08, 1.819079e-08, 1.802268e-08, 
    1.802481e-08, 1.808178e-08, 1.810879e-08, 1.790152e-08, 1.757937e-08, 
    1.699444e-08, 1.633328e-08, 1.583464e-08, 1.511631e-08, 1.472445e-08,
  1.882948e-08, 1.871412e-08, 1.854076e-08, 1.841544e-08, 1.824449e-08, 
    1.809991e-08, 1.802921e-08, 1.811687e-08, 1.821987e-08, 1.781593e-08, 
    1.721924e-08, 1.637416e-08, 1.561149e-08, 1.483419e-08, 1.433673e-08,
  1.925639e-08, 1.925613e-08, 1.922072e-08, 1.915931e-08, 1.900401e-08, 
    1.876336e-08, 1.844763e-08, 1.816498e-08, 1.804978e-08, 1.79791e-08, 
    1.747055e-08, 1.654482e-08, 1.560481e-08, 1.465591e-08, 1.400933e-08,
  2.017279e-08, 2.027717e-08, 2.02896e-08, 2.032108e-08, 2.021361e-08, 
    1.984578e-08, 1.947009e-08, 1.891388e-08, 1.839103e-08, 1.80957e-08, 
    1.773772e-08, 1.694434e-08, 1.584346e-08, 1.477923e-08, 1.383909e-08,
  2.088274e-08, 2.081954e-08, 2.084566e-08, 2.083878e-08, 2.088141e-08, 
    2.076809e-08, 2.050824e-08, 2.003342e-08, 1.916479e-08, 1.84125e-08, 
    1.790936e-08, 1.725514e-08, 1.62545e-08, 1.504086e-08, 1.386875e-08,
  2.136602e-08, 2.130293e-08, 2.126526e-08, 2.129094e-08, 2.130179e-08, 
    2.136247e-08, 2.121889e-08, 2.110387e-08, 2.058225e-08, 1.9569e-08, 
    1.859194e-08, 1.769052e-08, 1.679759e-08, 1.547338e-08, 1.395281e-08,
  2.184121e-08, 2.211069e-08, 2.214765e-08, 2.214627e-08, 2.211294e-08, 
    2.20713e-08, 2.195423e-08, 2.169693e-08, 2.151425e-08, 2.082034e-08, 
    1.950102e-08, 1.835805e-08, 1.727152e-08, 1.58743e-08, 1.409746e-08,
  2.023284e-08, 2.106599e-08, 2.144864e-08, 2.184564e-08, 2.222672e-08, 
    2.22923e-08, 2.17107e-08, 2.077699e-08, 1.994689e-08, 1.939481e-08, 
    1.929912e-08, 1.932404e-08, 1.950203e-08, 1.962279e-08, 1.955997e-08,
  2.101432e-08, 2.14641e-08, 2.217605e-08, 2.260356e-08, 2.278755e-08, 
    2.23316e-08, 2.125883e-08, 2.011071e-08, 1.919622e-08, 1.891035e-08, 
    1.904707e-08, 1.934744e-08, 1.954318e-08, 1.958591e-08, 1.933275e-08,
  2.249831e-08, 2.245949e-08, 2.254067e-08, 2.276361e-08, 2.257708e-08, 
    2.172826e-08, 2.077488e-08, 1.983533e-08, 1.926445e-08, 1.917379e-08, 
    1.92542e-08, 1.960104e-08, 1.957753e-08, 1.933854e-08, 1.886532e-08,
  2.31661e-08, 2.289587e-08, 2.247356e-08, 2.208501e-08, 2.136932e-08, 
    2.059046e-08, 2.008261e-08, 1.967905e-08, 1.951416e-08, 1.95764e-08, 
    1.975264e-08, 1.961611e-08, 1.928697e-08, 1.905698e-08, 1.852942e-08,
  2.28713e-08, 2.239734e-08, 2.151338e-08, 2.070081e-08, 2.01369e-08, 
    1.978204e-08, 1.970838e-08, 1.965364e-08, 1.96266e-08, 1.970619e-08, 
    1.971281e-08, 1.927359e-08, 1.905635e-08, 1.88495e-08, 1.837006e-08,
  2.206884e-08, 2.147399e-08, 2.079141e-08, 2.007548e-08, 1.956733e-08, 
    1.943466e-08, 1.948299e-08, 1.961022e-08, 1.976754e-08, 1.974431e-08, 
    1.944488e-08, 1.90981e-08, 1.896153e-08, 1.88171e-08, 1.852544e-08,
  2.161214e-08, 2.103499e-08, 2.05288e-08, 2.001788e-08, 1.970071e-08, 
    1.955979e-08, 1.952162e-08, 1.963048e-08, 1.975861e-08, 1.973301e-08, 
    1.93756e-08, 1.902055e-08, 1.871532e-08, 1.84751e-08, 1.839698e-08,
  2.150897e-08, 2.105389e-08, 2.064067e-08, 2.025439e-08, 1.995868e-08, 
    1.964328e-08, 1.956663e-08, 1.966696e-08, 1.978046e-08, 1.970333e-08, 
    1.939672e-08, 1.909626e-08, 1.858469e-08, 1.821446e-08, 1.825498e-08,
  2.11931e-08, 2.090722e-08, 2.062068e-08, 2.027135e-08, 1.995991e-08, 
    1.959583e-08, 1.953047e-08, 1.971413e-08, 1.979075e-08, 1.970817e-08, 
    1.933194e-08, 1.896531e-08, 1.861217e-08, 1.826223e-08, 1.817386e-08,
  2.075702e-08, 2.061569e-08, 2.040369e-08, 2.014015e-08, 1.989028e-08, 
    1.969627e-08, 1.968361e-08, 1.987713e-08, 1.996834e-08, 1.97911e-08, 
    1.954491e-08, 1.897234e-08, 1.864211e-08, 1.848301e-08, 1.824989e-08,
  1.196593e-08, 1.187916e-08, 1.194821e-08, 1.18961e-08, 1.210972e-08, 
    1.270477e-08, 1.399186e-08, 1.559391e-08, 1.73405e-08, 1.894666e-08, 
    2.040709e-08, 2.124287e-08, 2.13935e-08, 2.089856e-08, 2.044959e-08,
  1.210756e-08, 1.196218e-08, 1.207154e-08, 1.225899e-08, 1.26398e-08, 
    1.343598e-08, 1.492791e-08, 1.642783e-08, 1.789681e-08, 1.919385e-08, 
    2.037501e-08, 2.063713e-08, 2.035886e-08, 2.003215e-08, 1.976188e-08,
  1.297708e-08, 1.221826e-08, 1.214592e-08, 1.244313e-08, 1.312295e-08, 
    1.429763e-08, 1.573968e-08, 1.688864e-08, 1.783157e-08, 1.887748e-08, 
    1.965094e-08, 1.945955e-08, 1.955842e-08, 1.991712e-08, 1.990447e-08,
  1.507675e-08, 1.36753e-08, 1.314262e-08, 1.334462e-08, 1.415907e-08, 
    1.522912e-08, 1.616344e-08, 1.67439e-08, 1.754311e-08, 1.888575e-08, 
    1.980007e-08, 1.98568e-08, 2.030846e-08, 2.065278e-08, 2.068988e-08,
  1.698414e-08, 1.629968e-08, 1.558074e-08, 1.535844e-08, 1.560865e-08, 
    1.588374e-08, 1.624757e-08, 1.666572e-08, 1.782952e-08, 1.938227e-08, 
    2.037386e-08, 2.033303e-08, 2.055067e-08, 2.074032e-08, 2.074924e-08,
  1.887091e-08, 1.825017e-08, 1.778801e-08, 1.741373e-08, 1.717239e-08, 
    1.69682e-08, 1.693838e-08, 1.734925e-08, 1.866351e-08, 2.016705e-08, 
    2.101888e-08, 2.044976e-08, 2.062091e-08, 2.075336e-08, 2.086131e-08,
  1.973213e-08, 1.904955e-08, 1.881055e-08, 1.869319e-08, 1.837936e-08, 
    1.797299e-08, 1.784617e-08, 1.83478e-08, 1.950314e-08, 2.092717e-08, 
    2.119075e-08, 2.030989e-08, 2.060846e-08, 2.072802e-08, 2.091626e-08,
  2.227633e-08, 2.049252e-08, 1.917235e-08, 1.886777e-08, 1.905555e-08, 
    1.87524e-08, 1.877464e-08, 1.933586e-08, 2.038417e-08, 2.155323e-08, 
    2.103421e-08, 2.029682e-08, 2.071437e-08, 2.052579e-08, 2.07716e-08,
  2.316371e-08, 2.227225e-08, 2.134296e-08, 1.987405e-08, 1.926166e-08, 
    1.909955e-08, 1.927445e-08, 1.97463e-08, 2.062643e-08, 2.115639e-08, 
    2.023814e-08, 2.005936e-08, 2.055122e-08, 2.022731e-08, 2.04933e-08,
  2.606558e-08, 2.349464e-08, 2.23631e-08, 2.183384e-08, 2.108169e-08, 
    2.037461e-08, 2.010848e-08, 2.035454e-08, 2.074895e-08, 2.078269e-08, 
    2.010546e-08, 2.017111e-08, 2.040766e-08, 2.03232e-08, 2.021753e-08,
  1.55987e-08, 1.282881e-08, 1.051702e-08, 8.26592e-09, 6.590358e-09, 
    5.801077e-09, 5.646023e-09, 5.422764e-09, 5.062934e-09, 4.770754e-09, 
    4.804286e-09, 4.96565e-09, 5.86159e-09, 7.071605e-09, 8.136601e-09,
  1.586509e-08, 1.335875e-08, 1.080079e-08, 8.497741e-09, 6.805175e-09, 
    5.902993e-09, 5.630305e-09, 5.458312e-09, 5.167867e-09, 5.010087e-09, 
    5.118252e-09, 5.677474e-09, 6.873234e-09, 8.397301e-09, 9.611018e-09,
  1.602984e-08, 1.3786e-08, 1.116014e-08, 8.793134e-09, 7.122151e-09, 
    6.139865e-09, 5.882182e-09, 5.670421e-09, 5.473067e-09, 5.357238e-09, 
    5.60316e-09, 6.561921e-09, 7.937502e-09, 9.340834e-09, 1.058226e-08,
  1.650495e-08, 1.437787e-08, 1.16696e-08, 9.051164e-09, 7.40092e-09, 
    6.407034e-09, 6.109112e-09, 5.881219e-09, 5.762396e-09, 5.727804e-09, 
    6.118297e-09, 7.195299e-09, 8.596481e-09, 9.827911e-09, 1.137846e-08,
  1.692515e-08, 1.481939e-08, 1.235754e-08, 9.636142e-09, 7.721516e-09, 
    6.671614e-09, 6.329782e-09, 6.077464e-09, 5.9469e-09, 6.00606e-09, 
    6.47097e-09, 7.590758e-09, 8.787857e-09, 1.027308e-08, 1.232336e-08,
  1.854621e-08, 1.603789e-08, 1.338359e-08, 1.053946e-08, 8.393135e-09, 
    6.982806e-09, 6.464508e-09, 6.259266e-09, 6.162702e-09, 6.224895e-09, 
    6.729433e-09, 7.90669e-09, 9.098414e-09, 1.104394e-08, 1.360303e-08,
  1.976663e-08, 1.723288e-08, 1.452192e-08, 1.190008e-08, 9.605031e-09, 
    7.869112e-09, 7.018546e-09, 6.676464e-09, 6.493153e-09, 6.509812e-09, 
    7.215084e-09, 8.474909e-09, 9.629507e-09, 1.224957e-08, 1.506191e-08,
  2.199113e-08, 1.987189e-08, 1.682926e-08, 1.314138e-08, 1.082879e-08, 
    9.174401e-09, 8.023067e-09, 7.453095e-09, 7.103213e-09, 7.000649e-09, 
    7.73224e-09, 8.839545e-09, 1.0441e-08, 1.377133e-08, 1.642443e-08,
  2.192314e-08, 2.089018e-08, 1.961553e-08, 1.683881e-08, 1.316394e-08, 
    1.035869e-08, 8.874508e-09, 8.341926e-09, 8.083779e-09, 8.169338e-09, 
    9.095256e-09, 9.966574e-09, 1.234442e-08, 1.549745e-08, 1.737753e-08,
  2.316181e-08, 2.094729e-08, 1.961529e-08, 1.844153e-08, 1.677566e-08, 
    1.434496e-08, 1.136013e-08, 9.208224e-09, 8.67156e-09, 8.703463e-09, 
    9.952222e-09, 1.072495e-08, 1.361989e-08, 1.656151e-08, 1.737027e-08,
  1.759966e-08, 1.675786e-08, 1.610576e-08, 1.522453e-08, 1.407749e-08, 
    1.275918e-08, 1.185343e-08, 1.094425e-08, 9.237803e-09, 8.166749e-09, 
    9.093106e-09, 1.06714e-08, 1.151591e-08, 1.259453e-08, 1.330045e-08,
  1.82441e-08, 1.745845e-08, 1.672615e-08, 1.581074e-08, 1.469976e-08, 
    1.32544e-08, 1.213617e-08, 1.118218e-08, 9.288235e-09, 7.798802e-09, 
    8.387365e-09, 9.730052e-09, 1.052694e-08, 1.136051e-08, 1.21374e-08,
  1.902967e-08, 1.810184e-08, 1.733834e-08, 1.638866e-08, 1.524267e-08, 
    1.380474e-08, 1.249767e-08, 1.146048e-08, 9.458761e-09, 7.549846e-09, 
    7.859446e-09, 8.942748e-09, 9.629711e-09, 1.028074e-08, 1.103369e-08,
  1.983797e-08, 1.89918e-08, 1.799722e-08, 1.705178e-08, 1.594271e-08, 
    1.437493e-08, 1.294105e-08, 1.184652e-08, 9.747374e-09, 7.373949e-09, 
    7.30908e-09, 8.135018e-09, 8.827501e-09, 9.292106e-09, 1.003378e-08,
  2.033296e-08, 1.96014e-08, 1.86695e-08, 1.765292e-08, 1.659515e-08, 
    1.500989e-08, 1.342805e-08, 1.22226e-08, 1.008689e-08, 7.399736e-09, 
    6.977841e-09, 7.483779e-09, 8.138724e-09, 8.555888e-09, 9.128675e-09,
  2.08632e-08, 2.025243e-08, 1.934425e-08, 1.825753e-08, 1.720772e-08, 
    1.566775e-08, 1.391087e-08, 1.26671e-08, 1.044469e-08, 7.490229e-09, 
    6.64624e-09, 6.936562e-09, 7.544692e-09, 7.914955e-09, 8.37414e-09,
  2.100355e-08, 2.063268e-08, 1.995639e-08, 1.892787e-08, 1.786764e-08, 
    1.632633e-08, 1.444429e-08, 1.308701e-08, 1.090165e-08, 7.791155e-09, 
    6.522686e-09, 6.566959e-09, 7.040133e-09, 7.332241e-09, 7.705665e-09,
  2.147553e-08, 2.11705e-08, 2.03825e-08, 1.955888e-08, 1.852595e-08, 
    1.708702e-08, 1.502543e-08, 1.349778e-08, 1.129486e-08, 8.103962e-09, 
    6.420112e-09, 6.270183e-09, 6.633366e-09, 6.831212e-09, 7.152393e-09,
  2.193423e-08, 2.157861e-08, 2.102053e-08, 2.006778e-08, 1.910128e-08, 
    1.780638e-08, 1.576639e-08, 1.403227e-08, 1.176873e-08, 8.60228e-09, 
    6.490983e-09, 6.033535e-09, 6.260619e-09, 6.394871e-09, 6.780879e-09,
  2.282177e-08, 2.2327e-08, 2.156814e-08, 2.065429e-08, 1.960555e-08, 
    1.852099e-08, 1.648873e-08, 1.453153e-08, 1.220673e-08, 9.075353e-09, 
    6.609862e-09, 5.900146e-09, 5.941065e-09, 6.146664e-09, 6.735728e-09,
  1.995428e-08, 1.947461e-08, 1.878478e-08, 1.804822e-08, 1.723993e-08, 
    1.597077e-08, 1.450404e-08, 1.386215e-08, 1.341449e-08, 1.258248e-08, 
    1.227054e-08, 1.423466e-08, 1.817444e-08, 2.156938e-08, 2.216717e-08,
  2.095504e-08, 2.031118e-08, 1.941454e-08, 1.851543e-08, 1.758764e-08, 
    1.608923e-08, 1.461369e-08, 1.394294e-08, 1.358274e-08, 1.255858e-08, 
    1.193353e-08, 1.384723e-08, 1.788078e-08, 2.126325e-08, 2.17054e-08,
  2.182819e-08, 2.123044e-08, 2.034932e-08, 1.918251e-08, 1.809547e-08, 
    1.657376e-08, 1.479341e-08, 1.405069e-08, 1.376709e-08, 1.273923e-08, 
    1.177526e-08, 1.342965e-08, 1.743417e-08, 2.093233e-08, 2.126089e-08,
  2.292315e-08, 2.188156e-08, 2.113244e-08, 2.015276e-08, 1.880304e-08, 
    1.730549e-08, 1.533681e-08, 1.419396e-08, 1.381767e-08, 1.292261e-08, 
    1.172462e-08, 1.307594e-08, 1.680005e-08, 2.056169e-08, 2.084916e-08,
  2.36959e-08, 2.284676e-08, 2.171867e-08, 2.09774e-08, 1.974086e-08, 
    1.810522e-08, 1.60186e-08, 1.458882e-08, 1.399939e-08, 1.309837e-08, 
    1.177725e-08, 1.275737e-08, 1.604946e-08, 2.008824e-08, 2.046081e-08,
  2.435264e-08, 2.359643e-08, 2.254297e-08, 2.157107e-08, 2.062938e-08, 
    1.900251e-08, 1.690843e-08, 1.501525e-08, 1.413879e-08, 1.32538e-08, 
    1.185263e-08, 1.24973e-08, 1.530231e-08, 1.952736e-08, 2.007118e-08,
  2.47242e-08, 2.437347e-08, 2.321237e-08, 2.207891e-08, 2.124642e-08, 
    1.977871e-08, 1.761014e-08, 1.579829e-08, 1.457534e-08, 1.338078e-08, 
    1.196067e-08, 1.228748e-08, 1.460215e-08, 1.882819e-08, 1.970013e-08,
  2.453768e-08, 2.47748e-08, 2.431018e-08, 2.278554e-08, 2.163756e-08, 
    2.05841e-08, 1.837026e-08, 1.634723e-08, 1.505929e-08, 1.363187e-08, 
    1.201825e-08, 1.210808e-08, 1.402978e-08, 1.806469e-08, 1.923495e-08,
  2.392924e-08, 2.457721e-08, 2.458295e-08, 2.386963e-08, 2.233791e-08, 
    2.086163e-08, 1.902166e-08, 1.709848e-08, 1.563074e-08, 1.388433e-08, 
    1.210958e-08, 1.197013e-08, 1.358831e-08, 1.722244e-08, 1.873357e-08,
  2.319008e-08, 2.408684e-08, 2.442368e-08, 2.418599e-08, 2.321674e-08, 
    2.133024e-08, 1.924156e-08, 1.740834e-08, 1.600658e-08, 1.426408e-08, 
    1.218146e-08, 1.186569e-08, 1.331007e-08, 1.638374e-08, 1.813441e-08,
  1.876712e-08, 1.849555e-08, 1.80926e-08, 1.734652e-08, 1.714e-08, 
    1.721477e-08, 1.785466e-08, 1.744367e-08, 1.753799e-08, 1.693316e-08, 
    1.657278e-08, 1.562099e-08, 1.471638e-08, 1.455161e-08, 1.552369e-08,
  1.917351e-08, 1.914254e-08, 1.902215e-08, 1.82454e-08, 1.756146e-08, 
    1.711029e-08, 1.747469e-08, 1.753989e-08, 1.798124e-08, 1.701208e-08, 
    1.652669e-08, 1.540319e-08, 1.464397e-08, 1.475463e-08, 1.586345e-08,
  1.931294e-08, 1.983718e-08, 1.973267e-08, 1.917535e-08, 1.83815e-08, 
    1.769005e-08, 1.746061e-08, 1.757843e-08, 1.748714e-08, 1.740946e-08, 
    1.658869e-08, 1.529087e-08, 1.457851e-08, 1.498955e-08, 1.623614e-08,
  1.962651e-08, 2.006644e-08, 2.043133e-08, 2.014114e-08, 1.940112e-08, 
    1.850574e-08, 1.770421e-08, 1.751348e-08, 1.712395e-08, 1.78677e-08, 
    1.690798e-08, 1.538483e-08, 1.457286e-08, 1.522159e-08, 1.670027e-08,
  1.992679e-08, 2.026564e-08, 2.059855e-08, 2.102895e-08, 2.070013e-08, 
    1.98332e-08, 1.841499e-08, 1.760279e-08, 1.692748e-08, 1.744065e-08, 
    1.734496e-08, 1.580515e-08, 1.454692e-08, 1.540533e-08, 1.701324e-08,
  2.053702e-08, 2.057997e-08, 2.064299e-08, 2.106332e-08, 2.137582e-08, 
    2.097051e-08, 1.982773e-08, 1.824262e-08, 1.723815e-08, 1.66796e-08, 
    1.7707e-08, 1.624409e-08, 1.472253e-08, 1.5548e-08, 1.729742e-08,
  2.16546e-08, 2.159462e-08, 2.142061e-08, 2.141783e-08, 2.152894e-08, 
    2.139281e-08, 2.069808e-08, 1.92817e-08, 1.786758e-08, 1.682212e-08, 
    1.739398e-08, 1.679845e-08, 1.503754e-08, 1.56973e-08, 1.755015e-08,
  2.300446e-08, 2.320471e-08, 2.29528e-08, 2.264443e-08, 2.221154e-08, 
    2.192145e-08, 2.133635e-08, 2.02419e-08, 1.857368e-08, 1.74198e-08, 
    1.669449e-08, 1.70359e-08, 1.547094e-08, 1.581623e-08, 1.774263e-08,
  2.349076e-08, 2.414318e-08, 2.426628e-08, 2.382866e-08, 2.314823e-08, 
    2.264914e-08, 2.221058e-08, 2.139691e-08, 1.983561e-08, 1.828498e-08, 
    1.706404e-08, 1.690702e-08, 1.594461e-08, 1.59949e-08, 1.786298e-08,
  2.376007e-08, 2.433492e-08, 2.480519e-08, 2.483423e-08, 2.430222e-08, 
    2.356258e-08, 2.288603e-08, 2.227109e-08, 2.09228e-08, 1.937322e-08, 
    1.800031e-08, 1.663122e-08, 1.62382e-08, 1.633463e-08, 1.797563e-08,
  1.311343e-08, 1.206228e-08, 1.060201e-08, 9.814938e-09, 9.608898e-09, 
    1.00574e-08, 1.089835e-08, 1.204145e-08, 1.335915e-08, 1.406019e-08, 
    1.499795e-08, 1.608481e-08, 1.697169e-08, 1.747652e-08, 1.796818e-08,
  1.338386e-08, 1.267048e-08, 1.173537e-08, 1.087767e-08, 1.063285e-08, 
    1.073993e-08, 1.129342e-08, 1.204114e-08, 1.401996e-08, 1.465401e-08, 
    1.520372e-08, 1.639577e-08, 1.727417e-08, 1.770057e-08, 1.8296e-08,
  1.370518e-08, 1.311325e-08, 1.259994e-08, 1.176937e-08, 1.138499e-08, 
    1.121369e-08, 1.156203e-08, 1.217424e-08, 1.400175e-08, 1.500653e-08, 
    1.522444e-08, 1.639055e-08, 1.727631e-08, 1.776491e-08, 1.886555e-08,
  1.377873e-08, 1.346106e-08, 1.322425e-08, 1.253893e-08, 1.191402e-08, 
    1.160265e-08, 1.169999e-08, 1.238999e-08, 1.368889e-08, 1.558989e-08, 
    1.533451e-08, 1.616301e-08, 1.719317e-08, 1.794541e-08, 1.918059e-08,
  1.418198e-08, 1.350005e-08, 1.350585e-08, 1.309949e-08, 1.234993e-08, 
    1.191155e-08, 1.188037e-08, 1.240038e-08, 1.332648e-08, 1.581228e-08, 
    1.565192e-08, 1.612418e-08, 1.715303e-08, 1.810203e-08, 1.913391e-08,
  1.497595e-08, 1.375698e-08, 1.342994e-08, 1.335616e-08, 1.270428e-08, 
    1.22761e-08, 1.21729e-08, 1.251685e-08, 1.324673e-08, 1.561608e-08, 
    1.622839e-08, 1.602986e-08, 1.710475e-08, 1.802432e-08, 1.907924e-08,
  1.543004e-08, 1.412543e-08, 1.330312e-08, 1.329023e-08, 1.295339e-08, 
    1.269791e-08, 1.254307e-08, 1.27011e-08, 1.327906e-08, 1.507142e-08, 
    1.722531e-08, 1.638452e-08, 1.721282e-08, 1.797974e-08, 1.881497e-08,
  1.572411e-08, 1.450027e-08, 1.343222e-08, 1.315113e-08, 1.3241e-08, 
    1.313192e-08, 1.297184e-08, 1.294674e-08, 1.325183e-08, 1.438878e-08, 
    1.714259e-08, 1.712764e-08, 1.714463e-08, 1.801188e-08, 1.885141e-08,
  1.613811e-08, 1.501365e-08, 1.400724e-08, 1.350952e-08, 1.351864e-08, 
    1.374266e-08, 1.361135e-08, 1.361991e-08, 1.361439e-08, 1.440324e-08, 
    1.688908e-08, 1.812726e-08, 1.731437e-08, 1.792925e-08, 1.874071e-08,
  1.668139e-08, 1.563974e-08, 1.470953e-08, 1.405752e-08, 1.381988e-08, 
    1.400746e-08, 1.39357e-08, 1.399665e-08, 1.407162e-08, 1.473602e-08, 
    1.683405e-08, 1.841495e-08, 1.774006e-08, 1.789987e-08, 1.866719e-08,
  9.443408e-09, 8.777959e-09, 8.081415e-09, 7.34317e-09, 6.590207e-09, 
    5.710282e-09, 5.54072e-09, 5.514532e-09, 5.371754e-09, 5.536814e-09, 
    5.696727e-09, 5.982371e-09, 6.3357e-09, 6.961858e-09, 7.891266e-09,
  1.003695e-08, 9.186414e-09, 8.470073e-09, 7.659233e-09, 6.812325e-09, 
    5.985812e-09, 5.723699e-09, 5.646403e-09, 5.46633e-09, 5.66106e-09, 
    5.911398e-09, 6.134368e-09, 6.340332e-09, 6.721196e-09, 7.612348e-09,
  1.097824e-08, 9.715221e-09, 8.884054e-09, 7.954628e-09, 7.158733e-09, 
    6.411426e-09, 6.024669e-09, 5.886778e-09, 5.643782e-09, 5.735281e-09, 
    6.045215e-09, 6.286753e-09, 6.481998e-09, 6.671266e-09, 7.498501e-09,
  1.195013e-08, 1.039926e-08, 9.214008e-09, 8.242559e-09, 7.480931e-09, 
    6.895357e-09, 6.455209e-09, 6.161202e-09, 5.908601e-09, 5.853535e-09, 
    6.149093e-09, 6.450772e-09, 6.628443e-09, 6.741838e-09, 7.721242e-09,
  1.314529e-08, 1.131547e-08, 9.818657e-09, 8.51947e-09, 7.745979e-09, 
    7.236057e-09, 6.818292e-09, 6.445293e-09, 6.166057e-09, 6.07456e-09, 
    6.254757e-09, 6.525119e-09, 6.590005e-09, 6.795653e-09, 7.738249e-09,
  1.42906e-08, 1.246366e-08, 1.070561e-08, 9.127571e-09, 7.989688e-09, 
    7.503036e-09, 7.063335e-09, 6.696345e-09, 6.382926e-09, 6.332082e-09, 
    6.434626e-09, 6.566804e-09, 6.539805e-09, 6.757904e-09, 7.851828e-09,
  1.539793e-08, 1.350772e-08, 1.174758e-08, 1.002668e-08, 8.518659e-09, 
    7.719769e-09, 7.245183e-09, 6.877561e-09, 6.621835e-09, 6.572464e-09, 
    6.618887e-09, 6.690832e-09, 6.632297e-09, 6.878871e-09, 8.092168e-09,
  1.646324e-08, 1.437071e-08, 1.268318e-08, 1.101848e-08, 9.385505e-09, 
    8.122433e-09, 7.466461e-09, 6.968915e-09, 6.759301e-09, 6.777111e-09, 
    6.745474e-09, 6.803061e-09, 6.763535e-09, 7.028006e-09, 8.328435e-09,
  1.736877e-08, 1.534164e-08, 1.349062e-08, 1.179676e-08, 1.023287e-08, 
    8.829219e-09, 7.831959e-09, 7.231595e-09, 6.993671e-09, 6.974727e-09, 
    6.859055e-09, 6.892547e-09, 6.898238e-09, 7.241291e-09, 8.608713e-09,
  1.822934e-08, 1.628775e-08, 1.434354e-08, 1.259721e-08, 1.096356e-08, 
    9.608485e-09, 8.430384e-09, 7.859857e-09, 7.452838e-09, 7.218406e-09, 
    6.974623e-09, 6.949985e-09, 7.015966e-09, 7.420741e-09, 8.747092e-09,
  5.04994e-09, 5.100719e-09, 5.243437e-09, 5.440691e-09, 5.709371e-09, 
    6.15746e-09, 6.88933e-09, 7.394166e-09, 7.025426e-09, 6.914321e-09, 
    6.852413e-09, 6.008143e-09, 4.393002e-09, 3.961706e-09, 4.922465e-09,
  5.042424e-09, 5.092755e-09, 5.131785e-09, 5.351965e-09, 5.681618e-09, 
    5.993583e-09, 6.521154e-09, 7.416945e-09, 7.291135e-09, 7.178258e-09, 
    6.961868e-09, 6.730097e-09, 5.150191e-09, 4.104384e-09, 4.014872e-09,
  4.999137e-09, 5.13131e-09, 5.15995e-09, 5.296061e-09, 5.659599e-09, 
    5.844754e-09, 6.118043e-09, 7.152444e-09, 7.276754e-09, 7.366305e-09, 
    7.24959e-09, 7.034933e-09, 6.098438e-09, 4.843724e-09, 3.880422e-09,
  5.012534e-09, 5.221777e-09, 5.278828e-09, 5.342039e-09, 5.655749e-09, 
    5.782577e-09, 5.82079e-09, 6.601296e-09, 7.162058e-09, 7.334099e-09, 
    7.49549e-09, 7.208115e-09, 6.832977e-09, 5.675431e-09, 4.35821e-09,
  5.120213e-09, 5.338812e-09, 5.471383e-09, 5.476867e-09, 5.731365e-09, 
    5.861874e-09, 5.778718e-09, 6.188454e-09, 6.943456e-09, 6.981412e-09, 
    7.419097e-09, 7.326335e-09, 7.207328e-09, 6.481713e-09, 5.42665e-09,
  5.275632e-09, 5.459065e-09, 5.645412e-09, 5.659038e-09, 5.788775e-09, 
    6.006683e-09, 5.990365e-09, 6.124274e-09, 6.792117e-09, 6.902988e-09, 
    7.140545e-09, 7.266575e-09, 7.214695e-09, 6.990361e-09, 6.181051e-09,
  5.468372e-09, 5.60564e-09, 5.754278e-09, 5.865621e-09, 5.942343e-09, 
    6.178505e-09, 6.358903e-09, 6.334282e-09, 6.668672e-09, 6.998593e-09, 
    6.843316e-09, 7.330435e-09, 7.251003e-09, 7.442636e-09, 6.795765e-09,
  5.790185e-09, 5.81435e-09, 5.872346e-09, 5.999253e-09, 6.111134e-09, 
    6.380514e-09, 6.681869e-09, 6.808547e-09, 6.726698e-09, 7.09996e-09, 
    7.072507e-09, 7.046713e-09, 7.335759e-09, 7.38273e-09, 7.583616e-09,
  6.236721e-09, 6.057779e-09, 6.03546e-09, 6.105342e-09, 6.255274e-09, 
    6.543967e-09, 6.942761e-09, 7.189962e-09, 7.125888e-09, 7.237115e-09, 
    7.43869e-09, 7.08273e-09, 7.479895e-09, 7.403991e-09, 8.024993e-09,
  6.94793e-09, 6.448628e-09, 6.298159e-09, 6.180261e-09, 6.352349e-09, 
    6.624094e-09, 7.073707e-09, 7.503973e-09, 7.419673e-09, 7.606665e-09, 
    7.852527e-09, 7.627856e-09, 7.864516e-09, 7.8233e-09, 8.169095e-09,
  5.24889e-09, 5.959e-09, 6.715054e-09, 7.166097e-09, 7.444743e-09, 
    7.384039e-09, 7.135015e-09, 6.576125e-09, 5.855725e-09, 5.40761e-09, 
    5.988042e-09, 8.141397e-09, 1.07052e-08, 1.236789e-08, 1.318643e-08,
  5.192721e-09, 5.882357e-09, 6.611549e-09, 7.106539e-09, 7.357156e-09, 
    7.360987e-09, 7.20715e-09, 6.769283e-09, 6.154447e-09, 5.715393e-09, 
    5.874144e-09, 7.146914e-09, 9.283181e-09, 1.124314e-08, 1.2785e-08,
  5.111712e-09, 5.835617e-09, 6.548273e-09, 7.023986e-09, 7.26184e-09, 
    7.328115e-09, 7.274705e-09, 6.98776e-09, 6.522727e-09, 6.173523e-09, 
    5.937975e-09, 6.409103e-09, 7.901999e-09, 1.012172e-08, 1.184851e-08,
  5.061201e-09, 5.841768e-09, 6.518014e-09, 6.923896e-09, 7.12808e-09, 
    7.232368e-09, 7.305919e-09, 7.192408e-09, 6.958035e-09, 6.679175e-09, 
    6.394537e-09, 6.127255e-09, 6.851841e-09, 8.665236e-09, 1.036596e-08,
  5.046179e-09, 5.882158e-09, 6.511085e-09, 6.831289e-09, 7.011013e-09, 
    7.106106e-09, 7.227356e-09, 7.334338e-09, 7.25311e-09, 7.268198e-09, 
    7.131723e-09, 6.751261e-09, 6.613705e-09, 7.207529e-09, 8.743499e-09,
  5.084074e-09, 5.958319e-09, 6.527525e-09, 6.755546e-09, 6.899585e-09, 
    6.925002e-09, 7.031467e-09, 7.358367e-09, 7.502369e-09, 7.622355e-09, 
    7.757338e-09, 7.561051e-09, 7.080421e-09, 6.728702e-09, 7.435218e-09,
  5.126011e-09, 6.050395e-09, 6.559995e-09, 6.708842e-09, 6.778144e-09, 
    6.723932e-09, 6.780434e-09, 7.188662e-09, 7.491782e-09, 7.686601e-09, 
    7.961552e-09, 8.204122e-09, 7.94231e-09, 7.553308e-09, 7.121904e-09,
  5.195363e-09, 6.159241e-09, 6.582097e-09, 6.660129e-09, 6.644166e-09, 
    6.460543e-09, 6.480542e-09, 6.869559e-09, 7.282529e-09, 7.661338e-09, 
    7.817801e-09, 8.053566e-09, 8.347361e-09, 8.218463e-09, 7.852207e-09,
  5.265491e-09, 6.257684e-09, 6.589386e-09, 6.596957e-09, 6.490801e-09, 
    6.174843e-09, 6.198481e-09, 6.577077e-09, 6.773819e-09, 6.941435e-09, 
    6.912086e-09, 7.18015e-09, 7.792684e-09, 8.146534e-09, 8.736384e-09,
  5.333128e-09, 6.341272e-09, 6.563004e-09, 6.49806e-09, 6.326378e-09, 
    5.895122e-09, 5.951169e-09, 6.094469e-09, 5.937762e-09, 6.054246e-09, 
    6.399024e-09, 6.574394e-09, 7.041329e-09, 8.655259e-09, 8.801395e-09,
  6.80823e-09, 5.001108e-09, 4.042276e-09, 3.558124e-09, 4.045676e-09, 
    4.729962e-09, 5.719623e-09, 6.446354e-09, 5.591504e-09, 6.091113e-09, 
    9.88441e-09, 1.307446e-08, 1.385874e-08, 1.416656e-08, 1.474701e-08,
  8.604773e-09, 5.621646e-09, 4.398915e-09, 3.694091e-09, 4.003963e-09, 
    4.756202e-09, 5.733005e-09, 6.427857e-09, 5.640696e-09, 5.930469e-09, 
    9.056931e-09, 1.278872e-08, 1.370294e-08, 1.362272e-08, 1.451218e-08,
  1.084762e-08, 6.617194e-09, 4.81366e-09, 3.915232e-09, 3.974371e-09, 
    4.825167e-09, 5.853155e-09, 6.39572e-09, 5.652057e-09, 5.563033e-09, 
    7.987896e-09, 1.198769e-08, 1.352913e-08, 1.333055e-08, 1.413264e-08,
  1.290698e-08, 7.914637e-09, 5.343853e-09, 4.198529e-09, 4.053781e-09, 
    4.959326e-09, 5.973673e-09, 6.39916e-09, 5.748076e-09, 5.420923e-09, 
    6.84988e-09, 1.05323e-08, 1.316413e-08, 1.341192e-08, 1.368486e-08,
  1.379498e-08, 9.323506e-09, 6.013224e-09, 4.570514e-09, 4.224152e-09, 
    5.085766e-09, 6.053263e-09, 6.447976e-09, 5.909191e-09, 5.428487e-09, 
    6.114642e-09, 8.376115e-09, 1.197693e-08, 1.328627e-08, 1.305834e-08,
  1.43139e-08, 1.033073e-08, 6.764632e-09, 4.971803e-09, 4.523682e-09, 
    5.261369e-09, 6.13027e-09, 6.51078e-09, 6.184118e-09, 5.784035e-09, 
    6.054872e-09, 7.229067e-09, 9.813156e-09, 1.256988e-08, 1.297927e-08,
  1.450802e-08, 1.092063e-08, 7.481859e-09, 5.406674e-09, 4.86431e-09, 
    5.436954e-09, 6.227786e-09, 6.632592e-09, 6.481408e-09, 6.099578e-09, 
    6.386458e-09, 7.069986e-09, 8.073841e-09, 1.072787e-08, 1.272259e-08,
  1.444706e-08, 1.118527e-08, 8.051498e-09, 5.849142e-09, 5.242619e-09, 
    5.630938e-09, 6.319373e-09, 6.673724e-09, 6.752696e-09, 6.660782e-09, 
    6.974917e-09, 7.818341e-09, 8.024684e-09, 8.719611e-09, 1.105052e-08,
  1.428697e-08, 1.12316e-08, 8.291358e-09, 6.222407e-09, 5.604388e-09, 
    5.80423e-09, 6.385479e-09, 6.787153e-09, 7.101638e-09, 7.122968e-09, 
    7.415737e-09, 8.293168e-09, 8.301665e-09, 8.3194e-09, 8.887949e-09,
  1.400484e-08, 1.116915e-08, 8.369706e-09, 6.530268e-09, 5.921436e-09, 
    5.96759e-09, 6.46866e-09, 6.982114e-09, 7.305408e-09, 7.254113e-09, 
    7.737073e-09, 8.346429e-09, 8.531862e-09, 8.544262e-09, 8.424118e-09,
  6.558119e-09, 5.630391e-09, 5.355879e-09, 5.065357e-09, 4.238489e-09, 
    3.65774e-09, 3.376867e-09, 4.374778e-09, 6.435531e-09, 7.181389e-09, 
    1.037455e-08, 1.378069e-08, 1.441826e-08, 1.175447e-08, 8.233454e-09,
  7.302655e-09, 5.964375e-09, 5.384461e-09, 5.096651e-09, 4.525014e-09, 
    3.906313e-09, 3.497221e-09, 4.025521e-09, 5.957575e-09, 6.419975e-09, 
    8.661171e-09, 1.265218e-08, 1.423194e-08, 1.382473e-08, 1.042406e-08,
  9.067085e-09, 6.612153e-09, 5.579427e-09, 5.152448e-09, 4.651416e-09, 
    4.113894e-09, 3.587864e-09, 3.810817e-09, 5.691247e-09, 6.271456e-09, 
    7.831331e-09, 1.136696e-08, 1.425806e-08, 1.481727e-08, 1.244401e-08,
  1.266241e-08, 7.779173e-09, 5.978972e-09, 5.242269e-09, 4.6976e-09, 
    4.231344e-09, 3.707873e-09, 3.693564e-09, 5.320569e-09, 6.027315e-09, 
    6.838091e-09, 1.011892e-08, 1.361191e-08, 1.510792e-08, 1.401494e-08,
  1.646749e-08, 1.037199e-08, 6.87543e-09, 5.507161e-09, 4.773868e-09, 
    4.268166e-09, 3.825535e-09, 3.651471e-09, 4.968053e-09, 5.968837e-09, 
    6.450817e-09, 8.423475e-09, 1.183809e-08, 1.501395e-08, 1.505097e-08,
  2.049415e-08, 1.344821e-08, 8.464242e-09, 6.119421e-09, 4.919261e-09, 
    4.319035e-09, 3.894846e-09, 3.669633e-09, 4.669889e-09, 5.813114e-09, 
    6.178861e-09, 7.661361e-09, 1.003701e-08, 1.338753e-08, 1.517177e-08,
  2.38138e-08, 1.805704e-08, 1.119942e-08, 7.164926e-09, 5.293056e-09, 
    4.396009e-09, 3.966645e-09, 3.739574e-09, 4.477869e-09, 5.612881e-09, 
    6.057459e-09, 7.024715e-09, 8.969509e-09, 1.129912e-08, 1.47144e-08,
  2.434833e-08, 2.135402e-08, 1.500437e-08, 9.24525e-09, 6.079685e-09, 
    4.616299e-09, 4.029467e-09, 3.777536e-09, 4.402168e-09, 5.42309e-09, 
    6.026829e-09, 6.90581e-09, 8.145705e-09, 9.489699e-09, 1.223039e-08,
  2.394194e-08, 2.323152e-08, 1.882171e-08, 1.199774e-08, 7.349181e-09, 
    5.049162e-09, 4.205746e-09, 3.847139e-09, 4.353308e-09, 5.223137e-09, 
    5.927131e-09, 6.850263e-09, 7.931646e-09, 8.69494e-09, 1.033924e-08,
  2.199458e-08, 2.361475e-08, 2.149104e-08, 1.553424e-08, 9.387096e-09, 
    5.834241e-09, 4.467164e-09, 3.990615e-09, 4.440993e-09, 5.111829e-09, 
    5.867109e-09, 6.915901e-09, 7.835786e-09, 8.341186e-09, 8.824713e-09,
  8.917325e-09, 7.219623e-09, 5.330258e-09, 3.911727e-09, 3.475443e-09, 
    4.132942e-09, 5.388325e-09, 7.085736e-09, 9.10605e-09, 1.110488e-08, 
    1.344365e-08, 1.347288e-08, 9.569352e-09, 7.67638e-09, 8.096062e-09,
  9.050596e-09, 7.440913e-09, 5.643914e-09, 4.322548e-09, 3.727231e-09, 
    4.197703e-09, 4.853172e-09, 6.012262e-09, 7.878912e-09, 9.667624e-09, 
    1.248547e-08, 1.377114e-08, 1.180797e-08, 8.39144e-09, 7.881046e-09,
  9.257733e-09, 7.694437e-09, 5.991438e-09, 4.759405e-09, 4.092071e-09, 
    4.261403e-09, 4.717655e-09, 5.572334e-09, 7.371265e-09, 8.886616e-09, 
    1.150397e-08, 1.350888e-08, 1.302906e-08, 9.921633e-09, 7.910928e-09,
  9.675134e-09, 7.989224e-09, 6.330819e-09, 5.169835e-09, 4.484739e-09, 
    4.439773e-09, 4.559418e-09, 4.804436e-09, 6.378071e-09, 7.599781e-09, 
    9.877763e-09, 1.309688e-08, 1.376219e-08, 1.149762e-08, 8.680043e-09,
  1.0218e-08, 8.419199e-09, 6.716025e-09, 5.59086e-09, 4.88505e-09, 
    4.749344e-09, 4.651465e-09, 4.605962e-09, 5.82968e-09, 7.022571e-09, 
    8.09657e-09, 1.09481e-08, 1.354842e-08, 1.344547e-08, 1.017248e-08,
  1.114607e-08, 8.943379e-09, 7.146377e-09, 5.99675e-09, 5.259408e-09, 
    5.091958e-09, 4.834151e-09, 4.315115e-09, 4.95428e-09, 6.420974e-09, 
    7.279429e-09, 8.859602e-09, 1.176037e-08, 1.359803e-08, 1.171539e-08,
  1.228395e-08, 9.993593e-09, 7.772366e-09, 6.469221e-09, 5.627161e-09, 
    5.367921e-09, 5.108538e-09, 4.411181e-09, 4.403771e-09, 5.659567e-09, 
    6.691218e-09, 7.63062e-09, 9.747783e-09, 1.204441e-08, 1.352752e-08,
  1.340906e-08, 1.137785e-08, 8.74786e-09, 7.03383e-09, 6.034572e-09, 
    5.7006e-09, 5.424493e-09, 4.656423e-09, 4.207739e-09, 4.834916e-09, 
    6.181938e-09, 7.007861e-09, 8.095441e-09, 1.002273e-08, 1.249056e-08,
  1.416596e-08, 1.284039e-08, 1.049136e-08, 8.041934e-09, 6.527335e-09, 
    5.996409e-09, 5.72303e-09, 5.015565e-09, 4.266221e-09, 4.24728e-09, 
    5.339911e-09, 6.517597e-09, 7.478191e-09, 8.444148e-09, 1.058962e-08,
  1.428277e-08, 1.397502e-08, 1.221432e-08, 9.7674e-09, 7.467903e-09, 
    6.421945e-09, 5.982084e-09, 5.410543e-09, 4.510444e-09, 4.11954e-09, 
    4.569392e-09, 5.8507e-09, 6.854214e-09, 7.765483e-09, 9.076181e-09,
  1.069021e-08, 8.855539e-09, 7.017126e-09, 5.457113e-09, 6.339951e-09, 
    8.238114e-09, 9.060734e-09, 1.104477e-08, 1.193349e-08, 1.207501e-08, 
    1.139158e-08, 9.647784e-09, 8.842234e-09, 8.941328e-09, 9.532106e-09,
  9.826384e-09, 7.955619e-09, 5.889325e-09, 5.315223e-09, 7.304305e-09, 
    8.44135e-09, 9.861214e-09, 1.148745e-08, 1.198162e-08, 1.185654e-08, 
    1.111869e-08, 9.774431e-09, 9.119473e-09, 8.80365e-09, 9.391909e-09,
  8.919403e-09, 7.061428e-09, 5.337534e-09, 6.201582e-09, 8.045227e-09, 
    8.900107e-09, 1.024289e-08, 1.122077e-08, 1.165878e-08, 1.159123e-08, 
    1.094835e-08, 9.850001e-09, 9.142236e-09, 8.825981e-09, 9.021442e-09,
  8.380536e-09, 6.577268e-09, 5.919603e-09, 7.02904e-09, 7.817412e-09, 
    8.673299e-09, 9.55121e-09, 1.015963e-08, 1.080418e-08, 1.117319e-08, 
    1.101181e-08, 1.009228e-08, 9.169353e-09, 8.833655e-09, 8.639e-09,
  8.057727e-09, 6.881553e-09, 6.583902e-09, 6.915517e-09, 7.624413e-09, 
    8.277811e-09, 8.911045e-09, 9.413478e-09, 1.013732e-08, 1.061461e-08, 
    1.103401e-08, 1.049065e-08, 9.576755e-09, 8.87517e-09, 8.546309e-09,
  8.279257e-09, 7.129369e-09, 6.439549e-09, 6.480327e-09, 6.985435e-09, 
    7.413771e-09, 7.889676e-09, 8.457756e-09, 9.136713e-09, 9.649468e-09, 
    1.036843e-08, 1.050985e-08, 9.991023e-09, 8.941623e-09, 8.555119e-09,
  8.341527e-09, 6.979511e-09, 6.097339e-09, 5.97381e-09, 6.322654e-09, 
    6.684367e-09, 7.136648e-09, 7.694565e-09, 8.452266e-09, 9.037572e-09, 
    9.757147e-09, 1.02872e-08, 1.032131e-08, 9.74075e-09, 8.785592e-09,
  8.250188e-09, 6.881021e-09, 5.907812e-09, 5.558168e-09, 5.714735e-09, 
    5.999729e-09, 6.477896e-09, 6.899886e-09, 7.707303e-09, 8.444817e-09, 
    9.10141e-09, 9.618777e-09, 9.945686e-09, 9.841505e-09, 9.317419e-09,
  8.191868e-09, 6.876611e-09, 5.796195e-09, 5.245457e-09, 5.220997e-09, 
    5.508519e-09, 5.904667e-09, 6.288863e-09, 6.953886e-09, 7.861017e-09, 
    8.730233e-09, 9.391767e-09, 9.709693e-09, 9.818048e-09, 9.578236e-09,
  8.222699e-09, 6.948057e-09, 5.840808e-09, 5.078704e-09, 4.893026e-09, 
    5.054837e-09, 5.439752e-09, 5.871823e-09, 6.305627e-09, 7.192423e-09, 
    8.19974e-09, 9.075314e-09, 9.63565e-09, 9.711579e-09, 9.534807e-09,
  2.32999e-08, 2.195469e-08, 2.059089e-08, 1.896829e-08, 1.699714e-08, 
    1.479577e-08, 1.275317e-08, 1.084385e-08, 1.018075e-08, 1.005276e-08, 
    9.580088e-09, 9.441226e-09, 9.108843e-09, 9.149577e-09, 9.390255e-09,
  2.30215e-08, 2.128361e-08, 1.979139e-08, 1.80218e-08, 1.581979e-08, 
    1.35947e-08, 1.164412e-08, 1.036402e-08, 1.051811e-08, 9.829215e-09, 
    9.236037e-09, 9.378504e-09, 9.461237e-09, 9.674041e-09, 9.705922e-09,
  2.255031e-08, 2.059149e-08, 1.878467e-08, 1.68763e-08, 1.456858e-08, 
    1.249657e-08, 1.095192e-08, 1.079624e-08, 1.025773e-08, 9.361585e-09, 
    9.282531e-09, 9.686523e-09, 9.744664e-09, 9.775401e-09, 9.676365e-09,
  2.184171e-08, 1.968372e-08, 1.769107e-08, 1.561759e-08, 1.351813e-08, 
    1.174641e-08, 1.090297e-08, 1.071003e-08, 9.531081e-09, 9.070931e-09, 
    9.445324e-09, 9.664782e-09, 9.741634e-09, 9.713525e-09, 9.716207e-09,
  2.075464e-08, 1.856091e-08, 1.665315e-08, 1.450488e-08, 1.269909e-08, 
    1.139382e-08, 1.100019e-08, 9.990407e-09, 9.044625e-09, 9.233879e-09, 
    9.476354e-09, 9.587398e-09, 9.745659e-09, 9.758192e-09, 9.7585e-09,
  1.942658e-08, 1.748643e-08, 1.56182e-08, 1.355521e-08, 1.21504e-08, 
    1.119178e-08, 1.050208e-08, 9.318947e-09, 8.952255e-09, 9.300471e-09, 
    9.36337e-09, 9.431519e-09, 9.686682e-09, 9.813616e-09, 9.833721e-09,
  1.816899e-08, 1.637694e-08, 1.46221e-08, 1.28307e-08, 1.178832e-08, 
    1.088089e-08, 9.942877e-09, 9.098898e-09, 9.220621e-09, 9.201165e-09, 
    9.129097e-09, 9.270363e-09, 9.50408e-09, 9.68556e-09, 9.716056e-09,
  1.69249e-08, 1.532247e-08, 1.365149e-08, 1.22594e-08, 1.123969e-08, 
    1.046427e-08, 9.568152e-09, 9.152667e-09, 9.303225e-09, 9.09963e-09, 
    8.999861e-09, 9.072134e-09, 9.271661e-09, 9.47219e-09, 9.586416e-09,
  1.561966e-08, 1.411774e-08, 1.278136e-08, 1.155888e-08, 1.081911e-08, 
    1.007369e-08, 9.404361e-09, 9.434205e-09, 9.315584e-09, 9.100678e-09, 
    8.965439e-09, 8.875232e-09, 9.04268e-09, 9.194393e-09, 9.4319e-09,
  1.429024e-08, 1.297716e-08, 1.191171e-08, 1.098155e-08, 1.044055e-08, 
    9.727462e-09, 9.448536e-09, 9.524606e-09, 9.284827e-09, 9.048122e-09, 
    8.819511e-09, 8.62348e-09, 8.742302e-09, 8.929463e-09, 9.223688e-09,
  7.140104e-09, 7.879262e-09, 9.183748e-09, 1.19955e-08, 1.478543e-08, 
    2.003196e-08, 2.327637e-08, 2.079655e-08, 1.210633e-08, 9.613336e-09, 
    9.89989e-09, 1.006597e-08, 9.786651e-09, 9.593313e-09, 9.657218e-09,
  7.917101e-09, 8.507783e-09, 9.490679e-09, 1.378755e-08, 1.657117e-08, 
    2.141293e-08, 2.250515e-08, 1.803554e-08, 1.052915e-08, 9.774813e-09, 
    9.998163e-09, 1.019106e-08, 9.96717e-09, 9.999586e-09, 1.032555e-08,
  8.582979e-09, 9.1717e-09, 1.013503e-08, 1.434263e-08, 1.724874e-08, 
    2.136226e-08, 2.113454e-08, 1.475495e-08, 1.001486e-08, 9.94339e-09, 
    1.019388e-08, 1.016292e-08, 1.016079e-08, 1.043856e-08, 1.109538e-08,
  9.191496e-09, 9.977239e-09, 1.124323e-08, 1.520551e-08, 1.862822e-08, 
    2.119586e-08, 1.956853e-08, 1.275274e-08, 9.944784e-09, 1.003231e-08, 
    1.022546e-08, 1.011331e-08, 1.025466e-08, 1.064971e-08, 1.138592e-08,
  9.794767e-09, 1.069005e-08, 1.239867e-08, 1.601166e-08, 1.961114e-08, 
    2.062517e-08, 1.767398e-08, 1.116967e-08, 9.927518e-09, 1.016364e-08, 
    1.011509e-08, 1.015432e-08, 1.035266e-08, 1.085006e-08, 1.156002e-08,
  1.049931e-08, 1.145586e-08, 1.353619e-08, 1.692766e-08, 1.990625e-08, 
    1.972727e-08, 1.56743e-08, 1.038782e-08, 1.00455e-08, 1.017981e-08, 
    1.011319e-08, 1.02189e-08, 1.039187e-08, 1.106274e-08, 1.165558e-08,
  1.121148e-08, 1.213995e-08, 1.458658e-08, 1.739929e-08, 1.967072e-08, 
    1.845354e-08, 1.391236e-08, 1.008617e-08, 1.020414e-08, 1.010415e-08, 
    1.006571e-08, 1.01046e-08, 1.03735e-08, 1.103142e-08, 1.152638e-08,
  1.194854e-08, 1.294129e-08, 1.555591e-08, 1.783613e-08, 1.90145e-08, 
    1.698371e-08, 1.258026e-08, 1.009731e-08, 1.025401e-08, 9.96757e-09, 
    1.000569e-08, 9.984205e-09, 1.027662e-08, 1.081086e-08, 1.119148e-08,
  1.272306e-08, 1.386807e-08, 1.620307e-08, 1.809879e-08, 1.803396e-08, 
    1.581521e-08, 1.158156e-08, 1.016835e-08, 1.011597e-08, 9.91492e-09, 
    9.89766e-09, 9.873321e-09, 1.016602e-08, 1.059859e-08, 1.091106e-08,
  1.358186e-08, 1.470584e-08, 1.667658e-08, 1.796499e-08, 1.696175e-08, 
    1.468037e-08, 1.087439e-08, 1.01871e-08, 9.993086e-09, 9.877296e-09, 
    9.743023e-09, 9.770577e-09, 9.911776e-09, 1.026938e-08, 1.04792e-08,
  1.534885e-08, 1.368189e-08, 1.272725e-08, 1.150104e-08, 1.096987e-08, 
    1.069007e-08, 1.176344e-08, 1.294521e-08, 1.232277e-08, 1.144427e-08, 
    1.157483e-08, 1.168599e-08, 1.181559e-08, 1.201588e-08, 1.270016e-08,
  1.489691e-08, 1.328591e-08, 1.21395e-08, 1.08515e-08, 1.006141e-08, 
    1.134904e-08, 1.165959e-08, 1.286526e-08, 1.181963e-08, 1.202715e-08, 
    1.209564e-08, 1.183519e-08, 1.252458e-08, 1.374399e-08, 1.540088e-08,
  1.456005e-08, 1.281878e-08, 1.15942e-08, 1.007682e-08, 9.488364e-09, 
    1.108087e-08, 1.243405e-08, 1.167397e-08, 1.108006e-08, 1.18302e-08, 
    1.153309e-08, 1.278693e-08, 1.447295e-08, 1.577683e-08, 1.660966e-08,
  1.41955e-08, 1.238481e-08, 1.08581e-08, 9.25719e-09, 9.368322e-09, 
    1.110295e-08, 1.303603e-08, 1.207457e-08, 1.130609e-08, 1.109455e-08, 
    1.246408e-08, 1.471026e-08, 1.573538e-08, 1.620749e-08, 1.685928e-08,
  1.385498e-08, 1.175419e-08, 9.983482e-09, 8.490671e-09, 9.596576e-09, 
    1.158374e-08, 1.350752e-08, 1.183015e-08, 1.073257e-08, 1.208284e-08, 
    1.420043e-08, 1.520124e-08, 1.58219e-08, 1.657384e-08, 1.690614e-08,
  1.342223e-08, 1.100288e-08, 8.931178e-09, 8.065579e-09, 1.000502e-08, 
    1.222455e-08, 1.349112e-08, 1.089133e-08, 1.112231e-08, 1.319491e-08, 
    1.4465e-08, 1.519667e-08, 1.608751e-08, 1.651927e-08, 1.701612e-08,
  1.279864e-08, 9.982093e-09, 8.094077e-09, 8.284534e-09, 1.078173e-08, 
    1.302142e-08, 1.253399e-08, 1.066364e-08, 1.231364e-08, 1.344505e-08, 
    1.454627e-08, 1.52892e-08, 1.62628e-08, 1.662563e-08, 1.731023e-08,
  1.200091e-08, 9.046296e-09, 7.560557e-09, 8.768311e-09, 1.140567e-08, 
    1.344063e-08, 1.151357e-08, 1.085017e-08, 1.26085e-08, 1.342561e-08, 
    1.432275e-08, 1.506333e-08, 1.596181e-08, 1.663593e-08, 1.728167e-08,
  1.100967e-08, 8.153084e-09, 7.402994e-09, 9.500007e-09, 1.2407e-08, 
    1.295658e-08, 1.076041e-08, 1.140448e-08, 1.259794e-08, 1.341002e-08, 
    1.418157e-08, 1.517409e-08, 1.609826e-08, 1.719873e-08, 1.814258e-08,
  1.001557e-08, 7.582136e-09, 7.579669e-09, 9.95102e-09, 1.309048e-08, 
    1.238516e-08, 1.062502e-08, 1.179462e-08, 1.252479e-08, 1.350916e-08, 
    1.441786e-08, 1.557967e-08, 1.672297e-08, 1.815065e-08, 1.920565e-08,
  2.225372e-08, 2.058648e-08, 1.716568e-08, 1.45636e-08, 1.425526e-08, 
    1.418729e-08, 1.423011e-08, 1.392767e-08, 1.361094e-08, 1.352055e-08, 
    1.373194e-08, 1.425503e-08, 1.518305e-08, 1.654877e-08, 1.715988e-08,
  2.203807e-08, 2.126254e-08, 1.927589e-08, 1.629688e-08, 1.450892e-08, 
    1.442036e-08, 1.426112e-08, 1.404603e-08, 1.377096e-08, 1.362305e-08, 
    1.385754e-08, 1.43013e-08, 1.503293e-08, 1.634403e-08, 1.760618e-08,
  2.175211e-08, 2.096726e-08, 1.963259e-08, 1.796975e-08, 1.541686e-08, 
    1.451181e-08, 1.425075e-08, 1.403606e-08, 1.384204e-08, 1.385249e-08, 
    1.414982e-08, 1.454298e-08, 1.508433e-08, 1.610643e-08, 1.715703e-08,
  2.108635e-08, 2.045628e-08, 1.966995e-08, 1.86275e-08, 1.66544e-08, 
    1.494206e-08, 1.40635e-08, 1.38779e-08, 1.396355e-08, 1.40663e-08, 
    1.441252e-08, 1.463664e-08, 1.497411e-08, 1.563751e-08, 1.656498e-08,
  2.041388e-08, 1.982088e-08, 1.933635e-08, 1.871152e-08, 1.727356e-08, 
    1.561631e-08, 1.437838e-08, 1.39418e-08, 1.406275e-08, 1.400497e-08, 
    1.470403e-08, 1.484443e-08, 1.492573e-08, 1.553396e-08, 1.604076e-08,
  1.994711e-08, 1.96653e-08, 1.926243e-08, 1.851846e-08, 1.749772e-08, 
    1.59411e-08, 1.464853e-08, 1.426905e-08, 1.414845e-08, 1.467368e-08, 
    1.49209e-08, 1.514078e-08, 1.541511e-08, 1.557449e-08, 1.59973e-08,
  1.96342e-08, 1.953321e-08, 1.89609e-08, 1.810601e-08, 1.709957e-08, 
    1.567993e-08, 1.471566e-08, 1.418592e-08, 1.437793e-08, 1.509328e-08, 
    1.542352e-08, 1.571449e-08, 1.558742e-08, 1.608081e-08, 1.563037e-08,
  1.939458e-08, 1.906372e-08, 1.83931e-08, 1.72394e-08, 1.617937e-08, 
    1.501495e-08, 1.445787e-08, 1.432303e-08, 1.541091e-08, 1.569479e-08, 
    1.591157e-08, 1.576765e-08, 1.576133e-08, 1.570727e-08, 1.388977e-08,
  1.893356e-08, 1.840151e-08, 1.741255e-08, 1.615492e-08, 1.49977e-08, 
    1.440656e-08, 1.423771e-08, 1.48697e-08, 1.564524e-08, 1.572178e-08, 
    1.57383e-08, 1.555769e-08, 1.537791e-08, 1.422099e-08, 1.196617e-08,
  1.826742e-08, 1.745436e-08, 1.636878e-08, 1.492846e-08, 1.407391e-08, 
    1.391589e-08, 1.430784e-08, 1.539447e-08, 1.573417e-08, 1.574546e-08, 
    1.582095e-08, 1.521749e-08, 1.443634e-08, 1.297721e-08, 1.098474e-08,
  2.530511e-08, 2.323247e-08, 2.13817e-08, 1.770199e-08, 1.433412e-08, 
    1.108788e-08, 8.571496e-09, 7.089129e-09, 6.182774e-09, 5.478358e-09, 
    4.791881e-09, 4.18144e-09, 4.323803e-09, 5.499828e-09, 7.387685e-09,
  2.786779e-08, 2.421866e-08, 2.241596e-08, 1.987098e-08, 1.605695e-08, 
    1.265663e-08, 9.774064e-09, 7.77422e-09, 6.365194e-09, 5.46928e-09, 
    4.917709e-09, 4.339458e-09, 4.22286e-09, 5.563935e-09, 8.595451e-09,
  2.862063e-08, 2.617556e-08, 2.311387e-08, 2.118118e-08, 1.802359e-08, 
    1.426105e-08, 1.089809e-08, 8.40624e-09, 6.518804e-09, 5.551975e-09, 
    5.167046e-09, 4.531318e-09, 4.466636e-09, 6.351526e-09, 1.130496e-08,
  2.831423e-08, 2.682573e-08, 2.386939e-08, 2.14499e-08, 1.912279e-08, 
    1.557775e-08, 1.188871e-08, 8.887044e-09, 6.839147e-09, 6.035599e-09, 
    5.486443e-09, 4.879649e-09, 5.155337e-09, 7.727608e-09, 1.509065e-08,
  2.824635e-08, 2.61236e-08, 2.441176e-08, 2.160631e-08, 1.954058e-08, 
    1.61249e-08, 1.234627e-08, 9.352399e-09, 7.307142e-09, 6.29906e-09, 
    5.713345e-09, 5.185283e-09, 6.260061e-09, 9.513512e-09, 1.671488e-08,
  2.79783e-08, 2.517378e-08, 2.41654e-08, 2.150296e-08, 1.93683e-08, 
    1.671238e-08, 1.245449e-08, 9.378357e-09, 7.458381e-09, 6.38821e-09, 
    5.775105e-09, 5.585295e-09, 7.471075e-09, 1.29455e-08, 1.828214e-08,
  2.730709e-08, 2.450266e-08, 2.310849e-08, 2.119887e-08, 1.888904e-08, 
    1.649341e-08, 1.251164e-08, 9.366788e-09, 7.360626e-09, 6.349318e-09, 
    5.812973e-09, 6.197024e-09, 8.942083e-09, 1.57776e-08, 1.711315e-08,
  2.626371e-08, 2.347909e-08, 2.1961e-08, 2.024206e-08, 1.831236e-08, 
    1.582421e-08, 1.225042e-08, 9.145618e-09, 7.195278e-09, 6.197146e-09, 
    6.116538e-09, 7.360598e-09, 1.194029e-08, 1.725531e-08, 1.452881e-08,
  2.484645e-08, 2.216552e-08, 2.073006e-08, 1.90708e-08, 1.722459e-08, 
    1.498667e-08, 1.180293e-08, 8.890806e-09, 6.944186e-09, 6.3139e-09, 
    6.793624e-09, 9.269062e-09, 1.462717e-08, 1.658737e-08, 1.169487e-08,
  2.284363e-08, 2.092067e-08, 1.961581e-08, 1.780434e-08, 1.62955e-08, 
    1.391205e-08, 1.098924e-08, 8.510883e-09, 6.970165e-09, 6.705223e-09, 
    8.05812e-09, 1.152164e-08, 1.63374e-08, 1.439594e-08, 9.519352e-09,
  2.042867e-08, 1.936788e-08, 1.801046e-08, 1.59575e-08, 1.315147e-08, 
    1.065147e-08, 9.302665e-09, 8.914264e-09, 8.34806e-09, 7.53997e-09, 
    6.566339e-09, 5.492514e-09, 5.380127e-09, 6.392048e-09, 9.403956e-09,
  2.27741e-08, 2.119338e-08, 1.964743e-08, 1.790226e-08, 1.568655e-08, 
    1.304484e-08, 1.043775e-08, 9.201114e-09, 8.596718e-09, 7.886769e-09, 
    6.912011e-09, 5.787081e-09, 5.474308e-09, 6.037252e-09, 1.007112e-08,
  2.393946e-08, 2.324999e-08, 2.147071e-08, 1.987107e-08, 1.777853e-08, 
    1.542848e-08, 1.242662e-08, 1.017175e-08, 9.11122e-09, 8.379462e-09, 
    7.294238e-09, 6.004285e-09, 5.578492e-09, 5.699252e-09, 1.142461e-08,
  2.525235e-08, 2.417335e-08, 2.335688e-08, 2.135656e-08, 1.997215e-08, 
    1.767005e-08, 1.463705e-08, 1.155413e-08, 9.744673e-09, 8.789977e-09, 
    7.681265e-09, 6.220462e-09, 5.677808e-09, 6.091458e-09, 1.303664e-08,
  2.71996e-08, 2.536913e-08, 2.429803e-08, 2.299345e-08, 2.117857e-08, 
    1.998695e-08, 1.721483e-08, 1.358222e-08, 1.085524e-08, 9.331425e-09, 
    7.975019e-09, 6.357209e-09, 5.697106e-09, 6.980014e-09, 1.259066e-08,
  2.886445e-08, 2.761124e-08, 2.559519e-08, 2.437767e-08, 2.239382e-08, 
    2.112705e-08, 1.911786e-08, 1.539631e-08, 1.19706e-08, 9.83184e-09, 
    8.238276e-09, 6.508553e-09, 5.673918e-09, 8.699007e-09, 1.233543e-08,
  2.971903e-08, 2.900533e-08, 2.75494e-08, 2.552478e-08, 2.39286e-08, 
    2.228133e-08, 2.049653e-08, 1.687236e-08, 1.292721e-08, 1.012588e-08, 
    8.302011e-09, 6.524711e-09, 5.805014e-09, 1.009874e-08, 1.215013e-08,
  3.067846e-08, 2.956994e-08, 2.913705e-08, 2.698224e-08, 2.49883e-08, 
    2.354918e-08, 2.137087e-08, 1.793247e-08, 1.354613e-08, 1.015572e-08, 
    8.158898e-09, 6.488025e-09, 6.725823e-09, 1.118803e-08, 1.224102e-08,
  3.148342e-08, 3.001482e-08, 2.96924e-08, 2.821573e-08, 2.613243e-08, 
    2.457879e-08, 2.246999e-08, 1.851335e-08, 1.370849e-08, 9.978777e-09, 
    7.861022e-09, 6.439184e-09, 7.704957e-09, 1.169852e-08, 1.217543e-08,
  3.181454e-08, 2.975597e-08, 2.979369e-08, 2.905608e-08, 2.707218e-08, 
    2.541185e-08, 2.334392e-08, 1.894441e-08, 1.348735e-08, 9.653109e-09, 
    7.546669e-09, 6.75659e-09, 9.361274e-09, 1.214969e-08, 1.226654e-08,
  8.805364e-09, 7.96364e-09, 7.884833e-09, 7.949756e-09, 8.408833e-09, 
    8.586153e-09, 9.207591e-09, 9.995561e-09, 9.491713e-09, 8.874895e-09, 
    9.141351e-09, 9.672896e-09, 1.093809e-08, 1.184207e-08, 1.1692e-08,
  1.001748e-08, 8.670686e-09, 8.326354e-09, 8.37147e-09, 8.833103e-09, 
    9.318156e-09, 9.556071e-09, 1.02518e-08, 9.76529e-09, 8.969742e-09, 
    8.975001e-09, 9.558553e-09, 1.086987e-08, 1.190858e-08, 1.155934e-08,
  1.145508e-08, 9.60816e-09, 8.816832e-09, 8.77793e-09, 9.065026e-09, 
    9.751899e-09, 1.008396e-08, 1.065141e-08, 1.019093e-08, 9.275745e-09, 
    9.006262e-09, 9.616431e-09, 1.113624e-08, 1.199572e-08, 1.150043e-08,
  1.284397e-08, 1.102702e-08, 9.437323e-09, 9.057455e-09, 9.296057e-09, 
    9.923093e-09, 1.05151e-08, 1.098307e-08, 1.062393e-08, 9.560503e-09, 
    8.888187e-09, 9.670314e-09, 1.134188e-08, 1.20136e-08, 1.125238e-08,
  1.417375e-08, 1.24583e-08, 1.067742e-08, 9.575409e-09, 9.413329e-09, 
    9.901037e-09, 1.080702e-08, 1.130542e-08, 1.116959e-08, 9.950259e-09, 
    8.926683e-09, 9.704499e-09, 1.149532e-08, 1.211176e-08, 1.124235e-08,
  1.557117e-08, 1.388624e-08, 1.17853e-08, 1.049907e-08, 9.711884e-09, 
    1.003053e-08, 1.083931e-08, 1.156422e-08, 1.169943e-08, 1.04071e-08, 
    9.020785e-09, 9.707922e-09, 1.193735e-08, 1.216043e-08, 1.108344e-08,
  1.698362e-08, 1.56998e-08, 1.356436e-08, 1.140539e-08, 1.020241e-08, 
    1.003836e-08, 1.089188e-08, 1.170003e-08, 1.218985e-08, 1.09298e-08, 
    9.237513e-09, 9.669303e-09, 1.223956e-08, 1.212293e-08, 1.087051e-08,
  1.896795e-08, 1.728335e-08, 1.543714e-08, 1.315395e-08, 1.10479e-08, 
    1.021116e-08, 1.086935e-08, 1.179677e-08, 1.239014e-08, 1.154796e-08, 
    9.58027e-09, 9.663911e-09, 1.273912e-08, 1.180954e-08, 1.023002e-08,
  2.114145e-08, 1.966145e-08, 1.768825e-08, 1.504354e-08, 1.260769e-08, 
    1.066637e-08, 1.076907e-08, 1.185452e-08, 1.261456e-08, 1.209546e-08, 
    1.0007e-08, 9.761913e-09, 1.291523e-08, 1.133922e-08, 9.887251e-09,
  2.327389e-08, 2.151712e-08, 1.974138e-08, 1.761481e-08, 1.459376e-08, 
    1.185608e-08, 1.076603e-08, 1.174845e-08, 1.272088e-08, 1.257374e-08, 
    1.045848e-08, 9.890791e-09, 1.309963e-08, 1.084268e-08, 9.413816e-09,
  1.406004e-08, 1.331761e-08, 9.542956e-09, 6.684549e-09, 6.011802e-09, 
    5.760795e-09, 8.545436e-09, 1.083799e-08, 1.083822e-08, 1.052751e-08, 
    9.533554e-09, 9.058907e-09, 8.494029e-09, 9.11518e-09, 9.156239e-09,
  1.281608e-08, 1.498016e-08, 1.280675e-08, 8.826467e-09, 6.58527e-09, 
    5.724338e-09, 6.469721e-09, 1.00204e-08, 1.073011e-08, 1.075585e-08, 
    9.623871e-09, 9.314698e-09, 8.225465e-09, 8.592791e-09, 8.651027e-09,
  1.127073e-08, 1.386969e-08, 1.524609e-08, 1.231749e-08, 8.813605e-09, 
    6.133878e-09, 5.76817e-09, 8.219736e-09, 1.085059e-08, 1.095902e-08, 
    9.806085e-09, 9.563906e-09, 8.288859e-09, 8.270979e-09, 8.443471e-09,
  1.104574e-08, 1.19905e-08, 1.442895e-08, 1.455567e-08, 1.173099e-08, 
    8.27285e-09, 5.815397e-09, 6.992678e-09, 9.851477e-09, 1.117606e-08, 
    1.018979e-08, 9.669185e-09, 8.424617e-09, 7.952853e-09, 8.263136e-09,
  1.110044e-08, 1.156573e-08, 1.26465e-08, 1.43236e-08, 1.390083e-08, 
    1.105674e-08, 7.099023e-09, 6.341782e-09, 8.32818e-09, 1.095206e-08, 
    1.061145e-08, 9.54426e-09, 8.544019e-09, 7.847378e-09, 8.262364e-09,
  1.124902e-08, 1.151504e-08, 1.200456e-08, 1.288626e-08, 1.402913e-08, 
    1.337285e-08, 9.820232e-09, 6.808745e-09, 7.321568e-09, 9.83994e-09, 
    1.132098e-08, 9.583064e-09, 8.497531e-09, 7.842102e-09, 8.18341e-09,
  1.138571e-08, 1.173089e-08, 1.194715e-08, 1.226532e-08, 1.282024e-08, 
    1.388504e-08, 1.216169e-08, 8.65008e-09, 7.140709e-09, 8.402509e-09, 
    1.134878e-08, 9.983013e-09, 8.401621e-09, 7.938284e-09, 8.064992e-09,
  1.166233e-08, 1.186093e-08, 1.215875e-08, 1.228544e-08, 1.249793e-08, 
    1.297279e-08, 1.343346e-08, 1.078825e-08, 8.012164e-09, 7.921986e-09, 
    1.064036e-08, 1.043563e-08, 8.491904e-09, 7.971741e-09, 8.050369e-09,
  1.267783e-08, 1.267101e-08, 1.266908e-08, 1.280089e-08, 1.268419e-08, 
    1.269258e-08, 1.302794e-08, 1.238405e-08, 9.68603e-09, 7.970589e-09, 
    9.522177e-09, 1.103191e-08, 8.665799e-09, 7.970518e-09, 8.038795e-09,
  1.422257e-08, 1.39062e-08, 1.383119e-08, 1.38914e-08, 1.390548e-08, 
    1.336987e-08, 1.296015e-08, 1.263358e-08, 1.118703e-08, 9.009137e-09, 
    8.818232e-09, 1.110398e-08, 9.263943e-09, 8.02279e-09, 8.045132e-09,
  6.34512e-09, 5.7489e-09, 5.54943e-09, 5.870207e-09, 7.492385e-09, 
    1.000489e-08, 9.940452e-09, 8.911421e-09, 9.204141e-09, 9.839345e-09, 
    1.044974e-08, 1.092457e-08, 1.118105e-08, 1.126552e-08, 1.122313e-08,
  7.13503e-09, 6.508951e-09, 6.058327e-09, 5.764723e-09, 6.257463e-09, 
    8.639242e-09, 1.020069e-08, 9.368061e-09, 8.774378e-09, 9.395989e-09, 
    9.999756e-09, 1.058223e-08, 1.090535e-08, 1.092742e-08, 1.094121e-08,
  7.994484e-09, 7.273e-09, 6.934513e-09, 6.432139e-09, 6.055912e-09, 
    6.731964e-09, 9.390936e-09, 1.007904e-08, 9.033171e-09, 8.841811e-09, 
    9.589399e-09, 1.018e-08, 1.057602e-08, 1.080615e-08, 1.075398e-08,
  8.968559e-09, 8.143576e-09, 7.760701e-09, 7.398355e-09, 6.909288e-09, 
    6.330364e-09, 7.281503e-09, 1.025974e-08, 9.340504e-09, 8.834321e-09, 
    9.16749e-09, 9.659235e-09, 1.031617e-08, 1.072921e-08, 1.053122e-08,
  9.93755e-09, 8.953504e-09, 8.742536e-09, 8.47739e-09, 7.983298e-09, 
    7.165716e-09, 6.477868e-09, 8.865765e-09, 1.015444e-08, 9.009923e-09, 
    8.685691e-09, 9.381252e-09, 1.004219e-08, 1.054409e-08, 1.041077e-08,
  1.078671e-08, 9.701362e-09, 9.291421e-09, 9.470511e-09, 9.221289e-09, 
    8.609267e-09, 7.085094e-09, 7.103045e-09, 9.660909e-09, 9.303728e-09, 
    8.638503e-09, 9.129161e-09, 9.775743e-09, 1.024308e-08, 1.034823e-08,
  1.171714e-08, 1.037951e-08, 9.79761e-09, 9.851749e-09, 1.003684e-08, 
    1.003797e-08, 8.734002e-09, 7.11793e-09, 8.434543e-09, 9.740899e-09, 
    8.919686e-09, 8.783649e-09, 9.408662e-09, 1.003663e-08, 1.048551e-08,
  1.250971e-08, 1.10149e-08, 1.014684e-08, 1.008429e-08, 1.025932e-08, 
    1.08223e-08, 1.05728e-08, 8.465951e-09, 7.532502e-09, 9.243085e-09, 
    9.211763e-09, 8.58603e-09, 9.224551e-09, 1.007409e-08, 1.055538e-08,
  1.346434e-08, 1.161912e-08, 1.042422e-08, 1.01127e-08, 1.017911e-08, 
    1.07945e-08, 1.15689e-08, 1.059999e-08, 8.227962e-09, 8.539058e-09, 
    9.476283e-09, 8.629092e-09, 8.905264e-09, 1.006864e-08, 1.071495e-08,
  1.414071e-08, 1.237848e-08, 1.078638e-08, 1.014636e-08, 1.005753e-08, 
    1.038476e-08, 1.167181e-08, 1.207778e-08, 9.792593e-09, 8.326904e-09, 
    9.227398e-09, 8.816761e-09, 8.779753e-09, 1.002206e-08, 1.090672e-08,
  1.215311e-08, 1.167107e-08, 1.262437e-08, 1.061505e-08, 8.07411e-09, 
    9.474422e-09, 9.256116e-09, 1.058524e-08, 1.159573e-08, 1.163411e-08, 
    1.154176e-08, 1.092068e-08, 1.00344e-08, 9.594693e-09, 9.122826e-09,
  1.249282e-08, 1.165065e-08, 1.188506e-08, 1.193467e-08, 8.575119e-09, 
    8.75843e-09, 9.272442e-09, 9.517652e-09, 1.130728e-08, 1.178986e-08, 
    1.156316e-08, 1.117061e-08, 1.052422e-08, 9.957726e-09, 9.551631e-09,
  1.286159e-08, 1.208463e-08, 1.164432e-08, 1.23386e-08, 9.891501e-09, 
    7.794699e-09, 9.472187e-09, 8.798661e-09, 1.058278e-08, 1.143744e-08, 
    1.175129e-08, 1.129956e-08, 1.07676e-08, 1.019031e-08, 9.784733e-09,
  1.339456e-08, 1.250277e-08, 1.178816e-08, 1.196385e-08, 1.130068e-08, 
    7.619459e-09, 8.71982e-09, 9.144891e-09, 9.278018e-09, 1.113764e-08, 
    1.169518e-08, 1.147292e-08, 1.098985e-08, 1.038702e-08, 9.99907e-09,
  1.375129e-08, 1.316642e-08, 1.223491e-08, 1.191361e-08, 1.232685e-08, 
    8.929724e-09, 7.181796e-09, 9.462855e-09, 9.124184e-09, 1.046613e-08, 
    1.122287e-08, 1.163827e-08, 1.09974e-08, 1.055497e-08, 9.943104e-09,
  1.402008e-08, 1.385805e-08, 1.301057e-08, 1.2199e-08, 1.237209e-08, 
    1.061099e-08, 6.965885e-09, 8.676188e-09, 9.200575e-09, 9.459918e-09, 
    1.071787e-08, 1.134274e-08, 1.111314e-08, 1.055206e-08, 1.001481e-08,
  1.429991e-08, 1.43579e-08, 1.383412e-08, 1.287194e-08, 1.234504e-08, 
    1.196053e-08, 8.314025e-09, 7.228863e-09, 9.110023e-09, 9.187409e-09, 
    1.033626e-08, 1.105468e-08, 1.13349e-08, 1.053503e-08, 1.02751e-08,
  1.464113e-08, 1.496504e-08, 1.451823e-08, 1.374283e-08, 1.271426e-08, 
    1.251323e-08, 1.002427e-08, 6.977653e-09, 8.471116e-09, 9.086628e-09, 
    9.723848e-09, 1.067125e-08, 1.117286e-08, 1.075423e-08, 1.023466e-08,
  1.490755e-08, 1.540235e-08, 1.526604e-08, 1.465247e-08, 1.346028e-08, 
    1.279734e-08, 1.132978e-08, 7.934474e-09, 7.65113e-09, 8.870331e-09, 
    9.433673e-09, 1.035898e-08, 1.094862e-08, 1.090594e-08, 1.039031e-08,
  1.535167e-08, 1.588575e-08, 1.595156e-08, 1.553268e-08, 1.445629e-08, 
    1.319519e-08, 1.237211e-08, 9.296529e-09, 7.199506e-09, 8.594092e-09, 
    9.212525e-09, 9.968089e-09, 1.070706e-08, 1.093056e-08, 1.047989e-08,
  1.161868e-08, 1.209612e-08, 1.219313e-08, 1.133642e-08, 9.912814e-09, 
    9.65017e-09, 9.528972e-09, 8.71621e-09, 8.733519e-09, 9.060433e-09, 
    9.452538e-09, 9.77914e-09, 9.953998e-09, 1.019939e-08, 1.072165e-08,
  1.099717e-08, 1.18302e-08, 1.24867e-08, 1.272268e-08, 1.100043e-08, 
    9.688026e-09, 9.987551e-09, 9.355176e-09, 8.774201e-09, 9.084101e-09, 
    9.613171e-09, 1.003385e-08, 1.026806e-08, 1.038685e-08, 1.070934e-08,
  1.021268e-08, 1.154153e-08, 1.209845e-08, 1.316204e-08, 1.297108e-08, 
    9.990143e-09, 9.839179e-09, 1.004099e-08, 9.134711e-09, 9.052316e-09, 
    9.586705e-09, 1.040434e-08, 1.065955e-08, 1.072411e-08, 1.090042e-08,
  9.015363e-09, 1.076137e-08, 1.177358e-08, 1.283743e-08, 1.41278e-08, 
    1.246503e-08, 9.786203e-09, 1.040791e-08, 9.762295e-09, 9.068705e-09, 
    9.464952e-09, 1.034873e-08, 1.091959e-08, 1.11242e-08, 1.111671e-08,
  7.731873e-09, 9.579042e-09, 1.091796e-08, 1.217294e-08, 1.345334e-08, 
    1.453198e-08, 1.035655e-08, 9.900488e-09, 1.052776e-08, 9.624941e-09, 
    9.273704e-09, 1.003367e-08, 1.088829e-08, 1.135197e-08, 1.127871e-08,
  6.37093e-09, 8.17219e-09, 9.740273e-09, 1.124292e-08, 1.295773e-08, 
    1.536187e-08, 1.405937e-08, 9.591362e-09, 1.057614e-08, 1.010735e-08, 
    9.273618e-09, 9.637061e-09, 1.053997e-08, 1.115625e-08, 1.126256e-08,
  5.220715e-09, 6.793779e-09, 8.292888e-09, 9.657511e-09, 1.145837e-08, 
    1.397311e-08, 1.621682e-08, 1.154544e-08, 9.933455e-09, 1.052734e-08, 
    9.721703e-09, 9.834379e-09, 1.021318e-08, 1.088076e-08, 1.108753e-08,
  4.724737e-09, 5.838874e-09, 7.273172e-09, 8.349732e-09, 9.877932e-09, 
    1.208225e-08, 1.581487e-08, 1.547067e-08, 1.012757e-08, 1.049884e-08, 
    1.000992e-08, 9.753986e-09, 1.000058e-08, 1.044974e-08, 1.038813e-08,
  4.624263e-09, 5.395848e-09, 6.679403e-09, 7.638405e-09, 8.514432e-09, 
    1.008651e-08, 1.346023e-08, 1.693365e-08, 1.280984e-08, 1.00885e-08, 
    1.057459e-08, 9.932354e-09, 1.002617e-08, 9.799958e-09, 9.515136e-09,
  4.643509e-09, 5.483353e-09, 6.555937e-09, 7.518123e-09, 7.90792e-09, 
    8.728096e-09, 1.063644e-08, 1.542586e-08, 1.59437e-08, 1.127234e-08, 
    1.063187e-08, 1.007974e-08, 9.930196e-09, 9.281626e-09, 8.720589e-09,
  9.944768e-09, 1.020387e-08, 1.046789e-08, 1.086549e-08, 1.12689e-08, 
    1.169968e-08, 1.232009e-08, 1.302205e-08, 1.337678e-08, 1.365091e-08, 
    1.3872e-08, 1.387911e-08, 1.362953e-08, 1.34776e-08, 1.300065e-08,
  9.94152e-09, 1.017249e-08, 1.051281e-08, 1.078134e-08, 1.092186e-08, 
    1.14471e-08, 1.206383e-08, 1.271044e-08, 1.332798e-08, 1.363311e-08, 
    1.37564e-08, 1.387897e-08, 1.385937e-08, 1.371674e-08, 1.337851e-08,
  1.000297e-08, 1.019825e-08, 1.049688e-08, 1.066857e-08, 1.084332e-08, 
    1.115432e-08, 1.163449e-08, 1.235303e-08, 1.305421e-08, 1.327304e-08, 
    1.348722e-08, 1.35891e-08, 1.381718e-08, 1.383032e-08, 1.363754e-08,
  1.035007e-08, 1.031224e-08, 1.034317e-08, 1.041539e-08, 1.05963e-08, 
    1.093078e-08, 1.129497e-08, 1.17664e-08, 1.23957e-08, 1.304086e-08, 
    1.343484e-08, 1.372496e-08, 1.371059e-08, 1.360944e-08, 1.342178e-08,
  1.087747e-08, 1.067804e-08, 1.0476e-08, 1.037577e-08, 1.038941e-08, 
    1.066662e-08, 1.112469e-08, 1.153426e-08, 1.185444e-08, 1.2514e-08, 
    1.308906e-08, 1.349382e-08, 1.365184e-08, 1.3651e-08, 1.355493e-08,
  1.159708e-08, 1.139472e-08, 1.117226e-08, 1.082981e-08, 1.052025e-08, 
    1.044789e-08, 1.076193e-08, 1.127386e-08, 1.164163e-08, 1.190736e-08, 
    1.256833e-08, 1.315077e-08, 1.358153e-08, 1.369009e-08, 1.330814e-08,
  1.146308e-08, 1.147095e-08, 1.155628e-08, 1.1417e-08, 1.123021e-08, 
    1.099621e-08, 1.062819e-08, 1.075457e-08, 1.133272e-08, 1.177777e-08, 
    1.206236e-08, 1.276008e-08, 1.327874e-08, 1.324341e-08, 1.289281e-08,
  1.075201e-08, 1.075672e-08, 1.094955e-08, 1.131051e-08, 1.167696e-08, 
    1.154549e-08, 1.120387e-08, 1.078888e-08, 1.085594e-08, 1.13975e-08, 
    1.182427e-08, 1.204531e-08, 1.258612e-08, 1.273319e-08, 1.227057e-08,
  1.006626e-08, 1.001983e-08, 1.019096e-08, 1.043712e-08, 1.089657e-08, 
    1.140772e-08, 1.161531e-08, 1.146408e-08, 1.090644e-08, 1.103659e-08, 
    1.145021e-08, 1.169721e-08, 1.203334e-08, 1.227148e-08, 1.185437e-08,
  9.471707e-09, 9.46206e-09, 9.473741e-09, 9.593026e-09, 9.99843e-09, 
    1.038732e-08, 1.11755e-08, 1.14354e-08, 1.140005e-08, 1.091579e-08, 
    1.104025e-08, 1.144049e-08, 1.145865e-08, 1.162913e-08, 1.137882e-08,
  1.351252e-08, 1.373923e-08, 1.404002e-08, 1.433144e-08, 1.387083e-08, 
    1.357246e-08, 1.319351e-08, 1.271551e-08, 1.208062e-08, 1.18203e-08, 
    1.15184e-08, 1.109051e-08, 1.053915e-08, 1.01546e-08, 9.774909e-09,
  1.332836e-08, 1.363923e-08, 1.375369e-08, 1.398623e-08, 1.386566e-08, 
    1.383514e-08, 1.369481e-08, 1.355283e-08, 1.308764e-08, 1.242697e-08, 
    1.202315e-08, 1.154475e-08, 1.103869e-08, 1.071511e-08, 1.025664e-08,
  1.295237e-08, 1.319801e-08, 1.330778e-08, 1.358025e-08, 1.36595e-08, 
    1.387596e-08, 1.433018e-08, 1.427044e-08, 1.416967e-08, 1.358001e-08, 
    1.289065e-08, 1.236755e-08, 1.177754e-08, 1.125638e-08, 1.095223e-08,
  1.260019e-08, 1.276368e-08, 1.282273e-08, 1.304205e-08, 1.333242e-08, 
    1.376106e-08, 1.394466e-08, 1.460465e-08, 1.451424e-08, 1.410034e-08, 
    1.360101e-08, 1.306241e-08, 1.254762e-08, 1.21069e-08, 1.138363e-08,
  1.223741e-08, 1.235258e-08, 1.237239e-08, 1.255853e-08, 1.288689e-08, 
    1.327999e-08, 1.374456e-08, 1.413986e-08, 1.510058e-08, 1.510555e-08, 
    1.442086e-08, 1.365473e-08, 1.312788e-08, 1.258331e-08, 1.241068e-08,
  1.189073e-08, 1.192762e-08, 1.188735e-08, 1.202463e-08, 1.252051e-08, 
    1.295896e-08, 1.328356e-08, 1.358369e-08, 1.424858e-08, 1.481611e-08, 
    1.488078e-08, 1.45092e-08, 1.385527e-08, 1.289354e-08, 1.227967e-08,
  1.15543e-08, 1.15814e-08, 1.151719e-08, 1.163473e-08, 1.212547e-08, 
    1.255888e-08, 1.284397e-08, 1.302622e-08, 1.345602e-08, 1.403464e-08, 
    1.445102e-08, 1.442239e-08, 1.429322e-08, 1.365895e-08, 1.278274e-08,
  1.128769e-08, 1.127953e-08, 1.122476e-08, 1.127632e-08, 1.179727e-08, 
    1.210675e-08, 1.244932e-08, 1.266842e-08, 1.299067e-08, 1.347314e-08, 
    1.409722e-08, 1.436271e-08, 1.426525e-08, 1.376137e-08, 1.304333e-08,
  1.109674e-08, 1.105015e-08, 1.103657e-08, 1.101867e-08, 1.143238e-08, 
    1.178749e-08, 1.212586e-08, 1.241456e-08, 1.278357e-08, 1.304384e-08, 
    1.351514e-08, 1.390195e-08, 1.40977e-08, 1.363766e-08, 1.293102e-08,
  1.089771e-08, 1.087192e-08, 1.084006e-08, 1.083486e-08, 1.121161e-08, 
    1.156117e-08, 1.193721e-08, 1.215508e-08, 1.252703e-08, 1.275159e-08, 
    1.323584e-08, 1.386289e-08, 1.39911e-08, 1.342618e-08, 1.255154e-08,
  1.249607e-08, 1.1571e-08, 1.040488e-08, 1.001932e-08, 9.750242e-09, 
    9.838727e-09, 9.750736e-09, 9.445601e-09, 8.732999e-09, 8.173999e-09, 
    7.525351e-09, 6.893434e-09, 6.432255e-09, 5.881899e-09, 5.484156e-09,
  1.248914e-08, 1.257082e-08, 1.165972e-08, 1.057225e-08, 1.007607e-08, 
    9.887842e-09, 9.94532e-09, 1.006336e-08, 1.013316e-08, 9.428517e-09, 
    8.888662e-09, 7.809125e-09, 7.187798e-09, 6.365948e-09, 5.921019e-09,
  1.278562e-08, 1.260211e-08, 1.250279e-08, 1.191131e-08, 1.122951e-08, 
    1.058282e-08, 1.0339e-08, 1.044707e-08, 1.099522e-08, 1.124726e-08, 
    1.079378e-08, 9.563053e-09, 8.30628e-09, 7.219223e-09, 6.291228e-09,
  1.401064e-08, 1.262295e-08, 1.26604e-08, 1.273117e-08, 1.262353e-08, 
    1.262816e-08, 1.194785e-08, 1.117157e-08, 1.132604e-08, 1.167458e-08, 
    1.286329e-08, 1.197147e-08, 1.010433e-08, 8.541203e-09, 6.995804e-09,
  1.534523e-08, 1.334683e-08, 1.257387e-08, 1.283328e-08, 1.320419e-08, 
    1.358105e-08, 1.380865e-08, 1.336545e-08, 1.287734e-08, 1.243385e-08, 
    1.238172e-08, 1.316945e-08, 1.233058e-08, 1.012226e-08, 8.12961e-09,
  1.607894e-08, 1.438619e-08, 1.326923e-08, 1.289959e-08, 1.328213e-08, 
    1.369339e-08, 1.392569e-08, 1.387935e-08, 1.386208e-08, 1.370443e-08, 
    1.265346e-08, 1.264245e-08, 1.271574e-08, 1.161888e-08, 9.126538e-09,
  1.72534e-08, 1.495825e-08, 1.390123e-08, 1.339008e-08, 1.346169e-08, 
    1.369332e-08, 1.362248e-08, 1.377561e-08, 1.392292e-08, 1.457877e-08, 
    1.367233e-08, 1.253904e-08, 1.265768e-08, 1.204426e-08, 1.02988e-08,
  1.877852e-08, 1.632845e-08, 1.453199e-08, 1.396665e-08, 1.38158e-08, 
    1.380675e-08, 1.366895e-08, 1.372617e-08, 1.391145e-08, 1.470335e-08, 
    1.483654e-08, 1.334224e-08, 1.268622e-08, 1.192115e-08, 1.075079e-08,
  1.909775e-08, 1.761723e-08, 1.541312e-08, 1.441491e-08, 1.423933e-08, 
    1.388517e-08, 1.376818e-08, 1.356769e-08, 1.38201e-08, 1.450005e-08, 
    1.51103e-08, 1.397836e-08, 1.277454e-08, 1.179595e-08, 1.071503e-08,
  1.853378e-08, 1.830843e-08, 1.676302e-08, 1.496091e-08, 1.441548e-08, 
    1.392262e-08, 1.37229e-08, 1.347094e-08, 1.368291e-08, 1.430624e-08, 
    1.527882e-08, 1.433038e-08, 1.272096e-08, 1.139844e-08, 1.056189e-08,
  1.110481e-08, 9.715318e-09, 7.724287e-09, 6.421451e-09, 5.471677e-09, 
    4.740761e-09, 4.034209e-09, 3.644985e-09, 3.368065e-09, 3.324184e-09, 
    3.319133e-09, 3.312046e-09, 2.993089e-09, 2.668196e-09, 2.447403e-09,
  1.356731e-08, 1.218798e-08, 1.052417e-08, 8.740393e-09, 7.113414e-09, 
    6.004986e-09, 5.099882e-09, 4.448212e-09, 3.912409e-09, 3.634198e-09, 
    3.578119e-09, 3.565946e-09, 3.351847e-09, 2.973669e-09, 2.888847e-09,
  1.704961e-08, 1.506656e-08, 1.339094e-08, 1.183195e-08, 1.011765e-08, 
    8.36135e-09, 6.861175e-09, 5.793109e-09, 5.074477e-09, 4.543473e-09, 
    4.289087e-09, 3.954197e-09, 3.791682e-09, 3.412087e-09, 3.284092e-09,
  1.893474e-08, 1.763698e-08, 1.607694e-08, 1.439088e-08, 1.284722e-08, 
    1.142296e-08, 9.941202e-09, 8.38169e-09, 7.054313e-09, 6.097618e-09, 
    5.429341e-09, 4.993742e-09, 4.273323e-09, 3.779817e-09, 3.531023e-09,
  2.140131e-08, 2.147787e-08, 1.982401e-08, 1.748405e-08, 1.54367e-08, 
    1.376743e-08, 1.247774e-08, 1.145071e-08, 1.011865e-08, 9.041953e-09, 
    7.957682e-09, 7.238055e-09, 6.735394e-09, 5.417926e-09, 4.518467e-09,
  2.133561e-08, 2.306196e-08, 2.331068e-08, 2.125186e-08, 1.853259e-08, 
    1.61593e-08, 1.425427e-08, 1.311449e-08, 1.22966e-08, 1.143494e-08, 
    9.948953e-09, 8.96394e-09, 8.057357e-09, 7.70804e-09, 6.350579e-09,
  1.897821e-08, 2.205779e-08, 2.453493e-08, 2.425361e-08, 2.188795e-08, 
    1.916601e-08, 1.631833e-08, 1.415239e-08, 1.278995e-08, 1.213985e-08, 
    1.112464e-08, 9.996104e-09, 9.309637e-09, 8.762855e-09, 8.236375e-09,
  1.587992e-08, 1.966134e-08, 2.314551e-08, 2.421636e-08, 2.354966e-08, 
    2.212013e-08, 1.973899e-08, 1.674651e-08, 1.399789e-08, 1.252939e-08, 
    1.165309e-08, 1.077109e-08, 1.060357e-08, 1.028079e-08, 9.200512e-09,
  1.275799e-08, 1.672459e-08, 2.063434e-08, 2.24303e-08, 2.215198e-08, 
    2.143269e-08, 2.117925e-08, 1.962691e-08, 1.66876e-08, 1.382706e-08, 
    1.255115e-08, 1.180031e-08, 1.144533e-08, 1.137726e-08, 1.052397e-08,
  9.802809e-09, 1.37766e-08, 1.916426e-08, 2.166354e-08, 2.165245e-08, 
    1.964942e-08, 1.91421e-08, 1.941092e-08, 1.832541e-08, 1.609145e-08, 
    1.347122e-08, 1.265912e-08, 1.21575e-08, 1.196019e-08, 1.126071e-08,
  6.270447e-09, 5.342283e-09, 4.993634e-09, 4.589491e-09, 4.35765e-09, 
    4.11708e-09, 3.906889e-09, 3.615137e-09, 3.518793e-09, 3.548246e-09, 
    3.52525e-09, 3.6018e-09, 3.256247e-09, 3.052014e-09, 3.004141e-09,
  6.56691e-09, 5.453165e-09, 4.921268e-09, 4.490845e-09, 4.233474e-09, 
    3.935684e-09, 3.693242e-09, 3.376379e-09, 3.103199e-09, 3.035755e-09, 
    2.992835e-09, 3.286328e-09, 3.257579e-09, 3.161265e-09, 3.181481e-09,
  8.55179e-09, 7.948815e-09, 7.041165e-09, 5.987347e-09, 4.95206e-09, 
    4.258195e-09, 3.860662e-09, 3.570366e-09, 3.249201e-09, 2.98381e-09, 
    2.736927e-09, 2.737978e-09, 3.145346e-09, 3.504989e-09, 3.448449e-09,
  1.026601e-08, 1.063267e-08, 1.098124e-08, 1.055641e-08, 9.591867e-09, 
    7.827534e-09, 5.968732e-09, 4.460308e-09, 3.662451e-09, 3.225106e-09, 
    2.969603e-09, 2.726184e-09, 2.886708e-09, 3.486528e-09, 3.741942e-09,
  1.06684e-08, 1.174119e-08, 1.293426e-08, 1.41334e-08, 1.457151e-08, 
    1.417115e-08, 1.250177e-08, 9.873027e-09, 6.751345e-09, 4.391309e-09, 
    3.286301e-09, 2.973011e-09, 2.93286e-09, 3.396206e-09, 3.791846e-09,
  9.565038e-09, 1.010209e-08, 1.184482e-08, 1.475892e-08, 1.758929e-08, 
    1.950646e-08, 2.014612e-08, 1.865322e-08, 1.539868e-08, 1.07501e-08, 
    6.157845e-09, 3.533085e-09, 3.079686e-09, 3.34256e-09, 3.945766e-09,
  8.863134e-09, 9.536499e-09, 1.142217e-08, 1.473273e-08, 1.885688e-08, 
    2.183219e-08, 2.32534e-08, 2.361944e-08, 2.193889e-08, 1.872914e-08, 
    1.337961e-08, 7.339033e-09, 3.776963e-09, 3.461556e-09, 3.959841e-09,
  8.674376e-09, 9.377571e-09, 1.063547e-08, 1.331569e-08, 1.773007e-08, 
    1.9496e-08, 2.03732e-08, 2.10891e-08, 2.185948e-08, 2.193532e-08, 
    1.961164e-08, 1.245154e-08, 6.397169e-09, 4.009119e-09, 4.111167e-09,
  9.453218e-09, 1.012462e-08, 1.0465e-08, 1.180408e-08, 1.607675e-08, 
    1.772417e-08, 1.82446e-08, 1.945758e-08, 2.113411e-08, 2.260192e-08, 
    2.326987e-08, 1.78667e-08, 9.804585e-09, 5.006799e-09, 4.443326e-09,
  9.965643e-09, 1.031137e-08, 1.026179e-08, 1.116195e-08, 1.469894e-08, 
    1.655647e-08, 1.650927e-08, 1.733567e-08, 1.996439e-08, 2.199147e-08, 
    2.461723e-08, 2.155512e-08, 1.367631e-08, 6.427233e-09, 4.883635e-09,
  1.482213e-08, 1.449601e-08, 1.427772e-08, 1.295006e-08, 1.141651e-08, 
    1.048415e-08, 1.022544e-08, 9.537184e-09, 9.030249e-09, 8.040288e-09, 
    7.828272e-09, 7.935242e-09, 7.497721e-09, 6.579235e-09, 5.857772e-09,
  1.459977e-08, 1.425373e-08, 1.396776e-08, 1.282173e-08, 1.114207e-08, 
    9.894483e-09, 9.14883e-09, 8.494766e-09, 8.009489e-09, 7.637869e-09, 
    7.299419e-09, 7.098889e-09, 6.714585e-09, 5.891738e-09, 5.441927e-09,
  1.438178e-08, 1.374707e-08, 1.310899e-08, 1.185711e-08, 1.043972e-08, 
    9.186095e-09, 8.296982e-09, 7.752829e-09, 7.323327e-09, 7.169507e-09, 
    6.914191e-09, 6.62781e-09, 6.357682e-09, 5.565779e-09, 5.164544e-09,
  1.395401e-08, 1.327075e-08, 1.208756e-08, 1.049691e-08, 9.287027e-09, 
    8.227006e-09, 7.417129e-09, 6.782982e-09, 6.44096e-09, 6.249659e-09, 
    6.142928e-09, 6.056278e-09, 5.772681e-09, 5.322959e-09, 5.114729e-09,
  1.280057e-08, 1.206663e-08, 1.046042e-08, 8.927855e-09, 7.81037e-09, 
    7.41213e-09, 7.05659e-09, 6.622699e-09, 5.981311e-09, 5.422824e-09, 
    5.111562e-09, 5.455862e-09, 5.248172e-09, 4.871246e-09, 4.742779e-09,
  1.151587e-08, 1.074943e-08, 9.483526e-09, 8.379798e-09, 8.322474e-09, 
    8.836782e-09, 9.731424e-09, 1.016252e-08, 1.008257e-08, 8.999427e-09, 
    6.53511e-09, 4.972134e-09, 4.668509e-09, 4.468608e-09, 4.378009e-09,
  1.070931e-08, 1.011262e-08, 9.547418e-09, 9.303026e-09, 9.976199e-09, 
    1.129219e-08, 1.267628e-08, 1.410936e-08, 1.503474e-08, 1.49649e-08, 
    1.445622e-08, 9.466157e-09, 4.987446e-09, 4.029786e-09, 3.987377e-09,
  1.044634e-08, 1.003461e-08, 9.574999e-09, 9.806699e-09, 1.054506e-08, 
    1.214427e-08, 1.300787e-08, 1.329004e-08, 1.414623e-08, 1.454325e-08, 
    1.669971e-08, 1.670175e-08, 8.999281e-09, 4.357335e-09, 3.548347e-09,
  1.04138e-08, 1.005755e-08, 9.67173e-09, 1.009512e-08, 1.101079e-08, 
    1.260256e-08, 1.283564e-08, 1.319004e-08, 1.383835e-08, 1.48147e-08, 
    1.533503e-08, 2.025219e-08, 1.467851e-08, 6.747935e-09, 3.456437e-09,
  1.054599e-08, 1.008277e-08, 9.956945e-09, 1.044404e-08, 1.187149e-08, 
    1.297958e-08, 1.290411e-08, 1.325665e-08, 1.393979e-08, 1.584898e-08, 
    1.638008e-08, 2.072622e-08, 1.915908e-08, 9.451536e-09, 3.963246e-09,
  1.391679e-08, 1.536103e-08, 1.642012e-08, 1.450984e-08, 1.324043e-08, 
    1.256586e-08, 1.188798e-08, 1.172338e-08, 1.164397e-08, 1.122982e-08, 
    1.167577e-08, 1.18334e-08, 1.205699e-08, 1.19155e-08, 1.12478e-08,
  1.3021e-08, 1.495232e-08, 1.644679e-08, 1.524572e-08, 1.270566e-08, 
    1.222319e-08, 1.176553e-08, 1.083928e-08, 1.097658e-08, 1.078232e-08, 
    1.081932e-08, 1.097577e-08, 1.059371e-08, 9.399009e-09, 8.73483e-09,
  1.151591e-08, 1.426051e-08, 1.596917e-08, 1.537448e-08, 1.238319e-08, 
    1.117876e-08, 1.081432e-08, 9.856531e-09, 9.573325e-09, 9.83302e-09, 
    9.832034e-09, 9.563862e-09, 8.328703e-09, 7.451338e-09, 7.529888e-09,
  1.087578e-08, 1.329487e-08, 1.544099e-08, 1.55667e-08, 1.253055e-08, 
    1.015737e-08, 1.008386e-08, 9.629596e-09, 8.435515e-09, 8.70078e-09, 
    8.825785e-09, 8.077488e-09, 7.203371e-09, 6.93937e-09, 7.363042e-09,
  1.039357e-08, 1.242695e-08, 1.449667e-08, 1.500874e-08, 1.26079e-08, 
    1.017682e-08, 8.662946e-09, 8.832288e-09, 8.376388e-09, 7.678713e-09, 
    7.81723e-09, 7.369217e-09, 6.80746e-09, 6.560045e-09, 7.093968e-09,
  1.032604e-08, 1.194298e-08, 1.370759e-08, 1.464184e-08, 1.291132e-08, 
    1.074041e-08, 9.040122e-09, 8.146493e-09, 7.785806e-09, 7.444086e-09, 
    7.179433e-09, 6.85767e-09, 6.46802e-09, 6.137078e-09, 5.979016e-09,
  1.030217e-08, 1.159664e-08, 1.294565e-08, 1.370898e-08, 1.285556e-08, 
    1.139388e-08, 1.018392e-08, 1.02077e-08, 8.257805e-09, 7.376386e-09, 
    6.804943e-09, 6.502704e-09, 6.025873e-09, 5.423071e-09, 4.925121e-09,
  1.035187e-08, 1.137213e-08, 1.249389e-08, 1.319397e-08, 1.270853e-08, 
    1.179615e-08, 1.14246e-08, 1.118863e-08, 1.103597e-08, 8.711901e-09, 
    7.21117e-09, 6.32441e-09, 5.693033e-09, 5.002081e-09, 4.271413e-09,
  1.04176e-08, 1.126095e-08, 1.215465e-08, 1.256262e-08, 1.250611e-08, 
    1.216739e-08, 1.181377e-08, 1.186787e-08, 1.264343e-08, 1.124636e-08, 
    8.512883e-09, 6.913842e-09, 5.557802e-09, 4.675353e-09, 3.933125e-09,
  1.051597e-08, 1.123705e-08, 1.188706e-08, 1.216013e-08, 1.252311e-08, 
    1.236549e-08, 1.211048e-08, 1.254595e-08, 1.268023e-08, 1.341156e-08, 
    1.065798e-08, 8.140648e-09, 5.973478e-09, 4.645847e-09, 3.874807e-09,
  1.142785e-08, 1.172432e-08, 1.103096e-08, 9.965851e-09, 9.127549e-09, 
    9.603786e-09, 1.083964e-08, 1.159278e-08, 1.249749e-08, 1.345407e-08, 
    1.476089e-08, 1.636591e-08, 1.79356e-08, 1.848085e-08, 1.579823e-08,
  1.095419e-08, 1.216748e-08, 1.234514e-08, 1.131521e-08, 9.636303e-09, 
    8.789967e-09, 9.709101e-09, 1.078624e-08, 1.166956e-08, 1.250265e-08, 
    1.339977e-08, 1.449202e-08, 1.538765e-08, 1.60326e-08, 1.532447e-08,
  8.961317e-09, 1.123308e-08, 1.252924e-08, 1.218065e-08, 1.117283e-08, 
    9.156095e-09, 8.940465e-09, 9.869371e-09, 1.068766e-08, 1.132814e-08, 
    1.191044e-08, 1.270847e-08, 1.342144e-08, 1.374594e-08, 1.352866e-08,
  7.194816e-09, 9.145927e-09, 1.186474e-08, 1.26315e-08, 1.198476e-08, 
    1.0737e-08, 8.755972e-09, 9.236852e-09, 9.952861e-09, 1.070688e-08, 
    1.134341e-08, 1.204565e-08, 1.243142e-08, 1.276133e-08, 1.271051e-08,
  6.094422e-09, 7.064379e-09, 9.840925e-09, 1.214494e-08, 1.27654e-08, 
    1.20223e-08, 1.009975e-08, 8.784556e-09, 9.372803e-09, 9.900285e-09, 
    1.05082e-08, 1.083409e-08, 1.0957e-08, 1.093841e-08, 1.089898e-08,
  5.765719e-09, 6.079265e-09, 7.35498e-09, 1.062773e-08, 1.257905e-08, 
    1.270187e-08, 1.201655e-08, 9.372862e-09, 8.913711e-09, 9.352521e-09, 
    9.711646e-09, 9.651416e-09, 9.344717e-09, 8.950286e-09, 8.926429e-09,
  5.539883e-09, 5.756013e-09, 6.168891e-09, 8.387232e-09, 1.155813e-08, 
    1.292653e-08, 1.289535e-08, 1.123781e-08, 8.694976e-09, 8.840503e-09, 
    8.794782e-09, 8.424309e-09, 7.758223e-09, 7.120796e-09, 6.93831e-09,
  4.831032e-09, 5.465765e-09, 5.584629e-09, 6.663676e-09, 9.954526e-09, 
    1.206854e-08, 1.346922e-08, 1.302806e-08, 9.516027e-09, 8.398866e-09, 
    8.026327e-09, 7.226852e-09, 6.153703e-09, 5.440084e-09, 5.1318e-09,
  3.9845e-09, 4.614757e-09, 5.267251e-09, 5.89778e-09, 8.523299e-09, 
    1.123734e-08, 1.325345e-08, 1.452917e-08, 1.124354e-08, 8.721083e-09, 
    7.326662e-09, 6.002874e-09, 4.690986e-09, 4.169921e-09, 3.932529e-09,
  3.647416e-09, 3.59215e-09, 4.367332e-09, 5.502771e-09, 7.610033e-09, 
    1.033676e-08, 1.346458e-08, 1.745724e-08, 1.349352e-08, 9.340142e-09, 
    6.809734e-09, 5.072613e-09, 3.790282e-09, 3.409367e-09, 3.203538e-09,
  9.911061e-09, 1.064095e-08, 1.129915e-08, 1.22253e-08, 1.335021e-08, 
    1.463359e-08, 1.617951e-08, 1.772625e-08, 1.895285e-08, 1.899006e-08, 
    1.742932e-08, 1.473243e-08, 1.231638e-08, 1.112644e-08, 1.038726e-08,
  9.752626e-09, 1.044174e-08, 1.098067e-08, 1.157846e-08, 1.245756e-08, 
    1.347156e-08, 1.468335e-08, 1.600878e-08, 1.738893e-08, 1.804043e-08, 
    1.739477e-08, 1.538491e-08, 1.315702e-08, 1.104771e-08, 1.04849e-08,
  9.543102e-09, 1.032134e-08, 1.09618e-08, 1.143438e-08, 1.19301e-08, 
    1.258133e-08, 1.340204e-08, 1.421299e-08, 1.524524e-08, 1.573962e-08, 
    1.5659e-08, 1.453591e-08, 1.283026e-08, 1.154126e-08, 1.068108e-08,
  9.127592e-09, 9.90479e-09, 1.064176e-08, 1.114788e-08, 1.162607e-08, 
    1.171774e-08, 1.225977e-08, 1.261226e-08, 1.313923e-08, 1.34293e-08, 
    1.315356e-08, 1.265368e-08, 1.179539e-08, 1.105368e-08, 1.028238e-08,
  8.849939e-09, 9.430391e-09, 1.038304e-08, 1.097125e-08, 1.14658e-08, 
    1.154908e-08, 1.154479e-08, 1.162639e-08, 1.160758e-08, 1.154864e-08, 
    1.141454e-08, 1.104166e-08, 1.076905e-08, 1.042329e-08, 1.011775e-08,
  8.377e-09, 8.852093e-09, 9.903983e-09, 1.071578e-08, 1.129392e-08, 
    1.12856e-08, 1.121477e-08, 1.100951e-08, 1.085575e-08, 1.069793e-08, 
    1.053516e-08, 1.045186e-08, 1.04198e-08, 1.036699e-08, 1.035751e-08,
  7.93067e-09, 8.242254e-09, 9.433255e-09, 1.037695e-08, 1.124941e-08, 
    1.14138e-08, 1.09668e-08, 1.065701e-08, 1.019584e-08, 9.97616e-09, 
    9.7551e-09, 9.568026e-09, 9.506283e-09, 9.387739e-09, 9.273449e-09,
  7.699731e-09, 7.62634e-09, 8.991499e-09, 1.012724e-08, 1.108235e-08, 
    1.157232e-08, 1.086679e-08, 1.006701e-08, 9.095757e-09, 8.657423e-09, 
    8.169078e-09, 7.897774e-09, 7.684148e-09, 7.54903e-09, 7.425855e-09,
  7.583218e-09, 7.112614e-09, 8.275148e-09, 9.758813e-09, 1.112564e-08, 
    1.170624e-08, 1.101077e-08, 9.675265e-09, 8.201813e-09, 7.497352e-09, 
    6.928751e-09, 6.694175e-09, 6.618921e-09, 6.595205e-09, 6.649001e-09,
  7.59024e-09, 6.720804e-09, 7.35423e-09, 9.199312e-09, 1.10134e-08, 
    1.217776e-08, 1.158818e-08, 9.821171e-09, 7.617345e-09, 6.801081e-09, 
    6.246219e-09, 6.131308e-09, 6.090755e-09, 6.086725e-09, 6.149631e-09,
  1.381233e-08, 1.461093e-08, 1.55006e-08, 1.642627e-08, 1.695069e-08, 
    1.703983e-08, 1.659648e-08, 1.536722e-08, 1.390543e-08, 1.216654e-08, 
    1.064243e-08, 9.632682e-09, 8.515522e-09, 7.278821e-09, 6.366615e-09,
  1.279765e-08, 1.326422e-08, 1.37308e-08, 1.46425e-08, 1.515581e-08, 
    1.551643e-08, 1.527137e-08, 1.459717e-08, 1.363103e-08, 1.247536e-08, 
    1.098705e-08, 9.754189e-09, 8.587413e-09, 7.175552e-09, 6.411568e-09,
  1.187076e-08, 1.209487e-08, 1.225837e-08, 1.268602e-08, 1.304012e-08, 
    1.33446e-08, 1.335437e-08, 1.300482e-08, 1.255171e-08, 1.173403e-08, 
    1.063858e-08, 9.679058e-09, 8.828573e-09, 7.491834e-09, 6.55083e-09,
  1.14334e-08, 1.147729e-08, 1.142603e-08, 1.149696e-08, 1.162325e-08, 
    1.169362e-08, 1.178253e-08, 1.173539e-08, 1.167968e-08, 1.125011e-08, 
    1.060765e-08, 9.934402e-09, 8.927477e-09, 7.695784e-09, 6.798057e-09,
  1.102e-08, 1.107533e-08, 1.098461e-08, 1.101913e-08, 1.109621e-08, 
    1.106275e-08, 1.111152e-08, 1.110732e-08, 1.110596e-08, 1.074211e-08, 
    1.012364e-08, 9.451794e-09, 8.606971e-09, 7.642956e-09, 6.896824e-09,
  1.071874e-08, 1.076136e-08, 1.076194e-08, 1.086125e-08, 1.092403e-08, 
    1.087406e-08, 1.0847e-08, 1.074892e-08, 1.049156e-08, 1.008716e-08, 
    9.463895e-09, 8.87983e-09, 8.18532e-09, 7.445012e-09, 6.863073e-09,
  1.053759e-08, 1.059063e-08, 1.060938e-08, 1.077864e-08, 1.085106e-08, 
    1.078396e-08, 1.065326e-08, 1.041086e-08, 1.003609e-08, 9.531787e-09, 
    8.974563e-09, 8.492095e-09, 7.902626e-09, 7.396959e-09, 6.900969e-09,
  1.047473e-08, 1.04162e-08, 1.058158e-08, 1.068139e-08, 1.067936e-08, 
    1.048098e-08, 1.027224e-08, 9.870173e-09, 9.426648e-09, 8.941701e-09, 
    8.514497e-09, 8.146483e-09, 7.804004e-09, 7.560614e-09, 7.39375e-09,
  1.044707e-08, 1.043577e-08, 1.0571e-08, 1.055471e-08, 1.030819e-08, 
    9.993294e-09, 9.737051e-09, 9.327165e-09, 8.885376e-09, 8.555917e-09, 
    8.233474e-09, 8.090918e-09, 7.888586e-09, 7.846331e-09, 7.98862e-09,
  1.048736e-08, 1.038225e-08, 1.056547e-08, 1.043146e-08, 9.908667e-09, 
    9.450775e-09, 9.191549e-09, 8.808151e-09, 8.554728e-09, 8.289627e-09, 
    8.084647e-09, 8.043308e-09, 7.95295e-09, 8.092699e-09, 8.14189e-09,
  1.575157e-08, 1.53101e-08, 1.454718e-08, 1.328828e-08, 1.21275e-08, 
    1.122976e-08, 1.02101e-08, 8.888997e-09, 7.7916e-09, 7.000347e-09, 
    6.174735e-09, 5.580212e-09, 5.112775e-09, 4.924297e-09, 4.807801e-09,
  1.564674e-08, 1.565436e-08, 1.500093e-08, 1.383022e-08, 1.257024e-08, 
    1.141899e-08, 1.042374e-08, 9.075243e-09, 7.86388e-09, 6.97562e-09, 
    6.130832e-09, 5.533393e-09, 5.127266e-09, 5.006665e-09, 4.900152e-09,
  1.543443e-08, 1.572461e-08, 1.514806e-08, 1.40545e-08, 1.286063e-08, 
    1.170711e-08, 1.055842e-08, 9.224248e-09, 7.967439e-09, 6.887253e-09, 
    6.172681e-09, 5.530511e-09, 5.195325e-09, 5.024453e-09, 4.81884e-09,
  1.515373e-08, 1.554926e-08, 1.504289e-08, 1.40586e-08, 1.300934e-08, 
    1.18705e-08, 1.069594e-08, 9.384477e-09, 8.003564e-09, 6.873419e-09, 
    6.138073e-09, 5.480413e-09, 5.127458e-09, 4.914988e-09, 4.681291e-09,
  1.492459e-08, 1.526764e-08, 1.485159e-08, 1.396876e-08, 1.302761e-08, 
    1.193105e-08, 1.078565e-08, 9.436578e-09, 7.986308e-09, 6.845517e-09, 
    6.049024e-09, 5.497822e-09, 5.085487e-09, 4.835369e-09, 4.712702e-09,
  1.469818e-08, 1.502624e-08, 1.468188e-08, 1.380704e-08, 1.291837e-08, 
    1.194296e-08, 1.077082e-08, 9.38474e-09, 7.885888e-09, 6.714981e-09, 
    5.928192e-09, 5.395244e-09, 5.041257e-09, 4.861946e-09, 4.901958e-09,
  1.433471e-08, 1.472888e-08, 1.451341e-08, 1.357848e-08, 1.277607e-08, 
    1.185777e-08, 1.067029e-08, 9.194738e-09, 7.636804e-09, 6.556567e-09, 
    5.885763e-09, 5.399249e-09, 5.022925e-09, 4.959456e-09, 5.036816e-09,
  1.389504e-08, 1.439456e-08, 1.431452e-08, 1.346966e-08, 1.256477e-08, 
    1.164619e-08, 1.043364e-08, 8.822155e-09, 7.389014e-09, 6.406946e-09, 
    5.746782e-09, 5.253107e-09, 4.973046e-09, 5.092941e-09, 5.167488e-09,
  1.338063e-08, 1.396147e-08, 1.407074e-08, 1.331042e-08, 1.234279e-08, 
    1.129741e-08, 1.010854e-08, 8.465883e-09, 7.17443e-09, 6.245041e-09, 
    5.608146e-09, 5.150699e-09, 5.143636e-09, 5.324178e-09, 5.519078e-09,
  1.296842e-08, 1.350277e-08, 1.375192e-08, 1.316629e-08, 1.212365e-08, 
    1.093248e-08, 9.724575e-09, 8.144537e-09, 6.954892e-09, 6.037541e-09, 
    5.409846e-09, 5.201781e-09, 5.439365e-09, 5.826619e-09, 5.17765e-09,
  1.06366e-08, 8.699951e-09, 7.62868e-09, 6.828072e-09, 6.299866e-09, 
    5.954839e-09, 6.015954e-09, 6.05769e-09, 6.09947e-09, 6.166326e-09, 
    6.406154e-09, 6.674071e-09, 7.091622e-09, 7.458694e-09, 7.830576e-09,
  1.092684e-08, 8.943181e-09, 7.736932e-09, 6.830929e-09, 6.237133e-09, 
    6.012849e-09, 6.03826e-09, 5.893544e-09, 5.850415e-09, 5.965411e-09, 
    6.105403e-09, 6.285727e-09, 6.552868e-09, 6.926012e-09, 7.348716e-09,
  1.128994e-08, 9.290891e-09, 7.975824e-09, 6.998647e-09, 6.322499e-09, 
    6.169898e-09, 6.022439e-09, 5.706049e-09, 5.616647e-09, 5.588956e-09, 
    5.616343e-09, 5.799206e-09, 5.977265e-09, 6.321199e-09, 6.686671e-09,
  1.166547e-08, 9.68454e-09, 8.284845e-09, 7.270152e-09, 6.526052e-09, 
    6.349378e-09, 5.964425e-09, 5.476582e-09, 5.281287e-09, 5.311928e-09, 
    5.358833e-09, 5.497711e-09, 5.695574e-09, 5.966958e-09, 6.236572e-09,
  1.211206e-08, 1.011835e-08, 8.679868e-09, 7.596356e-09, 6.789469e-09, 
    6.514571e-09, 5.903943e-09, 5.25486e-09, 5.164011e-09, 5.220239e-09, 
    5.32245e-09, 5.600161e-09, 5.822225e-09, 6.075414e-09, 6.232564e-09,
  1.259145e-08, 1.058071e-08, 9.102735e-09, 7.981655e-09, 7.115996e-09, 
    6.675973e-09, 5.868401e-09, 5.170167e-09, 5.140462e-09, 5.237217e-09, 
    5.504475e-09, 5.696033e-09, 5.920652e-09, 6.067434e-09, 6.1133e-09,
  1.321839e-08, 1.107294e-08, 9.541775e-09, 8.367121e-09, 7.416364e-09, 
    6.843536e-09, 5.87626e-09, 5.17153e-09, 5.194021e-09, 5.363507e-09, 
    5.531467e-09, 5.637776e-09, 5.749018e-09, 5.743973e-09, 5.730773e-09,
  1.386865e-08, 1.160668e-08, 1.000449e-08, 8.762285e-09, 7.721509e-09, 
    7.043705e-09, 5.916226e-09, 5.243668e-09, 5.268524e-09, 5.426471e-09, 
    5.493695e-09, 5.566569e-09, 5.570117e-09, 5.456718e-09, 5.400368e-09,
  1.461988e-08, 1.222207e-08, 1.050684e-08, 9.154784e-09, 8.045232e-09, 
    7.266949e-09, 6.020803e-09, 5.317565e-09, 5.34425e-09, 5.438809e-09, 
    5.484149e-09, 5.435565e-09, 5.313374e-09, 5.106934e-09, 5.012739e-09,
  1.520162e-08, 1.296035e-08, 1.106255e-08, 9.564077e-09, 8.382193e-09, 
    7.521027e-09, 6.168492e-09, 5.403317e-09, 5.401067e-09, 5.474643e-09, 
    5.430597e-09, 5.29894e-09, 4.97693e-09, 4.60546e-09, 4.415981e-09 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
