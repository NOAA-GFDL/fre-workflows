netcdf \00010101.atmos_daily.tile4.pv350K {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pv350K(time, grid_yt, grid_xt) ;
		pv350K:_FillValue = -1.e+10f ;
		pv350K:missing_value = -1.e+10f ;
		pv350K:units = "(K m**2) / (kg s)" ;
		pv350K:long_name = "350-K potential vorticity; needs x350 scaling" ;
		pv350K:cell_methods = "time: mean" ;
		pv350K:time_avg_info = "average_T1,average_T2,average_DT" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:03 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile4.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile4.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.2466774, 0.6143242, 0.0668168, 0.2301621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.4924844, 0.2132108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.600569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1560082, 0,
  1, 1, 0.7132517, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02739768, 0,
  0.6230268, 0.6280472, 0.3043983, 0.08344039, 0, 0.3148882, 0.01188002, 0, 
    0, 0, 0, 0.08803581, 0, 0, 0,
  0, 0, 0, 0, 0.01144353, 0.8597386, 0.8205094, 0.5086318, 0.1258651, 
    0.08909279, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.291879, 0.6933324, 1, 0.9996726, 0.6666086, 0.08008575, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.611689, 0.7180831, 0.4623523, 0.2838529, 0.02767258, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0.002817577, 0.8915156, 0.5654301, 0.7485356, 0.3018697, 0, 0, 0, 
    0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pv350K =
  1.763946e-08, 1.320075e-08, 8.926571e-09, 5.418471e-09, 3.740519e-09, 
    3.104116e-09, 2.718356e-09, 2.333481e-09, 1.756542e-09, 1.226549e-09, 
    7.532366e-10, 4.061283e-10, 3.051805e-10, 5.073194e-10, 7.653645e-10,
  1.824778e-08, 1.424091e-08, 9.799625e-09, 5.916711e-09, 3.908095e-09, 
    3.196909e-09, 2.779213e-09, 2.374651e-09, 1.773806e-09, 1.188054e-09, 
    7.256077e-10, 3.669118e-10, 2.334334e-10, 4.040162e-10, 7.04689e-10,
  1.864193e-08, 1.527089e-08, 1.070404e-08, 6.436788e-09, 4.0715e-09, 
    3.249067e-09, 2.836499e-09, 2.43275e-09, 1.836753e-09, 1.211074e-09, 
    7.162912e-10, 3.757084e-10, 2.060561e-10, 3.499665e-10, 6.566421e-10,
  1.927314e-08, 1.609961e-08, 1.168845e-08, 7.057263e-09, 4.340741e-09, 
    3.39563e-09, 2.977395e-09, 2.51403e-09, 1.91984e-09, 1.256533e-09, 
    7.079829e-10, 3.866014e-10, 1.94463e-10, 3.177981e-10, 5.998343e-10,
  1.972093e-08, 1.684464e-08, 1.281462e-08, 7.827079e-09, 4.656465e-09, 
    3.494412e-09, 3.092937e-09, 2.595397e-09, 2.00835e-09, 1.332818e-09, 
    7.315407e-10, 3.84401e-10, 1.891533e-10, 2.579324e-10, 5.236017e-10,
  2.022448e-08, 1.743467e-08, 1.379317e-08, 8.614753e-09, 5.052078e-09, 
    3.638043e-09, 3.197948e-09, 2.656457e-09, 2.070883e-09, 1.390808e-09, 
    7.691425e-10, 3.889835e-10, 1.803502e-10, 1.828716e-10, 4.384595e-10,
  2.075666e-08, 1.804057e-08, 1.470475e-08, 9.594135e-09, 5.394694e-09, 
    3.65821e-09, 3.274986e-09, 2.822758e-09, 2.277065e-09, 1.53322e-09, 
    8.228013e-10, 3.91968e-10, 1.596345e-10, 1.164512e-10, 4.130951e-10,
  2.1193e-08, 1.869134e-08, 1.562117e-08, 1.063566e-08, 5.953062e-09, 
    3.819459e-09, 3.371765e-09, 3.076596e-09, 2.600721e-09, 1.701541e-09, 
    8.660221e-10, 3.908031e-10, 1.507199e-10, 1.075313e-10, 4.185763e-10,
  2.161422e-08, 1.924648e-08, 1.638756e-08, 1.164352e-08, 6.746177e-09, 
    4.391973e-09, 3.803409e-09, 3.287744e-09, 2.534304e-09, 1.673121e-09, 
    9.049457e-10, 4.049696e-10, 1.599935e-10, 1.496859e-10, 4.553197e-10,
  2.196286e-08, 1.979274e-08, 1.711542e-08, 1.281403e-08, 7.691031e-09, 
    4.623553e-09, 3.942348e-09, 3.450054e-09, 2.55892e-09, 1.707257e-09, 
    9.612952e-10, 4.492486e-10, 1.88149e-10, 2.172054e-10, 4.94964e-10,
  2.269588e-08, 2.089269e-08, 1.718123e-08, 1.278464e-08, 8.871353e-09, 
    5.755027e-09, 4.69296e-09, 4.377922e-09, 3.989816e-09, 3.324904e-09, 
    2.724384e-09, 2.250775e-09, 2.03023e-09, 2.108368e-09, 2.076416e-09,
  2.277233e-08, 2.103762e-08, 1.720567e-08, 1.281168e-08, 8.925277e-09, 
    5.836427e-09, 4.628537e-09, 4.231674e-09, 3.710839e-09, 2.896687e-09, 
    2.136425e-09, 1.640705e-09, 1.574583e-09, 1.798155e-09, 1.936154e-09,
  2.284275e-08, 2.113959e-08, 1.746594e-08, 1.313196e-08, 9.101597e-09, 
    5.735768e-09, 4.404141e-09, 3.999629e-09, 3.421764e-09, 2.521759e-09, 
    1.820478e-09, 1.475518e-09, 1.502671e-09, 1.893328e-09, 2.042296e-09,
  2.286018e-08, 2.141e-08, 1.753529e-08, 1.321902e-08, 9.17084e-09, 
    5.696355e-09, 4.297841e-09, 3.883023e-09, 3.270075e-09, 2.334719e-09, 
    1.618562e-09, 1.358551e-09, 1.592481e-09, 2.01693e-09, 2.134853e-09,
  2.278295e-08, 2.138682e-08, 1.779548e-08, 1.34546e-08, 9.258785e-09, 
    5.583954e-09, 4.104439e-09, 3.734705e-09, 3.115025e-09, 2.096456e-09, 
    1.373889e-09, 1.284177e-09, 1.693919e-09, 2.114059e-09, 2.065748e-09,
  2.262877e-08, 2.143886e-08, 1.784596e-08, 1.359923e-08, 9.38063e-09, 
    5.493945e-09, 3.880396e-09, 3.433309e-09, 2.784894e-09, 1.800319e-09, 
    1.191256e-09, 1.312874e-09, 1.842774e-09, 2.14586e-09, 1.920154e-09,
  2.282289e-08, 2.127486e-08, 1.775498e-08, 1.371868e-08, 9.295825e-09, 
    5.239225e-09, 3.673905e-09, 3.308708e-09, 2.825935e-09, 1.812189e-09, 
    1.194266e-09, 1.45604e-09, 1.963524e-09, 2.108141e-09, 1.726467e-09,
  2.284286e-08, 2.125535e-08, 1.770888e-08, 1.373235e-08, 9.213983e-09, 
    5.309701e-09, 3.924622e-09, 3.798605e-09, 3.31387e-09, 1.950773e-09, 
    1.220752e-09, 1.555876e-09, 2.008864e-09, 1.977436e-09, 1.496321e-09,
  2.285065e-08, 2.116632e-08, 1.759678e-08, 1.35591e-08, 9.403846e-09, 
    5.941212e-09, 4.492203e-09, 3.932854e-09, 2.881428e-09, 1.631943e-09, 
    1.20763e-09, 1.550208e-09, 1.894915e-09, 1.746492e-09, 1.281706e-09,
  2.287505e-08, 2.10893e-08, 1.750367e-08, 1.365604e-08, 9.593266e-09, 
    5.749145e-09, 4.207783e-09, 3.539842e-09, 2.481078e-09, 1.587075e-09, 
    1.270557e-09, 1.490563e-09, 1.67252e-09, 1.458946e-09, 1.115899e-09,
  2.286494e-08, 2.226209e-08, 2.138702e-08, 1.990592e-08, 1.733777e-08, 
    1.377608e-08, 1.044773e-08, 8.41049e-09, 6.955642e-09, 5.609991e-09, 
    4.477228e-09, 3.877827e-09, 3.477817e-09, 3.101498e-09, 2.706025e-09,
  2.308187e-08, 2.236201e-08, 2.131009e-08, 2.002667e-08, 1.756561e-08, 
    1.385386e-08, 1.030393e-08, 8.177484e-09, 6.662498e-09, 5.264491e-09, 
    4.16772e-09, 3.59118e-09, 3.222815e-09, 2.908466e-09, 2.48287e-09,
  2.305212e-08, 2.233755e-08, 2.141559e-08, 1.995294e-08, 1.743564e-08, 
    1.355448e-08, 9.910353e-09, 7.80483e-09, 6.318595e-09, 4.893472e-09, 
    3.822992e-09, 3.354001e-09, 3.094198e-09, 2.780643e-09, 2.257705e-09,
  2.312475e-08, 2.255729e-08, 2.146348e-08, 1.986616e-08, 1.725363e-08, 
    1.317413e-08, 9.430096e-09, 7.429403e-09, 6.005181e-09, 4.603863e-09, 
    3.642339e-09, 3.280005e-09, 3.045899e-09, 2.663321e-09, 1.990608e-09,
  2.312848e-08, 2.253759e-08, 2.138608e-08, 1.977121e-08, 1.68886e-08, 
    1.261108e-08, 8.946897e-09, 7.113315e-09, 5.710967e-09, 4.317654e-09, 
    3.452137e-09, 3.176255e-09, 2.919841e-09, 2.449831e-09, 1.735866e-09,
  2.297999e-08, 2.249326e-08, 2.118287e-08, 1.950943e-08, 1.671888e-08, 
    1.215884e-08, 8.37146e-09, 6.590921e-09, 5.264809e-09, 3.973718e-09, 
    3.286833e-09, 3.060606e-09, 2.790687e-09, 2.290686e-09, 1.533571e-09,
  2.28689e-08, 2.229891e-08, 2.081265e-08, 1.918308e-08, 1.60283e-08, 
    1.147779e-08, 7.94628e-09, 6.322079e-09, 5.055936e-09, 3.85787e-09, 
    3.235419e-09, 2.999281e-09, 2.67334e-09, 2.107431e-09, 1.440336e-09,
  2.30901e-08, 2.22631e-08, 2.061554e-08, 1.892759e-08, 1.562892e-08, 
    1.101469e-08, 7.859446e-09, 6.733269e-09, 5.476693e-09, 3.916935e-09, 
    3.193335e-09, 2.945334e-09, 2.563982e-09, 2.02266e-09, 1.342917e-09,
  2.292304e-08, 2.215018e-08, 2.039221e-08, 1.838703e-08, 1.530242e-08, 
    1.099684e-08, 8.080084e-09, 6.693834e-09, 4.932227e-09, 3.432319e-09, 
    2.988892e-09, 2.807892e-09, 2.486304e-09, 1.932882e-09, 1.270332e-09,
  2.288816e-08, 2.203889e-08, 2.011748e-08, 1.799961e-08, 1.466191e-08, 
    1.01547e-08, 7.536165e-09, 6.150404e-09, 4.314717e-09, 3.119848e-09, 
    2.842366e-09, 2.617996e-09, 2.309982e-09, 1.748742e-09, 1.285846e-09,
  2.414212e-08, 2.329332e-08, 2.317081e-08, 2.347766e-08, 2.242738e-08, 
    2.087308e-08, 1.886471e-08, 1.620482e-08, 1.331107e-08, 1.073018e-08, 
    8.640543e-09, 7.058105e-09, 5.849437e-09, 4.802568e-09, 3.891458e-09,
  2.43351e-08, 2.353276e-08, 2.321428e-08, 2.34816e-08, 2.240454e-08, 
    2.068159e-08, 1.83326e-08, 1.555411e-08, 1.265084e-08, 1.010828e-08, 
    8.129944e-09, 6.622287e-09, 5.456593e-09, 4.371139e-09, 3.573321e-09,
  2.444472e-08, 2.365312e-08, 2.315529e-08, 2.339207e-08, 2.220995e-08, 
    2.035857e-08, 1.7834e-08, 1.488551e-08, 1.185527e-08, 9.368831e-09, 
    7.564447e-09, 6.191118e-09, 5.023658e-09, 3.920001e-09, 3.326475e-09,
  2.423898e-08, 2.362652e-08, 2.326045e-08, 2.329763e-08, 2.199463e-08, 
    1.99825e-08, 1.718056e-08, 1.40646e-08, 1.106015e-08, 8.748334e-09, 
    7.114409e-09, 5.793839e-09, 4.596758e-09, 3.6257e-09, 3.207531e-09,
  2.446889e-08, 2.371812e-08, 2.327616e-08, 2.325987e-08, 2.169001e-08, 
    1.943062e-08, 1.658598e-08, 1.338124e-08, 1.0326e-08, 8.207789e-09, 
    6.672322e-09, 5.350222e-09, 4.181228e-09, 3.481801e-09, 3.096655e-09,
  2.401197e-08, 2.351557e-08, 2.321123e-08, 2.312387e-08, 2.151496e-08, 
    1.886701e-08, 1.557049e-08, 1.230603e-08, 9.465712e-09, 7.6721e-09, 
    6.182356e-09, 4.881599e-09, 3.859393e-09, 3.327193e-09, 2.942497e-09,
  2.413074e-08, 2.34822e-08, 2.311967e-08, 2.304316e-08, 2.108445e-08, 
    1.811583e-08, 1.493354e-08, 1.151326e-08, 8.856397e-09, 7.234745e-09, 
    5.683481e-09, 4.445947e-09, 3.577684e-09, 3.093608e-09, 2.726437e-09,
  2.407731e-08, 2.337962e-08, 2.307478e-08, 2.297299e-08, 2.066664e-08, 
    1.777302e-08, 1.463788e-08, 1.130955e-08, 8.704483e-09, 6.879266e-09, 
    5.227422e-09, 4.053181e-09, 3.27642e-09, 2.893623e-09, 2.534783e-09,
  2.410516e-08, 2.341106e-08, 2.319594e-08, 2.284609e-08, 2.078165e-08, 
    1.801796e-08, 1.416196e-08, 1.060453e-08, 8.093769e-09, 6.307019e-09, 
    4.809106e-09, 3.747814e-09, 3.052082e-09, 2.761094e-09, 2.286206e-09,
  2.406608e-08, 2.332521e-08, 2.31504e-08, 2.25042e-08, 2.043659e-08, 
    1.750773e-08, 1.32652e-08, 9.800364e-09, 7.386662e-09, 5.73816e-09, 
    4.403963e-09, 3.395725e-09, 2.879874e-09, 2.59487e-09, 2.034124e-09,
  2.466771e-08, 2.375221e-08, 2.293219e-08, 2.274246e-08, 2.248159e-08, 
    2.172123e-08, 2.051621e-08, 1.886127e-08, 1.702238e-08, 1.502517e-08, 
    1.271784e-08, 1.049325e-08, 8.801758e-09, 7.447712e-09, 6.228686e-09,
  2.48216e-08, 2.383948e-08, 2.295579e-08, 2.260928e-08, 2.227672e-08, 
    2.15057e-08, 2.012196e-08, 1.842665e-08, 1.652845e-08, 1.438527e-08, 
    1.197185e-08, 9.903204e-09, 8.364869e-09, 7.08719e-09, 5.87287e-09,
  2.502057e-08, 2.38729e-08, 2.284267e-08, 2.253433e-08, 2.210436e-08, 
    2.124146e-08, 1.970892e-08, 1.79326e-08, 1.589868e-08, 1.360992e-08, 
    1.121062e-08, 9.284801e-09, 7.882946e-09, 6.645515e-09, 5.449234e-09,
  2.484953e-08, 2.379793e-08, 2.286939e-08, 2.25672e-08, 2.209302e-08, 
    2.107658e-08, 1.929851e-08, 1.739499e-08, 1.53125e-08, 1.290957e-08, 
    1.05821e-08, 8.848667e-09, 7.503149e-09, 6.228211e-09, 5.020469e-09,
  2.516702e-08, 2.389968e-08, 2.272089e-08, 2.247312e-08, 2.191645e-08, 
    2.086362e-08, 1.900588e-08, 1.704303e-08, 1.478639e-08, 1.228781e-08, 
    1.008291e-08, 8.450193e-09, 7.057135e-09, 5.769149e-09, 4.599413e-09,
  2.468463e-08, 2.374553e-08, 2.274624e-08, 2.253834e-08, 2.193571e-08, 
    2.061413e-08, 1.85425e-08, 1.647642e-08, 1.414695e-08, 1.163688e-08, 
    9.54564e-09, 7.973752e-09, 6.535324e-09, 5.308131e-09, 4.195377e-09,
  2.474773e-08, 2.371318e-08, 2.269957e-08, 2.245516e-08, 2.159733e-08, 
    2.035769e-08, 1.813132e-08, 1.58612e-08, 1.344581e-08, 1.0928e-08, 
    8.959461e-09, 7.422716e-09, 6.051625e-09, 4.887833e-09, 3.850647e-09,
  2.469182e-08, 2.373323e-08, 2.267366e-08, 2.250628e-08, 2.145698e-08, 
    1.991655e-08, 1.771658e-08, 1.551579e-08, 1.290234e-08, 1.026213e-08, 
    8.384208e-09, 6.863987e-09, 5.647624e-09, 4.530526e-09, 3.574314e-09,
  2.472123e-08, 2.371221e-08, 2.261577e-08, 2.23508e-08, 2.134115e-08, 
    1.981814e-08, 1.73128e-08, 1.500561e-08, 1.200549e-08, 9.440825e-09, 
    7.786253e-09, 6.423245e-09, 5.2904e-09, 4.191885e-09, 3.270941e-09,
  2.47134e-08, 2.367634e-08, 2.256239e-08, 2.222446e-08, 2.097532e-08, 
    1.94147e-08, 1.636736e-08, 1.402963e-08, 1.093311e-08, 8.797485e-09, 
    7.297627e-09, 6.01402e-09, 4.939837e-09, 3.851878e-09, 2.983604e-09,
  2.425671e-08, 2.396548e-08, 2.285835e-08, 2.122296e-08, 2.001603e-08, 
    1.918768e-08, 1.944789e-08, 1.987802e-08, 1.828377e-08, 1.63598e-08, 
    1.460419e-08, 1.316287e-08, 1.156529e-08, 9.603888e-09, 7.551419e-09,
  2.423013e-08, 2.412532e-08, 2.319888e-08, 2.144269e-08, 2.033291e-08, 
    1.938425e-08, 1.950248e-08, 1.964203e-08, 1.797416e-08, 1.614826e-08, 
    1.444399e-08, 1.299462e-08, 1.138632e-08, 9.437243e-09, 7.411875e-09,
  2.438322e-08, 2.439915e-08, 2.345299e-08, 2.176881e-08, 2.054911e-08, 
    1.950487e-08, 1.963141e-08, 1.951411e-08, 1.770493e-08, 1.580476e-08, 
    1.414949e-08, 1.267176e-08, 1.105975e-08, 9.193389e-09, 7.226526e-09,
  2.398171e-08, 2.42029e-08, 2.368637e-08, 2.193624e-08, 2.075279e-08, 
    1.962182e-08, 1.97065e-08, 1.919238e-08, 1.729618e-08, 1.549701e-08, 
    1.391389e-08, 1.248143e-08, 1.090515e-08, 9.032802e-09, 7.115191e-09,
  2.396779e-08, 2.422503e-08, 2.371019e-08, 2.203292e-08, 2.07377e-08, 
    1.962855e-08, 1.979883e-08, 1.903887e-08, 1.7038e-08, 1.522983e-08, 
    1.37347e-08, 1.233635e-08, 1.070678e-08, 8.777508e-09, 6.924377e-09,
  2.410611e-08, 2.408699e-08, 2.361592e-08, 2.200467e-08, 2.07844e-08, 
    1.954013e-08, 1.963709e-08, 1.863158e-08, 1.663494e-08, 1.496205e-08, 
    1.356106e-08, 1.214134e-08, 1.041114e-08, 8.419765e-09, 6.673031e-09,
  2.370245e-08, 2.374205e-08, 2.338013e-08, 2.192424e-08, 2.057794e-08, 
    1.969066e-08, 1.987004e-08, 1.838661e-08, 1.626831e-08, 1.474e-08, 
    1.333845e-08, 1.18332e-08, 1.000948e-08, 8.01728e-09, 6.380438e-09,
  2.313408e-08, 2.350808e-08, 2.334077e-08, 2.187063e-08, 2.065667e-08, 
    1.963825e-08, 1.9706e-08, 1.846008e-08, 1.642941e-08, 1.462994e-08, 
    1.306498e-08, 1.147574e-08, 9.566453e-09, 7.600901e-09, 6.025715e-09,
  2.412026e-08, 2.444756e-08, 2.354623e-08, 2.178199e-08, 2.063289e-08, 
    2.007554e-08, 1.984104e-08, 1.826496e-08, 1.59468e-08, 1.405667e-08, 
    1.270275e-08, 1.103973e-08, 9.090004e-09, 7.147018e-09, 5.595839e-09,
  2.497775e-08, 2.467286e-08, 2.364951e-08, 2.171099e-08, 2.054847e-08, 
    1.999496e-08, 1.917131e-08, 1.736605e-08, 1.49806e-08, 1.366283e-08, 
    1.231474e-08, 1.051918e-08, 8.563549e-09, 6.637047e-09, 5.078894e-09,
  2.1163e-08, 1.991039e-08, 1.913269e-08, 1.862089e-08, 1.801729e-08, 
    1.75101e-08, 1.7198e-08, 1.690696e-08, 1.642827e-08, 1.608377e-08, 
    1.620847e-08, 1.553981e-08, 1.386857e-08, 1.20113e-08, 1.073345e-08,
  2.179669e-08, 2.039153e-08, 1.913793e-08, 1.85647e-08, 1.811521e-08, 
    1.770778e-08, 1.731532e-08, 1.703794e-08, 1.659906e-08, 1.618203e-08, 
    1.616668e-08, 1.58144e-08, 1.432509e-08, 1.245538e-08, 1.101214e-08,
  2.24212e-08, 2.116641e-08, 1.942874e-08, 1.866043e-08, 1.81518e-08, 
    1.780006e-08, 1.750933e-08, 1.720414e-08, 1.686003e-08, 1.632243e-08, 
    1.618914e-08, 1.600916e-08, 1.473708e-08, 1.286988e-08, 1.125692e-08,
  2.300161e-08, 2.132525e-08, 1.999604e-08, 1.896667e-08, 1.831973e-08, 
    1.798971e-08, 1.769086e-08, 1.751204e-08, 1.708129e-08, 1.647027e-08, 
    1.619708e-08, 1.608763e-08, 1.499551e-08, 1.31813e-08, 1.150423e-08,
  2.38304e-08, 2.173732e-08, 2.033155e-08, 1.914796e-08, 1.836357e-08, 
    1.793251e-08, 1.787508e-08, 1.78061e-08, 1.741806e-08, 1.659233e-08, 
    1.618047e-08, 1.612191e-08, 1.519574e-08, 1.342574e-08, 1.168724e-08,
  2.417709e-08, 2.2139e-08, 2.080679e-08, 1.933928e-08, 1.848836e-08, 
    1.809318e-08, 1.790015e-08, 1.807668e-08, 1.76842e-08, 1.673818e-08, 
    1.620464e-08, 1.608148e-08, 1.529573e-08, 1.360668e-08, 1.184514e-08,
  2.443345e-08, 2.255251e-08, 2.117168e-08, 1.953656e-08, 1.812587e-08, 
    1.774143e-08, 1.823781e-08, 1.866614e-08, 1.817675e-08, 1.688214e-08, 
    1.622814e-08, 1.601067e-08, 1.528466e-08, 1.367977e-08, 1.195352e-08,
  2.443525e-08, 2.282257e-08, 2.14396e-08, 1.978159e-08, 1.835417e-08, 
    1.755637e-08, 1.783831e-08, 1.841083e-08, 1.811143e-08, 1.690465e-08, 
    1.620649e-08, 1.584758e-08, 1.517981e-08, 1.367068e-08, 1.201081e-08,
  2.498759e-08, 2.37117e-08, 2.18166e-08, 1.974571e-08, 1.821082e-08, 
    1.745462e-08, 1.776317e-08, 1.833032e-08, 1.816257e-08, 1.707282e-08, 
    1.613383e-08, 1.565238e-08, 1.498221e-08, 1.355794e-08, 1.197012e-08,
  2.490937e-08, 2.357516e-08, 2.181554e-08, 1.974132e-08, 1.822511e-08, 
    1.740909e-08, 1.778343e-08, 1.872672e-08, 1.8474e-08, 1.717357e-08, 
    1.606548e-08, 1.547719e-08, 1.477519e-08, 1.340074e-08, 1.186493e-08,
  1.85626e-08, 1.771609e-08, 1.706006e-08, 1.663442e-08, 1.631472e-08, 
    1.586457e-08, 1.520311e-08, 1.395942e-08, 1.28461e-08, 1.199864e-08, 
    1.111307e-08, 9.937356e-09, 9.365159e-09, 8.904668e-09, 8.537681e-09,
  1.91931e-08, 1.804023e-08, 1.737181e-08, 1.678997e-08, 1.656666e-08, 
    1.621e-08, 1.588243e-08, 1.502979e-08, 1.381074e-08, 1.272346e-08, 
    1.196636e-08, 1.061308e-08, 9.673842e-09, 9.055956e-09, 8.790978e-09,
  2.003664e-08, 1.895199e-08, 1.793919e-08, 1.71724e-08, 1.678594e-08, 
    1.648218e-08, 1.618488e-08, 1.576711e-08, 1.478974e-08, 1.356041e-08, 
    1.271819e-08, 1.139021e-08, 1.011585e-08, 9.297454e-09, 8.884325e-09,
  2.069697e-08, 1.957307e-08, 1.854627e-08, 1.748083e-08, 1.703735e-08, 
    1.671935e-08, 1.645923e-08, 1.617189e-08, 1.559853e-08, 1.449632e-08, 
    1.347953e-08, 1.230291e-08, 1.078288e-08, 9.666889e-09, 8.99912e-09,
  2.269678e-08, 2.102355e-08, 1.937997e-08, 1.794038e-08, 1.729255e-08, 
    1.687617e-08, 1.658251e-08, 1.647138e-08, 1.619916e-08, 1.53794e-08, 
    1.433567e-08, 1.31942e-08, 1.160438e-08, 1.020804e-08, 9.236444e-09,
  2.337971e-08, 2.165471e-08, 2.036456e-08, 1.845622e-08, 1.756462e-08, 
    1.732842e-08, 1.688811e-08, 1.652418e-08, 1.64475e-08, 1.603296e-08, 
    1.523236e-08, 1.416612e-08, 1.262853e-08, 1.09624e-08, 9.663598e-09,
  2.439664e-08, 2.263193e-08, 2.108128e-08, 1.94639e-08, 1.770697e-08, 
    1.735346e-08, 1.738992e-08, 1.722779e-08, 1.690891e-08, 1.650714e-08, 
    1.59896e-08, 1.501509e-08, 1.367404e-08, 1.189561e-08, 1.029616e-08,
  2.523222e-08, 2.349978e-08, 2.198655e-08, 2.020154e-08, 1.870912e-08, 
    1.760191e-08, 1.740587e-08, 1.728039e-08, 1.714952e-08, 1.667069e-08, 
    1.650853e-08, 1.576093e-08, 1.466369e-08, 1.290424e-08, 1.111532e-08,
  2.637128e-08, 2.448746e-08, 2.293418e-08, 2.108946e-08, 1.935784e-08, 
    1.812455e-08, 1.76156e-08, 1.696994e-08, 1.683539e-08, 1.667761e-08, 
    1.675126e-08, 1.627138e-08, 1.545159e-08, 1.390782e-08, 1.200159e-08,
  2.685341e-08, 2.526727e-08, 2.385475e-08, 2.187647e-08, 2.023249e-08, 
    1.855496e-08, 1.776417e-08, 1.719212e-08, 1.689841e-08, 1.663344e-08, 
    1.682785e-08, 1.667864e-08, 1.602952e-08, 1.480806e-08, 1.28845e-08,
  1.687999e-08, 1.603202e-08, 1.517854e-08, 1.481401e-08, 1.479895e-08, 
    1.528723e-08, 1.581327e-08, 1.603963e-08, 1.564645e-08, 1.486295e-08, 
    1.34212e-08, 1.173199e-08, 9.651024e-09, 7.736131e-09, 6.220466e-09,
  1.707622e-08, 1.626982e-08, 1.574323e-08, 1.515921e-08, 1.489826e-08, 
    1.523991e-08, 1.554264e-08, 1.572395e-08, 1.562157e-08, 1.522513e-08, 
    1.430382e-08, 1.261829e-08, 1.097908e-08, 8.957135e-09, 7.377071e-09,
  1.684e-08, 1.652844e-08, 1.607192e-08, 1.548841e-08, 1.48555e-08, 
    1.478813e-08, 1.507195e-08, 1.520025e-08, 1.504315e-08, 1.479734e-08, 
    1.478065e-08, 1.340359e-08, 1.188974e-08, 1.022476e-08, 8.495293e-09,
  1.741401e-08, 1.720168e-08, 1.660722e-08, 1.576557e-08, 1.502108e-08, 
    1.457125e-08, 1.459018e-08, 1.465372e-08, 1.454664e-08, 1.400612e-08, 
    1.438174e-08, 1.382897e-08, 1.264264e-08, 1.128769e-08, 9.655862e-09,
  1.882193e-08, 1.80363e-08, 1.733127e-08, 1.623835e-08, 1.531461e-08, 
    1.457035e-08, 1.444257e-08, 1.446125e-08, 1.457017e-08, 1.419914e-08, 
    1.449571e-08, 1.420988e-08, 1.31901e-08, 1.19968e-08, 1.050311e-08,
  1.9982e-08, 1.909489e-08, 1.794083e-08, 1.662143e-08, 1.578534e-08, 
    1.49262e-08, 1.448431e-08, 1.405542e-08, 1.457172e-08, 1.454973e-08, 
    1.443602e-08, 1.423767e-08, 1.330003e-08, 1.230495e-08, 1.084774e-08,
  1.96797e-08, 1.889377e-08, 1.80576e-08, 1.695325e-08, 1.591245e-08, 
    1.494349e-08, 1.456121e-08, 1.388178e-08, 1.417609e-08, 1.451112e-08, 
    1.431316e-08, 1.398097e-08, 1.32008e-08, 1.243812e-08, 1.086674e-08,
  1.975185e-08, 1.904136e-08, 1.839201e-08, 1.734603e-08, 1.60142e-08, 
    1.518282e-08, 1.504929e-08, 1.50957e-08, 1.510765e-08, 1.453105e-08, 
    1.422482e-08, 1.350477e-08, 1.318028e-08, 1.273278e-08, 1.101247e-08,
  2.094226e-08, 1.968756e-08, 1.875162e-08, 1.749001e-08, 1.649734e-08, 
    1.636089e-08, 1.609636e-08, 1.597397e-08, 1.521136e-08, 1.433525e-08, 
    1.430694e-08, 1.348873e-08, 1.300445e-08, 1.29928e-08, 1.148062e-08,
  2.186929e-08, 2.025863e-08, 1.924417e-08, 1.80383e-08, 1.75267e-08, 
    1.702765e-08, 1.648357e-08, 1.610831e-08, 1.513042e-08, 1.414804e-08, 
    1.413786e-08, 1.384537e-08, 1.284908e-08, 1.268213e-08, 1.215075e-08,
  2.329322e-08, 2.348377e-08, 2.323724e-08, 2.244256e-08, 2.117794e-08, 
    1.964606e-08, 1.781792e-08, 1.594618e-08, 1.38426e-08, 1.089925e-08, 
    7.546633e-09, 4.997555e-09, 3.730394e-09, 3.396969e-09, 3.382506e-09,
  2.368098e-08, 2.373866e-08, 2.35639e-08, 2.298708e-08, 2.189527e-08, 
    2.066148e-08, 1.903043e-08, 1.733786e-08, 1.530426e-08, 1.261395e-08, 
    9.788232e-09, 6.826188e-09, 4.682878e-09, 3.697522e-09, 3.598035e-09,
  2.286101e-08, 2.290098e-08, 2.36941e-08, 2.361974e-08, 2.279191e-08, 
    2.164546e-08, 1.997513e-08, 1.827956e-08, 1.651773e-08, 1.414085e-08, 
    1.144168e-08, 8.714061e-09, 6.059722e-09, 4.507793e-09, 3.702428e-09,
  2.199478e-08, 2.27592e-08, 2.338202e-08, 2.375923e-08, 2.322152e-08, 
    2.217124e-08, 2.107035e-08, 1.939559e-08, 1.762633e-08, 1.56424e-08, 
    1.308115e-08, 1.056372e-08, 7.799388e-09, 5.693103e-09, 4.420307e-09,
  2.226721e-08, 2.288508e-08, 2.333037e-08, 2.371085e-08, 2.348931e-08, 
    2.291642e-08, 2.162556e-08, 2.02526e-08, 1.861218e-08, 1.675341e-08, 
    1.421081e-08, 1.213835e-08, 9.677393e-09, 7.13237e-09, 5.514613e-09,
  2.349565e-08, 2.43726e-08, 2.445959e-08, 2.383086e-08, 2.272516e-08, 
    2.23235e-08, 2.177199e-08, 2.049856e-08, 1.917215e-08, 1.769807e-08, 
    1.525734e-08, 1.306104e-08, 1.114917e-08, 8.869282e-09, 6.794846e-09,
  2.409557e-08, 2.395138e-08, 2.365725e-08, 2.362025e-08, 2.291478e-08, 
    2.259706e-08, 2.148505e-08, 2.074735e-08, 1.995646e-08, 1.860849e-08, 
    1.637053e-08, 1.421511e-08, 1.237689e-08, 1.029134e-08, 8.320879e-09,
  2.283538e-08, 2.242624e-08, 2.379383e-08, 2.33328e-08, 2.077209e-08, 
    2.107104e-08, 2.146461e-08, 2.176315e-08, 2.094266e-08, 1.962323e-08, 
    1.773192e-08, 1.567751e-08, 1.323213e-08, 1.140788e-08, 9.617836e-09,
  2.179686e-08, 2.078589e-08, 2.310449e-08, 2.060826e-08, 1.866214e-08, 
    2.110685e-08, 2.103128e-08, 2.200234e-08, 2.101223e-08, 1.959729e-08, 
    1.812015e-08, 1.653665e-08, 1.458611e-08, 1.253281e-08, 1.052995e-08,
  1.948198e-08, 1.894576e-08, 2.115857e-08, 1.796762e-08, 1.797407e-08, 
    1.889816e-08, 1.9152e-08, 2.051657e-08, 1.975316e-08, 1.905598e-08, 
    1.811203e-08, 1.696258e-08, 1.616559e-08, 1.40783e-08, 1.105192e-08,
  2.17344e-08, 2.140255e-08, 2.182217e-08, 2.311466e-08, 2.231089e-08, 
    2.069071e-08, 1.843199e-08, 1.55586e-08, 1.214467e-08, 7.488945e-09, 
    4.863254e-09, 3.218999e-09, 2.476627e-09, 2.089793e-09, 1.780629e-09,
  2.207265e-08, 2.163965e-08, 2.170799e-08, 2.258718e-08, 2.251641e-08, 
    2.137444e-08, 1.957801e-08, 1.688569e-08, 1.384819e-08, 9.573872e-09, 
    5.802047e-09, 3.734872e-09, 2.70412e-09, 2.122515e-09, 1.846406e-09,
  2.240854e-08, 2.174439e-08, 2.182586e-08, 2.164291e-08, 2.253183e-08, 
    2.188992e-08, 2.029925e-08, 1.795673e-08, 1.527882e-08, 1.15575e-08, 
    7.316068e-09, 4.438816e-09, 2.864519e-09, 2.301969e-09, 1.897705e-09,
  2.295402e-08, 2.19533e-08, 2.191087e-08, 2.16868e-08, 2.222216e-08, 
    2.231843e-08, 2.101432e-08, 1.885228e-08, 1.625588e-08, 1.300162e-08, 
    8.973758e-09, 5.328801e-09, 3.316362e-09, 2.496403e-09, 2.004764e-09,
  2.301808e-08, 2.244791e-08, 2.237969e-08, 2.197299e-08, 2.211681e-08, 
    2.214819e-08, 2.152171e-08, 1.969105e-08, 1.740858e-08, 1.43779e-08, 
    1.064868e-08, 6.573665e-09, 3.976021e-09, 2.692427e-09, 2.147393e-09,
  2.396119e-08, 2.301907e-08, 2.307253e-08, 2.209167e-08, 2.204812e-08, 
    2.22098e-08, 2.165412e-08, 1.998317e-08, 1.800398e-08, 1.528672e-08, 
    1.19732e-08, 7.824394e-09, 4.688668e-09, 2.968735e-09, 2.33622e-09,
  2.506255e-08, 2.350824e-08, 2.350839e-08, 2.269391e-08, 2.251136e-08, 
    2.196786e-08, 2.184655e-08, 2.064465e-08, 1.879019e-08, 1.623039e-08, 
    1.314853e-08, 9.14856e-09, 5.480623e-09, 3.382274e-09, 2.544256e-09,
  2.419921e-08, 2.39161e-08, 2.418133e-08, 2.335882e-08, 2.279904e-08, 
    2.230334e-08, 2.19098e-08, 2.072807e-08, 1.919762e-08, 1.682206e-08, 
    1.408542e-08, 1.041166e-08, 6.424572e-09, 3.957448e-09, 2.77612e-09,
  2.447149e-08, 2.400308e-08, 2.407474e-08, 2.351376e-08, 2.279784e-08, 
    2.221486e-08, 2.162454e-08, 2.062205e-08, 1.933466e-08, 1.729592e-08, 
    1.484085e-08, 1.162893e-08, 7.442878e-09, 4.596952e-09, 3.079583e-09,
  2.451352e-08, 2.402407e-08, 2.443377e-08, 2.350703e-08, 2.30489e-08, 
    2.202058e-08, 2.08558e-08, 2.041229e-08, 1.952931e-08, 1.768584e-08, 
    1.543296e-08, 1.264287e-08, 8.522171e-09, 5.336116e-09, 3.443633e-09,
  2.05912e-08, 2.172386e-08, 2.340936e-08, 2.32381e-08, 2.144601e-08, 
    1.860394e-08, 1.508431e-08, 1.012638e-08, 4.728969e-09, 1.992569e-09, 
    1.00374e-09, 8.120583e-10, 7.343025e-10, 5.590401e-10, 3.464558e-10,
  1.970464e-08, 2.091012e-08, 2.267219e-08, 2.359703e-08, 2.274994e-08, 
    2.047303e-08, 1.735493e-08, 1.328542e-08, 7.348551e-09, 3.218094e-09, 
    1.338079e-09, 1.02018e-09, 7.543055e-10, 6.630778e-10, 4.397681e-10,
  1.900079e-08, 1.969922e-08, 2.143404e-08, 2.317102e-08, 2.356889e-08, 
    2.194184e-08, 1.930531e-08, 1.595043e-08, 1.050362e-08, 5.079515e-09, 
    2.103393e-09, 1.068004e-09, 8.406563e-10, 7.117913e-10, 5.206662e-10,
  1.881942e-08, 1.930397e-08, 2.036794e-08, 2.247154e-08, 2.350977e-08, 
    2.327409e-08, 2.087935e-08, 1.798854e-08, 1.359569e-08, 7.518055e-09, 
    3.220432e-09, 1.324145e-09, 1.036468e-09, 7.558803e-10, 5.987976e-10,
  1.889475e-08, 1.842431e-08, 1.924944e-08, 2.130085e-08, 2.300331e-08, 
    2.371775e-08, 2.231813e-08, 1.986995e-08, 1.616062e-08, 1.062507e-08, 
    4.984879e-09, 1.965973e-09, 1.134155e-09, 8.147946e-10, 6.550398e-10,
  1.964625e-08, 1.892736e-08, 1.862222e-08, 2.028286e-08, 2.241142e-08, 
    2.383011e-08, 2.331326e-08, 2.120926e-08, 1.821613e-08, 1.361855e-08, 
    7.331867e-09, 2.973463e-09, 1.196701e-09, 9.861579e-10, 7.255355e-10,
  2.076442e-08, 1.933933e-08, 1.854578e-08, 1.939334e-08, 2.134482e-08, 
    2.321176e-08, 2.412907e-08, 2.245898e-08, 1.96836e-08, 1.592139e-08, 
    1.008585e-08, 4.483244e-09, 1.676712e-09, 1.152005e-09, 7.769845e-10,
  2.197988e-08, 2.000712e-08, 1.883916e-08, 1.896255e-08, 2.05557e-08, 
    2.251795e-08, 2.39915e-08, 2.379547e-08, 2.152719e-08, 1.793489e-08, 
    1.281111e-08, 6.446639e-09, 2.433171e-09, 1.268436e-09, 8.369649e-10,
  2.223424e-08, 2.035294e-08, 1.924413e-08, 1.885564e-08, 1.986246e-08, 
    2.169798e-08, 2.402982e-08, 2.422768e-08, 2.23994e-08, 1.923502e-08, 
    1.500157e-08, 8.815452e-09, 3.583068e-09, 1.399473e-09, 1.025068e-09,
  2.247595e-08, 2.078028e-08, 1.950701e-08, 1.880438e-08, 1.951331e-08, 
    2.122274e-08, 2.28903e-08, 2.428025e-08, 2.316248e-08, 2.050775e-08, 
    1.676893e-08, 1.113478e-08, 5.127315e-09, 1.782059e-09, 1.204443e-09,
  2.305244e-08, 2.161965e-08, 1.968311e-08, 1.74436e-08, 1.494563e-08, 
    1.122976e-08, 7.270035e-09, 4.313391e-09, 2.892731e-09, 2.057959e-09, 
    1.299468e-09, 1.056442e-09, 7.202761e-10, 4.300082e-10, 3.054845e-10,
  2.337341e-08, 2.278576e-08, 2.133134e-08, 1.903597e-08, 1.658916e-08, 
    1.366983e-08, 9.794762e-09, 6.089268e-09, 3.625017e-09, 2.670179e-09, 
    1.766373e-09, 1.225982e-09, 9.360994e-10, 5.624042e-10, 3.507144e-10,
  2.381951e-08, 2.315538e-08, 2.244242e-08, 2.067572e-08, 1.833935e-08, 
    1.576462e-08, 1.237253e-08, 8.33129e-09, 4.834679e-09, 3.13187e-09, 
    2.309925e-09, 1.488505e-09, 1.143628e-09, 7.440547e-10, 4.294014e-10,
  2.381834e-08, 2.342655e-08, 2.306775e-08, 2.18119e-08, 2.009034e-08, 
    1.752707e-08, 1.477444e-08, 1.086264e-08, 6.810145e-09, 3.833855e-09, 
    2.722633e-09, 1.919625e-09, 1.344394e-09, 9.804614e-10, 5.66811e-10,
  2.323277e-08, 2.340371e-08, 2.346787e-08, 2.271643e-08, 2.151374e-08, 
    1.925016e-08, 1.646645e-08, 1.338496e-08, 9.277825e-09, 5.475934e-09, 
    3.184968e-09, 2.366096e-09, 1.661258e-09, 1.19379e-09, 7.756731e-10,
  2.231788e-08, 2.306166e-08, 2.369531e-08, 2.312148e-08, 2.255691e-08, 
    2.084091e-08, 1.823961e-08, 1.510888e-08, 1.124484e-08, 7.335121e-09, 
    4.184274e-09, 2.702834e-09, 2.030748e-09, 1.437464e-09, 1.003368e-09,
  2.236765e-08, 2.237021e-08, 2.32404e-08, 2.34175e-08, 2.301744e-08, 
    2.203066e-08, 2.021996e-08, 1.727585e-08, 1.393539e-08, 9.513964e-09, 
    5.714448e-09, 3.302259e-09, 2.337098e-09, 1.731378e-09, 1.21511e-09,
  2.236526e-08, 2.217967e-08, 2.27948e-08, 2.308767e-08, 2.350808e-08, 
    2.25293e-08, 2.142875e-08, 1.893339e-08, 1.555419e-08, 1.184136e-08, 
    7.461233e-09, 4.376586e-09, 2.733118e-09, 2.019563e-09, 1.42531e-09,
  2.255605e-08, 2.182479e-08, 2.227453e-08, 2.29392e-08, 2.347346e-08, 
    2.306749e-08, 2.252038e-08, 2.05288e-08, 1.731322e-08, 1.353795e-08, 
    9.46899e-09, 5.787624e-09, 3.360633e-09, 2.308738e-09, 1.669519e-09,
  2.230047e-08, 2.171137e-08, 2.173455e-08, 2.275578e-08, 2.321186e-08, 
    2.300072e-08, 2.28388e-08, 2.175269e-08, 1.90218e-08, 1.563691e-08, 
    1.180423e-08, 7.514288e-09, 4.438566e-09, 2.721658e-09, 1.917142e-09,
  2.128055e-08, 1.786698e-08, 1.459363e-08, 1.175562e-08, 8.591649e-09, 
    5.563647e-09, 2.997669e-09, 1.497914e-09, 9.063282e-10, 7.33869e-10, 
    7.047277e-10, 6.093632e-10, 4.798636e-10, 4.027997e-10, 3.487756e-10,
  2.24518e-08, 1.991426e-08, 1.641597e-08, 1.323994e-08, 1.021287e-08, 
    7.019752e-09, 4.084062e-09, 2.053631e-09, 1.116794e-09, 8.135151e-10, 
    7.482545e-10, 6.797907e-10, 5.429312e-10, 4.498931e-10, 3.886566e-10,
  2.348231e-08, 2.157467e-08, 1.840796e-08, 1.487966e-08, 1.17754e-08, 
    8.629789e-09, 5.39767e-09, 2.820719e-09, 1.427167e-09, 9.360818e-10, 
    8.007525e-10, 7.370384e-10, 6.189682e-10, 4.964472e-10, 4.243643e-10,
  2.416775e-08, 2.294438e-08, 2.025915e-08, 1.674452e-08, 1.342963e-08, 
    1.036284e-08, 6.987687e-09, 3.932004e-09, 1.873183e-09, 1.078446e-09, 
    8.611414e-10, 7.828823e-10, 6.794555e-10, 5.540108e-10, 4.496351e-10,
  2.449844e-08, 2.356756e-08, 2.208977e-08, 1.875151e-08, 1.524241e-08, 
    1.202708e-08, 8.728765e-09, 5.446577e-09, 2.773438e-09, 1.348391e-09, 
    9.524782e-10, 8.354401e-10, 7.291663e-10, 6.138529e-10, 4.778611e-10,
  2.462466e-08, 2.384815e-08, 2.298185e-08, 2.062576e-08, 1.724664e-08, 
    1.39917e-08, 1.061603e-08, 7.042579e-09, 3.8693e-09, 1.823e-09, 
    1.072667e-09, 8.873962e-10, 7.746939e-10, 6.675664e-10, 5.310561e-10,
  2.512905e-08, 2.445488e-08, 2.364015e-08, 2.201508e-08, 1.90179e-08, 
    1.570703e-08, 1.253151e-08, 9.108477e-09, 5.527006e-09, 2.665694e-09, 
    1.270916e-09, 9.703873e-10, 8.268128e-10, 7.173289e-10, 5.948596e-10,
  2.558759e-08, 2.497193e-08, 2.42423e-08, 2.309761e-08, 2.089511e-08, 
    1.759277e-08, 1.408196e-08, 1.087036e-08, 7.61729e-09, 4.076413e-09, 
    1.68744e-09, 1.081666e-09, 8.987721e-10, 7.729331e-10, 6.545146e-10,
  2.555918e-08, 2.533653e-08, 2.472393e-08, 2.374905e-08, 2.240482e-08, 
    1.973992e-08, 1.6422e-08, 1.271513e-08, 9.002681e-09, 5.494331e-09, 
    2.544245e-09, 1.254155e-09, 9.858734e-10, 8.352307e-10, 7.150812e-10,
  2.611e-08, 2.55191e-08, 2.531698e-08, 2.468697e-08, 2.327295e-08, 
    2.143271e-08, 1.841526e-08, 1.47563e-08, 1.085745e-08, 7.275404e-09, 
    3.90567e-09, 1.716669e-09, 1.098509e-09, 9.100057e-10, 7.82532e-10,
  2.379919e-08, 2.259736e-08, 2.178818e-08, 2.068292e-08, 1.842812e-08, 
    1.472234e-08, 1.015678e-08, 5.842598e-09, 2.642107e-09, 9.952983e-10, 
    6.159777e-10, 6.605974e-10, 5.970938e-10, 4.501445e-10, 2.761973e-10,
  2.37996e-08, 2.284104e-08, 2.200123e-08, 2.09376e-08, 1.901521e-08, 
    1.57143e-08, 1.151666e-08, 7.091927e-09, 3.552642e-09, 1.380601e-09, 
    6.728488e-10, 6.27487e-10, 5.977965e-10, 4.954638e-10, 3.275072e-10,
  2.400469e-08, 2.286628e-08, 2.199086e-08, 2.113452e-08, 1.949682e-08, 
    1.652366e-08, 1.264144e-08, 8.314781e-09, 4.477855e-09, 1.903684e-09, 
    8.011067e-10, 6.083337e-10, 5.962866e-10, 5.004104e-10, 3.750498e-10,
  2.409407e-08, 2.299538e-08, 2.220428e-08, 2.123508e-08, 1.985541e-08, 
    1.717726e-08, 1.363501e-08, 9.430875e-09, 5.341247e-09, 2.46717e-09, 
    9.893308e-10, 6.42308e-10, 5.947989e-10, 4.945966e-10, 4.245697e-10,
  2.452942e-08, 2.347117e-08, 2.254983e-08, 2.142626e-08, 1.9984e-08, 
    1.762187e-08, 1.439219e-08, 1.053159e-08, 6.324831e-09, 3.117812e-09, 
    1.268187e-09, 7.039657e-10, 6.052711e-10, 4.944498e-10, 4.633548e-10,
  2.459615e-08, 2.360255e-08, 2.282165e-08, 2.166867e-08, 2.038635e-08, 
    1.80815e-08, 1.496251e-08, 1.135195e-08, 7.235863e-09, 3.799482e-09, 
    1.603372e-09, 7.960059e-10, 6.210303e-10, 5.014513e-10, 4.885231e-10,
  2.466904e-08, 2.376841e-08, 2.288649e-08, 2.182697e-08, 2.026814e-08, 
    1.835474e-08, 1.543347e-08, 1.201667e-08, 8.226045e-09, 4.552294e-09, 
    1.98328e-09, 8.940435e-10, 6.340697e-10, 5.08859e-10, 5.043423e-10,
  2.437268e-08, 2.357519e-08, 2.29207e-08, 2.187282e-08, 2.053265e-08, 
    1.853748e-08, 1.598282e-08, 1.296258e-08, 9.342846e-09, 5.385111e-09, 
    2.393901e-09, 1.008347e-09, 6.691127e-10, 5.175239e-10, 5.187003e-10,
  2.421748e-08, 2.357642e-08, 2.294006e-08, 2.194181e-08, 2.068084e-08, 
    1.911815e-08, 1.689684e-08, 1.389251e-08, 9.941369e-09, 6.070919e-09, 
    2.834173e-09, 1.156793e-09, 7.236305e-10, 5.494432e-10, 5.357457e-10,
  2.414744e-08, 2.360508e-08, 2.297277e-08, 2.219844e-08, 2.122245e-08, 
    1.950788e-08, 1.728483e-08, 1.431665e-08, 1.049748e-08, 6.805273e-09, 
    3.413243e-09, 1.381426e-09, 8.076341e-10, 5.984994e-10, 5.423911e-10,
  2.448744e-08, 2.365156e-08, 2.220861e-08, 1.868735e-08, 1.403247e-08, 
    9.179168e-09, 5.491718e-09, 3.131263e-09, 1.757172e-09, 1.244388e-09, 
    1.046463e-09, 8.573719e-10, 5.589481e-10, 3.593293e-10, 2.415933e-10,
  2.554749e-08, 2.460218e-08, 2.35081e-08, 2.124987e-08, 1.751612e-08, 
    1.223064e-08, 7.569516e-09, 4.302217e-09, 2.308338e-09, 1.353079e-09, 
    1.061967e-09, 9.282602e-10, 6.703132e-10, 4.330354e-10, 2.613639e-10,
  2.586742e-08, 2.521383e-08, 2.426245e-08, 2.307201e-08, 2.024856e-08, 
    1.517331e-08, 9.93596e-09, 5.946132e-09, 3.135674e-09, 1.642698e-09, 
    1.123622e-09, 9.800107e-10, 7.587304e-10, 5.119479e-10, 2.988036e-10,
  2.484975e-08, 2.489903e-08, 2.432999e-08, 2.390928e-08, 2.234115e-08, 
    1.814703e-08, 1.255466e-08, 7.701526e-09, 4.258672e-09, 2.144701e-09, 
    1.254871e-09, 1.04874e-09, 8.439991e-10, 5.900628e-10, 3.554405e-10,
  2.339417e-08, 2.489068e-08, 2.485924e-08, 2.447802e-08, 2.346319e-08, 
    2.072952e-08, 1.531581e-08, 9.742112e-09, 5.631871e-09, 2.867096e-09, 
    1.477918e-09, 1.123294e-09, 9.198379e-10, 6.698663e-10, 4.146365e-10,
  2.259934e-08, 2.349002e-08, 2.485863e-08, 2.516277e-08, 2.4358e-08, 
    2.281214e-08, 1.811371e-08, 1.219014e-08, 7.162814e-09, 3.79587e-09, 
    1.856075e-09, 1.221907e-09, 9.933723e-10, 7.532059e-10, 4.738529e-10,
  2.371464e-08, 2.339328e-08, 2.424438e-08, 2.555491e-08, 2.483103e-08, 
    2.408647e-08, 2.078832e-08, 1.526873e-08, 9.179969e-09, 4.882288e-09, 
    2.401774e-09, 1.354658e-09, 1.06713e-09, 8.401504e-10, 5.335085e-10,
  2.451029e-08, 2.365401e-08, 2.363207e-08, 2.501561e-08, 2.59534e-08, 
    2.495598e-08, 2.239673e-08, 1.727093e-08, 1.076505e-08, 5.922964e-09, 
    2.981316e-09, 1.528332e-09, 1.139399e-09, 9.275785e-10, 6.050755e-10,
  2.52878e-08, 2.393971e-08, 2.326517e-08, 2.457747e-08, 2.573396e-08, 
    2.540251e-08, 2.387314e-08, 1.915128e-08, 1.263717e-08, 7.069942e-09, 
    3.541079e-09, 1.71708e-09, 1.184786e-09, 1.006732e-09, 6.803248e-10,
  2.635547e-08, 2.485926e-08, 2.375474e-08, 2.411887e-08, 2.51944e-08, 
    2.507695e-08, 2.411376e-08, 2.084009e-08, 1.490818e-08, 8.41225e-09, 
    4.146278e-09, 1.916083e-09, 1.224204e-09, 1.077494e-09, 7.553427e-10,
  1.81515e-08, 1.358833e-08, 8.525696e-09, 4.274792e-09, 2.183171e-09, 
    1.59246e-09, 1.119902e-09, 8.83476e-10, 7.864164e-10, 7.741307e-10, 
    6.560701e-10, 5.367142e-10, 4.77952e-10, 4.659239e-10, 4.218502e-10,
  2.037503e-08, 1.692347e-08, 1.181394e-08, 6.578878e-09, 3.155377e-09, 
    1.89958e-09, 1.320605e-09, 9.534727e-10, 7.924346e-10, 7.580731e-10, 
    6.593562e-10, 5.342582e-10, 4.469288e-10, 4.362078e-10, 4.030509e-10,
  2.227688e-08, 1.915617e-08, 1.499051e-08, 9.562026e-09, 4.819268e-09, 
    2.475492e-09, 1.601495e-09, 1.099369e-09, 8.401814e-10, 7.668001e-10, 
    7.032866e-10, 5.77964e-10, 4.67865e-10, 4.2474e-10, 4.093202e-10,
  2.275275e-08, 2.095865e-08, 1.77679e-08, 1.296311e-08, 7.348543e-09, 
    3.6071e-09, 2.08558e-09, 1.345116e-09, 9.455732e-10, 7.873479e-10, 
    7.509934e-10, 6.41743e-10, 5.018581e-10, 3.976018e-10, 4.051406e-10,
  2.273694e-08, 2.230213e-08, 2.006335e-08, 1.628378e-08, 1.065398e-08, 
    5.533643e-09, 2.844759e-09, 1.747328e-09, 1.157212e-09, 8.469923e-10, 
    7.63983e-10, 6.898327e-10, 5.39679e-10, 3.75874e-10, 3.844176e-10,
  2.286195e-08, 2.329864e-08, 2.179148e-08, 1.900447e-08, 1.422261e-08, 
    8.56333e-09, 4.368303e-09, 2.392408e-09, 1.473453e-09, 9.72657e-10, 
    7.825108e-10, 7.343439e-10, 5.835333e-10, 3.909129e-10, 3.631005e-10,
  2.300564e-08, 2.36935e-08, 2.328153e-08, 2.083408e-08, 1.728074e-08, 
    1.181326e-08, 6.766654e-09, 3.614539e-09, 2.028024e-09, 1.206525e-09, 
    8.373384e-10, 7.716573e-10, 6.388255e-10, 4.311921e-10, 3.402361e-10,
  2.297561e-08, 2.330326e-08, 2.394079e-08, 2.281528e-08, 1.994863e-08, 
    1.522954e-08, 9.1583e-09, 4.721659e-09, 2.447878e-09, 1.450469e-09, 
    9.381081e-10, 7.910487e-10, 6.837675e-10, 4.821658e-10, 3.195338e-10,
  2.339389e-08, 2.299958e-08, 2.382014e-08, 2.371635e-08, 2.206826e-08, 
    1.793554e-08, 1.203495e-08, 6.331716e-09, 3.083495e-09, 1.737215e-09, 
    1.055073e-09, 7.903706e-10, 7.161239e-10, 5.341655e-10, 3.092844e-10,
  2.372018e-08, 2.305315e-08, 2.324284e-08, 2.420472e-08, 2.304745e-08, 
    2.01387e-08, 1.524167e-08, 8.961725e-09, 4.538859e-09, 2.329543e-09, 
    1.262701e-09, 8.229126e-10, 7.477216e-10, 5.773e-10, 3.100713e-10,
  1.633318e-08, 1.233416e-08, 7.394197e-09, 3.012179e-09, 1.085886e-09, 
    7.921033e-10, 7.698273e-10, 8.151539e-10, 8.617765e-10, 7.15192e-10, 
    6.775992e-10, 5.938179e-10, 5.240075e-10, 5.01951e-10, 6.461635e-10,
  1.812835e-08, 1.500413e-08, 1.03396e-08, 5.104553e-09, 1.769752e-09, 
    8.71527e-10, 7.838983e-10, 7.871937e-10, 8.528383e-10, 7.683824e-10, 
    6.744684e-10, 6.716184e-10, 6.604195e-10, 6.037128e-10, 7.239782e-10,
  1.948198e-08, 1.675835e-08, 1.303649e-08, 7.929145e-09, 3.146457e-09, 
    1.121148e-09, 8.185786e-10, 8.006464e-10, 8.310297e-10, 8.242007e-10, 
    6.629644e-10, 6.971928e-10, 6.334558e-10, 5.687517e-10, 6.444272e-10,
  2.072017e-08, 1.834886e-08, 1.545747e-08, 1.103414e-08, 5.398739e-09, 
    1.80515e-09, 8.913076e-10, 8.236392e-10, 8.204481e-10, 8.768664e-10, 
    6.629312e-10, 7.159121e-10, 5.603248e-10, 5.252475e-10, 5.829127e-10,
  2.095584e-08, 1.961592e-08, 1.757135e-08, 1.39519e-08, 8.268388e-09, 
    3.183276e-09, 1.120471e-09, 8.288075e-10, 8.154586e-10, 8.863277e-10, 
    6.957878e-10, 7.196356e-10, 5.611232e-10, 5.014204e-10, 5.600908e-10,
  2.220954e-08, 2.077484e-08, 1.910864e-08, 1.626857e-08, 1.128174e-08, 
    5.404996e-09, 1.771003e-09, 8.951544e-10, 8.471513e-10, 8.678726e-10, 
    7.632062e-10, 7.087803e-10, 6.138862e-10, 5.044585e-10, 5.458581e-10,
  2.383775e-08, 2.227136e-08, 2.028427e-08, 1.83357e-08, 1.410076e-08, 
    8.34095e-09, 3.156547e-09, 1.150857e-09, 9.176774e-10, 8.760018e-10, 
    8.437582e-10, 6.820559e-10, 6.807931e-10, 5.114872e-10, 5.399193e-10,
  2.457053e-08, 2.313891e-08, 2.120166e-08, 1.960899e-08, 1.694908e-08, 
    1.158866e-08, 5.155943e-09, 1.580804e-09, 9.257196e-10, 9.201674e-10, 
    8.980436e-10, 6.780198e-10, 7.245894e-10, 5.139423e-10, 5.252729e-10,
  2.498363e-08, 2.405553e-08, 2.213937e-08, 2.082718e-08, 1.906677e-08, 
    1.442565e-08, 7.838563e-09, 2.642444e-09, 9.729929e-10, 9.169547e-10, 
    9.143306e-10, 7.285513e-10, 7.336411e-10, 5.140831e-10, 5.076115e-10,
  2.55075e-08, 2.476521e-08, 2.319695e-08, 2.164089e-08, 2.017712e-08, 
    1.700268e-08, 1.093112e-08, 4.699023e-09, 1.388163e-09, 9.201104e-10, 
    9.144173e-10, 7.95054e-10, 7.13872e-10, 5.305641e-10, 4.836676e-10,
  1.906165e-08, 1.559086e-08, 1.126389e-08, 6.909842e-09, 3.332058e-09, 
    1.569853e-09, 1.044517e-09, 9.342944e-10, 7.453049e-10, 5.059448e-10, 
    3.49228e-10, 3.188641e-10, 6.484341e-10, 8.738822e-10, 7.963653e-10,
  1.998517e-08, 1.686755e-08, 1.252298e-08, 8.000178e-09, 4.039156e-09, 
    1.78097e-09, 1.080721e-09, 9.646777e-10, 8.397347e-10, 6.252366e-10, 
    4.299064e-10, 3.837049e-10, 6.678618e-10, 8.914989e-10, 8.010786e-10,
  2.068672e-08, 1.770342e-08, 1.384841e-08, 9.242979e-09, 4.896054e-09, 
    2.094169e-09, 1.154101e-09, 9.923297e-10, 9.000998e-10, 6.751242e-10, 
    4.456282e-10, 4.043708e-10, 6.472091e-10, 8.947816e-10, 7.639198e-10,
  2.113277e-08, 1.841836e-08, 1.489664e-08, 1.044792e-08, 5.860634e-09, 
    2.511497e-09, 1.252252e-09, 1.021584e-09, 9.539077e-10, 7.291454e-10, 
    4.566972e-10, 4.293509e-10, 6.404406e-10, 8.951465e-10, 7.198181e-10,
  2.14401e-08, 1.930863e-08, 1.604442e-08, 1.174437e-08, 6.897238e-09, 
    3.014717e-09, 1.35539e-09, 1.040565e-09, 1.010886e-09, 8.254658e-10, 
    4.914569e-10, 4.701919e-10, 6.691149e-10, 9.007318e-10, 6.739789e-10,
  2.167891e-08, 1.998006e-08, 1.707129e-08, 1.302476e-08, 8.016483e-09, 
    3.701553e-09, 1.498809e-09, 1.072743e-09, 1.036337e-09, 9.070647e-10, 
    5.268507e-10, 4.774059e-10, 7.089611e-10, 8.886152e-10, 6.240105e-10,
  2.240397e-08, 2.074671e-08, 1.810588e-08, 1.428288e-08, 9.196468e-09, 
    4.535472e-09, 1.755853e-09, 1.147186e-09, 1.080938e-09, 9.989906e-10, 
    5.617317e-10, 4.642257e-10, 7.347379e-10, 8.632825e-10, 5.76148e-10,
  2.312179e-08, 2.164957e-08, 1.900318e-08, 1.545927e-08, 1.055302e-08, 
    5.436804e-09, 2.006144e-09, 1.133308e-09, 1.083835e-09, 1.090237e-09, 
    6.160334e-10, 4.494674e-10, 7.588816e-10, 8.3267e-10, 5.391116e-10,
  2.297901e-08, 2.173867e-08, 1.965718e-08, 1.66329e-08, 1.196423e-08, 
    6.279913e-09, 2.406025e-09, 1.163807e-09, 1.077515e-09, 1.102588e-09, 
    6.984939e-10, 4.370823e-10, 7.792998e-10, 8.205619e-10, 5.226082e-10,
  2.358623e-08, 2.246355e-08, 2.03788e-08, 1.771507e-08, 1.323091e-08, 
    7.446588e-09, 3.002147e-09, 1.298654e-09, 1.129289e-09, 1.092158e-09, 
    7.832856e-10, 4.312153e-10, 7.838324e-10, 8.262633e-10, 5.208959e-10,
  1.932483e-08, 1.848075e-08, 1.742696e-08, 1.659094e-08, 1.477207e-08, 
    1.075936e-08, 6.061979e-09, 2.491522e-09, 1.24369e-09, 1.03859e-09, 
    1.02914e-09, 9.915261e-10, 6.428941e-10, 8.194394e-11, 1.119521e-10,
  2.012096e-08, 1.896311e-08, 1.773463e-08, 1.67851e-08, 1.576713e-08, 
    1.241219e-08, 7.658943e-09, 3.340974e-09, 1.381651e-09, 1.066249e-09, 
    1.034295e-09, 9.908273e-10, 6.06189e-10, -1.739642e-11, 1.933679e-12,
  2.03757e-08, 1.954441e-08, 1.807204e-08, 1.711908e-08, 1.64361e-08, 
    1.390928e-08, 9.310293e-09, 4.467927e-09, 1.625762e-09, 1.108861e-09, 
    1.052957e-09, 1.013059e-09, 5.709488e-10, -8.235543e-11, -7.817045e-11,
  1.937297e-08, 1.915393e-08, 1.816255e-08, 1.746578e-08, 1.675358e-08, 
    1.504721e-08, 1.087233e-08, 5.752091e-09, 2.128202e-09, 1.149385e-09, 
    1.072947e-09, 1.036005e-09, 5.355552e-10, -1.536126e-10, -1.622733e-10,
  1.89895e-08, 1.880727e-08, 1.819497e-08, 1.804983e-08, 1.714855e-08, 
    1.586402e-08, 1.241786e-08, 7.119078e-09, 2.833675e-09, 1.194438e-09, 
    1.090492e-09, 1.067936e-09, 5.099687e-10, -2.405784e-10, -2.542202e-10,
  1.925519e-08, 1.875897e-08, 1.863108e-08, 1.842489e-08, 1.746811e-08, 
    1.645791e-08, 1.357548e-08, 8.405515e-09, 3.609967e-09, 1.330028e-09, 
    1.100671e-09, 1.09895e-09, 4.94018e-10, -2.730966e-10, -3.110256e-10,
  1.997369e-08, 1.977178e-08, 1.931819e-08, 1.897957e-08, 1.785469e-08, 
    1.693065e-08, 1.461299e-08, 9.65574e-09, 4.371414e-09, 1.559517e-09, 
    1.11567e-09, 1.121606e-09, 4.866413e-10, -2.593801e-10, -3.567065e-10,
  2.052128e-08, 2.060992e-08, 1.968419e-08, 1.92861e-08, 1.821892e-08, 
    1.724431e-08, 1.525354e-08, 1.048343e-08, 4.863704e-09, 1.760259e-09, 
    1.155285e-09, 1.142641e-09, 4.774895e-10, -2.402621e-10, -3.584414e-10,
  2.048928e-08, 2.038889e-08, 1.986342e-08, 1.953122e-08, 1.861973e-08, 
    1.72342e-08, 1.574537e-08, 1.130815e-08, 5.639169e-09, 2.04278e-09, 
    1.194907e-09, 1.166137e-09, 4.607123e-10, -2.18836e-10, -3.256783e-10,
  2.06934e-08, 2.051191e-08, 2.012788e-08, 1.963781e-08, 1.894895e-08, 
    1.782331e-08, 1.602137e-08, 1.204936e-08, 6.43407e-09, 2.340353e-09, 
    1.220914e-09, 1.182733e-09, 4.304031e-10, -2.102937e-10, -2.734484e-10,
  1.887217e-08, 1.846986e-08, 1.807654e-08, 1.654508e-08, 1.381309e-08, 
    1.047089e-08, 7.199545e-09, 4.075426e-09, 1.796548e-09, 1.104247e-09, 
    8.93803e-10, 7.551184e-10, 5.324495e-10, 1.903641e-10, 3.942664e-10,
  1.917222e-08, 1.89069e-08, 1.846086e-08, 1.747826e-08, 1.529803e-08, 
    1.215441e-08, 8.720498e-09, 5.312028e-09, 2.333036e-09, 1.22997e-09, 
    9.469531e-10, 7.86589e-10, 5.739129e-10, 1.750494e-10, 3.323066e-10,
  1.930012e-08, 1.917008e-08, 1.875201e-08, 1.811467e-08, 1.65231e-08, 
    1.369143e-08, 1.029623e-08, 6.669449e-09, 3.198512e-09, 1.41405e-09, 
    1.009185e-09, 8.163873e-10, 6.16955e-10, 1.848643e-10, 3.467431e-10,
  1.907957e-08, 1.934707e-08, 1.90121e-08, 1.836902e-08, 1.75319e-08, 
    1.507524e-08, 1.182078e-08, 8.104753e-09, 4.26405e-09, 1.679777e-09, 
    1.076001e-09, 8.508725e-10, 6.52576e-10, 2.099102e-10, 3.611414e-10,
  1.896066e-08, 1.918161e-08, 1.905044e-08, 1.86294e-08, 1.820078e-08, 
    1.63769e-08, 1.334241e-08, 9.619748e-09, 5.510556e-09, 2.147665e-09, 
    1.161448e-09, 8.920873e-10, 6.784346e-10, 2.384559e-10, 3.718111e-10,
  1.936182e-08, 1.894122e-08, 1.92645e-08, 1.884156e-08, 1.861598e-08, 
    1.74668e-08, 1.46545e-08, 1.105919e-08, 6.833556e-09, 2.886034e-09, 
    1.26714e-09, 9.374882e-10, 7.061807e-10, 2.64305e-10, 3.726938e-10,
  2.005642e-08, 1.890143e-08, 1.922694e-08, 1.910619e-08, 1.876488e-08, 
    1.814607e-08, 1.598109e-08, 1.263717e-08, 8.183433e-09, 3.780701e-09, 
    1.412948e-09, 9.793336e-10, 7.365139e-10, 2.866568e-10, 3.452204e-10,
  2.091294e-08, 1.957418e-08, 1.899393e-08, 1.91061e-08, 1.911198e-08, 
    1.86598e-08, 1.675887e-08, 1.365548e-08, 9.230904e-09, 4.735836e-09, 
    1.646075e-09, 1.018586e-09, 7.670965e-10, 3.242032e-10, 3.14187e-10,
  2.15778e-08, 2.025911e-08, 1.900315e-08, 1.87856e-08, 1.89063e-08, 
    1.886961e-08, 1.721268e-08, 1.462428e-08, 1.075664e-08, 5.991224e-09, 
    2.046406e-09, 1.060215e-09, 7.960473e-10, 3.7419e-10, 2.932331e-10,
  2.20999e-08, 2.080136e-08, 1.953579e-08, 1.865915e-08, 1.848675e-08, 
    1.875769e-08, 1.777188e-08, 1.562844e-08, 1.202813e-08, 7.223333e-09, 
    2.576009e-09, 1.109646e-09, 8.257839e-10, 4.224888e-10, 2.657404e-10,
  1.937581e-08, 1.838781e-08, 1.752104e-08, 1.603255e-08, 1.336011e-08, 
    1.008348e-08, 8.223248e-09, 6.916084e-09, 5.662739e-09, 3.842214e-09, 
    1.747347e-09, 7.729419e-10, 8.900691e-10, 8.455519e-10, 5.673439e-10,
  2.078232e-08, 1.942595e-08, 1.844899e-08, 1.734794e-08, 1.540199e-08, 
    1.268164e-08, 9.539168e-09, 7.682786e-09, 6.373752e-09, 4.662124e-09, 
    2.61685e-09, 8.885628e-10, 8.6795e-10, 8.386274e-10, 5.263077e-10,
  2.209028e-08, 2.042591e-08, 1.934749e-08, 1.832528e-08, 1.68741e-08, 
    1.459414e-08, 1.174129e-08, 8.718082e-09, 7.116291e-09, 5.455678e-09, 
    3.53736e-09, 1.333202e-09, 8.250813e-10, 8.700113e-10, 5.867375e-10,
  2.239072e-08, 2.119962e-08, 1.980143e-08, 1.901063e-08, 1.813489e-08, 
    1.628518e-08, 1.408833e-08, 1.069683e-08, 8.245519e-09, 6.555194e-09, 
    4.808554e-09, 2.074187e-09, 7.595718e-10, 8.997612e-10, 6.506142e-10,
  2.235067e-08, 2.202352e-08, 2.074831e-08, 1.990511e-08, 1.910118e-08, 
    1.757338e-08, 1.575557e-08, 1.304769e-08, 1.001014e-08, 7.810208e-09, 
    5.967811e-09, 3.164448e-09, 8.651035e-10, 9.012417e-10, 6.998569e-10,
  2.268482e-08, 2.241655e-08, 2.155621e-08, 2.071383e-08, 1.997417e-08, 
    1.892261e-08, 1.717436e-08, 1.472849e-08, 1.140789e-08, 8.805626e-09, 
    6.874834e-09, 4.182282e-09, 1.194195e-09, 8.758687e-10, 7.473235e-10,
  2.330314e-08, 2.311056e-08, 2.206607e-08, 2.125238e-08, 2.053883e-08, 
    1.962371e-08, 1.846576e-08, 1.670451e-08, 1.348293e-08, 9.828153e-09, 
    7.560943e-09, 4.998094e-09, 1.70864e-09, 8.417047e-10, 7.814756e-10,
  2.354708e-08, 2.347924e-08, 2.263024e-08, 2.14233e-08, 2.105914e-08, 
    2.017349e-08, 1.881966e-08, 1.719044e-08, 1.473645e-08, 1.099724e-08, 
    8.227579e-09, 5.590299e-09, 2.250614e-09, 8.228865e-10, 7.921507e-10,
  2.375156e-08, 2.349865e-08, 2.296587e-08, 2.186814e-08, 2.130824e-08, 
    2.068575e-08, 1.934507e-08, 1.750523e-08, 1.584113e-08, 1.240009e-08, 
    9.188394e-09, 6.343364e-09, 2.890022e-09, 8.883162e-10, 7.905812e-10,
  2.41428e-08, 2.364668e-08, 2.324817e-08, 2.232736e-08, 2.11021e-08, 
    2.058168e-08, 1.987156e-08, 1.849262e-08, 1.726914e-08, 1.41288e-08, 
    1.039495e-08, 7.234194e-09, 3.619679e-09, 1.095087e-09, 7.80599e-10,
  1.706598e-08, 1.501969e-08, 1.248239e-08, 8.684378e-09, 5.771094e-09, 
    4.06157e-09, 3.159703e-09, 2.331153e-09, 1.806829e-09, 1.505586e-09, 
    1.176935e-09, 1.005863e-09, 9.448773e-10, 9.752888e-10, 9.253334e-10,
  1.832655e-08, 1.648281e-08, 1.451589e-08, 1.131032e-08, 7.419117e-09, 
    5.062365e-09, 3.759875e-09, 2.905726e-09, 2.123251e-09, 1.742909e-09, 
    1.306167e-09, 1.063931e-09, 9.472484e-10, 9.880928e-10, 1.003157e-09,
  1.971778e-08, 1.757295e-08, 1.58214e-08, 1.346345e-08, 9.773842e-09, 
    6.341484e-09, 4.472823e-09, 3.427035e-09, 2.59579e-09, 2.033932e-09, 
    1.540917e-09, 1.17984e-09, 9.524191e-10, 9.770328e-10, 1.03815e-09,
  2.098538e-08, 1.890849e-08, 1.697478e-08, 1.508059e-08, 1.203346e-08, 
    8.207316e-09, 5.602718e-09, 4.1167e-09, 3.101069e-09, 2.435429e-09, 
    1.883282e-09, 1.380768e-09, 9.959231e-10, 9.621089e-10, 1.0459e-09,
  2.166967e-08, 2.015813e-08, 1.852552e-08, 1.647791e-08, 1.396318e-08, 
    1.030776e-08, 7.031459e-09, 5.03221e-09, 3.725448e-09, 2.856145e-09, 
    2.266803e-09, 1.666323e-09, 1.126168e-09, 9.456803e-10, 1.041848e-09,
  2.300421e-08, 2.120456e-08, 1.969144e-08, 1.775373e-08, 1.568097e-08, 
    1.245574e-08, 8.722218e-09, 6.090474e-09, 4.406928e-09, 3.311756e-09, 
    2.679153e-09, 2.012988e-09, 1.343176e-09, 9.425765e-10, 1.037669e-09,
  2.361979e-08, 2.244797e-08, 2.058331e-08, 1.88682e-08, 1.708187e-08, 
    1.436945e-08, 1.077001e-08, 7.623205e-09, 5.495878e-09, 3.824581e-09, 
    3.017226e-09, 2.369268e-09, 1.613473e-09, 1.018555e-09, 1.016689e-09,
  2.402909e-08, 2.318533e-08, 2.17832e-08, 1.986379e-08, 1.834517e-08, 
    1.61505e-08, 1.280073e-08, 9.141105e-09, 6.554567e-09, 4.623772e-09, 
    3.4688e-09, 2.769365e-09, 1.911271e-09, 1.17881e-09, 9.841937e-10,
  2.424271e-08, 2.37277e-08, 2.255581e-08, 2.094632e-08, 1.939166e-08, 
    1.747221e-08, 1.482348e-08, 1.105493e-08, 7.884402e-09, 5.664124e-09, 
    4.091522e-09, 3.251848e-09, 2.289676e-09, 1.407556e-09, 9.448886e-10,
  2.449708e-08, 2.405717e-08, 2.313202e-08, 2.181435e-08, 2.046656e-08, 
    1.873433e-08, 1.638419e-08, 1.279327e-08, 9.232009e-09, 6.74667e-09, 
    4.861589e-09, 3.717397e-09, 2.74322e-09, 1.700356e-09, 9.525597e-10,
  1.884561e-08, 1.695338e-08, 1.442519e-08, 1.091857e-08, 5.982939e-09, 
    2.845258e-09, 1.524434e-09, 9.755474e-10, 7.084028e-10, 4.775795e-10, 
    3.205714e-10, 1.806501e-10, 1.147808e-10, 1.473539e-10, 1.987378e-10,
  2.005114e-08, 1.836746e-08, 1.620546e-08, 1.318357e-08, 8.482354e-09, 
    3.894728e-09, 1.908992e-09, 1.064998e-09, 7.436212e-10, 5.298902e-10, 
    3.66188e-10, 2.278676e-10, 1.291678e-10, 1.512946e-10, 2.092678e-10,
  2.1904e-08, 1.955823e-08, 1.748876e-08, 1.510022e-08, 1.109566e-08, 
    5.619734e-09, 2.533548e-09, 1.310988e-09, 8.330239e-10, 6.033995e-10, 
    4.141936e-10, 2.783345e-10, 1.472711e-10, 1.464426e-10, 2.191487e-10,
  2.312231e-08, 2.064511e-08, 1.859669e-08, 1.673518e-08, 1.343486e-08, 
    8.112123e-09, 3.565685e-09, 1.682433e-09, 9.614217e-10, 6.682049e-10, 
    4.519027e-10, 3.308241e-10, 1.760677e-10, 1.40567e-10, 2.315891e-10,
  2.431951e-08, 2.207437e-08, 1.959747e-08, 1.792755e-08, 1.548751e-08, 
    1.091528e-08, 5.15843e-09, 2.34254e-09, 1.187623e-09, 7.55694e-10, 
    5.079216e-10, 3.784836e-10, 2.256576e-10, 1.549693e-10, 2.369551e-10,
  2.501604e-08, 2.348348e-08, 2.084007e-08, 1.895087e-08, 1.720369e-08, 
    1.354682e-08, 7.362834e-09, 3.170534e-09, 1.473255e-09, 8.701082e-10, 
    5.92502e-10, 4.256794e-10, 2.682653e-10, 1.9584e-10, 2.453013e-10,
  2.609247e-08, 2.468937e-08, 2.228137e-08, 1.998603e-08, 1.837198e-08, 
    1.569202e-08, 1.020486e-08, 4.533954e-09, 1.993129e-09, 1.006817e-09, 
    6.582122e-10, 4.566345e-10, 2.960139e-10, 2.336878e-10, 2.504326e-10,
  2.672956e-08, 2.580651e-08, 2.384576e-08, 2.100137e-08, 1.93285e-08, 
    1.737855e-08, 1.258363e-08, 6.018638e-09, 2.606207e-09, 1.200717e-09, 
    7.186891e-10, 4.918801e-10, 3.275627e-10, 2.400959e-10, 2.443796e-10,
  2.630657e-08, 2.633715e-08, 2.49541e-08, 2.233928e-08, 2.000406e-08, 
    1.854548e-08, 1.474932e-08, 8.141762e-09, 3.451198e-09, 1.46434e-09, 
    7.93781e-10, 5.41142e-10, 3.465906e-10, 2.572987e-10, 2.455897e-10,
  2.590955e-08, 2.65752e-08, 2.573154e-08, 2.353714e-08, 2.076827e-08, 
    1.93232e-08, 1.648701e-08, 1.069212e-08, 4.809634e-09, 1.941472e-09, 
    9.334018e-10, 6.067304e-10, 3.852635e-10, 2.674949e-10, 2.52656e-10,
  1.394308e-08, 1.167153e-08, 9.756072e-09, 8.511109e-09, 7.473016e-09, 
    5.480177e-09, 3.786686e-09, 2.780371e-09, 2.21696e-09, 1.925577e-09, 
    1.588744e-09, 9.744716e-10, 2.775656e-10, 3.613117e-11, 8.070768e-11,
  1.516318e-08, 1.315279e-08, 1.085115e-08, 9.295503e-09, 8.16374e-09, 
    6.447363e-09, 4.529499e-09, 3.226572e-09, 2.441159e-09, 2.054109e-09, 
    1.734872e-09, 1.210648e-09, 4.554884e-10, 7.50013e-11, 6.208568e-11,
  1.639331e-08, 1.474826e-08, 1.224782e-08, 1.004191e-08, 8.765564e-09, 
    7.414099e-09, 5.296624e-09, 3.715848e-09, 2.785124e-09, 2.176771e-09, 
    1.845821e-09, 1.430469e-09, 6.626866e-10, 1.235523e-10, 3.968161e-11,
  1.771658e-08, 1.624882e-08, 1.397749e-08, 1.096308e-08, 9.461107e-09, 
    8.309827e-09, 6.240619e-09, 4.316709e-09, 3.118461e-09, 2.335753e-09, 
    1.941823e-09, 1.621014e-09, 8.924436e-10, 2.246598e-10, 3.709489e-11,
  1.929942e-08, 1.763703e-08, 1.547753e-08, 1.226692e-08, 1.021143e-08, 
    8.91247e-09, 7.173062e-09, 5.13704e-09, 3.594406e-09, 2.638949e-09, 
    2.049161e-09, 1.771381e-09, 1.142303e-09, 3.507128e-10, 5.903202e-11,
  2.011448e-08, 1.85771e-08, 1.668048e-08, 1.377265e-08, 1.116931e-08, 
    9.687226e-09, 8.103229e-09, 5.88921e-09, 4.064947e-09, 2.933769e-09, 
    2.120062e-09, 1.849601e-09, 1.356624e-09, 5.167038e-10, 9.628096e-11,
  2.146234e-08, 1.94799e-08, 1.763402e-08, 1.526664e-08, 1.236676e-08, 
    1.041035e-08, 8.959554e-09, 6.889001e-09, 4.858524e-09, 3.335632e-09, 
    2.212724e-09, 1.861752e-09, 1.532431e-09, 7.107426e-10, 1.554353e-10,
  2.276149e-08, 2.063497e-08, 1.878972e-08, 1.663697e-08, 1.400283e-08, 
    1.146438e-08, 9.74736e-09, 7.737317e-09, 5.720615e-09, 3.833418e-09, 
    2.350133e-09, 1.818294e-09, 1.642772e-09, 9.357604e-10, 2.517282e-10,
  2.335583e-08, 2.164846e-08, 1.966212e-08, 1.77824e-08, 1.541505e-08, 
    1.274035e-08, 1.077306e-08, 8.846524e-09, 6.484704e-09, 4.320215e-09, 
    2.579373e-09, 1.822863e-09, 1.73027e-09, 1.146602e-09, 3.855803e-10,
  2.35881e-08, 2.254641e-08, 2.050762e-08, 1.87433e-08, 1.680432e-08, 
    1.422089e-08, 1.17754e-08, 9.789442e-09, 7.239341e-09, 5.142955e-09, 
    3.02399e-09, 1.929495e-09, 1.804672e-09, 1.336593e-09, 5.596802e-10,
  9.116494e-09, 8.289496e-09, 7.017746e-09, 5.360684e-09, 3.80756e-09, 
    2.506705e-09, 1.849461e-09, 1.627532e-09, 1.482752e-09, 1.426558e-09, 
    1.273767e-09, 9.492175e-10, 5.246009e-10, 2.850565e-10, 3.438374e-10,
  9.611529e-09, 8.92419e-09, 7.898495e-09, 6.320034e-09, 4.65273e-09, 
    3.132101e-09, 2.161863e-09, 1.783242e-09, 1.617092e-09, 1.507161e-09, 
    1.397057e-09, 1.107716e-09, 6.2747e-10, 3.236916e-10, 2.888676e-10,
  1.033118e-08, 9.482148e-09, 8.693967e-09, 7.238896e-09, 5.553412e-09, 
    3.891094e-09, 2.577205e-09, 1.999338e-09, 1.774631e-09, 1.62031e-09, 
    1.493838e-09, 1.290139e-09, 7.756683e-10, 3.806101e-10, 2.626241e-10,
  1.095386e-08, 1.011053e-08, 9.281065e-09, 8.09059e-09, 6.504257e-09, 
    4.837611e-09, 3.213694e-09, 2.259955e-09, 1.868917e-09, 1.717839e-09, 
    1.566643e-09, 1.448387e-09, 9.894597e-10, 4.623997e-10, 2.631308e-10,
  1.19559e-08, 1.086544e-08, 9.845824e-09, 8.860992e-09, 7.437196e-09, 
    5.795465e-09, 4.006131e-09, 2.747765e-09, 2.099132e-09, 1.812565e-09, 
    1.631287e-09, 1.544784e-09, 1.228206e-09, 5.868572e-10, 2.820116e-10,
  1.318401e-08, 1.161812e-08, 1.050402e-08, 9.496174e-09, 8.280641e-09, 
    6.837621e-09, 4.984026e-09, 3.257387e-09, 2.285304e-09, 1.877852e-09, 
    1.670567e-09, 1.592122e-09, 1.437389e-09, 7.709229e-10, 3.262527e-10,
  1.515896e-08, 1.247524e-08, 1.109715e-08, 1.013962e-08, 9.050465e-09, 
    7.583948e-09, 5.979956e-09, 4.172657e-09, 2.804202e-09, 2.079616e-09, 
    1.750308e-09, 1.626337e-09, 1.57184e-09, 1.013369e-09, 4.066877e-10,
  1.729283e-08, 1.428604e-08, 1.190434e-08, 1.071532e-08, 9.76144e-09, 
    8.449209e-09, 6.819314e-09, 4.995996e-09, 3.452217e-09, 2.409366e-09, 
    1.845251e-09, 1.66832e-09, 1.642459e-09, 1.281701e-09, 5.337287e-10,
  1.894528e-08, 1.653245e-08, 1.345161e-08, 1.142936e-08, 1.03621e-08, 
    9.370031e-09, 8.069867e-09, 6.151952e-09, 4.090747e-09, 2.719252e-09, 
    1.996614e-09, 1.708006e-09, 1.65618e-09, 1.505415e-09, 7.195526e-10,
  2.050122e-08, 1.855909e-08, 1.551586e-08, 1.268586e-08, 1.109866e-08, 
    1.022064e-08, 8.933884e-09, 7.068692e-09, 4.919006e-09, 3.334933e-09, 
    2.336402e-09, 1.755452e-09, 1.633821e-09, 1.645622e-09, 9.547028e-10,
  6.234702e-09, 5.212128e-09, 4.075177e-09, 3.045429e-09, 2.387926e-09, 
    2.04359e-09, 1.86279e-09, 1.873444e-09, 1.92945e-09, 1.804413e-09, 
    1.45012e-09, 9.137062e-10, 4.086503e-10, 1.962618e-10, 2.310359e-10,
  6.250158e-09, 5.50244e-09, 4.5336e-09, 3.360061e-09, 2.431146e-09, 
    1.970566e-09, 1.812317e-09, 1.861874e-09, 1.945609e-09, 1.843431e-09, 
    1.511886e-09, 9.738393e-10, 4.65675e-10, 3.034186e-10, 3.880979e-10,
  6.470568e-09, 5.851974e-09, 4.996082e-09, 3.694956e-09, 2.589361e-09, 
    2.019124e-09, 1.856949e-09, 1.880394e-09, 1.983913e-09, 1.914419e-09, 
    1.606861e-09, 1.084059e-09, 5.523471e-10, 3.777096e-10, 4.354225e-10,
  6.862612e-09, 6.286727e-09, 5.448867e-09, 4.181939e-09, 3.040833e-09, 
    2.275208e-09, 1.961879e-09, 1.876164e-09, 1.932458e-09, 1.928122e-09, 
    1.713793e-09, 1.240516e-09, 6.73552e-10, 4.14765e-10, 3.816955e-10,
  7.814995e-09, 6.860756e-09, 5.857736e-09, 4.725058e-09, 3.5844e-09, 
    2.606371e-09, 2.078351e-09, 1.819976e-09, 1.796838e-09, 1.850523e-09, 
    1.775124e-09, 1.410588e-09, 8.095907e-10, 4.085298e-10, 2.56683e-10,
  8.585768e-09, 7.419894e-09, 6.249192e-09, 5.079682e-09, 4.084985e-09, 
    3.038221e-09, 2.284486e-09, 1.732011e-09, 1.572567e-09, 1.731701e-09, 
    1.821488e-09, 1.563865e-09, 9.698703e-10, 4.300886e-10, 1.765858e-10,
  8.705635e-09, 7.660257e-09, 6.538075e-09, 5.501803e-09, 4.388866e-09, 
    3.230329e-09, 2.36875e-09, 1.793325e-09, 1.576728e-09, 1.732308e-09, 
    1.922286e-09, 1.697952e-09, 1.136202e-09, 5.3134e-10, 1.869769e-10,
  9.40634e-09, 8.242942e-09, 7.027425e-09, 5.797819e-09, 4.721345e-09, 
    3.492944e-09, 2.502529e-09, 1.918822e-09, 1.804378e-09, 1.848844e-09, 
    1.995177e-09, 1.81308e-09, 1.273506e-09, 6.770437e-10, 2.836635e-10,
  1.056618e-08, 8.912562e-09, 7.664209e-09, 6.017487e-09, 5.073256e-09, 
    4.241447e-09, 3.141913e-09, 2.188287e-09, 1.780108e-09, 1.801888e-09, 
    1.998597e-09, 1.8481e-09, 1.356479e-09, 8.150955e-10, 4.062096e-10,
  1.253415e-08, 9.90256e-09, 8.367529e-09, 6.702611e-09, 5.549418e-09, 
    4.736335e-09, 3.702006e-09, 2.532355e-09, 1.891217e-09, 1.834438e-09, 
    2.002033e-09, 1.921918e-09, 1.445104e-09, 9.415683e-10, 5.387697e-10,
  1.471912e-08, 1.345085e-08, 1.260175e-08, 1.18007e-08, 1.055912e-08, 
    9.301526e-09, 8.101148e-09, 7.05237e-09, 6.22705e-09, 5.40584e-09, 
    4.738173e-09, 4.417998e-09, 3.962121e-09, 3.592027e-09, 3.000502e-09,
  1.448984e-08, 1.350616e-08, 1.27079e-08, 1.179729e-08, 1.0457e-08, 
    9.157536e-09, 7.937342e-09, 6.908876e-09, 6.082428e-09, 5.251559e-09, 
    4.660619e-09, 4.33175e-09, 3.828725e-09, 3.451036e-09, 2.902522e-09,
  1.425321e-08, 1.343813e-08, 1.270511e-08, 1.167094e-08, 1.020474e-08, 
    8.891021e-09, 7.739972e-09, 6.794662e-09, 5.999473e-09, 5.166268e-09, 
    4.572324e-09, 4.220025e-09, 3.679559e-09, 3.278569e-09, 2.8135e-09,
  1.440961e-08, 1.378854e-08, 1.293285e-08, 1.161318e-08, 1.006529e-08, 
    8.704656e-09, 7.603152e-09, 6.692124e-09, 5.923378e-09, 5.138111e-09, 
    4.513145e-09, 4.137425e-09, 3.560306e-09, 3.193723e-09, 2.824519e-09,
  1.502095e-08, 1.415517e-08, 1.311423e-08, 1.159873e-08, 9.889519e-09, 
    8.550289e-09, 7.572978e-09, 6.703949e-09, 5.941623e-09, 5.132201e-09, 
    4.479833e-09, 4.097157e-09, 3.494514e-09, 3.143601e-09, 2.821709e-09,
  1.584317e-08, 1.453445e-08, 1.305789e-08, 1.146843e-08, 9.904609e-09, 
    8.460041e-09, 7.448858e-09, 6.514389e-09, 5.782192e-09, 5.084997e-09, 
    4.49035e-09, 4.080685e-09, 3.442105e-09, 3.116705e-09, 2.810549e-09,
  1.575466e-08, 1.399812e-08, 1.266437e-08, 1.128464e-08, 9.611686e-09, 
    8.262365e-09, 7.347503e-09, 6.421157e-09, 5.743261e-09, 5.107281e-09, 
    4.477066e-09, 4.005101e-09, 3.367502e-09, 3.094153e-09, 2.773718e-09,
  1.554718e-08, 1.393851e-08, 1.262969e-08, 1.108571e-08, 9.366895e-09, 
    8.085054e-09, 7.312155e-09, 6.530924e-09, 5.908525e-09, 5.175098e-09, 
    4.43662e-09, 3.869501e-09, 3.247143e-09, 3.050136e-09, 2.717823e-09,
  1.587111e-08, 1.417003e-08, 1.261025e-08, 1.07452e-08, 9.183685e-09, 
    8.409067e-09, 7.575713e-09, 6.617528e-09, 5.779536e-09, 5.082233e-09, 
    4.399694e-09, 3.745914e-09, 3.104149e-09, 2.980483e-09, 2.639619e-09,
  1.625854e-08, 1.452994e-08, 1.255716e-08, 1.06891e-08, 9.340215e-09, 
    8.430137e-09, 7.589924e-09, 6.499258e-09, 5.465802e-09, 4.904712e-09, 
    4.378934e-09, 3.657432e-09, 2.966896e-09, 2.889921e-09, 2.532674e-09,
  2.476609e-08, 2.190546e-08, 1.942233e-08, 1.690175e-08, 1.401477e-08, 
    1.121471e-08, 8.829619e-09, 6.836276e-09, 5.301947e-09, 3.80903e-09, 
    2.899191e-09, 2.505362e-09, 2.246853e-09, 1.817627e-09, 1.35211e-09,
  2.533842e-08, 2.316494e-08, 2.022748e-08, 1.759187e-08, 1.480539e-08, 
    1.192282e-08, 9.349468e-09, 7.2355e-09, 5.630743e-09, 4.065055e-09, 
    3.035623e-09, 2.579764e-09, 2.361029e-09, 1.969544e-09, 1.500425e-09,
  2.560982e-08, 2.3973e-08, 2.11723e-08, 1.832934e-08, 1.54882e-08, 
    1.261679e-08, 9.920193e-09, 7.676831e-09, 5.984509e-09, 4.329704e-09, 
    3.175927e-09, 2.654819e-09, 2.458606e-09, 2.080175e-09, 1.55581e-09,
  2.573458e-08, 2.437205e-08, 2.203072e-08, 1.912588e-08, 1.618576e-08, 
    1.329283e-08, 1.047524e-08, 8.084474e-09, 6.324001e-09, 4.619511e-09, 
    3.353282e-09, 2.763605e-09, 2.576747e-09, 2.219368e-09, 1.672981e-09,
  2.525628e-08, 2.453607e-08, 2.272523e-08, 1.99295e-08, 1.683603e-08, 
    1.383565e-08, 1.106171e-08, 8.569783e-09, 6.718963e-09, 4.939584e-09, 
    3.571769e-09, 2.884511e-09, 2.683574e-09, 2.378243e-09, 1.810633e-09,
  2.443666e-08, 2.432036e-08, 2.307844e-08, 2.071701e-08, 1.760621e-08, 
    1.447984e-08, 1.146777e-08, 8.9302e-09, 7.064757e-09, 5.26419e-09, 
    3.765977e-09, 2.96748e-09, 2.749897e-09, 2.529304e-09, 1.967935e-09,
  2.423994e-08, 2.445903e-08, 2.35215e-08, 2.136631e-08, 1.820864e-08, 
    1.501336e-08, 1.207037e-08, 9.353093e-09, 7.379257e-09, 5.569616e-09, 
    3.949309e-09, 3.034684e-09, 2.793214e-09, 2.662738e-09, 2.139732e-09,
  2.414349e-08, 2.435114e-08, 2.372136e-08, 2.193161e-08, 1.905026e-08, 
    1.557579e-08, 1.243399e-08, 9.781972e-09, 7.872631e-09, 5.924439e-09, 
    4.121041e-09, 3.088712e-09, 2.830479e-09, 2.797787e-09, 2.30007e-09,
  2.381026e-08, 2.408049e-08, 2.372048e-08, 2.236827e-08, 1.960925e-08, 
    1.633539e-08, 1.313986e-08, 1.022851e-08, 8.133149e-09, 6.096014e-09, 
    4.307333e-09, 3.192145e-09, 2.914342e-09, 2.940001e-09, 2.451393e-09,
  2.358059e-08, 2.380061e-08, 2.362237e-08, 2.267255e-08, 2.014178e-08, 
    1.702444e-08, 1.367027e-08, 1.058419e-08, 8.297145e-09, 6.371088e-09, 
    4.602812e-09, 3.331437e-09, 3.043173e-09, 3.105183e-09, 2.624286e-09,
  1.968398e-08, 1.653058e-08, 1.372076e-08, 1.143323e-08, 9.710058e-09, 
    8.127416e-09, 6.50848e-09, 4.992852e-09, 3.910879e-09, 3.001855e-09, 
    2.201565e-09, 1.554942e-09, 9.346905e-10, 6.943512e-10, 5.273352e-10,
  2.037381e-08, 1.754346e-08, 1.439656e-08, 1.189963e-08, 1.006538e-08, 
    8.496873e-09, 6.853492e-09, 5.254296e-09, 4.081736e-09, 3.1453e-09, 
    2.305108e-09, 1.643263e-09, 9.815229e-10, 7.18928e-10, 5.693898e-10,
  2.100859e-08, 1.835125e-08, 1.514164e-08, 1.236069e-08, 1.039829e-08, 
    8.79926e-09, 7.177627e-09, 5.520193e-09, 4.248648e-09, 3.28564e-09, 
    2.402559e-09, 1.721732e-09, 1.024614e-09, 7.368158e-10, 5.989595e-10,
  2.197924e-08, 1.925236e-08, 1.607241e-08, 1.291929e-08, 1.076313e-08, 
    9.142697e-09, 7.505668e-09, 5.784036e-09, 4.435336e-09, 3.438672e-09, 
    2.51668e-09, 1.806123e-09, 1.084604e-09, 7.574234e-10, 6.412634e-10,
  2.315732e-08, 2.015116e-08, 1.696889e-08, 1.362985e-08, 1.113918e-08, 
    9.422339e-09, 7.864126e-09, 6.159497e-09, 4.707665e-09, 3.647756e-09, 
    2.66735e-09, 1.896332e-09, 1.164733e-09, 7.857306e-10, 6.85576e-10,
  2.420889e-08, 2.101125e-08, 1.790363e-08, 1.436411e-08, 1.164295e-08, 
    9.775729e-09, 8.183785e-09, 6.461189e-09, 4.922917e-09, 3.815539e-09, 
    2.769961e-09, 1.965965e-09, 1.231728e-09, 8.145291e-10, 7.166515e-10,
  2.502975e-08, 2.182936e-08, 1.864029e-08, 1.520998e-08, 1.208544e-08, 
    1.00663e-08, 8.496548e-09, 6.796906e-09, 5.186124e-09, 4.021441e-09, 
    2.871369e-09, 2.02297e-09, 1.296857e-09, 8.44674e-10, 7.308362e-10,
  2.563327e-08, 2.276185e-08, 1.952642e-08, 1.604975e-08, 1.283362e-08, 
    1.036032e-08, 8.789935e-09, 7.205878e-09, 5.601144e-09, 4.277314e-09, 
    2.999915e-09, 2.102083e-09, 1.3835e-09, 8.934596e-10, 7.612543e-10,
  2.633856e-08, 2.373927e-08, 2.042607e-08, 1.691547e-08, 1.354734e-08, 
    1.090276e-08, 9.329104e-09, 7.659558e-09, 5.897294e-09, 4.430849e-09, 
    3.125501e-09, 2.187002e-09, 1.473803e-09, 9.54867e-10, 8.078866e-10,
  2.658956e-08, 2.484426e-08, 2.143285e-08, 1.788056e-08, 1.441342e-08, 
    1.137921e-08, 9.644987e-09, 7.986453e-09, 6.129364e-09, 4.593599e-09, 
    3.253895e-09, 2.263392e-09, 1.568872e-09, 1.027914e-09, 8.588586e-10,
  2.374435e-08, 2.237984e-08, 2.097856e-08, 1.979354e-08, 1.807732e-08, 
    1.609334e-08, 1.398632e-08, 1.10167e-08, 7.591197e-09, 5.031903e-09, 
    3.752922e-09, 2.620715e-09, 1.71598e-09, 1.289064e-09, 1.092194e-09,
  2.414943e-08, 2.30091e-08, 2.146916e-08, 2.022654e-08, 1.874502e-08, 
    1.678573e-08, 1.472102e-08, 1.208658e-08, 8.691977e-09, 5.671558e-09, 
    4.094924e-09, 2.972632e-09, 2.008891e-09, 1.439525e-09, 1.172162e-09,
  2.463012e-08, 2.337221e-08, 2.184062e-08, 2.048669e-08, 1.923702e-08, 
    1.7341e-08, 1.541616e-08, 1.293218e-08, 9.796262e-09, 6.41356e-09, 
    4.450289e-09, 3.273056e-09, 2.246058e-09, 1.577633e-09, 1.236639e-09,
  2.46304e-08, 2.376994e-08, 2.233943e-08, 2.086157e-08, 1.960763e-08, 
    1.783062e-08, 1.594097e-08, 1.364861e-08, 1.070959e-08, 7.299729e-09, 
    4.861988e-09, 3.565109e-09, 2.476303e-09, 1.722678e-09, 1.296465e-09,
  2.487947e-08, 2.419109e-08, 2.283892e-08, 2.106373e-08, 1.981269e-08, 
    1.811945e-08, 1.640436e-08, 1.424312e-08, 1.152971e-08, 8.173076e-09, 
    5.323673e-09, 3.874589e-09, 2.708668e-09, 1.882943e-09, 1.369666e-09,
  2.444992e-08, 2.426882e-08, 2.327561e-08, 2.148921e-08, 2.005449e-08, 
    1.846948e-08, 1.658757e-08, 1.45725e-08, 1.202308e-08, 8.975809e-09, 
    5.866905e-09, 4.206747e-09, 2.928661e-09, 2.043116e-09, 1.461068e-09,
  2.376652e-08, 2.404934e-08, 2.343895e-08, 2.181821e-08, 2.023449e-08, 
    1.873738e-08, 1.711986e-08, 1.518305e-08, 1.270284e-08, 9.666286e-09, 
    6.51895e-09, 4.53984e-09, 3.169338e-09, 2.195645e-09, 1.566492e-09,
  2.325995e-08, 2.394128e-08, 2.371629e-08, 2.21726e-08, 2.061074e-08, 
    1.905167e-08, 1.73341e-08, 1.533794e-08, 1.304587e-08, 1.026047e-08, 
    7.22618e-09, 4.903126e-09, 3.435323e-09, 2.351412e-09, 1.668116e-09,
  2.272088e-08, 2.377459e-08, 2.384413e-08, 2.24331e-08, 2.084051e-08, 
    1.913527e-08, 1.747168e-08, 1.573296e-08, 1.36221e-08, 1.088073e-08, 
    7.844539e-09, 5.307115e-09, 3.716801e-09, 2.500622e-09, 1.753901e-09,
  2.220496e-08, 2.362001e-08, 2.395786e-08, 2.27175e-08, 2.122205e-08, 
    1.948531e-08, 1.75293e-08, 1.583212e-08, 1.39175e-08, 1.134958e-08, 
    8.375569e-09, 5.721845e-09, 3.97979e-09, 2.656356e-09, 1.823995e-09,
  1.989038e-08, 1.840118e-08, 1.69144e-08, 1.491984e-08, 1.247527e-08, 
    1.010652e-08, 8.266106e-09, 6.57556e-09, 4.972443e-09, 3.706846e-09, 
    2.918705e-09, 2.278669e-09, 1.71733e-09, 1.303818e-09, 1.074336e-09,
  2.078528e-08, 1.95966e-08, 1.811276e-08, 1.623945e-08, 1.413148e-08, 
    1.163065e-08, 9.521431e-09, 7.670084e-09, 5.858377e-09, 4.298858e-09, 
    3.277294e-09, 2.554301e-09, 1.922126e-09, 1.414361e-09, 1.122038e-09,
  2.157065e-08, 2.060999e-08, 1.925415e-08, 1.739754e-08, 1.534478e-08, 
    1.312952e-08, 1.081235e-08, 8.79301e-09, 6.916719e-09, 5.096174e-09, 
    3.779356e-09, 2.882934e-09, 2.146826e-09, 1.58413e-09, 1.233183e-09,
  2.253436e-08, 2.159385e-08, 2.019817e-08, 1.85283e-08, 1.671871e-08, 
    1.44716e-08, 1.226573e-08, 1.001092e-08, 7.962565e-09, 5.934321e-09, 
    4.349541e-09, 3.273331e-09, 2.415275e-09, 1.788043e-09, 1.362338e-09,
  2.303739e-08, 2.23571e-08, 2.098907e-08, 1.945894e-08, 1.794507e-08, 
    1.582926e-08, 1.355221e-08, 1.135574e-08, 9.25935e-09, 7.038426e-09, 
    5.045307e-09, 3.704559e-09, 2.73252e-09, 2.018661e-09, 1.498937e-09,
  2.326226e-08, 2.271001e-08, 2.190873e-08, 2.039493e-08, 1.895118e-08, 
    1.733861e-08, 1.502394e-08, 1.258246e-08, 1.025528e-08, 8.058954e-09, 
    5.839514e-09, 4.193359e-09, 3.078602e-09, 2.289199e-09, 1.686257e-09,
  2.368462e-08, 2.29655e-08, 2.243877e-08, 2.144007e-08, 1.978508e-08, 
    1.834011e-08, 1.652393e-08, 1.432791e-08, 1.179828e-08, 9.318119e-09, 
    6.829456e-09, 4.796171e-09, 3.461231e-09, 2.564378e-09, 1.935422e-09,
  2.36001e-08, 2.325826e-08, 2.27931e-08, 2.215179e-08, 2.097107e-08, 
    1.928959e-08, 1.74216e-08, 1.520538e-08, 1.294254e-08, 1.052261e-08, 
    7.966982e-09, 5.557752e-09, 3.924429e-09, 2.851163e-09, 2.198229e-09,
  2.355508e-08, 2.348446e-08, 2.300225e-08, 2.247478e-08, 2.178175e-08, 
    2.047883e-08, 1.864004e-08, 1.63564e-08, 1.408907e-08, 1.167459e-08, 
    9.130694e-09, 6.466768e-09, 4.460277e-09, 3.174975e-09, 2.431436e-09,
  2.323755e-08, 2.350674e-08, 2.326032e-08, 2.274828e-08, 2.200894e-08, 
    2.107602e-08, 1.964544e-08, 1.762916e-08, 1.542432e-08, 1.290839e-08, 
    1.029943e-08, 7.475757e-09, 5.106345e-09, 3.53094e-09, 2.639723e-09,
  1.404288e-08, 1.13823e-08, 9.123327e-09, 6.433266e-09, 4.420617e-09, 
    3.177488e-09, 2.527274e-09, 2.17666e-09, 1.773064e-09, 1.280586e-09, 
    9.249361e-10, 7.799595e-10, 7.448858e-10, 7.955119e-10, 8.141158e-10,
  1.496233e-08, 1.260309e-08, 1.020657e-08, 7.614334e-09, 5.332212e-09, 
    3.67291e-09, 2.795959e-09, 2.309622e-09, 1.92166e-09, 1.419363e-09, 
    9.48117e-10, 7.519479e-10, 7.637433e-10, 8.482838e-10, 8.385493e-10,
  1.622354e-08, 1.40394e-08, 1.13844e-08, 8.628048e-09, 6.325634e-09, 
    4.420768e-09, 3.217624e-09, 2.51341e-09, 2.019225e-09, 1.540373e-09, 
    1.074552e-09, 8.190483e-10, 8.474252e-10, 9.347615e-10, 8.848567e-10,
  1.757175e-08, 1.554787e-08, 1.27618e-08, 9.690266e-09, 7.333572e-09, 
    5.263209e-09, 3.811178e-09, 2.801967e-09, 2.127889e-09, 1.651088e-09, 
    1.273828e-09, 1.013803e-09, 9.789574e-10, 9.994811e-10, 8.924366e-10,
  1.915507e-08, 1.700871e-08, 1.400385e-08, 1.109879e-08, 8.396739e-09, 
    6.016524e-09, 4.305484e-09, 3.160086e-09, 2.331639e-09, 1.810543e-09, 
    1.459833e-09, 1.195837e-09, 1.089143e-09, 1.018845e-09, 8.777442e-10,
  2.033956e-08, 1.833416e-08, 1.556598e-08, 1.251539e-08, 9.708469e-09, 
    7.263896e-09, 5.133695e-09, 3.674523e-09, 2.653464e-09, 2.013509e-09, 
    1.58968e-09, 1.320754e-09, 1.157972e-09, 1.032718e-09, 8.722218e-10,
  2.081418e-08, 1.932284e-08, 1.692599e-08, 1.420476e-08, 1.116305e-08, 
    8.356671e-09, 6.103206e-09, 4.537684e-09, 3.274437e-09, 2.338419e-09, 
    1.739702e-09, 1.415333e-09, 1.196437e-09, 1.051804e-09, 8.860803e-10,
  2.172525e-08, 2.028877e-08, 1.826499e-08, 1.563093e-08, 1.285651e-08, 
    9.856368e-09, 6.901871e-09, 4.866651e-09, 3.676202e-09, 2.677536e-09, 
    1.91988e-09, 1.515243e-09, 1.25427e-09, 1.07718e-09, 9.140533e-10,
  2.301355e-08, 2.142846e-08, 1.942798e-08, 1.671862e-08, 1.430119e-08, 
    1.160952e-08, 8.375072e-09, 5.573657e-09, 3.950453e-09, 3.000232e-09, 
    2.133922e-09, 1.609026e-09, 1.299228e-09, 1.098389e-09, 9.433894e-10,
  2.32723e-08, 2.229917e-08, 2.030767e-08, 1.767981e-08, 1.563256e-08, 
    1.317048e-08, 1.005779e-08, 6.832353e-09, 4.700111e-09, 3.444901e-09, 
    2.41762e-09, 1.745663e-09, 1.34122e-09, 1.114403e-09, 9.685619e-10,
  1.952623e-08, 1.717696e-08, 1.343928e-08, 8.640034e-09, 5.00873e-09, 
    3.230556e-09, 2.227217e-09, 1.488839e-09, 9.971565e-10, 7.463918e-10, 
    6.169689e-10, 5.736862e-10, 6.022688e-10, 5.734775e-10, 5.634497e-10,
  2.011312e-08, 1.822129e-08, 1.47293e-08, 1.008345e-08, 5.778163e-09, 
    3.519818e-09, 2.378986e-09, 1.567108e-09, 1.03602e-09, 7.513887e-10, 
    6.115214e-10, 5.510209e-10, 5.564318e-10, 5.002916e-10, 4.639751e-10,
  2.064326e-08, 1.892874e-08, 1.591361e-08, 1.159027e-08, 6.810505e-09, 
    3.944199e-09, 2.572836e-09, 1.684913e-09, 1.100757e-09, 7.685867e-10, 
    6.265305e-10, 5.54513e-10, 5.520248e-10, 4.957463e-10, 4.780401e-10,
  2.099874e-08, 1.928486e-08, 1.691532e-08, 1.306815e-08, 8.06972e-09, 
    4.536392e-09, 2.828722e-09, 1.829906e-09, 1.189933e-09, 8.066899e-10, 
    6.41671e-10, 5.606128e-10, 5.571552e-10, 5.084341e-10, 5.086355e-10,
  2.171827e-08, 1.987399e-08, 1.772962e-08, 1.439998e-08, 9.525702e-09, 
    5.290375e-09, 3.146726e-09, 1.997887e-09, 1.286636e-09, 8.520396e-10, 
    6.576837e-10, 5.696835e-10, 5.71196e-10, 5.163872e-10, 5.075845e-10,
  2.188749e-08, 2.01375e-08, 1.843469e-08, 1.564431e-08, 1.109716e-08, 
    6.382185e-09, 3.605302e-09, 2.253405e-09, 1.419847e-09, 9.087017e-10, 
    6.730624e-10, 5.785216e-10, 5.818179e-10, 5.112556e-10, 4.698598e-10,
  2.296122e-08, 2.090917e-08, 1.916345e-08, 1.677545e-08, 1.261997e-08, 
    7.753634e-09, 4.356939e-09, 2.6648e-09, 1.60869e-09, 9.928729e-10, 
    7.073641e-10, 5.875028e-10, 5.888598e-10, 5.015438e-10, 4.290894e-10,
  2.360838e-08, 2.140258e-08, 1.972533e-08, 1.776702e-08, 1.431662e-08, 
    9.302796e-09, 5.02024e-09, 2.778603e-09, 1.677642e-09, 1.055786e-09, 
    7.464977e-10, 6.01676e-10, 5.964899e-10, 4.938224e-10, 3.964809e-10,
  2.399771e-08, 2.209157e-08, 2.027983e-08, 1.864106e-08, 1.559694e-08, 
    1.033452e-08, 5.65749e-09, 2.955584e-09, 1.767518e-09, 1.122685e-09, 
    7.762083e-10, 6.151383e-10, 6.063596e-10, 4.878022e-10, 3.709578e-10,
  2.413346e-08, 2.281917e-08, 2.089265e-08, 1.919354e-08, 1.680015e-08, 
    1.172887e-08, 6.740855e-09, 3.506962e-09, 2.04209e-09, 1.234574e-09, 
    8.223576e-10, 6.380003e-10, 6.23836e-10, 4.886356e-10, 3.594807e-10,
  1.886021e-08, 1.711825e-08, 1.58206e-08, 1.422768e-08, 1.189428e-08, 
    9.091763e-09, 6.636881e-09, 4.65708e-09, 2.953968e-09, 1.648841e-09, 
    1.001005e-09, 8.273839e-10, 8.003956e-10, 5.115016e-10, -6.548859e-11,
  2.003324e-08, 1.80643e-08, 1.62848e-08, 1.490536e-08, 1.265901e-08, 
    9.809784e-09, 7.113396e-09, 4.963312e-09, 3.173794e-09, 1.772623e-09, 
    1.033531e-09, 8.126954e-10, 7.832472e-10, 4.813586e-10, -1.068507e-10,
  2.173291e-08, 1.935384e-08, 1.695243e-08, 1.535062e-08, 1.34575e-08, 
    1.065135e-08, 7.688021e-09, 5.364783e-09, 3.440576e-09, 1.923338e-09, 
    1.087204e-09, 8.189738e-10, 7.722384e-10, 4.926747e-10, -2.047336e-10,
  2.34533e-08, 2.033856e-08, 1.789078e-08, 1.582456e-08, 1.41668e-08, 
    1.152932e-08, 8.316643e-09, 5.729012e-09, 3.716097e-09, 2.099306e-09, 
    1.156732e-09, 8.363033e-10, 7.618625e-10, 4.700033e-10, -1.653497e-10,
  2.497505e-08, 2.218045e-08, 1.882995e-08, 1.658273e-08, 1.4775e-08, 
    1.237799e-08, 9.18371e-09, 6.260937e-09, 4.019412e-09, 2.297926e-09, 
    1.244064e-09, 8.593969e-10, 7.582701e-10, 4.413971e-10, -5.811773e-11,
  2.455773e-08, 2.286123e-08, 1.996582e-08, 1.742113e-08, 1.535662e-08, 
    1.326316e-08, 1.002766e-08, 6.815002e-09, 4.430175e-09, 2.53896e-09, 
    1.34732e-09, 8.90268e-10, 7.602243e-10, 4.152641e-10, -1.062441e-10,
  2.422908e-08, 2.351216e-08, 2.128381e-08, 1.830759e-08, 1.593659e-08, 
    1.394957e-08, 1.105502e-08, 7.644951e-09, 4.916719e-09, 2.797019e-09, 
    1.443693e-09, 9.159626e-10, 7.650197e-10, 3.941842e-10, -1.18805e-10,
  2.448079e-08, 2.401102e-08, 2.21531e-08, 1.927151e-08, 1.674876e-08, 
    1.456257e-08, 1.189132e-08, 8.396854e-09, 5.212124e-09, 3.020645e-09, 
    1.536805e-09, 9.309438e-10, 7.696982e-10, 3.683909e-10, -1.37304e-10,
  2.447668e-08, 2.436209e-08, 2.275701e-08, 2.02831e-08, 1.754585e-08, 
    1.511265e-08, 1.265866e-08, 9.345952e-09, 5.843904e-09, 3.39421e-09, 
    1.672558e-09, 9.53715e-10, 7.770974e-10, 3.518947e-10, -1.584065e-10,
  2.399466e-08, 2.435495e-08, 2.351836e-08, 2.114966e-08, 1.827555e-08, 
    1.582225e-08, 1.35102e-08, 1.018712e-08, 6.582138e-09, 3.80065e-09, 
    1.8379e-09, 9.855977e-10, 7.875071e-10, 3.795091e-10, -1.849618e-10,
  1.875223e-08, 1.706619e-08, 1.510545e-08, 1.281433e-08, 1.019156e-08, 
    7.48809e-09, 5.023337e-09, 3.122621e-09, 1.758604e-09, 1.013345e-09, 
    6.986048e-10, 6.750504e-10, 6.197273e-10, 6.906912e-10, 8.377694e-10,
  1.902582e-08, 1.809629e-08, 1.595506e-08, 1.376607e-08, 1.118837e-08, 
    8.421648e-09, 5.757013e-09, 3.588863e-09, 2.035333e-09, 1.120671e-09, 
    7.106615e-10, 6.224425e-10, 5.743396e-10, 6.34078e-10, 6.553876e-10,
  1.943523e-08, 1.874638e-08, 1.696327e-08, 1.467516e-08, 1.21912e-08, 
    9.399139e-09, 6.551651e-09, 4.168928e-09, 2.410116e-09, 1.26365e-09, 
    7.694057e-10, 6.262926e-10, 5.764839e-10, 6.302705e-10, 5.993593e-10,
  1.954956e-08, 1.906042e-08, 1.788247e-08, 1.565133e-08, 1.317503e-08, 
    1.045809e-08, 7.42443e-09, 4.785821e-09, 2.812104e-09, 1.455244e-09, 
    8.325797e-10, 6.223042e-10, 5.697579e-10, 6.379416e-10, 5.943496e-10,
  2.040986e-08, 1.962348e-08, 1.842244e-08, 1.663282e-08, 1.423095e-08, 
    1.146361e-08, 8.414588e-09, 5.560495e-09, 3.303323e-09, 1.701542e-09, 
    9.079832e-10, 6.492274e-10, 6.113137e-10, 6.671294e-10, 6.245693e-10,
  2.03851e-08, 1.974723e-08, 1.876006e-08, 1.73147e-08, 1.523856e-08, 
    1.257217e-08, 9.3958e-09, 6.311909e-09, 3.847194e-09, 2.001968e-09, 
    1.009389e-09, 6.782443e-10, 6.445148e-10, 6.907828e-10, 6.249721e-10,
  2.078835e-08, 2.005976e-08, 1.925899e-08, 1.792687e-08, 1.6093e-08, 
    1.362219e-08, 1.055714e-08, 7.292097e-09, 4.486241e-09, 2.33739e-09, 
    1.149317e-09, 7.042197e-10, 6.475619e-10, 6.933929e-10, 6.147231e-10,
  2.129201e-08, 2.043698e-08, 1.957933e-08, 1.846118e-08, 1.687036e-08, 
    1.46915e-08, 1.156282e-08, 8.206078e-09, 5.121381e-09, 2.705396e-09, 
    1.318171e-09, 7.373862e-10, 6.462501e-10, 6.954142e-10, 5.891314e-10,
  2.19782e-08, 2.090708e-08, 1.994308e-08, 1.884455e-08, 1.737952e-08, 
    1.542669e-08, 1.26918e-08, 9.334425e-09, 6.030814e-09, 3.203633e-09, 
    1.511411e-09, 7.788674e-10, 6.435829e-10, 6.980848e-10, 5.990924e-10,
  2.248804e-08, 2.139881e-08, 2.033946e-08, 1.925015e-08, 1.789523e-08, 
    1.62034e-08, 1.378628e-08, 1.030753e-08, 6.927013e-09, 3.754126e-09, 
    1.743832e-09, 8.396744e-10, 6.484526e-10, 7.023671e-10, 6.023468e-10,
  2.192286e-08, 2.021479e-08, 1.814607e-08, 1.576004e-08, 1.248942e-08, 
    9.039113e-09, 5.770802e-09, 3.270602e-09, 1.642262e-09, 5.744318e-10, 
    5.858424e-10, 5.482789e-10, 4.491446e-10, 6.20112e-10, 8.967529e-10,
  2.219089e-08, 2.103067e-08, 1.901654e-08, 1.669393e-08, 1.359751e-08, 
    1.001674e-08, 6.576634e-09, 3.680668e-09, 1.833153e-09, 6.380301e-10, 
    5.62093e-10, 5.54409e-10, 4.149295e-10, 4.849255e-10, 7.607326e-10,
  2.267654e-08, 2.16634e-08, 1.988123e-08, 1.760285e-08, 1.463756e-08, 
    1.101103e-08, 7.412163e-09, 4.212566e-09, 2.062228e-09, 7.406405e-10, 
    5.520776e-10, 6.449253e-10, 5.106088e-10, 4.406248e-10, 6.235849e-10,
  2.27008e-08, 2.233352e-08, 2.057781e-08, 1.850183e-08, 1.566066e-08, 
    1.208916e-08, 8.27033e-09, 4.816092e-09, 2.293118e-09, 8.410507e-10, 
    4.970001e-10, 6.810964e-10, 5.033514e-10, 4.018156e-10, 6.696128e-10,
  2.332338e-08, 2.306905e-08, 2.13252e-08, 1.926167e-08, 1.665944e-08, 
    1.312395e-08, 9.201523e-09, 5.50114e-09, 2.579705e-09, 9.601473e-10, 
    4.841754e-10, 6.493488e-10, 3.803088e-10, 3.727186e-10, 6.192613e-10,
  2.31351e-08, 2.316063e-08, 2.190868e-08, 1.981566e-08, 1.761143e-08, 
    1.422794e-08, 1.015364e-08, 6.222655e-09, 2.943254e-09, 1.10223e-09, 
    5.055568e-10, 6.515127e-10, 3.839e-10, 3.286053e-10, 5.484451e-10,
  2.246945e-08, 2.30079e-08, 2.22327e-08, 2.038659e-08, 1.832036e-08, 
    1.520613e-08, 1.130445e-08, 7.172801e-09, 3.434276e-09, 1.267804e-09, 
    5.393856e-10, 6.517781e-10, 5.020393e-10, 3.840316e-10, 4.955507e-10,
  2.212076e-08, 2.274825e-08, 2.254131e-08, 2.08707e-08, 1.899809e-08, 
    1.621245e-08, 1.230724e-08, 8.024472e-09, 3.897314e-09, 1.409511e-09, 
    5.585106e-10, 5.886606e-10, 5.778413e-10, 5.224792e-10, 4.508157e-10,
  2.200202e-08, 2.25083e-08, 2.261045e-08, 2.115846e-08, 1.945664e-08, 
    1.728692e-08, 1.349689e-08, 9.197405e-09, 4.697304e-09, 1.644449e-09, 
    5.92135e-10, 5.499213e-10, 6.515502e-10, 6.383933e-10, 3.910218e-10,
  2.177175e-08, 2.2166e-08, 2.258504e-08, 2.155371e-08, 2.002697e-08, 
    1.822461e-08, 1.456857e-08, 1.027097e-08, 5.490672e-09, 1.976805e-09, 
    6.445469e-10, 4.981742e-10, 6.867966e-10, 6.332488e-10, 3.430667e-10,
  2.441067e-08, 2.353662e-08, 2.097527e-08, 1.847961e-08, 1.527964e-08, 
    1.085609e-08, 6.29119e-09, 3.622852e-09, 2.760648e-09, 1.404323e-09, 
    6.107406e-10, 3.211781e-10, 3.306633e-10, 3.831603e-10, 2.022e-10,
  2.383047e-08, 2.415209e-08, 2.215518e-08, 1.959723e-08, 1.671667e-08, 
    1.277997e-08, 8.001576e-09, 4.410374e-09, 3.103687e-09, 1.851808e-09, 
    7.510095e-10, 3.522735e-10, 3.034751e-10, 2.842352e-10, 1.322982e-10,
  2.348829e-08, 2.432762e-08, 2.313877e-08, 2.059276e-08, 1.797447e-08, 
    1.441654e-08, 9.757106e-09, 5.491811e-09, 3.425645e-09, 2.349592e-09, 
    9.663812e-10, 3.972763e-10, 2.905101e-10, 2.332516e-10, 8.572933e-11,
  2.29989e-08, 2.439464e-08, 2.385316e-08, 2.161218e-08, 1.904471e-08, 
    1.586526e-08, 1.148154e-08, 6.789532e-09, 3.928838e-09, 2.772687e-09, 
    1.259886e-09, 4.660322e-10, 2.929049e-10, 1.752751e-10, 6.878127e-11,
  2.33554e-08, 2.431005e-08, 2.431675e-08, 2.248926e-08, 1.999854e-08, 
    1.703979e-08, 1.311498e-08, 8.319806e-09, 4.695068e-09, 3.215439e-09, 
    1.580579e-09, 5.679355e-10, 3.081266e-10, 1.503666e-10, 1.998008e-11,
  2.378878e-08, 2.414168e-08, 2.456184e-08, 2.309209e-08, 2.091279e-08, 
    1.819058e-08, 1.441185e-08, 9.683911e-09, 5.654912e-09, 3.622746e-09, 
    1.926568e-09, 7.109478e-10, 3.212984e-10, 1.312965e-10, 1.662194e-12,
  2.358573e-08, 2.372984e-08, 2.436449e-08, 2.357758e-08, 2.154684e-08, 
    1.908933e-08, 1.585108e-08, 1.122068e-08, 6.772342e-09, 4.153702e-09, 
    2.316709e-09, 8.956356e-10, 3.523082e-10, 1.264755e-10, -2.763822e-11,
  2.348498e-08, 2.345929e-08, 2.42855e-08, 2.379006e-08, 2.226878e-08, 
    1.994607e-08, 1.686027e-08, 1.247452e-08, 7.810067e-09, 4.776954e-09, 
    2.752991e-09, 1.134041e-09, 4.035517e-10, 1.451963e-10, -6.54903e-11,
  2.361328e-08, 2.34571e-08, 2.39627e-08, 2.370508e-08, 2.245834e-08, 
    2.071766e-08, 1.779784e-08, 1.38294e-08, 9.133927e-09, 5.52093e-09, 
    3.231138e-09, 1.397301e-09, 4.739346e-10, 1.632721e-10, -5.635493e-11,
  2.350607e-08, 2.33907e-08, 2.377305e-08, 2.374134e-08, 2.292098e-08, 
    2.136729e-08, 1.851736e-08, 1.467563e-08, 1.021346e-08, 6.361739e-09, 
    3.775436e-09, 1.682524e-09, 5.728895e-10, 1.893092e-10, -6.189355e-11,
  2.282597e-08, 2.209315e-08, 2.070486e-08, 1.810356e-08, 1.423657e-08, 
    1.011394e-08, 6.094997e-09, 4.070731e-09, 2.819006e-09, 1.938675e-09, 
    1.536698e-09, 1.207484e-09, 1.056178e-09, 8.873966e-10, 6.886649e-10,
  2.26865e-08, 2.286412e-08, 2.192493e-08, 1.987082e-08, 1.666184e-08, 
    1.247661e-08, 8.074582e-09, 4.903096e-09, 3.376642e-09, 2.270291e-09, 
    1.725045e-09, 1.361368e-09, 1.111465e-09, 9.002022e-10, 6.507632e-10,
  2.316362e-08, 2.297789e-08, 2.265744e-08, 2.126962e-08, 1.857578e-08, 
    1.495356e-08, 1.021009e-08, 6.160703e-09, 3.96385e-09, 2.708494e-09, 
    1.962617e-09, 1.520308e-09, 1.207146e-09, 9.419148e-10, 6.673514e-10,
  2.363921e-08, 2.325748e-08, 2.307214e-08, 2.225229e-08, 2.015767e-08, 
    1.710326e-08, 1.258163e-08, 7.942882e-09, 4.714448e-09, 3.127868e-09, 
    2.239242e-09, 1.700359e-09, 1.309633e-09, 9.986287e-10, 7.085675e-10,
  2.324135e-08, 2.319698e-08, 2.344293e-08, 2.296858e-08, 2.144438e-08, 
    1.880001e-08, 1.481102e-08, 1.002303e-08, 5.987728e-09, 3.614849e-09, 
    2.481741e-09, 1.871528e-09, 1.412062e-09, 1.06114e-09, 7.730321e-10,
  2.300342e-08, 2.332329e-08, 2.345198e-08, 2.341789e-08, 2.242296e-08, 
    2.023619e-08, 1.688085e-08, 1.201678e-08, 7.395811e-09, 4.36244e-09, 
    2.736652e-09, 1.995676e-09, 1.491961e-09, 1.131283e-09, 8.268791e-10,
  2.269788e-08, 2.321656e-08, 2.34957e-08, 2.372489e-08, 2.312763e-08, 
    2.136071e-08, 1.875739e-08, 1.419915e-08, 9.349845e-09, 5.373204e-09, 
    3.094302e-09, 2.109262e-09, 1.571472e-09, 1.186176e-09, 8.730605e-10,
  2.287371e-08, 2.304602e-08, 2.33867e-08, 2.367502e-08, 2.380989e-08, 
    2.210139e-08, 1.975766e-08, 1.585655e-08, 1.098439e-08, 6.544828e-09, 
    3.67367e-09, 2.238091e-09, 1.64935e-09, 1.238855e-09, 9.073176e-10,
  2.288546e-08, 2.286732e-08, 2.322226e-08, 2.3697e-08, 2.427812e-08, 
    2.304388e-08, 2.074801e-08, 1.736302e-08, 1.257485e-08, 7.718207e-09, 
    4.414704e-09, 2.548459e-09, 1.759489e-09, 1.304611e-09, 9.493062e-10,
  2.303239e-08, 2.277642e-08, 2.308046e-08, 2.359027e-08, 2.419151e-08, 
    2.347105e-08, 2.152356e-08, 1.861805e-08, 1.404307e-08, 9.040249e-09, 
    5.188809e-09, 2.951303e-09, 1.893594e-09, 1.388742e-09, 9.977033e-10,
  1.902738e-08, 1.617413e-08, 1.290705e-08, 9.195071e-09, 6.303416e-09, 
    4.546806e-09, 3.116954e-09, 2.094419e-09, 1.292894e-09, 1.112608e-09, 
    9.958429e-10, 7.040694e-10, 5.038654e-10, 4.746348e-10, 4.96985e-10,
  2.011233e-08, 1.806728e-08, 1.520102e-08, 1.156716e-08, 8.043545e-09, 
    5.640322e-09, 3.90204e-09, 2.692228e-09, 1.674464e-09, 1.177357e-09, 
    1.092978e-09, 8.687532e-10, 5.635318e-10, 4.869802e-10, 4.985292e-10,
  2.100893e-08, 1.942892e-08, 1.710528e-08, 1.399139e-08, 1.020615e-08, 
    7.076908e-09, 4.954685e-09, 3.309996e-09, 2.276839e-09, 1.405985e-09, 
    1.200075e-09, 1.00183e-09, 6.631727e-10, 5.061159e-10, 4.910493e-10,
  2.152134e-08, 2.0706e-08, 1.876237e-08, 1.604655e-08, 1.254427e-08, 
    8.989192e-09, 6.163984e-09, 4.211473e-09, 2.846063e-09, 1.859192e-09, 
    1.387487e-09, 1.155218e-09, 7.892386e-10, 5.479486e-10, 4.89652e-10,
  2.19441e-08, 2.136727e-08, 2.027316e-08, 1.802289e-08, 1.495482e-08, 
    1.116389e-08, 7.756403e-09, 5.32204e-09, 3.530548e-09, 2.432384e-09, 
    1.677315e-09, 1.335528e-09, 9.259813e-10, 6.134563e-10, 5.02567e-10,
  2.270302e-08, 2.181303e-08, 2.110921e-08, 1.938155e-08, 1.706979e-08, 
    1.368661e-08, 9.81432e-09, 6.625265e-09, 4.470167e-09, 2.970372e-09, 
    2.058863e-09, 1.56642e-09, 1.052775e-09, 7.06153e-10, 5.320323e-10,
  2.284819e-08, 2.245458e-08, 2.176119e-08, 2.067137e-08, 1.864425e-08, 
    1.588197e-08, 1.229652e-08, 8.529448e-09, 5.722372e-09, 3.813299e-09, 
    2.572364e-09, 1.88549e-09, 1.226575e-09, 8.104634e-10, 5.76013e-10,
  2.268405e-08, 2.291308e-08, 2.241347e-08, 2.151716e-08, 2.004266e-08, 
    1.776746e-08, 1.453021e-08, 1.039148e-08, 7.132185e-09, 4.63396e-09, 
    3.182588e-09, 2.228579e-09, 1.50412e-09, 9.03307e-10, 6.373169e-10,
  2.286808e-08, 2.319528e-08, 2.296735e-08, 2.217826e-08, 2.123459e-08, 
    1.9372e-08, 1.679632e-08, 1.284972e-08, 8.713849e-09, 5.602469e-09, 
    3.758764e-09, 2.588889e-09, 1.841238e-09, 1.00097e-09, 7.085524e-10,
  2.283326e-08, 2.303968e-08, 2.332838e-08, 2.296403e-08, 2.189624e-08, 
    2.060915e-08, 1.861025e-08, 1.512232e-08, 1.077331e-08, 7.001059e-09, 
    4.387627e-09, 3.060583e-09, 2.104527e-09, 1.135651e-09, 7.858967e-10,
  6.144459e-09, 3.696313e-09, 2.098414e-09, 1.243342e-09, 9.00447e-10, 
    7.020686e-10, 5.309411e-10, 5.224238e-10, 5.622992e-10, 7.28616e-10, 
    8.2793e-10, 9.470084e-10, 1.012585e-09, 8.160244e-10, 4.892945e-10,
  7.898856e-09, 4.952907e-09, 2.863141e-09, 1.571628e-09, 1.027833e-09, 
    8.001544e-10, 5.927931e-10, 5.329683e-10, 5.691747e-10, 6.593523e-10, 
    7.919276e-10, 8.939079e-10, 1.00933e-09, 8.796061e-10, 5.705479e-10,
  9.710774e-09, 6.489967e-09, 3.960496e-09, 2.093187e-09, 1.242654e-09, 
    9.163781e-10, 6.818197e-10, 5.499471e-10, 5.49896e-10, 5.939162e-10, 
    7.280301e-10, 8.381736e-10, 9.777722e-10, 9.214883e-10, 6.561948e-10,
  1.183864e-08, 8.390777e-09, 5.364603e-09, 2.961139e-09, 1.603381e-09, 
    1.077667e-09, 8.088838e-10, 6.189589e-10, 5.303524e-10, 5.485538e-10, 
    6.755326e-10, 7.859771e-10, 9.119163e-10, 9.245273e-10, 7.636958e-10,
  1.34584e-08, 1.031439e-08, 7.05156e-09, 4.209217e-09, 2.202277e-09, 
    1.289134e-09, 9.436684e-10, 7.381008e-10, 5.573049e-10, 5.04785e-10, 
    6.298717e-10, 7.428776e-10, 8.397241e-10, 9.179147e-10, 8.553745e-10,
  1.536303e-08, 1.233759e-08, 8.981366e-09, 5.746389e-09, 3.203937e-09, 
    1.699621e-09, 1.155598e-09, 9.157536e-10, 7.073933e-10, 5.550819e-10, 
    5.848515e-10, 7.159906e-10, 7.584605e-10, 8.720339e-10, 9.033859e-10,
  1.650653e-08, 1.3908e-08, 1.080204e-08, 7.553202e-09, 4.51352e-09, 
    2.380172e-09, 1.427275e-09, 1.147192e-09, 9.100908e-10, 6.734155e-10, 
    5.913745e-10, 6.838282e-10, 7.071684e-10, 8.247695e-10, 9.19071e-10,
  1.783794e-08, 1.561927e-08, 1.267318e-08, 9.41101e-09, 6.168245e-09, 
    3.494209e-09, 1.822235e-09, 1.224648e-09, 9.907618e-10, 7.779925e-10, 
    6.35881e-10, 6.357737e-10, 6.678653e-10, 7.864193e-10, 9.13677e-10,
  1.905271e-08, 1.710431e-08, 1.446373e-08, 1.113971e-08, 8.018666e-09, 
    5.121065e-09, 2.779546e-09, 1.513606e-09, 1.037656e-09, 8.604226e-10, 
    6.968793e-10, 5.818678e-10, 6.24063e-10, 7.478567e-10, 8.961126e-10,
  2.024663e-08, 1.844444e-08, 1.620082e-08, 1.30086e-08, 1.007972e-08, 
    6.961636e-09, 4.113117e-09, 2.256299e-09, 1.329393e-09, 9.985806e-10, 
    7.986949e-10, 6.020688e-10, 5.771565e-10, 6.967159e-10, 8.603164e-10,
  6.207944e-09, 3.623537e-09, 1.783918e-09, 1.073703e-09, 1.001419e-09, 
    9.269942e-10, 7.853436e-10, 5.960306e-10, 4.864202e-10, 3.826404e-10, 
    3.023161e-10, 3.969708e-10, 4.871974e-10, 4.952404e-10, 5.007025e-10,
  7.078302e-09, 4.45303e-09, 2.368525e-09, 1.22834e-09, 1.016783e-09, 
    9.575648e-10, 8.15388e-10, 6.454831e-10, 5.067346e-10, 3.758218e-10, 
    2.724015e-10, 3.619518e-10, 4.631162e-10, 4.700327e-10, 4.663217e-10,
  8.43175e-09, 5.581878e-09, 3.1329e-09, 1.461233e-09, 1.087001e-09, 
    9.868641e-10, 8.461872e-10, 6.849039e-10, 5.296678e-10, 3.820532e-10, 
    2.668271e-10, 3.532374e-10, 4.618286e-10, 4.483531e-10, 4.565216e-10,
  1.005272e-08, 6.825837e-09, 4.044213e-09, 1.863554e-09, 1.220688e-09, 
    1.035096e-09, 9.046949e-10, 7.309395e-10, 5.577274e-10, 3.984525e-10, 
    2.689835e-10, 3.480381e-10, 4.571036e-10, 4.627979e-10, 4.661376e-10,
  1.149603e-08, 8.121091e-09, 5.047181e-09, 2.497419e-09, 1.417431e-09, 
    1.113074e-09, 9.452394e-10, 7.965332e-10, 6.10218e-10, 4.331987e-10, 
    2.784728e-10, 3.31544e-10, 4.454876e-10, 4.755484e-10, 4.536871e-10,
  1.270824e-08, 9.467562e-09, 6.200224e-09, 3.263391e-09, 1.696333e-09, 
    1.265997e-09, 1.017022e-09, 8.411464e-10, 6.162437e-10, 4.508742e-10, 
    2.953317e-10, 3.245813e-10, 4.260703e-10, 4.744465e-10, 4.369071e-10,
  1.375979e-08, 1.043844e-08, 7.238008e-09, 4.242291e-09, 2.089869e-09, 
    1.386817e-09, 1.106457e-09, 9.362224e-10, 6.857765e-10, 4.857152e-10, 
    3.154202e-10, 3.282597e-10, 4.030356e-10, 4.558757e-10, 4.12741e-10,
  1.470334e-08, 1.180353e-08, 8.445933e-09, 5.278309e-09, 2.724651e-09, 
    1.592016e-09, 1.170689e-09, 9.878882e-10, 8.170338e-10, 5.882165e-10, 
    3.515616e-10, 3.597653e-10, 4.003211e-10, 4.222999e-10, 3.953128e-10,
  1.558037e-08, 1.299237e-08, 9.626419e-09, 6.283852e-09, 3.501309e-09, 
    2.126844e-09, 1.439239e-09, 1.019674e-09, 8.404787e-10, 6.20926e-10, 
    3.962902e-10, 3.928216e-10, 4.280022e-10, 4.022388e-10, 3.924015e-10,
  1.643145e-08, 1.403471e-08, 1.081096e-08, 7.516726e-09, 4.439196e-09, 
    2.623161e-09, 1.778696e-09, 1.188175e-09, 8.818831e-10, 6.414099e-10, 
    4.229281e-10, 3.832047e-10, 4.47195e-10, 4.174048e-10, 4.195044e-10,
  1.156567e-08, 6.853178e-09, 3.402703e-09, 1.890669e-09, 1.62724e-09, 
    1.440626e-09, 1.225881e-09, 1.061165e-09, 9.299882e-10, 9.22696e-10, 
    9.719957e-10, 8.341138e-10, 5.6609e-10, 4.587176e-10, 4.242821e-10,
  1.304773e-08, 8.500566e-09, 4.445907e-09, 2.166024e-09, 1.672993e-09, 
    1.487328e-09, 1.288968e-09, 1.126989e-09, 9.683586e-10, 9.124935e-10, 
    9.305298e-10, 8.1377e-10, 5.089797e-10, 4.131024e-10, 3.588514e-10,
  1.463135e-08, 1.021317e-08, 5.775318e-09, 2.665947e-09, 1.756019e-09, 
    1.555953e-09, 1.364283e-09, 1.168887e-09, 9.979989e-10, 8.916572e-10, 
    9.036408e-10, 8.281493e-10, 4.938854e-10, 5.215597e-10, 5.240643e-10,
  1.629831e-08, 1.181089e-08, 7.238108e-09, 3.465036e-09, 1.932986e-09, 
    1.645184e-09, 1.45179e-09, 1.201725e-09, 1.028343e-09, 8.826358e-10, 
    8.791242e-10, 8.372927e-10, 4.868166e-10, 4.821362e-10, 7.050898e-10,
  1.753907e-08, 1.327209e-08, 8.785197e-09, 4.501301e-09, 2.223289e-09, 
    1.764444e-09, 1.527696e-09, 1.263413e-09, 1.103759e-09, 9.129256e-10, 
    8.668201e-10, 8.544166e-10, 4.983723e-10, 3.625813e-10, 8.337939e-10,
  1.875287e-08, 1.480278e-08, 1.037953e-08, 5.665508e-09, 2.693802e-09, 
    1.93079e-09, 1.663653e-09, 1.318781e-09, 1.145961e-09, 9.610976e-10, 
    8.780004e-10, 8.745595e-10, 5.137585e-10, 2.925178e-10, 7.822885e-10,
  1.973309e-08, 1.60295e-08, 1.179144e-08, 7.033786e-09, 3.281196e-09, 
    2.020335e-09, 1.823633e-09, 1.465025e-09, 1.240229e-09, 1.06304e-09, 
    9.054415e-10, 9.098191e-10, 5.422398e-10, 2.513424e-10, 6.651208e-10,
  2.055514e-08, 1.731086e-08, 1.329741e-08, 8.463479e-09, 4.161258e-09, 
    2.14403e-09, 1.757936e-09, 1.51374e-09, 1.333099e-09, 1.18174e-09, 
    9.306168e-10, 9.615587e-10, 5.968652e-10, 2.529073e-10, 5.556213e-10,
  2.096628e-08, 1.813894e-08, 1.460092e-08, 9.804466e-09, 5.169489e-09, 
    2.599771e-09, 1.922451e-09, 1.557192e-09, 1.320138e-09, 1.178301e-09, 
    9.446863e-10, 1.022223e-09, 6.823169e-10, 2.786797e-10, 4.846253e-10,
  2.127204e-08, 1.904296e-08, 1.574282e-08, 1.12758e-08, 6.286784e-09, 
    3.003249e-09, 2.077322e-09, 1.738537e-09, 1.328582e-09, 1.20097e-09, 
    9.829005e-10, 1.047013e-09, 7.816918e-10, 3.288473e-10, 4.539291e-10,
  7.290604e-09, 3.788042e-09, 1.988455e-09, 1.689936e-09, 1.386621e-09, 
    9.888964e-10, 8.110285e-10, 8.795582e-10, 1.010284e-09, 7.585683e-10, 
    5.999042e-10, 9.461313e-10, 1.20864e-09, 1.230983e-09, 1.041372e-09,
  9.163019e-09, 4.775302e-09, 2.258242e-09, 1.711672e-09, 1.463193e-09, 
    1.072987e-09, 8.442593e-10, 8.722779e-10, 9.50181e-10, 7.764626e-10, 
    6.107497e-10, 9.051039e-10, 1.120111e-09, 1.11562e-09, 9.906873e-10,
  1.113296e-08, 5.97504e-09, 2.721782e-09, 1.770178e-09, 1.527192e-09, 
    1.158551e-09, 8.701959e-10, 8.776667e-10, 9.421317e-10, 8.258162e-10, 
    6.614143e-10, 8.724561e-10, 1.065803e-09, 1.081302e-09, 9.984741e-10,
  1.349554e-08, 7.279324e-09, 3.374374e-09, 1.857018e-09, 1.583072e-09, 
    1.25693e-09, 9.067507e-10, 8.896882e-10, 9.595574e-10, 8.210607e-10, 
    7.169862e-10, 8.075091e-10, 1.056119e-09, 1.058029e-09, 9.521262e-10,
  1.585769e-08, 8.639035e-09, 4.252131e-09, 2.041721e-09, 1.635176e-09, 
    1.35195e-09, 9.627455e-10, 9.199397e-10, 9.650534e-10, 7.838458e-10, 
    7.710245e-10, 7.315782e-10, 9.6617e-10, 1.086999e-09, 8.477246e-10,
  1.795539e-08, 1.060765e-08, 5.388078e-09, 2.387221e-09, 1.683185e-09, 
    1.490038e-09, 1.052143e-09, 9.411122e-10, 9.575766e-10, 7.514005e-10, 
    7.940023e-10, 6.368787e-10, 8.768518e-10, 1.055626e-09, 6.692888e-10,
  2.047608e-08, 1.287051e-08, 6.923116e-09, 3.037565e-09, 1.779665e-09, 
    1.577777e-09, 1.191715e-09, 1.022226e-09, 9.91726e-10, 7.592725e-10, 
    8.115237e-10, 5.451652e-10, 7.806737e-10, 9.531196e-10, 5.203772e-10,
  2.218471e-08, 1.528278e-08, 8.575205e-09, 3.881759e-09, 2.063256e-09, 
    1.677863e-09, 1.204303e-09, 9.8177e-10, 9.599438e-10, 7.950985e-10, 
    7.890777e-10, 4.552457e-10, 6.796997e-10, 8.085027e-10, 4.171628e-10,
  2.304559e-08, 1.764389e-08, 1.046821e-08, 4.911077e-09, 2.316803e-09, 
    1.83438e-09, 1.312094e-09, 9.336416e-10, 9.253145e-10, 8.703677e-10, 
    7.668433e-10, 4.085585e-10, 5.820007e-10, 7.185792e-10, 3.183162e-10,
  2.362646e-08, 1.954323e-08, 1.25292e-08, 6.168306e-09, 2.587253e-09, 
    1.921263e-09, 1.511587e-09, 1.071524e-09, 9.739586e-10, 9.036901e-10, 
    8.255596e-10, 3.798016e-10, 5.038439e-10, 6.685153e-10, 2.393399e-10,
  1.607583e-08, 1.248059e-08, 8.365871e-09, 4.177164e-09, 1.857687e-09, 
    1.130764e-09, 8.066348e-10, 6.239885e-10, 5.507523e-10, 6.185421e-10, 
    8.345428e-10, 8.244332e-10, 9.865307e-10, 1.167844e-09, 8.502122e-10,
  1.828858e-08, 1.409475e-08, 9.783741e-09, 5.365115e-09, 2.319263e-09, 
    1.278673e-09, 8.904857e-10, 6.469761e-10, 5.927037e-10, 6.161806e-10, 
    7.907449e-10, 8.865477e-10, 1.040859e-09, 1.19088e-09, 8.034869e-10,
  1.991979e-08, 1.552435e-08, 1.124722e-08, 6.847203e-09, 3.050795e-09, 
    1.47842e-09, 9.812262e-10, 7.177025e-10, 6.26277e-10, 6.427932e-10, 
    7.431942e-10, 9.293278e-10, 1.024022e-09, 1.145894e-09, 8.000205e-10,
  2.127714e-08, 1.684969e-08, 1.280191e-08, 8.49501e-09, 4.059085e-09, 
    1.785813e-09, 1.067295e-09, 7.622115e-10, 6.006254e-10, 6.378652e-10, 
    6.581144e-10, 8.960959e-10, 9.846057e-10, 1.107066e-09, 7.621028e-10,
  2.236994e-08, 1.846056e-08, 1.449008e-08, 1.011686e-08, 5.356923e-09, 
    2.274865e-09, 1.181e-09, 8.440615e-10, 6.326039e-10, 6.520118e-10, 
    6.270213e-10, 8.137813e-10, 9.858834e-10, 1.078071e-09, 7.38402e-10,
  2.308139e-08, 2.000209e-08, 1.626945e-08, 1.195128e-08, 6.885144e-09, 
    3.02241e-09, 1.401561e-09, 9.152206e-10, 6.625862e-10, 6.431154e-10, 
    6.283346e-10, 7.34957e-10, 1.046791e-09, 9.904889e-10, 7.012171e-10,
  2.479485e-08, 2.160019e-08, 1.781165e-08, 1.361597e-08, 8.479742e-09, 
    3.9596e-09, 1.771137e-09, 1.013681e-09, 7.439849e-10, 6.460458e-10, 
    6.665016e-10, 7.37269e-10, 1.116692e-09, 9.511151e-10, 6.505064e-10,
  2.513403e-08, 2.274657e-08, 1.911053e-08, 1.499005e-08, 1.011047e-08, 
    4.970209e-09, 2.120603e-09, 1.15475e-09, 8.215099e-10, 6.865806e-10, 
    6.757357e-10, 7.253116e-10, 1.158271e-09, 9.823116e-10, 5.918575e-10,
  2.504427e-08, 2.375013e-08, 2.044933e-08, 1.663551e-08, 1.171341e-08, 
    6.021208e-09, 2.552786e-09, 1.308264e-09, 8.602007e-10, 6.41162e-10, 
    6.292941e-10, 6.361052e-10, 1.122311e-09, 1.040939e-09, 5.509758e-10,
  2.461401e-08, 2.438326e-08, 2.170916e-08, 1.801225e-08, 1.289422e-08, 
    7.253446e-09, 3.146254e-09, 1.539829e-09, 8.95482e-10, 6.426412e-10, 
    6.280327e-10, 6.072122e-10, 1.073427e-09, 1.093965e-09, 5.429315e-10,
  1.407916e-08, 1.043465e-08, 7.148159e-09, 4.019677e-09, 2.274669e-09, 
    1.413407e-09, 1.086832e-09, 1.132038e-09, 1.199803e-09, 1.097421e-09, 
    1.058632e-09, 1.110487e-09, 1.053025e-09, 4.338238e-10, 1.769542e-10,
  1.585623e-08, 1.254316e-08, 9.106673e-09, 5.51293e-09, 3.006163e-09, 
    1.742675e-09, 1.194601e-09, 1.135789e-09, 1.266958e-09, 1.2473e-09, 
    1.175817e-09, 1.180132e-09, 1.067098e-09, 3.139103e-10, -4.159711e-11,
  1.759374e-08, 1.459631e-08, 1.129524e-08, 7.344944e-09, 4.068884e-09, 
    2.226773e-09, 1.373709e-09, 1.159416e-09, 1.292591e-09, 1.352888e-09, 
    1.2685e-09, 1.20665e-09, 9.475928e-10, 7.318724e-11, -2.066471e-10,
  1.914165e-08, 1.657568e-08, 1.331903e-08, 9.520064e-09, 5.595469e-09, 
    2.960806e-09, 1.657547e-09, 1.208964e-09, 1.272167e-09, 1.397163e-09, 
    1.339309e-09, 1.168887e-09, 7.788992e-10, -3.36663e-11, -1.736086e-10,
  2.061401e-08, 1.840089e-08, 1.528501e-08, 1.179693e-08, 7.613209e-09, 
    4.099198e-09, 2.108668e-09, 1.352844e-09, 1.248172e-09, 1.400337e-09, 
    1.370906e-09, 1.15405e-09, 7.164587e-10, 1.349048e-11, -8.194755e-11,
  2.219304e-08, 1.981417e-08, 1.708671e-08, 1.38587e-08, 9.920138e-09, 
    5.782892e-09, 2.938963e-09, 1.641661e-09, 1.288472e-09, 1.404762e-09, 
    1.383171e-09, 1.162552e-09, 7.413229e-10, 1.585611e-10, -4.610068e-11,
  2.306885e-08, 2.134647e-08, 1.879342e-08, 1.580618e-08, 1.216755e-08, 
    7.706482e-09, 4.116552e-09, 2.185415e-09, 1.517704e-09, 1.468881e-09, 
    1.441892e-09, 1.236423e-09, 8.424381e-10, 2.777845e-10, -6.886626e-11,
  2.39647e-08, 2.273467e-08, 2.053089e-08, 1.754546e-08, 1.424492e-08, 
    1.008416e-08, 5.570883e-09, 2.818649e-09, 1.721323e-09, 1.497819e-09, 
    1.477238e-09, 1.315582e-09, 9.524878e-10, 4.0805e-10, -4.184447e-11,
  2.430068e-08, 2.390115e-08, 2.204472e-08, 1.91896e-08, 1.613613e-08, 
    1.244925e-08, 7.752633e-09, 3.903802e-09, 2.036493e-09, 1.513626e-09, 
    1.456585e-09, 1.37125e-09, 1.058287e-09, 5.334038e-10, 1.73166e-11,
  2.451805e-08, 2.454327e-08, 2.350902e-08, 2.090137e-08, 1.798282e-08, 
    1.456133e-08, 1.019211e-08, 5.451538e-09, 2.671171e-09, 1.726621e-09, 
    1.496145e-09, 1.413503e-09, 1.156881e-09, 6.618493e-10, 1.179095e-10,
  9.845542e-09, 7.636107e-09, 5.775201e-09, 4.009605e-09, 2.860054e-09, 
    2.198926e-09, 1.828751e-09, 1.686078e-09, 1.704218e-09, 1.883629e-09, 
    1.958511e-09, 1.839916e-09, 1.628155e-09, 1.371412e-09, 9.963554e-10,
  1.100161e-08, 8.681764e-09, 6.673302e-09, 4.710043e-09, 3.303811e-09, 
    2.444616e-09, 1.965789e-09, 1.729427e-09, 1.642708e-09, 1.800443e-09, 
    1.978584e-09, 1.942231e-09, 1.726976e-09, 1.412637e-09, 1.000734e-09,
  1.268565e-08, 1.018522e-08, 7.719031e-09, 5.407873e-09, 3.845438e-09, 
    2.812001e-09, 2.182398e-09, 1.851742e-09, 1.704019e-09, 1.749492e-09, 
    1.969896e-09, 2.03479e-09, 1.812162e-09, 1.464903e-09, 1.047362e-09,
  1.423443e-08, 1.185564e-08, 8.881205e-09, 6.13617e-09, 4.389924e-09, 
    3.212521e-09, 2.441154e-09, 2.006707e-09, 1.804611e-09, 1.760574e-09, 
    1.923179e-09, 2.06772e-09, 1.903943e-09, 1.571437e-09, 1.165423e-09,
  1.563759e-08, 1.340964e-08, 1.020254e-08, 7.237464e-09, 5.00013e-09, 
    3.559141e-09, 2.589724e-09, 2.05664e-09, 1.811427e-09, 1.74659e-09, 
    1.828427e-09, 2.03354e-09, 1.956455e-09, 1.685692e-09, 1.299749e-09,
  1.728422e-08, 1.464735e-08, 1.174156e-08, 8.590851e-09, 5.905813e-09, 
    4.178941e-09, 2.964867e-09, 2.232445e-09, 1.836907e-09, 1.710926e-09, 
    1.716085e-09, 1.931138e-09, 1.96735e-09, 1.778713e-09, 1.425903e-09,
  1.81324e-08, 1.587131e-08, 1.307365e-08, 1.027312e-08, 7.175937e-09, 
    4.823479e-09, 3.444436e-09, 2.653981e-09, 2.142372e-09, 1.815013e-09, 
    1.690615e-09, 1.813782e-09, 1.977911e-09, 1.841603e-09, 1.534031e-09,
  1.928288e-08, 1.739582e-08, 1.468243e-08, 1.173842e-08, 8.775215e-09, 
    5.934648e-09, 3.825795e-09, 2.573285e-09, 2.137451e-09, 1.909843e-09, 
    1.741002e-09, 1.747341e-09, 1.957414e-09, 1.888528e-09, 1.637568e-09,
  2.02869e-08, 1.868577e-08, 1.613117e-08, 1.289845e-08, 1.023467e-08, 
    7.522326e-09, 4.832565e-09, 2.863202e-09, 2.082669e-09, 1.955131e-09, 
    1.759617e-09, 1.708517e-09, 1.918945e-09, 1.926374e-09, 1.718445e-09,
  2.148264e-08, 1.981251e-08, 1.745516e-08, 1.426765e-08, 1.169545e-08, 
    9.080972e-09, 6.179628e-09, 3.812313e-09, 2.601243e-09, 2.141801e-09, 
    1.793159e-09, 1.655595e-09, 1.838727e-09, 1.945676e-09, 1.801683e-09,
  1.62142e-08, 1.42299e-08, 1.206952e-08, 1.00544e-08, 8.038018e-09, 
    6.199772e-09, 4.327268e-09, 3.036711e-09, 2.355462e-09, 1.829075e-09, 
    1.355982e-09, 1.010312e-09, 8.753831e-10, 9.000037e-10, 7.541042e-10,
  1.713334e-08, 1.53955e-08, 1.312356e-08, 1.099126e-08, 8.906531e-09, 
    7.012209e-09, 5.070227e-09, 3.469635e-09, 2.534191e-09, 1.978146e-09, 
    1.50434e-09, 1.115941e-09, 9.019901e-10, 9.140552e-10, 7.895007e-10,
  1.790396e-08, 1.628141e-08, 1.422192e-08, 1.193775e-08, 9.775036e-09, 
    7.782985e-09, 5.828868e-09, 4.01708e-09, 2.824108e-09, 2.140565e-09, 
    1.655195e-09, 1.236247e-09, 9.556118e-10, 9.419796e-10, 8.508814e-10,
  1.899254e-08, 1.714995e-08, 1.517341e-08, 1.287295e-08, 1.067255e-08, 
    8.624856e-09, 6.603302e-09, 4.661961e-09, 3.168626e-09, 2.302446e-09, 
    1.789377e-09, 1.354212e-09, 1.028663e-09, 9.729364e-10, 9.131141e-10,
  1.953914e-08, 1.771556e-08, 1.617221e-08, 1.385473e-08, 1.15686e-08, 
    9.421533e-09, 7.342712e-09, 5.427002e-09, 3.714959e-09, 2.542988e-09, 
    1.905845e-09, 1.441656e-09, 1.095098e-09, 9.948622e-10, 9.67424e-10,
  2.053298e-08, 1.85568e-08, 1.692403e-08, 1.478786e-08, 1.250277e-08, 
    1.034103e-08, 8.157873e-09, 6.049611e-09, 4.21154e-09, 2.833259e-09, 
    2.030791e-09, 1.505589e-09, 1.136695e-09, 1.003619e-09, 1.009185e-09,
  2.147103e-08, 1.964279e-08, 1.772988e-08, 1.56807e-08, 1.333875e-08, 
    1.110287e-08, 9.003857e-09, 6.93222e-09, 4.9788e-09, 3.303077e-09, 
    2.23604e-09, 1.600553e-09, 1.183954e-09, 1.003123e-09, 1.03206e-09,
  2.221914e-08, 2.035451e-08, 1.840302e-08, 1.651496e-08, 1.43477e-08, 
    1.187093e-08, 9.621033e-09, 7.569465e-09, 5.665371e-09, 3.894484e-09, 
    2.578636e-09, 1.805901e-09, 1.283151e-09, 1.022338e-09, 1.037295e-09,
  2.248948e-08, 2.09716e-08, 1.924601e-08, 1.714029e-08, 1.52536e-08, 
    1.29526e-08, 1.051869e-08, 8.184877e-09, 5.970867e-09, 4.284717e-09, 
    2.927952e-09, 2.04566e-09, 1.425429e-09, 1.058739e-09, 1.027594e-09,
  2.29653e-08, 2.148514e-08, 2.00248e-08, 1.803897e-08, 1.572065e-08, 
    1.360261e-08, 1.133801e-08, 8.924308e-09, 6.594692e-09, 4.726725e-09, 
    3.259968e-09, 2.260048e-09, 1.577515e-09, 1.101606e-09, 1.006161e-09,
  1.791726e-08, 1.68252e-08, 1.530534e-08, 1.292532e-08, 1.031307e-08, 
    7.687182e-09, 5.252822e-09, 3.516721e-09, 2.617499e-09, 2.078363e-09, 
    1.463589e-09, 9.824815e-10, 7.682134e-10, 6.907399e-10, 7.519099e-10,
  1.81558e-08, 1.754925e-08, 1.631969e-08, 1.428275e-08, 1.17395e-08, 
    9.118407e-09, 6.424041e-09, 4.259284e-09, 2.906349e-09, 2.286192e-09, 
    1.695613e-09, 1.10256e-09, 7.819992e-10, 6.586786e-10, 6.566102e-10,
  1.858426e-08, 1.797804e-08, 1.723611e-08, 1.546907e-08, 1.309162e-08, 
    1.039462e-08, 7.734908e-09, 5.15623e-09, 3.393507e-09, 2.539159e-09, 
    1.922488e-09, 1.284422e-09, 8.510505e-10, 6.914201e-10, 6.306137e-10,
  1.895784e-08, 1.859032e-08, 1.779469e-08, 1.651628e-08, 1.438482e-08, 
    1.17576e-08, 9.059555e-09, 6.207566e-09, 4.000515e-09, 2.804526e-09, 
    2.162482e-09, 1.513254e-09, 9.606264e-10, 7.431554e-10, 6.318691e-10,
  1.973819e-08, 1.896533e-08, 1.814476e-08, 1.712891e-08, 1.558075e-08, 
    1.302821e-08, 1.031558e-08, 7.549946e-09, 4.938216e-09, 3.226709e-09, 
    2.40465e-09, 1.723933e-09, 1.094648e-09, 7.980392e-10, 6.390673e-10,
  2.008985e-08, 1.924138e-08, 1.846352e-08, 1.753379e-08, 1.651778e-08, 
    1.442352e-08, 1.158613e-08, 8.730613e-09, 5.812297e-09, 3.810112e-09, 
    2.690727e-09, 1.947333e-09, 1.264687e-09, 8.577155e-10, 6.469275e-10,
  2.075745e-08, 1.962879e-08, 1.865736e-08, 1.785142e-08, 1.708497e-08, 
    1.546699e-08, 1.303552e-08, 1.01312e-08, 7.114676e-09, 4.547169e-09, 
    3.061849e-09, 2.215482e-09, 1.451641e-09, 9.466713e-10, 6.686301e-10,
  2.195634e-08, 2.032729e-08, 1.915622e-08, 1.825845e-08, 1.770359e-08, 
    1.645806e-08, 1.404134e-08, 1.136132e-08, 8.43075e-09, 5.435667e-09, 
    3.482233e-09, 2.488812e-09, 1.652824e-09, 1.075792e-09, 7.170703e-10,
  2.267023e-08, 2.098805e-08, 1.960098e-08, 1.864898e-08, 1.814319e-08, 
    1.735937e-08, 1.538899e-08, 1.256515e-08, 9.619404e-09, 6.213641e-09, 
    3.941147e-09, 2.758732e-09, 1.858046e-09, 1.222326e-09, 7.884028e-10,
  2.338078e-08, 2.169998e-08, 2.008692e-08, 1.891448e-08, 1.841065e-08, 
    1.780174e-08, 1.637019e-08, 1.375045e-08, 1.0758e-08, 7.361138e-09, 
    4.542012e-09, 3.086414e-09, 2.081773e-09, 1.363307e-09, 8.739064e-10,
  1.850907e-08, 1.660398e-08, 1.426927e-08, 1.147379e-08, 8.56015e-09, 
    5.973785e-09, 4.092561e-09, 2.998701e-09, 2.287449e-09, 1.683382e-09, 
    1.257537e-09, 1.14318e-09, 1.101185e-09, 1.121176e-09, 9.137894e-10,
  1.896094e-08, 1.741573e-08, 1.534785e-08, 1.259042e-08, 9.662986e-09, 
    6.880424e-09, 4.686409e-09, 3.272035e-09, 2.432283e-09, 1.82983e-09, 
    1.347534e-09, 1.166405e-09, 1.113577e-09, 1.114952e-09, 9.608907e-10,
  1.939286e-08, 1.818362e-08, 1.629154e-08, 1.362437e-08, 1.080658e-08, 
    7.882421e-09, 5.40689e-09, 3.70127e-09, 2.664276e-09, 2.004584e-09, 
    1.470155e-09, 1.210108e-09, 1.133655e-09, 1.139042e-09, 1.029653e-09,
  1.965858e-08, 1.886074e-08, 1.719884e-08, 1.460351e-08, 1.187125e-08, 
    8.983947e-09, 6.257022e-09, 4.218328e-09, 2.912222e-09, 2.172133e-09, 
    1.597358e-09, 1.262036e-09, 1.148083e-09, 1.16291e-09, 1.073162e-09,
  2.006643e-08, 1.94296e-08, 1.792139e-08, 1.561832e-08, 1.2892e-08, 
    1.005521e-08, 7.202646e-09, 4.875065e-09, 3.242499e-09, 2.337757e-09, 
    1.724802e-09, 1.314612e-09, 1.159839e-09, 1.183949e-09, 1.104616e-09,
  2.01703e-08, 1.962892e-08, 1.840421e-08, 1.642484e-08, 1.397108e-08, 
    1.121599e-08, 8.212984e-09, 5.592181e-09, 3.65376e-09, 2.56739e-09, 
    1.88452e-09, 1.383531e-09, 1.187819e-09, 1.221014e-09, 1.123198e-09,
  1.979665e-08, 1.965727e-08, 1.873738e-08, 1.718145e-08, 1.481004e-08, 
    1.2165e-08, 9.385273e-09, 6.59692e-09, 4.263141e-09, 2.886162e-09, 
    2.100132e-09, 1.48148e-09, 1.227272e-09, 1.254418e-09, 1.129942e-09,
  2.01353e-08, 1.997862e-08, 1.908738e-08, 1.763427e-08, 1.571576e-08, 
    1.314556e-08, 1.042323e-08, 7.47614e-09, 4.852403e-09, 3.237702e-09, 
    2.32871e-09, 1.61547e-09, 1.267815e-09, 1.279029e-09, 1.130418e-09,
  2.066269e-08, 2.024619e-08, 1.934452e-08, 1.78426e-08, 1.63467e-08, 
    1.426157e-08, 1.14683e-08, 8.428731e-09, 5.585005e-09, 3.678277e-09, 
    2.557695e-09, 1.770994e-09, 1.315144e-09, 1.298066e-09, 1.131445e-09,
  2.124955e-08, 2.047626e-08, 1.947492e-08, 1.814391e-08, 1.679763e-08, 
    1.516232e-08, 1.247977e-08, 9.483731e-09, 6.491493e-09, 4.261407e-09, 
    2.83532e-09, 1.942231e-09, 1.370524e-09, 1.314755e-09, 1.135829e-09,
  2.341591e-08, 2.329124e-08, 2.22807e-08, 1.941345e-08, 1.484958e-08, 
    1.0003e-08, 6.010928e-09, 3.320804e-09, 2.121953e-09, 1.367968e-09, 
    8.197116e-10, 6.610754e-10, 7.000364e-10, 7.759524e-10, 6.708624e-10,
  2.344094e-08, 2.34476e-08, 2.287157e-08, 2.057061e-08, 1.644765e-08, 
    1.149718e-08, 7.039965e-09, 3.870483e-09, 2.327956e-09, 1.499216e-09, 
    8.738408e-10, 6.599022e-10, 7.017078e-10, 7.856238e-10, 6.680911e-10,
  2.345952e-08, 2.328295e-08, 2.314229e-08, 2.156287e-08, 1.78906e-08, 
    1.294703e-08, 8.16866e-09, 4.593857e-09, 2.702558e-09, 1.74752e-09, 
    1.014947e-09, 7.134318e-10, 7.308442e-10, 8.077922e-10, 6.822521e-10,
  2.351926e-08, 2.313973e-08, 2.31026e-08, 2.215569e-08, 1.909475e-08, 
    1.441481e-08, 9.326619e-09, 5.297966e-09, 3.085348e-09, 2.009265e-09, 
    1.172093e-09, 7.546306e-10, 7.377948e-10, 7.873489e-10, 6.532005e-10,
  2.340422e-08, 2.315236e-08, 2.313303e-08, 2.276287e-08, 2.002035e-08, 
    1.570004e-08, 1.059142e-08, 6.108842e-09, 3.50295e-09, 2.236197e-09, 
    1.303861e-09, 7.815072e-10, 7.27799e-10, 7.577053e-10, 6.195821e-10,
  2.350519e-08, 2.300703e-08, 2.281859e-08, 2.287196e-08, 2.091023e-08, 
    1.685386e-08, 1.169406e-08, 6.843326e-09, 3.875706e-09, 2.430767e-09, 
    1.392825e-09, 8.069806e-10, 7.287254e-10, 7.473491e-10, 6.034462e-10,
  2.384167e-08, 2.320806e-08, 2.279998e-08, 2.289785e-08, 2.132514e-08, 
    1.775423e-08, 1.290954e-08, 7.77746e-09, 4.275365e-09, 2.458138e-09, 
    1.390098e-09, 8.159094e-10, 7.386736e-10, 7.493623e-10, 5.967146e-10,
  2.419546e-08, 2.333909e-08, 2.275878e-08, 2.273426e-08, 2.190226e-08, 
    1.835429e-08, 1.373912e-08, 8.367122e-09, 4.404895e-09, 2.411595e-09, 
    1.341971e-09, 8.042693e-10, 7.476081e-10, 7.572761e-10, 5.978117e-10,
  2.424805e-08, 2.350075e-08, 2.277091e-08, 2.25409e-08, 2.221418e-08, 
    1.895839e-08, 1.43996e-08, 8.791102e-09, 4.584602e-09, 2.557964e-09, 
    1.360511e-09, 8.080868e-10, 7.560734e-10, 7.555666e-10, 6.049607e-10,
  2.431944e-08, 2.360894e-08, 2.284219e-08, 2.239839e-08, 2.193776e-08, 
    1.917527e-08, 1.508136e-08, 9.385856e-09, 5.01205e-09, 2.727155e-09, 
    1.409877e-09, 8.301146e-10, 7.641282e-10, 7.477874e-10, 6.040662e-10,
  2.583466e-08, 2.513889e-08, 2.242754e-08, 1.871009e-08, 1.263458e-08, 
    6.807408e-09, 2.589053e-09, 6.696451e-10, 6.344602e-10, 8.693496e-10, 
    9.899649e-10, 7.823451e-10, 4.99551e-10, 3.685474e-10, 3.069793e-10,
  2.543838e-08, 2.617702e-08, 2.363793e-08, 2.03314e-08, 1.473178e-08, 
    8.471305e-09, 3.44575e-09, 7.873484e-10, 6.19812e-10, 8.088649e-10, 
    9.736287e-10, 7.839427e-10, 4.996781e-10, 3.459518e-10, 2.531206e-10,
  2.391411e-08, 2.605107e-08, 2.475454e-08, 2.198167e-08, 1.684222e-08, 
    1.032719e-08, 4.490551e-09, 1.173962e-09, 5.969833e-10, 7.721274e-10, 
    9.769702e-10, 8.045579e-10, 5.219674e-10, 3.677562e-10, 2.375614e-10,
  2.293922e-08, 2.500714e-08, 2.546412e-08, 2.346561e-08, 1.888991e-08, 
    1.239244e-08, 5.728094e-09, 1.707358e-09, 5.734026e-10, 7.411758e-10, 
    9.688093e-10, 8.17057e-10, 5.326801e-10, 3.608836e-10, 2.170981e-10,
  2.259831e-08, 2.417271e-08, 2.577718e-08, 2.477959e-08, 2.069712e-08, 
    1.440608e-08, 7.187155e-09, 2.347069e-09, 5.689015e-10, 7.09475e-10, 
    9.583024e-10, 8.259226e-10, 5.402061e-10, 3.481185e-10, 2.117583e-10,
  2.295956e-08, 2.310454e-08, 2.516699e-08, 2.57106e-08, 2.249922e-08, 
    1.644043e-08, 8.684392e-09, 2.990127e-09, 6.352279e-10, 6.848592e-10, 
    9.509595e-10, 8.349696e-10, 5.527428e-10, 3.527166e-10, 2.105214e-10,
  2.354534e-08, 2.316278e-08, 2.424145e-08, 2.604259e-08, 2.376308e-08, 
    1.821605e-08, 1.030519e-08, 3.769709e-09, 8.238778e-10, 6.711733e-10, 
    9.45045e-10, 8.395731e-10, 5.553479e-10, 3.434157e-10, 2.070579e-10,
  2.393996e-08, 2.335081e-08, 2.346986e-08, 2.584055e-08, 2.550856e-08, 
    1.974766e-08, 1.16841e-08, 4.335636e-09, 9.785994e-10, 6.935289e-10, 
    9.370472e-10, 8.386343e-10, 5.420371e-10, 3.266694e-10, 2.02349e-10,
  2.405645e-08, 2.362895e-08, 2.319801e-08, 2.546979e-08, 2.643819e-08, 
    2.036132e-08, 1.259987e-08, 4.811145e-09, 1.159464e-09, 6.970526e-10, 
    9.311789e-10, 8.36009e-10, 5.198553e-10, 3.042132e-10, 1.968266e-10,
  2.405595e-08, 2.383293e-08, 2.317084e-08, 2.474523e-08, 2.625933e-08, 
    2.116221e-08, 1.364282e-08, 5.533716e-09, 1.343063e-09, 6.85987e-10, 
    9.261826e-10, 8.385432e-10, 5.042531e-10, 2.90965e-10, 2.037106e-10,
  2.464531e-08, 2.287436e-08, 1.987317e-08, 1.585296e-08, 1.089471e-08, 
    6.25953e-09, 2.893682e-09, 1.618274e-09, 1.163984e-09, 9.405379e-10, 
    7.678123e-10, 5.657438e-10, 4.00484e-10, 3.740007e-10, 3.963359e-10,
  2.515349e-08, 2.414587e-08, 2.140639e-08, 1.774411e-08, 1.292512e-08, 
    7.865857e-09, 3.703206e-09, 1.77635e-09, 1.21929e-09, 9.720442e-10, 
    8.02408e-10, 5.792811e-10, 3.856168e-10, 3.419551e-10, 3.628289e-10,
  2.520611e-08, 2.473828e-08, 2.272907e-08, 1.958194e-08, 1.493854e-08, 
    9.652256e-09, 4.833921e-09, 2.054685e-09, 1.307509e-09, 1.00491e-09, 
    8.496306e-10, 6.064853e-10, 3.89086e-10, 3.262183e-10, 3.37371e-10,
  2.490511e-08, 2.509278e-08, 2.37301e-08, 2.130259e-08, 1.691769e-08, 
    1.162882e-08, 6.231375e-09, 2.61937e-09, 1.385315e-09, 1.035298e-09, 
    8.888307e-10, 6.39482e-10, 4.017408e-10, 3.162953e-10, 3.177547e-10,
  2.420283e-08, 2.533161e-08, 2.470026e-08, 2.269002e-08, 1.876405e-08, 
    1.355955e-08, 7.858085e-09, 3.387269e-09, 1.498968e-09, 1.063088e-09, 
    9.171757e-10, 6.737664e-10, 4.197357e-10, 3.113488e-10, 3.057312e-10,
  2.275782e-08, 2.476362e-08, 2.509026e-08, 2.384333e-08, 2.05704e-08, 
    1.551522e-08, 9.596953e-09, 4.353528e-09, 1.722764e-09, 1.089532e-09, 
    9.356659e-10, 6.99903e-10, 4.358273e-10, 3.064959e-10, 2.933133e-10,
  2.235559e-08, 2.434324e-08, 2.526659e-08, 2.46729e-08, 2.199722e-08, 
    1.736847e-08, 1.17105e-08, 5.754071e-09, 2.115043e-09, 1.132515e-09, 
    9.504957e-10, 7.195122e-10, 4.440254e-10, 2.990121e-10, 2.802615e-10,
  2.201366e-08, 2.352182e-08, 2.494406e-08, 2.507938e-08, 2.377641e-08, 
    1.905211e-08, 1.358158e-08, 6.820807e-09, 2.39616e-09, 1.187483e-09, 
    9.661633e-10, 7.343616e-10, 4.443819e-10, 2.889296e-10, 2.670051e-10,
  2.177236e-08, 2.286385e-08, 2.449315e-08, 2.539795e-08, 2.482427e-08, 
    2.015822e-08, 1.50489e-08, 8.120959e-09, 2.966323e-09, 1.2707e-09, 
    9.906811e-10, 7.465701e-10, 4.448553e-10, 2.766057e-10, 2.548246e-10,
  2.179537e-08, 2.241372e-08, 2.394853e-08, 2.528141e-08, 2.532148e-08, 
    2.140566e-08, 1.678568e-08, 9.714875e-09, 3.808738e-09, 1.364869e-09, 
    1.017007e-09, 7.584084e-10, 4.45093e-10, 2.644515e-10, 2.392508e-10,
  2.22759e-08, 2.117527e-08, 1.90824e-08, 1.514035e-08, 1.032738e-08, 
    5.916037e-09, 2.882389e-09, 1.786624e-09, 1.341156e-09, 1.203516e-09, 
    1.102181e-09, 9.581287e-10, 7.696769e-10, 7.186441e-10, 7.904257e-10,
  2.251957e-08, 2.160994e-08, 1.974458e-08, 1.617096e-08, 1.128272e-08, 
    6.57319e-09, 3.136055e-09, 1.820317e-09, 1.384009e-09, 1.214423e-09, 
    1.128669e-09, 9.925367e-10, 8.229691e-10, 7.584111e-10, 8.109289e-10,
  2.285397e-08, 2.176413e-08, 2.023039e-08, 1.713333e-08, 1.232363e-08, 
    7.36192e-09, 3.557202e-09, 1.899447e-09, 1.426358e-09, 1.211692e-09, 
    1.154438e-09, 1.031464e-09, 8.531072e-10, 7.602768e-10, 7.87058e-10,
  2.309927e-08, 2.183168e-08, 2.064235e-08, 1.800916e-08, 1.331551e-08, 
    8.218892e-09, 4.038585e-09, 1.972174e-09, 1.45583e-09, 1.199861e-09, 
    1.169856e-09, 1.059063e-09, 8.831e-10, 7.680327e-10, 7.637976e-10,
  2.297459e-08, 2.220044e-08, 2.128333e-08, 1.885667e-08, 1.433698e-08, 
    9.056935e-09, 4.58378e-09, 2.065331e-09, 1.490267e-09, 1.196945e-09, 
    1.195522e-09, 1.091885e-09, 9.237288e-10, 7.890606e-10, 7.51458e-10,
  2.268716e-08, 2.225637e-08, 2.155508e-08, 1.959694e-08, 1.53927e-08, 
    9.974511e-09, 5.111158e-09, 2.19348e-09, 1.500745e-09, 1.205657e-09, 
    1.203098e-09, 1.128024e-09, 9.754021e-10, 8.083609e-10, 7.319775e-10,
  2.293971e-08, 2.267724e-08, 2.196644e-08, 2.012211e-08, 1.634352e-08, 
    1.095177e-08, 5.794808e-09, 2.441155e-09, 1.52354e-09, 1.239472e-09, 
    1.210857e-09, 1.166963e-09, 1.019839e-09, 8.258974e-10, 7.15292e-10,
  2.292357e-08, 2.288403e-08, 2.227004e-08, 2.057019e-08, 1.7333e-08, 
    1.182404e-08, 6.245734e-09, 2.566794e-09, 1.598773e-09, 1.318111e-09, 
    1.210314e-09, 1.190958e-09, 1.041594e-09, 8.461336e-10, 6.985005e-10,
  2.257673e-08, 2.275525e-08, 2.242458e-08, 2.109691e-08, 1.804909e-08, 
    1.221283e-08, 6.465801e-09, 2.656187e-09, 1.627449e-09, 1.311536e-09, 
    1.177526e-09, 1.191119e-09, 1.049626e-09, 8.655936e-10, 6.970073e-10,
  2.23767e-08, 2.287607e-08, 2.266153e-08, 2.150236e-08, 1.863836e-08, 
    1.290677e-08, 6.905781e-09, 2.881137e-09, 1.617715e-09, 1.296701e-09, 
    1.174112e-09, 1.186741e-09, 1.050719e-09, 8.605089e-10, 6.960597e-10,
  2.235508e-08, 2.237299e-08, 2.200089e-08, 2.013137e-08, 1.620358e-08, 
    1.111278e-08, 6.564372e-09, 3.609985e-09, 1.98542e-09, 1.088508e-09, 
    8.076296e-10, 6.498567e-10, 5.66734e-10, 5.758042e-10, 5.521502e-10,
  2.254232e-08, 2.267552e-08, 2.232673e-08, 2.133187e-08, 1.783406e-08, 
    1.288511e-08, 7.628201e-09, 4.07609e-09, 2.18451e-09, 1.147571e-09, 
    8.423254e-10, 6.765028e-10, 5.67328e-10, 5.387814e-10, 4.998618e-10,
  2.282159e-08, 2.25218e-08, 2.227637e-08, 2.205972e-08, 1.925556e-08, 
    1.467397e-08, 8.969329e-09, 4.777259e-09, 2.460879e-09, 1.248795e-09, 
    8.731079e-10, 7.098072e-10, 5.86528e-10, 5.48648e-10, 4.915395e-10,
  2.300673e-08, 2.220851e-08, 2.227432e-08, 2.261653e-08, 2.054698e-08, 
    1.63801e-08, 1.048244e-08, 5.566064e-09, 2.757118e-09, 1.353174e-09, 
    9.018207e-10, 7.357086e-10, 6.073019e-10, 5.625928e-10, 4.632286e-10,
  2.291593e-08, 2.206907e-08, 2.232421e-08, 2.2907e-08, 2.165222e-08, 
    1.780907e-08, 1.212518e-08, 6.526945e-09, 3.13974e-09, 1.449736e-09, 
    9.360814e-10, 7.544254e-10, 6.226406e-10, 5.733997e-10, 4.416084e-10,
  2.286187e-08, 2.227785e-08, 2.231896e-08, 2.300136e-08, 2.264018e-08, 
    1.92642e-08, 1.351728e-08, 7.431473e-09, 3.568761e-09, 1.549358e-09, 
    9.821953e-10, 7.74248e-10, 6.329116e-10, 5.799131e-10, 4.298944e-10,
  2.377922e-08, 2.277516e-08, 2.235928e-08, 2.296394e-08, 2.314315e-08, 
    2.047581e-08, 1.516644e-08, 8.561096e-09, 3.994211e-09, 1.654608e-09, 
    1.022219e-09, 7.980966e-10, 6.424877e-10, 5.776085e-10, 4.189518e-10,
  2.396533e-08, 2.289204e-08, 2.222506e-08, 2.266432e-08, 2.38235e-08, 
    2.133766e-08, 1.612102e-08, 9.231851e-09, 4.199385e-09, 1.778832e-09, 
    1.062548e-09, 8.117212e-10, 6.457184e-10, 5.690814e-10, 4.050354e-10,
  2.414988e-08, 2.307783e-08, 2.22905e-08, 2.268474e-08, 2.390439e-08, 
    2.173983e-08, 1.67761e-08, 9.809888e-09, 4.598304e-09, 1.921547e-09, 
    1.084263e-09, 8.145402e-10, 6.575203e-10, 5.63766e-10, 3.942548e-10,
  2.432928e-08, 2.337243e-08, 2.26236e-08, 2.270917e-08, 2.327578e-08, 
    2.207726e-08, 1.772721e-08, 1.077725e-08, 5.151937e-09, 2.027114e-09, 
    1.109901e-09, 8.205618e-10, 6.812555e-10, 5.635599e-10, 3.94148e-10,
  2.292393e-08, 1.903213e-08, 1.275902e-08, 6.530487e-09, 3.643813e-09, 
    2.342817e-09, 1.587027e-09, 1.058962e-09, 7.754353e-10, 7.061702e-10, 
    8.078568e-10, 9.176978e-10, 7.227191e-10, -4.019717e-11, 1.288842e-10,
  2.395264e-08, 2.066185e-08, 1.515774e-08, 8.161361e-09, 4.330526e-09, 
    2.646696e-09, 1.739354e-09, 1.158161e-09, 8.234998e-10, 7.198272e-10, 
    8.245895e-10, 9.326458e-10, 5.031431e-10, -1.116663e-10, 1.766442e-10,
  2.457321e-08, 2.22965e-08, 1.73471e-08, 1.018036e-08, 5.268008e-09, 
    3.067541e-09, 1.920807e-09, 1.27432e-09, 8.869712e-10, 7.484575e-10, 
    8.392587e-10, 9.479328e-10, 3.705817e-10, -6.287065e-11, 2.675627e-10,
  2.42247e-08, 2.351925e-08, 1.937179e-08, 1.25703e-08, 6.506344e-09, 
    3.67486e-09, 2.174123e-09, 1.394059e-09, 9.627601e-10, 7.789446e-10, 
    8.530986e-10, 9.460468e-10, 2.60138e-10, -1.677185e-11, 3.506072e-10,
  2.434401e-08, 2.411285e-08, 2.118786e-08, 1.498585e-08, 8.178141e-09, 
    4.454766e-09, 2.539722e-09, 1.547754e-09, 1.05027e-09, 8.236102e-10, 
    8.653363e-10, 9.305348e-10, 1.613017e-10, 5.491961e-11, 4.337441e-10,
  2.366851e-08, 2.42721e-08, 2.251575e-08, 1.737332e-08, 1.026721e-08, 
    5.574746e-09, 3.042668e-09, 1.712045e-09, 1.124836e-09, 8.724756e-10, 
    8.854212e-10, 9.086985e-10, 8.724425e-11, 1.227037e-10, 4.661134e-10,
  2.325104e-08, 2.40337e-08, 2.346523e-08, 1.969703e-08, 1.257715e-08, 
    6.937611e-09, 3.758468e-09, 1.998243e-09, 1.234283e-09, 9.32503e-10, 
    9.129253e-10, 8.936359e-10, 4.286424e-11, 1.62784e-10, 4.326213e-10,
  2.285967e-08, 2.400238e-08, 2.398935e-08, 2.158876e-08, 1.523814e-08, 
    8.53822e-09, 4.511417e-09, 2.290793e-09, 1.36265e-09, 9.959052e-10, 
    9.430348e-10, 8.867821e-10, 2.447252e-11, 1.767667e-10, 3.594404e-10,
  2.265564e-08, 2.352922e-08, 2.395772e-08, 2.286325e-08, 1.749772e-08, 
    1.016064e-08, 5.441486e-09, 2.671668e-09, 1.455494e-09, 1.016407e-09, 
    9.594319e-10, 8.891225e-10, 2.796574e-11, 1.747492e-10, 2.946097e-10,
  2.269712e-08, 2.339653e-08, 2.375988e-08, 2.332055e-08, 1.936253e-08, 
    1.211251e-08, 6.664792e-09, 3.265815e-09, 1.629955e-09, 1.054198e-09, 
    9.695718e-10, 8.906739e-10, 5.877315e-11, 1.896881e-10, 2.601173e-10,
  2.062374e-08, 1.61724e-08, 1.013148e-08, 5.520785e-09, 3.314332e-09, 
    1.985788e-09, 1.342183e-09, 1.142744e-09, 1.116051e-09, 1.261751e-09, 
    1.391688e-09, 1.212482e-09, 9.450722e-10, 6.598387e-10, 5.241414e-10,
  2.145774e-08, 1.763899e-08, 1.141243e-08, 6.094715e-09, 3.513634e-09, 
    2.079172e-09, 1.368812e-09, 1.141611e-09, 1.090574e-09, 1.241444e-09, 
    1.363327e-09, 1.112156e-09, 7.423977e-10, 4.786382e-10, 3.909804e-10,
  2.232382e-08, 1.876932e-08, 1.284051e-08, 6.768705e-09, 3.769549e-09, 
    2.154551e-09, 1.373228e-09, 1.137856e-09, 1.100572e-09, 1.270169e-09, 
    1.37689e-09, 1.050958e-09, 6.256355e-10, 4.182169e-10, 4.063794e-10,
  2.302642e-08, 2.005708e-08, 1.433484e-08, 7.638038e-09, 4.113346e-09, 
    2.280922e-09, 1.391585e-09, 1.126833e-09, 1.118763e-09, 1.293592e-09, 
    1.365478e-09, 9.760297e-10, 5.049658e-10, 3.742014e-10, 4.595631e-10,
  2.387561e-08, 2.123317e-08, 1.578158e-08, 8.718671e-09, 4.50167e-09, 
    2.408594e-09, 1.437069e-09, 1.138352e-09, 1.124306e-09, 1.287314e-09, 
    1.333439e-09, 9.093735e-10, 4.189136e-10, 3.900914e-10, 4.850221e-10,
  2.39704e-08, 2.218579e-08, 1.728006e-08, 1.000534e-08, 5.04586e-09, 
    2.607009e-09, 1.484425e-09, 1.135857e-09, 1.106584e-09, 1.270935e-09, 
    1.281494e-09, 8.195045e-10, 3.599792e-10, 4.102958e-10, 4.817098e-10,
  2.346475e-08, 2.264724e-08, 1.853211e-08, 1.153363e-08, 5.673061e-09, 
    2.812682e-09, 1.56858e-09, 1.163379e-09, 1.125507e-09, 1.263506e-09, 
    1.236687e-09, 7.249673e-10, 3.224138e-10, 4.194724e-10, 4.655235e-10,
  2.284439e-08, 2.305979e-08, 2.008874e-08, 1.318735e-08, 6.598373e-09, 
    3.109952e-09, 1.712473e-09, 1.201338e-09, 1.081869e-09, 1.247121e-09, 
    1.191789e-09, 6.555595e-10, 3.085968e-10, 4.178092e-10, 4.339707e-10,
  2.280043e-08, 2.345928e-08, 2.14481e-08, 1.495119e-08, 7.59935e-09, 
    3.512278e-09, 1.932983e-09, 1.2629e-09, 1.047527e-09, 1.237134e-09, 
    1.137824e-09, 5.869748e-10, 3.124189e-10, 4.050524e-10, 3.941255e-10,
  2.274055e-08, 2.363998e-08, 2.230573e-08, 1.669502e-08, 8.967912e-09, 
    4.008832e-09, 2.020464e-09, 1.291236e-09, 1.053416e-09, 1.241386e-09, 
    1.09246e-09, 5.217904e-10, 3.181508e-10, 4.018935e-10, 3.558243e-10,
  2.201125e-08, 1.944972e-08, 1.418486e-08, 1.052754e-08, 8.597803e-09, 
    6.514345e-09, 4.431433e-09, 2.647076e-09, 1.491497e-09, 8.997816e-10, 
    6.326696e-10, 5.412387e-10, 4.413956e-10, 3.282027e-10, 1.906126e-10,
  2.261037e-08, 2.066679e-08, 1.554697e-08, 1.103399e-08, 8.833339e-09, 
    6.675471e-09, 4.49934e-09, 2.63357e-09, 1.496022e-09, 9.059057e-10, 
    6.491372e-10, 5.466856e-10, 3.977435e-10, 2.46854e-10, 1.02616e-10,
  2.29704e-08, 2.173574e-08, 1.701596e-08, 1.170927e-08, 9.024457e-09, 
    6.857656e-09, 4.62407e-09, 2.652454e-09, 1.47334e-09, 8.844969e-10, 
    6.52503e-10, 5.494332e-10, 3.689903e-10, 2.235562e-10, 9.090022e-11,
  2.231475e-08, 2.242352e-08, 1.852438e-08, 1.264256e-08, 9.403167e-09, 
    7.130068e-09, 4.754474e-09, 2.685937e-09, 1.474264e-09, 8.889857e-10, 
    6.638921e-10, 5.490094e-10, 3.480585e-10, 2.055337e-10, 5.173217e-11,
  2.231326e-08, 2.289556e-08, 1.988932e-08, 1.38487e-08, 9.834056e-09, 
    7.394924e-09, 4.937852e-09, 2.778818e-09, 1.518704e-09, 9.170723e-10, 
    6.835216e-10, 5.50729e-10, 3.280755e-10, 1.689797e-10, -1.259951e-11,
  2.155242e-08, 2.291344e-08, 2.118528e-08, 1.526044e-08, 1.050171e-08, 
    7.723643e-09, 5.171388e-09, 2.876884e-09, 1.552014e-09, 9.387615e-10, 
    6.980446e-10, 5.478536e-10, 3.165468e-10, 1.125833e-10, -3.35291e-11,
  2.119454e-08, 2.235496e-08, 2.217357e-08, 1.678993e-08, 1.115352e-08, 
    8.083479e-09, 5.500567e-09, 2.964264e-09, 1.559529e-09, 9.411097e-10, 
    7.082353e-10, 5.413011e-10, 3.095231e-10, 6.211225e-11, -1.779907e-10,
  2.112957e-08, 2.192332e-08, 2.314519e-08, 1.837929e-08, 1.21261e-08, 
    8.488402e-09, 5.901549e-09, 3.167129e-09, 1.652747e-09, 9.319315e-10, 
    7.075672e-10, 5.281093e-10, 2.888785e-10, -4.595796e-11, -2.450311e-10,
  2.14515e-08, 2.171808e-08, 2.344433e-08, 1.964026e-08, 1.2969e-08, 
    8.91229e-09, 6.314729e-09, 3.477191e-09, 1.721417e-09, 8.813725e-10, 
    7.434554e-10, 5.280488e-10, 2.617722e-10, -1.367238e-10, -4.058964e-11,
  2.159961e-08, 2.154009e-08, 2.351448e-08, 2.079186e-08, 1.428557e-08, 
    9.495086e-09, 6.651962e-09, 3.551979e-09, 1.658513e-09, 9.193785e-10, 
    8.111236e-10, 5.382486e-10, 2.446657e-10, -1.461509e-10, 4.944955e-11,
  2.018057e-08, 1.939024e-08, 1.841837e-08, 1.664002e-08, 1.431917e-08, 
    1.23749e-08, 9.932893e-09, 7.071621e-09, 4.531342e-09, 2.380323e-09, 
    5.540762e-10, 1.681598e-10, 1.884314e-10, 4.408251e-10, 7.167612e-10,
  2.055384e-08, 1.96955e-08, 1.862911e-08, 1.714101e-08, 1.466999e-08, 
    1.25434e-08, 9.998684e-09, 7.04749e-09, 4.420451e-09, 2.233069e-09, 
    4.854495e-10, 1.702558e-10, 2.028245e-10, 5.019162e-10, 7.025365e-10,
  2.115635e-08, 2.019367e-08, 1.884718e-08, 1.734114e-08, 1.514213e-08, 
    1.280533e-08, 1.021667e-08, 7.158866e-09, 4.368967e-09, 2.093381e-09, 
    4.324514e-10, 1.723804e-10, 2.291853e-10, 5.521885e-10, 6.365989e-10,
  2.169962e-08, 2.03089e-08, 1.920255e-08, 1.77597e-08, 1.56515e-08, 
    1.314514e-08, 1.041487e-08, 7.210357e-09, 4.287742e-09, 1.936831e-09, 
    3.897093e-10, 1.88404e-10, 2.796685e-10, 5.820214e-10, 6.084706e-10,
  2.283139e-08, 2.078585e-08, 1.948917e-08, 1.80205e-08, 1.61287e-08, 
    1.343709e-08, 1.068894e-08, 7.271079e-09, 4.164708e-09, 1.792608e-09, 
    3.625702e-10, 2.019554e-10, 3.28002e-10, 5.688351e-10, 5.955808e-10,
  2.290855e-08, 2.108743e-08, 1.984613e-08, 1.827344e-08, 1.670881e-08, 
    1.387076e-08, 1.077466e-08, 7.209088e-09, 4.089392e-09, 1.708177e-09, 
    3.425679e-10, 2.045496e-10, 3.694624e-10, 5.322454e-10, 6.142351e-10,
  2.291368e-08, 2.159613e-08, 2.03136e-08, 1.863446e-08, 1.70018e-08, 
    1.42935e-08, 1.115464e-08, 7.317059e-09, 4.026489e-09, 1.677293e-09, 
    3.281134e-10, 2.110309e-10, 4.288375e-10, 4.899155e-10, 6.448665e-10,
  2.280791e-08, 2.194412e-08, 2.077255e-08, 1.901127e-08, 1.75382e-08, 
    1.480614e-08, 1.141907e-08, 7.454387e-09, 3.958491e-09, 1.654354e-09, 
    3.062979e-10, 2.259207e-10, 4.628208e-10, 4.663474e-10, 6.450227e-10,
  2.293376e-08, 2.21976e-08, 2.113843e-08, 1.937526e-08, 1.768427e-08, 
    1.516019e-08, 1.150382e-08, 7.512054e-09, 4.138048e-09, 1.727363e-09, 
    3.012733e-10, 2.419484e-10, 4.608779e-10, 4.408376e-10, 6.134757e-10,
  2.295437e-08, 2.219589e-08, 2.153756e-08, 1.972756e-08, 1.788621e-08, 
    1.548241e-08, 1.182214e-08, 7.713069e-09, 4.258263e-09, 1.745497e-09, 
    3.045602e-10, 2.598158e-10, 4.306068e-10, 3.915012e-10, 5.669854e-10,
  2.082696e-08, 2.061993e-08, 2.067492e-08, 1.974686e-08, 1.824976e-08, 
    1.709216e-08, 1.589246e-08, 1.389004e-08, 1.100111e-08, 7.540612e-09, 
    4.305853e-09, 1.969335e-09, 8.973746e-10, 5.012568e-10, 2.132867e-10,
  2.131473e-08, 2.079764e-08, 2.054889e-08, 2.004333e-08, 1.864855e-08, 
    1.738933e-08, 1.614612e-08, 1.417636e-08, 1.126278e-08, 7.675856e-09, 
    4.310774e-09, 1.941472e-09, 8.314112e-10, 3.949598e-10, 1.068899e-10,
  2.181681e-08, 2.17216e-08, 2.088878e-08, 2.008257e-08, 1.904374e-08, 
    1.76635e-08, 1.641063e-08, 1.452781e-08, 1.148316e-08, 7.813944e-09, 
    4.387587e-09, 1.980337e-09, 8.321233e-10, 3.442371e-10, 6.318776e-11,
  2.214433e-08, 2.191398e-08, 2.127699e-08, 2.031585e-08, 1.934369e-08, 
    1.811577e-08, 1.668245e-08, 1.477066e-08, 1.167372e-08, 7.905387e-09, 
    4.419393e-09, 1.98374e-09, 8.212994e-10, 3.04501e-10, 5.551348e-11,
  2.363726e-08, 2.261143e-08, 2.171516e-08, 2.057047e-08, 1.972818e-08, 
    1.846725e-08, 1.709743e-08, 1.504837e-08, 1.181759e-08, 7.947558e-09, 
    4.443532e-09, 1.97141e-09, 8.098213e-10, 2.748031e-10, 5.688193e-11,
  2.366042e-08, 2.25629e-08, 2.195747e-08, 2.071982e-08, 2.006616e-08, 
    1.907095e-08, 1.733212e-08, 1.520229e-08, 1.203557e-08, 8.057911e-09, 
    4.511903e-09, 1.959954e-09, 7.926406e-10, 2.499113e-10, 6.138407e-11,
  2.297414e-08, 2.262856e-08, 2.199416e-08, 2.117149e-08, 2.019268e-08, 
    1.945449e-08, 1.815843e-08, 1.568055e-08, 1.228743e-08, 8.199438e-09, 
    4.594072e-09, 1.968808e-09, 7.807202e-10, 2.478291e-10, 8.681909e-11,
  2.254126e-08, 2.276196e-08, 2.219679e-08, 2.139977e-08, 2.095188e-08, 
    1.991887e-08, 1.861249e-08, 1.585728e-08, 1.219735e-08, 8.268019e-09, 
    4.661537e-09, 1.967382e-09, 7.767799e-10, 2.723089e-10, 1.160235e-10,
  2.229734e-08, 2.278884e-08, 2.219111e-08, 2.167818e-08, 2.093709e-08, 
    2.005949e-08, 1.833271e-08, 1.58777e-08, 1.265869e-08, 8.581035e-09, 
    4.716258e-09, 1.948997e-09, 7.740928e-10, 3.023264e-10, 1.299716e-10,
  2.196365e-08, 2.277915e-08, 2.236154e-08, 2.190484e-08, 2.068592e-08, 
    2.009402e-08, 1.898125e-08, 1.623103e-08, 1.294215e-08, 8.779528e-09, 
    4.747429e-09, 1.944197e-09, 7.719955e-10, 3.24261e-10, 1.226342e-10,
  2.121885e-08, 1.99551e-08, 1.849251e-08, 1.808408e-08, 1.917235e-08, 
    1.885266e-08, 1.643477e-08, 1.295605e-08, 9.037359e-09, 4.936812e-09, 
    1.867572e-09, 7.716287e-10, 4.648012e-10, 2.932387e-10, 1.12922e-10,
  2.172196e-08, 2.058926e-08, 1.89275e-08, 1.816255e-08, 1.882589e-08, 
    1.915316e-08, 1.709638e-08, 1.383289e-08, 9.920567e-09, 5.676498e-09, 
    2.254742e-09, 8.527276e-10, 4.730155e-10, 2.643625e-10, 9.630702e-11,
  2.189207e-08, 2.135818e-08, 1.966353e-08, 1.839111e-08, 1.85429e-08, 
    1.918307e-08, 1.766265e-08, 1.466524e-08, 1.075519e-08, 6.419124e-09, 
    2.75531e-09, 9.585023e-10, 4.80108e-10, 2.538229e-10, 6.928021e-11,
  2.155262e-08, 2.174115e-08, 2.043308e-08, 1.878704e-08, 1.843034e-08, 
    1.920402e-08, 1.81275e-08, 1.53491e-08, 1.150958e-08, 7.130503e-09, 
    3.292705e-09, 1.089597e-09, 4.890635e-10, 2.437861e-10, 6.902529e-11,
  2.250037e-08, 2.218905e-08, 2.11233e-08, 1.937448e-08, 1.847248e-08, 
    1.890642e-08, 1.854889e-08, 1.621921e-08, 1.233975e-08, 7.869263e-09, 
    3.88303e-09, 1.247385e-09, 5.051925e-10, 2.329232e-10, 3.499218e-11,
  2.257696e-08, 2.215582e-08, 2.144991e-08, 1.992695e-08, 1.871105e-08, 
    1.894371e-08, 1.84614e-08, 1.65796e-08, 1.299712e-08, 8.599177e-09, 
    4.480505e-09, 1.418118e-09, 5.199628e-10, 2.169915e-10, 5.287292e-12,
  2.249311e-08, 2.220154e-08, 2.158406e-08, 2.040075e-08, 1.895312e-08, 
    1.884973e-08, 1.874313e-08, 1.728054e-08, 1.378052e-08, 9.355327e-09, 
    5.004015e-09, 1.606863e-09, 5.253217e-10, 2.051664e-10, -3.311619e-12,
  2.205298e-08, 2.220177e-08, 2.189267e-08, 2.075321e-08, 1.953961e-08, 
    1.885742e-08, 1.865484e-08, 1.76631e-08, 1.45865e-08, 1.001244e-08, 
    5.445691e-09, 1.773223e-09, 5.243045e-10, 1.983504e-10, 1.527878e-11,
  2.192923e-08, 2.226724e-08, 2.201698e-08, 2.100739e-08, 1.97929e-08, 
    1.909154e-08, 1.884147e-08, 1.824844e-08, 1.559405e-08, 1.092912e-08, 
    5.885854e-09, 1.92263e-09, 5.303701e-10, 2.028118e-10, 3.966811e-11,
  2.148389e-08, 2.205188e-08, 2.206705e-08, 2.147423e-08, 2.027771e-08, 
    1.937904e-08, 1.883934e-08, 1.816085e-08, 1.601275e-08, 1.167208e-08, 
    6.290152e-09, 2.084929e-09, 5.643819e-10, 2.199166e-10, 7.119055e-11,
  2.176054e-08, 2.04561e-08, 1.863186e-08, 1.809539e-08, 1.952075e-08, 
    1.980653e-08, 1.654105e-08, 1.186961e-08, 6.94487e-09, 2.98845e-09, 
    1.309433e-09, 8.252297e-10, 6.924935e-10, 5.614003e-10, 4.442292e-10,
  2.252164e-08, 2.123145e-08, 1.912294e-08, 1.803705e-08, 1.912719e-08, 
    2.009568e-08, 1.720002e-08, 1.251892e-08, 7.460537e-09, 3.184247e-09, 
    1.383661e-09, 8.310743e-10, 6.350815e-10, 4.489778e-10, 3.495025e-10,
  2.285481e-08, 2.146789e-08, 1.948746e-08, 1.80526e-08, 1.866099e-08, 
    2.009896e-08, 1.773896e-08, 1.314517e-08, 7.922815e-09, 3.385825e-09, 
    1.436484e-09, 8.057796e-10, 5.794052e-10, 3.477311e-10, 3.60996e-10,
  2.310673e-08, 2.158372e-08, 1.992607e-08, 1.831106e-08, 1.838925e-08, 
    2.018567e-08, 1.816951e-08, 1.360573e-08, 8.388925e-09, 3.573757e-09, 
    1.438992e-09, 7.544591e-10, 4.986416e-10, 2.711135e-10, 3.633145e-10,
  2.296776e-08, 2.205559e-08, 2.042928e-08, 1.849263e-08, 1.810977e-08, 
    1.993404e-08, 1.855738e-08, 1.407555e-08, 8.721732e-09, 3.650894e-09, 
    1.387081e-09, 6.847412e-10, 4.327095e-10, 2.267676e-10, 3.512705e-10,
  2.223669e-08, 2.192345e-08, 2.070982e-08, 1.878542e-08, 1.811673e-08, 
    1.986366e-08, 1.853928e-08, 1.418606e-08, 8.874749e-09, 3.64553e-09, 
    1.320184e-09, 6.360541e-10, 3.963072e-10, 2.107086e-10, 2.900182e-10,
  2.250749e-08, 2.266814e-08, 2.12437e-08, 1.907691e-08, 1.794945e-08, 
    1.961164e-08, 1.882604e-08, 1.441564e-08, 8.995067e-09, 3.643374e-09, 
    1.293627e-09, 6.121345e-10, 3.750715e-10, 2.161018e-10, 2.18809e-10,
  2.245876e-08, 2.285454e-08, 2.158994e-08, 1.92685e-08, 1.812749e-08, 
    1.937993e-08, 1.896525e-08, 1.457514e-08, 9.09395e-09, 3.671363e-09, 
    1.31289e-09, 6.01715e-10, 3.514973e-10, 2.235782e-10, 1.61331e-10,
  2.244372e-08, 2.296525e-08, 2.187594e-08, 1.965547e-08, 1.818322e-08, 
    1.919867e-08, 1.901117e-08, 1.477205e-08, 9.164027e-09, 3.715255e-09, 
    1.30576e-09, 5.820689e-10, 3.203338e-10, 2.185686e-10, 8.610414e-11,
  2.245529e-08, 2.29852e-08, 2.212901e-08, 1.98766e-08, 1.822576e-08, 
    1.905657e-08, 1.89675e-08, 1.472867e-08, 9.079416e-09, 3.709406e-09, 
    1.261132e-09, 5.331255e-10, 2.721679e-10, 1.121176e-10, 7.290263e-12,
  1.842719e-08, 1.882328e-08, 1.967138e-08, 2.040672e-08, 2.080611e-08, 
    1.989047e-08, 1.753408e-08, 1.41566e-08, 1.080014e-08, 7.44057e-09, 
    5.320394e-09, 4.1894e-09, 3.146894e-09, 2.154322e-09, 1.265145e-09,
  1.857397e-08, 1.870657e-08, 1.950118e-08, 2.011488e-08, 2.074044e-08, 
    2.032547e-08, 1.81896e-08, 1.485085e-08, 1.14258e-08, 7.871869e-09, 
    5.471916e-09, 4.210623e-09, 3.100186e-09, 2.017257e-09, 1.03503e-09,
  1.877057e-08, 1.865093e-08, 1.91289e-08, 1.97748e-08, 2.059219e-08, 
    2.053597e-08, 1.885594e-08, 1.555806e-08, 1.199211e-08, 8.240025e-09, 
    5.589111e-09, 4.232328e-09, 3.097961e-09, 1.934525e-09, 9.134912e-10,
  1.885961e-08, 1.837945e-08, 1.906083e-08, 1.950839e-08, 2.036874e-08, 
    2.077714e-08, 1.925243e-08, 1.599311e-08, 1.239821e-08, 8.514134e-09, 
    5.661156e-09, 4.219843e-09, 3.05892e-09, 1.837575e-09, 7.889307e-10,
  1.898628e-08, 1.830019e-08, 1.865254e-08, 1.926029e-08, 2.007489e-08, 
    2.075365e-08, 1.985684e-08, 1.657242e-08, 1.280221e-08, 8.748446e-09, 
    5.689927e-09, 4.172287e-09, 2.986985e-09, 1.676187e-09, 6.278728e-10,
  1.881442e-08, 1.820509e-08, 1.848565e-08, 1.898835e-08, 1.995399e-08, 
    2.093961e-08, 1.995641e-08, 1.674117e-08, 1.301049e-08, 8.836349e-09, 
    5.667944e-09, 4.097565e-09, 2.852816e-09, 1.537177e-09, 5.033694e-10,
  1.907495e-08, 1.840008e-08, 1.84234e-08, 1.884695e-08, 1.961261e-08, 
    2.092516e-08, 2.069016e-08, 1.736774e-08, 1.326207e-08, 8.883506e-09, 
    5.6158e-09, 4.00864e-09, 2.719824e-09, 1.338635e-09, 4.382166e-10,
  1.952448e-08, 1.870656e-08, 1.846811e-08, 1.866528e-08, 1.987173e-08, 
    2.101966e-08, 2.093756e-08, 1.739721e-08, 1.324723e-08, 8.831742e-09, 
    5.549689e-09, 3.913466e-09, 2.575122e-09, 1.088299e-09, 3.709814e-10,
  1.98227e-08, 1.885752e-08, 1.846898e-08, 1.86719e-08, 1.960366e-08, 
    2.093105e-08, 2.08134e-08, 1.712888e-08, 1.306718e-08, 8.746669e-09, 
    5.451847e-09, 3.788148e-09, 2.373689e-09, 8.179841e-10, 3.055336e-10,
  1.991635e-08, 1.893958e-08, 1.847071e-08, 1.853076e-08, 1.932454e-08, 
    2.109909e-08, 2.113394e-08, 1.727157e-08, 1.31279e-08, 8.602157e-09, 
    5.276655e-09, 3.621025e-09, 2.085852e-09, 6.13987e-10, 2.329989e-10,
  2.519632e-08, 2.487283e-08, 2.361583e-08, 2.255772e-08, 2.131959e-08, 
    1.914342e-08, 1.629083e-08, 1.393737e-08, 1.16744e-08, 9.097693e-09, 
    6.512525e-09, 4.214051e-09, 2.436004e-09, 1.209509e-09, 5.948153e-10,
  2.556198e-08, 2.491199e-08, 2.380093e-08, 2.26736e-08, 2.154705e-08, 
    1.964366e-08, 1.676401e-08, 1.420595e-08, 1.191781e-08, 9.359537e-09, 
    6.687473e-09, 4.177972e-09, 2.347064e-09, 1.109394e-09, 4.85004e-10,
  2.57952e-08, 2.501176e-08, 2.387972e-08, 2.277848e-08, 2.195122e-08, 
    2.009215e-08, 1.721789e-08, 1.450925e-08, 1.215375e-08, 9.546469e-09, 
    6.770977e-09, 4.13704e-09, 2.263721e-09, 9.723027e-10, 3.531082e-10,
  2.531712e-08, 2.441097e-08, 2.399501e-08, 2.313221e-08, 2.22214e-08, 
    2.048984e-08, 1.753667e-08, 1.466353e-08, 1.223304e-08, 9.648313e-09, 
    6.738807e-09, 4.015881e-09, 2.137555e-09, 8.248257e-10, 3.096109e-10,
  2.526011e-08, 2.442919e-08, 2.387902e-08, 2.312792e-08, 2.24258e-08, 
    2.07179e-08, 1.787571e-08, 1.489027e-08, 1.236994e-08, 9.650456e-09, 
    6.585402e-09, 3.770384e-09, 1.969558e-09, 7.13861e-10, 2.423924e-10,
  2.419133e-08, 2.378831e-08, 2.374776e-08, 2.323679e-08, 2.262335e-08, 
    2.099357e-08, 1.794568e-08, 1.485521e-08, 1.220358e-08, 9.561199e-09, 
    6.334095e-09, 3.430925e-09, 1.754783e-09, 6.076775e-10, 1.770462e-10,
  2.443386e-08, 2.371843e-08, 2.351343e-08, 2.299496e-08, 2.26035e-08, 
    2.104076e-08, 1.822899e-08, 1.506248e-08, 1.224236e-08, 9.256531e-09, 
    5.957136e-09, 3.015421e-09, 1.503171e-09, 4.670034e-10, 1.716591e-10,
  2.438382e-08, 2.367302e-08, 2.321953e-08, 2.301714e-08, 2.273581e-08, 
    2.108894e-08, 1.817018e-08, 1.477115e-08, 1.172322e-08, 8.747146e-09, 
    5.437036e-09, 2.666766e-09, 1.239901e-09, 2.917104e-10, 1.880095e-10,
  2.430823e-08, 2.343369e-08, 2.292701e-08, 2.28957e-08, 2.274072e-08, 
    2.081338e-08, 1.758417e-08, 1.404092e-08, 1.112741e-08, 8.235872e-09, 
    4.797846e-09, 2.335067e-09, 1.004492e-09, 1.591591e-10, 2.149509e-10,
  2.45525e-08, 2.347316e-08, 2.276882e-08, 2.285697e-08, 2.246782e-08, 
    2.064647e-08, 1.750548e-08, 1.392837e-08, 1.093687e-08, 7.672722e-09, 
    4.108741e-09, 1.993355e-09, 7.729377e-10, 1.299349e-10, 2.6409e-10,
  2.212017e-08, 2.165269e-08, 2.11602e-08, 2.061371e-08, 1.947529e-08, 
    1.77944e-08, 1.511795e-08, 1.205231e-08, 8.092882e-09, 4.631985e-09, 
    2.274303e-09, 1.548028e-09, 1.43919e-09, 1.006658e-09, 4.530076e-10,
  2.277926e-08, 2.230997e-08, 2.154789e-08, 2.102245e-08, 1.996458e-08, 
    1.863153e-08, 1.629152e-08, 1.345262e-08, 9.459403e-09, 5.661009e-09, 
    2.743731e-09, 1.630263e-09, 1.497441e-09, 1.084338e-09, 4.781714e-10,
  2.321511e-08, 2.249063e-08, 2.167781e-08, 2.13071e-08, 2.049653e-08, 
    1.928515e-08, 1.726604e-08, 1.47933e-08, 1.09315e-08, 6.718631e-09, 
    3.341984e-09, 1.747724e-09, 1.536137e-09, 1.131156e-09, 4.733112e-10,
  2.347509e-08, 2.267113e-08, 2.219815e-08, 2.181088e-08, 2.094764e-08, 
    1.989443e-08, 1.809958e-08, 1.580826e-08, 1.225444e-08, 7.790693e-09, 
    3.993995e-09, 1.892635e-09, 1.573797e-09, 1.171637e-09, 4.615777e-10,
  2.364683e-08, 2.299658e-08, 2.252444e-08, 2.214851e-08, 2.128536e-08, 
    2.024238e-08, 1.877916e-08, 1.689564e-08, 1.359765e-08, 8.882841e-09, 
    4.671822e-09, 2.083308e-09, 1.615612e-09, 1.192578e-09, 4.282165e-10,
  2.338665e-08, 2.347907e-08, 2.328276e-08, 2.271458e-08, 2.174197e-08, 
    2.087342e-08, 1.913112e-08, 1.738006e-08, 1.463045e-08, 9.950798e-09, 
    5.298609e-09, 2.292711e-09, 1.651173e-09, 1.196714e-09, 3.767252e-10,
  2.370872e-08, 2.39813e-08, 2.367361e-08, 2.290008e-08, 2.17867e-08, 
    2.108667e-08, 1.988571e-08, 1.833007e-08, 1.569759e-08, 1.09378e-08, 
    5.884785e-09, 2.476345e-09, 1.665718e-09, 1.177513e-09, 3.481496e-10,
  2.391682e-08, 2.413828e-08, 2.355181e-08, 2.296136e-08, 2.231828e-08, 
    2.132756e-08, 2.015813e-08, 1.863167e-08, 1.634949e-08, 1.179302e-08, 
    6.404304e-09, 2.616056e-09, 1.68135e-09, 1.128228e-09, 3.633293e-10,
  2.395426e-08, 2.399889e-08, 2.363647e-08, 2.334806e-08, 2.274424e-08, 
    2.112762e-08, 2.008708e-08, 1.88718e-08, 1.713781e-08, 1.269131e-08, 
    6.831895e-09, 2.705145e-09, 1.673897e-09, 1.036853e-09, 3.789126e-10,
  2.417991e-08, 2.400827e-08, 2.386058e-08, 2.376496e-08, 2.290866e-08, 
    2.133663e-08, 2.049471e-08, 1.910117e-08, 1.761183e-08, 1.330943e-08, 
    7.18108e-09, 2.714182e-09, 1.641274e-09, 9.29987e-10, 3.81195e-10,
  2.248656e-08, 2.1731e-08, 1.979e-08, 1.677135e-08, 1.241061e-08, 
    8.435056e-09, 5.154929e-09, 3.003567e-09, 1.82356e-09, 1.301128e-09, 
    1.117349e-09, 9.862088e-10, 8.504937e-10, 8.144155e-10, 7.139414e-10,
  2.241958e-08, 2.241402e-08, 2.086106e-08, 1.83049e-08, 1.435761e-08, 
    1.006828e-08, 6.297411e-09, 3.681058e-09, 2.113444e-09, 1.410959e-09, 
    1.126649e-09, 9.985851e-10, 8.753689e-10, 8.466131e-10, 7.330933e-10,
  2.209333e-08, 2.2461e-08, 2.164128e-08, 1.951421e-08, 1.608736e-08, 
    1.18079e-08, 7.630972e-09, 4.521026e-09, 2.558169e-09, 1.589026e-09, 
    1.171559e-09, 9.980659e-10, 8.867327e-10, 8.613049e-10, 7.38011e-10,
  2.183082e-08, 2.225316e-08, 2.210518e-08, 2.064107e-08, 1.764406e-08, 
    1.357997e-08, 9.09762e-09, 5.485934e-09, 3.079422e-09, 1.807269e-09, 
    1.255577e-09, 1.006059e-09, 8.997953e-10, 8.7796e-10, 7.481722e-10,
  2.155315e-08, 2.178534e-08, 2.236909e-08, 2.13559e-08, 1.891864e-08, 
    1.524607e-08, 1.07568e-08, 6.631439e-09, 3.79122e-09, 2.098954e-09, 
    1.36602e-09, 1.031428e-09, 9.110872e-10, 8.947144e-10, 7.575687e-10,
  2.18139e-08, 2.153139e-08, 2.222345e-08, 2.190832e-08, 2.01021e-08, 
    1.687146e-08, 1.240485e-08, 7.843389e-09, 4.536938e-09, 2.443013e-09, 
    1.496202e-09, 1.063645e-09, 9.213597e-10, 9.144568e-10, 7.715486e-10,
  2.220736e-08, 2.173035e-08, 2.191708e-08, 2.218225e-08, 2.084486e-08, 
    1.824728e-08, 1.431239e-08, 9.485332e-09, 5.560553e-09, 2.92192e-09, 
    1.661616e-09, 1.110479e-09, 9.34351e-10, 9.358677e-10, 7.864823e-10,
  2.296054e-08, 2.193537e-08, 2.174697e-08, 2.228253e-08, 2.167074e-08, 
    1.9211e-08, 1.54849e-08, 1.062185e-08, 6.459256e-09, 3.433511e-09, 
    1.837479e-09, 1.16014e-09, 9.504105e-10, 9.626888e-10, 8.057521e-10,
  2.354455e-08, 2.223954e-08, 2.180086e-08, 2.2275e-08, 2.217912e-08, 
    2.005386e-08, 1.679219e-08, 1.196208e-08, 7.342224e-09, 3.950168e-09, 
    2.011212e-09, 1.198617e-09, 9.668603e-10, 9.911438e-10, 8.255086e-10,
  2.399801e-08, 2.264426e-08, 2.194623e-08, 2.222474e-08, 2.208812e-08, 
    2.041524e-08, 1.773402e-08, 1.335021e-08, 8.544595e-09, 4.647035e-09, 
    2.237701e-09, 1.244153e-09, 9.804378e-10, 1.017635e-09, 8.442468e-10,
  2.447914e-08, 2.249191e-08, 2.003214e-08, 1.725417e-08, 1.422881e-08, 
    1.101941e-08, 7.283855e-09, 4.806996e-09, 2.94474e-09, 1.923553e-09, 
    1.396295e-09, 1.054606e-09, 8.405912e-10, 7.253239e-10, 6.084671e-10,
  2.516648e-08, 2.376034e-08, 2.130807e-08, 1.855713e-08, 1.560677e-08, 
    1.234059e-08, 8.402758e-09, 5.373843e-09, 3.318484e-09, 2.076546e-09, 
    1.458675e-09, 1.090669e-09, 8.679911e-10, 7.543582e-10, 6.111234e-10,
  2.524833e-08, 2.432869e-08, 2.236115e-08, 1.987497e-08, 1.690244e-08, 
    1.370889e-08, 9.749937e-09, 6.05831e-09, 3.787294e-09, 2.281388e-09, 
    1.554592e-09, 1.126109e-09, 8.965103e-10, 7.725343e-10, 5.9771e-10,
  2.49121e-08, 2.451403e-08, 2.323551e-08, 2.111971e-08, 1.821954e-08, 
    1.51382e-08, 1.116369e-08, 6.899178e-09, 4.263526e-09, 2.510927e-09, 
    1.660001e-09, 1.153637e-09, 9.274808e-10, 7.945329e-10, 5.884333e-10,
  2.484565e-08, 2.496756e-08, 2.400064e-08, 2.218319e-08, 1.935991e-08, 
    1.64398e-08, 1.257041e-08, 8.044825e-09, 4.846356e-09, 2.7665e-09, 
    1.750622e-09, 1.17882e-09, 9.583084e-10, 8.157641e-10, 5.753555e-10,
  2.427094e-08, 2.465262e-08, 2.449466e-08, 2.302052e-08, 2.057311e-08, 
    1.773921e-08, 1.388175e-08, 9.189898e-09, 5.371384e-09, 3.052026e-09, 
    1.841312e-09, 1.199818e-09, 9.801745e-10, 8.374557e-10, 5.653488e-10,
  2.430241e-08, 2.464508e-08, 2.470365e-08, 2.372481e-08, 2.144518e-08, 
    1.891262e-08, 1.548198e-08, 1.07411e-08, 6.223563e-09, 3.404031e-09, 
    1.94537e-09, 1.241428e-09, 9.922131e-10, 8.625599e-10, 5.630356e-10,
  2.38948e-08, 2.444758e-08, 2.466055e-08, 2.418522e-08, 2.272339e-08, 
    1.993562e-08, 1.652645e-08, 1.176045e-08, 6.928233e-09, 3.758225e-09, 
    2.074173e-09, 1.29913e-09, 9.900508e-10, 8.796941e-10, 5.615621e-10,
  2.359426e-08, 2.434104e-08, 2.462363e-08, 2.45877e-08, 2.355437e-08, 
    2.074595e-08, 1.742639e-08, 1.285029e-08, 7.684819e-09, 4.132664e-09, 
    2.218711e-09, 1.362758e-09, 9.800517e-10, 8.975749e-10, 5.639709e-10,
  2.355082e-08, 2.409874e-08, 2.44915e-08, 2.482296e-08, 2.387187e-08, 
    2.134291e-08, 1.836715e-08, 1.429341e-08, 8.975196e-09, 4.59364e-09, 
    2.329281e-09, 1.412893e-09, 9.800809e-10, 9.112948e-10, 5.77166e-10,
  2.242466e-08, 2.047102e-08, 1.783643e-08, 1.404367e-08, 1.079708e-08, 
    8.611862e-09, 6.584063e-09, 4.65409e-09, 3.428477e-09, 2.608983e-09, 
    1.839798e-09, 1.223833e-09, 4.866844e-10, 4.622026e-11, 4.146134e-11,
  2.354739e-08, 2.203388e-08, 1.974007e-08, 1.636937e-08, 1.248224e-08, 
    9.741655e-09, 7.565574e-09, 5.391224e-09, 3.817461e-09, 2.910783e-09, 
    2.169271e-09, 1.465723e-09, 6.990357e-10, 8.971997e-11, 7.513724e-12,
  2.498081e-08, 2.3127e-08, 2.120547e-08, 1.844616e-08, 1.451446e-08, 
    1.102314e-08, 8.592765e-09, 6.297815e-09, 4.390106e-09, 3.293309e-09, 
    2.490857e-09, 1.637335e-09, 8.691692e-10, 1.294044e-10, -1.238659e-11,
  2.589588e-08, 2.409016e-08, 2.236907e-08, 2.025289e-08, 1.678893e-08, 
    1.270445e-08, 9.822358e-09, 7.258857e-09, 4.983248e-09, 3.630375e-09, 
    2.793968e-09, 1.832936e-09, 1.033041e-09, 1.875005e-10, 5.958674e-12,
  2.614021e-08, 2.537077e-08, 2.36578e-08, 2.181732e-08, 1.889328e-08, 
    1.470572e-08, 1.116368e-08, 8.531265e-09, 5.899636e-09, 4.079902e-09, 
    3.1075e-09, 2.090667e-09, 1.202795e-09, 2.617271e-10, 2.180683e-11,
  2.565233e-08, 2.561537e-08, 2.493133e-08, 2.313844e-08, 2.079863e-08, 
    1.698134e-08, 1.274171e-08, 9.662278e-09, 6.800132e-09, 4.568333e-09, 
    3.390803e-09, 2.377925e-09, 1.330543e-09, 3.546466e-10, 2.933032e-11,
  2.557744e-08, 2.612603e-08, 2.575793e-08, 2.434743e-08, 2.227982e-08, 
    1.888413e-08, 1.480432e-08, 1.132847e-08, 8.078361e-09, 5.213878e-09, 
    3.671409e-09, 2.643918e-09, 1.462068e-09, 4.595065e-10, 3.457461e-11,
  2.536239e-08, 2.600983e-08, 2.606891e-08, 2.504208e-08, 2.391117e-08, 
    2.089516e-08, 1.65405e-08, 1.273474e-08, 9.318291e-09, 5.991299e-09, 
    3.995913e-09, 2.898706e-09, 1.619283e-09, 5.689013e-10, 5.210176e-11,
  2.575875e-08, 2.565549e-08, 2.602336e-08, 2.569292e-08, 2.459458e-08, 
    2.228681e-08, 1.846583e-08, 1.433206e-08, 1.073091e-08, 6.93423e-09, 
    4.399716e-09, 3.190483e-09, 1.863421e-09, 6.603274e-10, 7.482701e-11,
  2.616069e-08, 2.561375e-08, 2.577966e-08, 2.590347e-08, 2.498783e-08, 
    2.348139e-08, 2.025743e-08, 1.604427e-08, 1.234228e-08, 8.236023e-09, 
    4.97523e-09, 3.545917e-09, 2.159468e-09, 7.461831e-10, 1.179768e-10,
  1.912205e-08, 1.594887e-08, 1.197241e-08, 8.401376e-09, 6.047833e-09, 
    4.334102e-09, 3.128402e-09, 2.679811e-09, 2.213366e-09, 1.799962e-09, 
    1.458104e-09, 8.908692e-10, 2.946109e-10, 1.39393e-10, 1.211738e-10,
  2.078528e-08, 1.762745e-08, 1.406003e-08, 1.002182e-08, 6.949449e-09, 
    5.022834e-09, 3.628732e-09, 2.819974e-09, 2.36191e-09, 1.939417e-09, 
    1.661793e-09, 1.201406e-09, 4.290806e-10, 1.619372e-10, 1.216225e-10,
  2.201579e-08, 1.96646e-08, 1.606871e-08, 1.186372e-08, 8.179581e-09, 
    5.774066e-09, 4.200977e-09, 3.143434e-09, 2.590075e-09, 2.147593e-09, 
    1.863125e-09, 1.475172e-09, 6.067015e-10, 1.992798e-10, 1.320038e-10,
  2.240428e-08, 2.14562e-08, 1.808832e-08, 1.398334e-08, 9.770389e-09, 
    6.834632e-09, 4.906586e-09, 3.562674e-09, 2.726904e-09, 2.31599e-09, 
    2.056976e-09, 1.692799e-09, 8.298953e-10, 2.386164e-10, 1.435767e-10,
  2.359998e-08, 2.266302e-08, 2.010167e-08, 1.617641e-08, 1.172599e-08, 
    7.978167e-09, 5.718188e-09, 4.22622e-09, 3.132291e-09, 2.592714e-09, 
    2.252043e-09, 1.869943e-09, 1.107958e-09, 2.945741e-10, 1.55251e-10,
  2.401364e-08, 2.308952e-08, 2.171225e-08, 1.829274e-08, 1.403757e-08, 
    9.621461e-09, 6.729208e-09, 4.62492e-09, 3.312813e-09, 2.774337e-09, 
    2.43072e-09, 2.039087e-09, 1.391653e-09, 3.719349e-10, 1.541786e-10,
  2.453951e-08, 2.334786e-08, 2.231873e-08, 2.050023e-08, 1.63124e-08, 
    1.144207e-08, 7.974478e-09, 5.44384e-09, 3.872056e-09, 3.089463e-09, 
    2.605655e-09, 2.207914e-09, 1.63143e-09, 4.900012e-10, 1.537039e-10,
  2.513915e-08, 2.432561e-08, 2.287984e-08, 2.173469e-08, 1.873003e-08, 
    1.379636e-08, 9.454915e-09, 6.607065e-09, 4.795418e-09, 3.550802e-09, 
    2.780016e-09, 2.37765e-09, 1.73439e-09, 6.570329e-10, 1.66266e-10,
  2.589232e-08, 2.523158e-08, 2.348375e-08, 2.225495e-08, 2.061791e-08, 
    1.635182e-08, 1.160422e-08, 7.996626e-09, 5.397455e-09, 3.74455e-09, 
    2.944364e-09, 2.546933e-09, 1.746376e-09, 8.871224e-10, 2.188802e-10,
  2.632213e-08, 2.584873e-08, 2.44199e-08, 2.276042e-08, 2.188194e-08, 
    1.881041e-08, 1.37904e-08, 9.417166e-09, 6.271546e-09, 4.167708e-09, 
    3.13195e-09, 2.661416e-09, 1.882256e-09, 1.141516e-09, 3.125023e-10,
  2.12914e-08, 1.861487e-08, 1.461888e-08, 1.005562e-08, 6.427801e-09, 
    4.349691e-09, 3.271701e-09, 2.759943e-09, 2.456564e-09, 1.981441e-09, 
    1.527611e-09, 1.104943e-09, 6.182184e-10, 3.98005e-10, 5.730555e-10,
  2.211753e-08, 1.995611e-08, 1.639214e-08, 1.163195e-08, 7.525725e-09, 
    4.91827e-09, 3.55476e-09, 2.89123e-09, 2.527292e-09, 2.006836e-09, 
    1.538168e-09, 1.188684e-09, 7.083302e-10, 4.337298e-10, 5.846539e-10,
  2.255611e-08, 2.121998e-08, 1.80034e-08, 1.327922e-08, 8.743957e-09, 
    5.546128e-09, 3.82714e-09, 3.015607e-09, 2.61457e-09, 2.074295e-09, 
    1.57649e-09, 1.297051e-09, 8.222224e-10, 4.623217e-10, 5.652961e-10,
  2.271228e-08, 2.187515e-08, 1.937021e-08, 1.503672e-08, 1.017271e-08, 
    6.420182e-09, 4.196361e-09, 3.135521e-09, 2.691763e-09, 2.175053e-09, 
    1.636604e-09, 1.365594e-09, 9.03604e-10, 4.754686e-10, 5.394747e-10,
  2.338335e-08, 2.250597e-08, 2.042438e-08, 1.665681e-08, 1.177289e-08, 
    7.380673e-09, 4.688738e-09, 3.374695e-09, 2.84446e-09, 2.308653e-09, 
    1.703487e-09, 1.41563e-09, 9.949244e-10, 4.914201e-10, 5.438609e-10,
  2.365674e-08, 2.277162e-08, 2.133015e-08, 1.808787e-08, 1.34023e-08, 
    8.678574e-09, 5.289324e-09, 3.496166e-09, 2.850217e-09, 2.372273e-09, 
    1.752812e-09, 1.477847e-09, 1.082074e-09, 5.217733e-10, 5.713183e-10,
  2.396488e-08, 2.315095e-08, 2.199658e-08, 1.945018e-08, 1.49451e-08, 
    9.880175e-09, 6.077063e-09, 3.770292e-09, 2.940978e-09, 2.475075e-09, 
    1.785688e-09, 1.467846e-09, 1.149243e-09, 5.510286e-10, 5.942457e-10,
  2.406123e-08, 2.360592e-08, 2.2481e-08, 2.052444e-08, 1.663321e-08, 
    1.136435e-08, 6.908523e-09, 4.290599e-09, 3.303015e-09, 2.739181e-09, 
    1.822194e-09, 1.45003e-09, 1.202431e-09, 5.783159e-10, 6.34025e-10,
  2.467706e-08, 2.408464e-08, 2.285633e-08, 2.123337e-08, 1.800896e-08, 
    1.309856e-08, 8.184957e-09, 4.945077e-09, 3.404607e-09, 2.745013e-09, 
    1.888711e-09, 1.459815e-09, 1.239979e-09, 5.824651e-10, 6.753116e-10,
  2.529638e-08, 2.448203e-08, 2.328164e-08, 2.184528e-08, 1.927107e-08, 
    1.479011e-08, 9.42668e-09, 5.499456e-09, 3.550187e-09, 2.86048e-09, 
    2.019298e-09, 1.457407e-09, 1.223931e-09, 5.513867e-10, 7.162738e-10,
  2.020531e-08, 1.90268e-08, 1.711423e-08, 1.442433e-08, 1.040763e-08, 
    6.63872e-09, 4.330819e-09, 2.936377e-09, 2.230741e-09, 1.96852e-09, 
    1.751081e-09, 1.414517e-09, 1.115403e-09, 9.141349e-10, 7.758568e-10,
  2.109485e-08, 1.974174e-08, 1.805145e-08, 1.555095e-08, 1.199682e-08, 
    7.747206e-09, 4.983776e-09, 3.253897e-09, 2.373399e-09, 2.065116e-09, 
    1.869055e-09, 1.50105e-09, 1.141906e-09, 9.133429e-10, 8.043098e-10,
  2.180306e-08, 2.04701e-08, 1.894026e-08, 1.659295e-08, 1.341236e-08, 
    9.025626e-09, 5.760542e-09, 3.670407e-09, 2.576945e-09, 2.188447e-09, 
    1.972806e-09, 1.56348e-09, 1.136033e-09, 8.912763e-10, 8.278995e-10,
  2.220003e-08, 2.094824e-08, 1.955755e-08, 1.768016e-08, 1.470457e-08, 
    1.048534e-08, 6.66329e-09, 4.141472e-09, 2.79649e-09, 2.297857e-09, 
    2.034789e-09, 1.565578e-09, 1.103699e-09, 8.794263e-10, 8.478978e-10,
  2.29879e-08, 2.187425e-08, 2.023818e-08, 1.852366e-08, 1.584429e-08, 
    1.193858e-08, 7.761845e-09, 4.854914e-09, 3.128051e-09, 2.434484e-09, 
    2.081058e-09, 1.549249e-09, 1.082348e-09, 9.123924e-10, 8.92011e-10,
  2.332774e-08, 2.229051e-08, 2.102159e-08, 1.940174e-08, 1.696676e-08, 
    1.338101e-08, 8.923407e-09, 5.51917e-09, 3.432365e-09, 2.541829e-09, 
    2.08983e-09, 1.52761e-09, 1.091049e-09, 9.704725e-10, 9.528105e-10,
  2.331406e-08, 2.298213e-08, 2.175486e-08, 2.013972e-08, 1.787311e-08, 
    1.457827e-08, 1.03716e-08, 6.433949e-09, 3.848546e-09, 2.685589e-09, 
    2.10368e-09, 1.520424e-09, 1.130759e-09, 1.050915e-09, 1.024847e-09,
  2.314562e-08, 2.365692e-08, 2.257359e-08, 2.103919e-08, 1.904403e-08, 
    1.573079e-08, 1.159423e-08, 7.442951e-09, 4.603411e-09, 2.933704e-09, 
    2.131732e-09, 1.541309e-09, 1.192843e-09, 1.123701e-09, 1.08648e-09,
  2.300245e-08, 2.361388e-08, 2.303821e-08, 2.176921e-08, 1.987912e-08, 
    1.683864e-08, 1.293614e-08, 8.574437e-09, 5.137911e-09, 3.028999e-09, 
    2.192444e-09, 1.596589e-09, 1.248028e-09, 1.170977e-09, 1.124685e-09,
  2.314494e-08, 2.3527e-08, 2.358521e-08, 2.242366e-08, 2.083423e-08, 
    1.783093e-08, 1.399676e-08, 9.539611e-09, 5.790216e-09, 3.34342e-09, 
    2.355784e-09, 1.682392e-09, 1.29238e-09, 1.182623e-09, 1.146795e-09,
  1.883678e-08, 1.751097e-08, 1.6727e-08, 1.579649e-08, 1.342319e-08, 
    1.001465e-08, 6.696355e-09, 3.795444e-09, 2.306991e-09, 1.79129e-09, 
    1.716986e-09, 1.60603e-09, 1.396293e-09, 1.351081e-09, 1.265861e-09,
  1.997419e-08, 1.841239e-08, 1.718116e-08, 1.635281e-08, 1.470905e-08, 
    1.162706e-08, 8.218084e-09, 4.909448e-09, 2.763103e-09, 1.964271e-09, 
    1.805576e-09, 1.729793e-09, 1.438814e-09, 1.310917e-09, 1.236334e-09,
  2.125381e-08, 1.93998e-08, 1.785946e-08, 1.68217e-08, 1.568124e-08, 
    1.310669e-08, 9.722098e-09, 6.267163e-09, 3.501103e-09, 2.286709e-09, 
    1.895717e-09, 1.750458e-09, 1.413277e-09, 1.195794e-09, 1.289757e-09,
  2.188943e-08, 2.044993e-08, 1.866352e-08, 1.722384e-08, 1.639233e-08, 
    1.444995e-08, 1.122958e-08, 7.702785e-09, 4.392023e-09, 2.663896e-09, 
    1.972844e-09, 1.685094e-09, 1.347242e-09, 1.198477e-09, 1.466888e-09,
  2.218815e-08, 2.161429e-08, 1.983658e-08, 1.786888e-08, 1.690579e-08, 
    1.54542e-08, 1.265675e-08, 9.214182e-09, 5.693355e-09, 3.199323e-09, 
    2.114841e-09, 1.639962e-09, 1.396543e-09, 1.397266e-09, 1.668445e-09,
  2.128012e-08, 2.153333e-08, 2.08186e-08, 1.873002e-08, 1.738446e-08, 
    1.639126e-08, 1.400851e-08, 1.044959e-08, 6.935637e-09, 3.904053e-09, 
    2.330004e-09, 1.674298e-09, 1.507626e-09, 1.604114e-09, 1.813054e-09,
  2.097274e-08, 2.139426e-08, 2.131266e-08, 1.981648e-08, 1.791873e-08, 
    1.686093e-08, 1.528709e-08, 1.202539e-08, 8.257719e-09, 4.796072e-09, 
    2.641774e-09, 1.752786e-09, 1.618753e-09, 1.774304e-09, 1.875238e-09,
  2.112759e-08, 2.1212e-08, 2.156154e-08, 2.064545e-08, 1.894181e-08, 
    1.7477e-08, 1.620629e-08, 1.337659e-08, 9.692467e-09, 5.980428e-09, 
    3.117609e-09, 1.930243e-09, 1.768883e-09, 1.917129e-09, 1.915966e-09,
  2.162704e-08, 2.118127e-08, 2.135776e-08, 2.129606e-08, 1.967495e-08, 
    1.805241e-08, 1.688762e-08, 1.474422e-08, 1.101531e-08, 7.150944e-09, 
    3.836617e-09, 2.217131e-09, 1.936892e-09, 2.04016e-09, 1.954469e-09,
  2.206968e-08, 2.143454e-08, 2.111735e-08, 2.154602e-08, 2.058147e-08, 
    1.888673e-08, 1.750491e-08, 1.546198e-08, 1.209053e-08, 8.399407e-09, 
    4.79819e-09, 2.607164e-09, 2.110903e-09, 2.115031e-09, 1.991976e-09,
  2.057278e-08, 1.834224e-08, 1.538179e-08, 1.203598e-08, 7.413977e-09, 
    3.747156e-09, 2.092782e-09, 1.859501e-09, 1.553855e-09, 1.216256e-09, 
    7.966857e-10, 6.530283e-10, 7.58362e-10, 1.08301e-09, 1.235069e-09,
  2.165474e-08, 1.995145e-08, 1.742309e-08, 1.413191e-08, 1.013195e-08, 
    5.779206e-09, 2.852261e-09, 1.914859e-09, 1.730913e-09, 1.358461e-09, 
    9.751102e-10, 7.237994e-10, 7.930769e-10, 1.08051e-09, 1.282863e-09,
  2.19791e-08, 2.089111e-08, 1.910102e-08, 1.620591e-08, 1.26268e-08, 
    8.062125e-09, 4.147025e-09, 2.139879e-09, 1.806111e-09, 1.535602e-09, 
    1.184223e-09, 8.479598e-10, 8.272493e-10, 1.025192e-09, 1.259293e-09,
  2.271475e-08, 2.116187e-08, 2.023629e-08, 1.802727e-08, 1.490536e-08, 
    1.052861e-08, 6.200371e-09, 2.941314e-09, 1.843305e-09, 1.633431e-09, 
    1.391379e-09, 9.875801e-10, 8.660901e-10, 9.63766e-10, 1.223219e-09,
  2.256898e-08, 2.195019e-08, 2.116092e-08, 1.951876e-08, 1.702166e-08, 
    1.300248e-08, 8.404046e-09, 4.501663e-09, 2.313295e-09, 1.752879e-09, 
    1.521085e-09, 1.166277e-09, 9.180504e-10, 9.23301e-10, 1.159807e-09,
  2.191845e-08, 2.183179e-08, 2.158202e-08, 2.060392e-08, 1.872626e-08, 
    1.553085e-08, 1.080454e-08, 6.34158e-09, 3.03702e-09, 1.803947e-09, 
    1.608998e-09, 1.27209e-09, 9.744887e-10, 9.141833e-10, 1.110416e-09,
  2.191368e-08, 2.22768e-08, 2.196428e-08, 2.139691e-08, 2.00417e-08, 
    1.772367e-08, 1.322076e-08, 8.722744e-09, 4.747457e-09, 2.307691e-09, 
    1.709245e-09, 1.398072e-09, 1.007426e-09, 9.281626e-10, 1.076753e-09,
  2.199647e-08, 2.218862e-08, 2.220334e-08, 2.170326e-08, 2.110994e-08, 
    1.948086e-08, 1.544502e-08, 1.064108e-08, 6.744916e-09, 3.381906e-09, 
    1.919282e-09, 1.53685e-09, 1.08634e-09, 9.531008e-10, 1.066695e-09,
  2.231294e-08, 2.208282e-08, 2.221724e-08, 2.229107e-08, 2.177867e-08, 
    2.050207e-08, 1.806156e-08, 1.281348e-08, 8.446952e-09, 4.628788e-09, 
    2.36971e-09, 1.718564e-09, 1.199333e-09, 9.770028e-10, 1.023499e-09,
  2.312201e-08, 2.207579e-08, 2.222662e-08, 2.232387e-08, 2.236674e-08, 
    2.131075e-08, 1.993577e-08, 1.510901e-08, 1.033574e-08, 6.353946e-09, 
    3.217843e-09, 1.97517e-09, 1.322979e-09, 1.000526e-09, 9.501572e-10,
  1.834763e-08, 1.445435e-08, 1.095507e-08, 8.49619e-09, 6.405906e-09, 
    4.781954e-09, 3.630855e-09, 2.627328e-09, 1.832307e-09, 1.210424e-09, 
    9.184619e-10, 8.239563e-10, 7.146326e-10, 7.1645e-10, 7.541984e-10,
  1.940646e-08, 1.609804e-08, 1.209798e-08, 9.268128e-09, 7.027641e-09, 
    5.236691e-09, 3.937481e-09, 2.859174e-09, 1.978843e-09, 1.280632e-09, 
    8.991012e-10, 7.797355e-10, 6.95931e-10, 7.057419e-10, 7.60427e-10,
  2.046579e-08, 1.750501e-08, 1.356529e-08, 1.015047e-08, 7.68882e-09, 
    5.735652e-09, 4.272332e-09, 3.098391e-09, 2.170183e-09, 1.407951e-09, 
    9.545016e-10, 7.899096e-10, 6.923719e-10, 6.914055e-10, 7.605111e-10,
  2.150414e-08, 1.882605e-08, 1.490097e-08, 1.124362e-08, 8.421114e-09, 
    6.339387e-09, 4.697478e-09, 3.350408e-09, 2.348704e-09, 1.56037e-09, 
    1.040128e-09, 8.066491e-10, 6.818697e-10, 6.602529e-10, 7.31527e-10,
  2.199025e-08, 2.015877e-08, 1.642603e-08, 1.253797e-08, 9.30117e-09, 
    6.927622e-09, 5.143682e-09, 3.677836e-09, 2.601298e-09, 1.730215e-09, 
    1.130193e-09, 8.426844e-10, 6.637022e-10, 6.32036e-10, 6.858445e-10,
  2.175918e-08, 2.071268e-08, 1.77716e-08, 1.392427e-08, 1.044857e-08, 
    7.825224e-09, 5.769282e-09, 4.033745e-09, 2.804305e-09, 1.879753e-09, 
    1.201622e-09, 8.397279e-10, 6.273301e-10, 5.989531e-10, 6.427082e-10,
  2.176635e-08, 2.142933e-08, 1.928928e-08, 1.557038e-08, 1.172218e-08, 
    8.638023e-09, 6.513331e-09, 4.668544e-09, 3.236421e-09, 2.130444e-09, 
    1.332394e-09, 8.924583e-10, 6.095008e-10, 5.572261e-10, 5.93956e-10,
  2.182231e-08, 2.157595e-08, 2.042222e-08, 1.710419e-08, 1.341451e-08, 
    9.847665e-09, 7.171892e-09, 5.155689e-09, 3.626646e-09, 2.448416e-09, 
    1.564252e-09, 1.061609e-09, 6.953634e-10, 5.431329e-10, 5.510981e-10,
  2.269793e-08, 2.191774e-08, 2.113434e-08, 1.869009e-08, 1.4964e-08, 
    1.140682e-08, 8.309632e-09, 5.830935e-09, 3.896457e-09, 2.591219e-09, 
    1.760218e-09, 1.251392e-09, 8.589281e-10, 6.01982e-10, 5.295374e-10,
  2.317101e-08, 2.23953e-08, 2.152344e-08, 1.998162e-08, 1.641934e-08, 
    1.303142e-08, 9.703122e-09, 6.837737e-09, 4.540845e-09, 2.894313e-09, 
    1.906567e-09, 1.407581e-09, 1.024883e-09, 6.724324e-10, 5.24925e-10,
  2.224292e-08, 1.960255e-08, 1.811159e-08, 1.563193e-08, 1.275535e-08, 
    9.953756e-09, 7.867402e-09, 6.117825e-09, 4.647685e-09, 3.269885e-09, 
    2.526545e-09, 2.184271e-09, 1.818273e-09, 1.614811e-09, 1.508754e-09,
  2.187125e-08, 1.995397e-08, 1.835473e-08, 1.591593e-08, 1.295724e-08, 
    1.017781e-08, 8.048186e-09, 6.233482e-09, 4.654741e-09, 3.270937e-09, 
    2.491451e-09, 2.212369e-09, 1.941812e-09, 1.70188e-09, 1.493689e-09,
  2.200495e-08, 2.049846e-08, 1.869335e-08, 1.622427e-08, 1.318464e-08, 
    1.033188e-08, 8.093833e-09, 6.322491e-09, 4.659995e-09, 3.324771e-09, 
    2.525319e-09, 2.226252e-09, 2.015754e-09, 1.774575e-09, 1.503565e-09,
  2.232033e-08, 2.127582e-08, 1.919076e-08, 1.646376e-08, 1.349617e-08, 
    1.057922e-08, 8.164051e-09, 6.368563e-09, 4.654209e-09, 3.465502e-09, 
    2.653123e-09, 2.253084e-09, 2.06067e-09, 1.82911e-09, 1.491916e-09,
  2.311437e-08, 2.173524e-08, 1.961841e-08, 1.689143e-08, 1.380179e-08, 
    1.075115e-08, 8.204068e-09, 6.462593e-09, 4.819389e-09, 3.710936e-09, 
    2.874788e-09, 2.313615e-09, 2.071747e-09, 1.869955e-09, 1.507011e-09,
  2.349136e-08, 2.211442e-08, 2.01979e-08, 1.733822e-08, 1.421695e-08, 
    1.109225e-08, 8.325712e-09, 6.334652e-09, 4.831298e-09, 3.923641e-09, 
    3.070444e-09, 2.366815e-09, 2.062262e-09, 1.879781e-09, 1.485319e-09,
  2.329448e-08, 2.219177e-08, 2.036842e-08, 1.789858e-08, 1.44493e-08, 
    1.115599e-08, 8.300952e-09, 6.359478e-09, 5.217553e-09, 4.281269e-09, 
    3.270781e-09, 2.384062e-09, 2.000295e-09, 1.840976e-09, 1.447153e-09,
  2.360849e-08, 2.26841e-08, 2.090626e-08, 1.853504e-08, 1.482408e-08, 
    1.145722e-08, 8.659941e-09, 6.732104e-09, 5.755534e-09, 4.65023e-09, 
    3.442308e-09, 2.462881e-09, 1.97363e-09, 1.789664e-09, 1.392147e-09,
  2.345871e-08, 2.309013e-08, 2.144848e-08, 1.891093e-08, 1.540828e-08, 
    1.234235e-08, 9.417109e-09, 7.02468e-09, 5.601024e-09, 4.611428e-09, 
    3.570259e-09, 2.577979e-09, 2.008472e-09, 1.758748e-09, 1.329406e-09,
  2.347336e-08, 2.323192e-08, 2.194684e-08, 1.954078e-08, 1.628086e-08, 
    1.297902e-08, 9.84461e-09, 7.073981e-09, 5.342494e-09, 4.540424e-09, 
    3.665036e-09, 2.732495e-09, 2.126178e-09, 1.785802e-09, 1.300256e-09,
  2.487683e-08, 2.484312e-08, 2.498072e-08, 2.405084e-08, 2.245504e-08, 
    1.985936e-08, 1.714316e-08, 1.475237e-08, 1.202095e-08, 9.085145e-09, 
    6.227201e-09, 4.351669e-09, 3.557239e-09, 3.007858e-09, 2.549696e-09,
  2.540276e-08, 2.52822e-08, 2.509346e-08, 2.399548e-08, 2.234548e-08, 
    1.97043e-08, 1.69008e-08, 1.446809e-08, 1.172814e-08, 8.694678e-09, 
    5.876029e-09, 4.202272e-09, 3.50677e-09, 2.922465e-09, 2.447384e-09,
  2.557405e-08, 2.537709e-08, 2.517285e-08, 2.408076e-08, 2.231868e-08, 
    1.957243e-08, 1.676493e-08, 1.419712e-08, 1.12879e-08, 8.153847e-09, 
    5.423857e-09, 3.954124e-09, 3.3332e-09, 2.754302e-09, 2.315683e-09,
  2.577579e-08, 2.576792e-08, 2.539977e-08, 2.414626e-08, 2.235971e-08, 
    1.949005e-08, 1.652711e-08, 1.383055e-08, 1.08562e-08, 7.663541e-09, 
    5.084484e-09, 3.805086e-09, 3.215941e-09, 2.635286e-09, 2.223035e-09,
  2.574061e-08, 2.567109e-08, 2.542816e-08, 2.427128e-08, 2.234439e-08, 
    1.93546e-08, 1.642029e-08, 1.360114e-08, 1.049966e-08, 7.263482e-09, 
    4.827946e-09, 3.684191e-09, 3.090662e-09, 2.521545e-09, 2.147303e-09,
  2.561716e-08, 2.548771e-08, 2.526723e-08, 2.42951e-08, 2.247344e-08, 
    1.920351e-08, 1.608075e-08, 1.308998e-08, 1.001778e-08, 6.826621e-09, 
    4.560054e-09, 3.54716e-09, 2.941367e-09, 2.406054e-09, 2.10818e-09,
  2.514198e-08, 2.524152e-08, 2.507097e-08, 2.426155e-08, 2.219499e-08, 
    1.894445e-08, 1.579268e-08, 1.271003e-08, 9.589041e-09, 6.457598e-09, 
    4.327183e-09, 3.421726e-09, 2.796041e-09, 2.301612e-09, 2.068304e-09,
  2.512965e-08, 2.526927e-08, 2.511524e-08, 2.424619e-08, 2.199987e-08, 
    1.857401e-08, 1.566006e-08, 1.258673e-08, 9.412114e-09, 6.132275e-09, 
    4.097675e-09, 3.260011e-09, 2.608515e-09, 2.211467e-09, 1.966948e-09,
  2.49593e-08, 2.534909e-08, 2.52196e-08, 2.405118e-08, 2.175205e-08, 
    1.858598e-08, 1.562078e-08, 1.227337e-08, 8.831343e-09, 5.58473e-09, 
    3.912636e-09, 3.116638e-09, 2.440586e-09, 2.137553e-09, 1.823341e-09,
  2.488732e-08, 2.546187e-08, 2.530858e-08, 2.400378e-08, 2.187806e-08, 
    1.850944e-08, 1.524317e-08, 1.171161e-08, 8.152826e-09, 5.24689e-09, 
    3.823831e-09, 2.990747e-09, 2.310915e-09, 2.088439e-09, 1.675046e-09,
  2.495205e-08, 2.494339e-08, 2.512559e-08, 2.522269e-08, 2.418195e-08, 
    2.280044e-08, 2.085083e-08, 1.781245e-08, 1.463086e-08, 1.188379e-08, 
    9.535902e-09, 7.222699e-09, 5.606842e-09, 4.198195e-09, 2.94607e-09,
  2.554786e-08, 2.542066e-08, 2.487933e-08, 2.478231e-08, 2.420983e-08, 
    2.296248e-08, 2.127904e-08, 1.840174e-08, 1.499604e-08, 1.211072e-08, 
    9.651994e-09, 7.298431e-09, 5.681396e-09, 4.218421e-09, 2.933962e-09,
  2.52776e-08, 2.579166e-08, 2.520582e-08, 2.47647e-08, 2.434103e-08, 
    2.323854e-08, 2.172629e-08, 1.896334e-08, 1.536063e-08, 1.226496e-08, 
    9.696996e-09, 7.308183e-09, 5.688913e-09, 4.106938e-09, 2.794435e-09,
  2.498765e-08, 2.551441e-08, 2.529693e-08, 2.500526e-08, 2.460784e-08, 
    2.362601e-08, 2.195341e-08, 1.935653e-08, 1.56084e-08, 1.239103e-08, 
    9.71791e-09, 7.296129e-09, 5.641534e-09, 3.919904e-09, 2.664362e-09,
  2.478514e-08, 2.536456e-08, 2.526904e-08, 2.509968e-08, 2.47969e-08, 
    2.38467e-08, 2.223201e-08, 1.996578e-08, 1.604123e-08, 1.245742e-08, 
    9.65979e-09, 7.223143e-09, 5.533185e-09, 3.694476e-09, 2.552754e-09,
  2.430424e-08, 2.508517e-08, 2.529356e-08, 2.511146e-08, 2.489129e-08, 
    2.416871e-08, 2.222762e-08, 1.998531e-08, 1.613205e-08, 1.249187e-08, 
    9.521378e-09, 7.111813e-09, 5.365041e-09, 3.495221e-09, 2.510641e-09,
  2.429198e-08, 2.477324e-08, 2.511277e-08, 2.536203e-08, 2.487187e-08, 
    2.424032e-08, 2.265326e-08, 2.034136e-08, 1.649117e-08, 1.241244e-08, 
    9.333472e-09, 6.950652e-09, 5.152083e-09, 3.342985e-09, 2.523202e-09,
  2.412483e-08, 2.450787e-08, 2.516871e-08, 2.534165e-08, 2.487943e-08, 
    2.4193e-08, 2.27141e-08, 2.051655e-08, 1.661111e-08, 1.238691e-08, 
    9.149902e-09, 6.803284e-09, 4.909107e-09, 3.236593e-09, 2.59225e-09,
  2.426357e-08, 2.461637e-08, 2.500587e-08, 2.505812e-08, 2.476581e-08, 
    2.448684e-08, 2.317023e-08, 2.049669e-08, 1.649604e-08, 1.212408e-08, 
    8.917847e-09, 6.597263e-09, 4.681305e-09, 3.17243e-09, 2.652847e-09,
  2.435996e-08, 2.468599e-08, 2.486504e-08, 2.473035e-08, 2.467803e-08, 
    2.446773e-08, 2.318031e-08, 2.04678e-08, 1.621784e-08, 1.17973e-08, 
    8.664707e-09, 6.331526e-09, 4.473755e-09, 3.128856e-09, 2.677705e-09,
  2.47522e-08, 2.482837e-08, 2.41272e-08, 2.238158e-08, 2.074273e-08, 
    1.887635e-08, 1.388308e-08, 1.026551e-08, 8.267572e-09, 6.787907e-09, 
    5.248551e-09, 3.656514e-09, 2.557206e-09, 2.065203e-09, 1.874325e-09,
  2.466325e-08, 2.493569e-08, 2.477882e-08, 2.317969e-08, 2.163374e-08, 
    1.986048e-08, 1.433958e-08, 1.028237e-08, 8.381214e-09, 6.923178e-09, 
    5.291714e-09, 3.696207e-09, 2.593198e-09, 2.084473e-09, 1.899473e-09,
  2.499534e-08, 2.562365e-08, 2.53215e-08, 2.394541e-08, 2.256467e-08, 
    2.099282e-08, 1.493076e-08, 1.033993e-08, 8.417485e-09, 7.004312e-09, 
    5.327495e-09, 3.705931e-09, 2.593697e-09, 2.066253e-09, 1.896818e-09,
  2.478738e-08, 2.57735e-08, 2.572415e-08, 2.494147e-08, 2.354076e-08, 
    2.240543e-08, 1.554631e-08, 1.040799e-08, 8.488238e-09, 7.103294e-09, 
    5.386499e-09, 3.709618e-09, 2.589734e-09, 2.054079e-09, 1.911024e-09,
  2.688362e-08, 2.579349e-08, 2.524541e-08, 2.549101e-08, 2.456806e-08, 
    2.359366e-08, 1.628576e-08, 1.063476e-08, 8.611187e-09, 7.191214e-09, 
    5.416715e-09, 3.698207e-09, 2.581664e-09, 2.054851e-09, 1.931815e-09,
  2.704605e-08, 2.55433e-08, 2.46645e-08, 2.518278e-08, 2.551499e-08, 
    2.50958e-08, 1.691755e-08, 1.087408e-08, 8.732652e-09, 7.282837e-09, 
    5.447308e-09, 3.695748e-09, 2.578013e-09, 2.061336e-09, 1.94065e-09,
  2.621573e-08, 2.53484e-08, 2.424254e-08, 2.538462e-08, 2.607896e-08, 
    2.622271e-08, 1.81108e-08, 1.130529e-08, 8.796942e-09, 7.305378e-09, 
    5.457431e-09, 3.683855e-09, 2.569271e-09, 2.068914e-09, 1.9523e-09,
  2.600224e-08, 2.640137e-08, 2.535553e-08, 2.558004e-08, 2.717329e-08, 
    2.739146e-08, 1.88459e-08, 1.182197e-08, 8.818184e-09, 7.295905e-09, 
    5.474215e-09, 3.677328e-09, 2.560319e-09, 2.07926e-09, 1.971756e-09,
  2.636903e-08, 2.7129e-08, 2.601328e-08, 2.544747e-08, 2.656466e-08, 
    2.833084e-08, 1.964204e-08, 1.242355e-08, 9.13897e-09, 7.396975e-09, 
    5.476402e-09, 3.656675e-09, 2.556279e-09, 2.097416e-09, 2.004903e-09,
  2.641337e-08, 2.702209e-08, 2.597393e-08, 2.556946e-08, 2.552466e-08, 
    2.831723e-08, 2.056452e-08, 1.294093e-08, 9.349082e-09, 7.431732e-09, 
    5.468107e-09, 3.640896e-09, 2.550784e-09, 2.127969e-09, 2.055933e-09,
  2.280213e-08, 2.436978e-08, 2.559421e-08, 2.511562e-08, 2.341293e-08, 
    1.920377e-08, 1.452571e-08, 1.113624e-08, 8.771605e-09, 6.939335e-09, 
    5.818441e-09, 4.480807e-09, 3.299245e-09, 2.354914e-09, 1.570133e-09,
  2.285445e-08, 2.417712e-08, 2.528459e-08, 2.520588e-08, 2.317498e-08, 
    1.965746e-08, 1.472757e-08, 1.092629e-08, 8.609703e-09, 6.852495e-09, 
    5.66961e-09, 4.311411e-09, 3.148129e-09, 2.209231e-09, 1.497521e-09,
  2.296301e-08, 2.389779e-08, 2.506402e-08, 2.475514e-08, 2.288971e-08, 
    1.991622e-08, 1.496059e-08, 1.088921e-08, 8.532017e-09, 6.765137e-09, 
    5.491019e-09, 4.076093e-09, 2.951299e-09, 2.051091e-09, 1.400594e-09,
  2.318907e-08, 2.410593e-08, 2.489246e-08, 2.426766e-08, 2.27114e-08, 
    1.981211e-08, 1.504769e-08, 1.074032e-08, 8.348955e-09, 6.658983e-09, 
    5.309731e-09, 3.858118e-09, 2.774491e-09, 1.905026e-09, 1.304462e-09,
  2.369049e-08, 2.430601e-08, 2.476093e-08, 2.429612e-08, 2.242551e-08, 
    1.962157e-08, 1.499441e-08, 1.059408e-08, 8.218707e-09, 6.511173e-09, 
    5.116882e-09, 3.656946e-09, 2.607379e-09, 1.767602e-09, 1.208566e-09,
  2.449637e-08, 2.446815e-08, 2.487865e-08, 2.424294e-08, 2.241049e-08, 
    1.944041e-08, 1.467357e-08, 1.029202e-08, 8.062479e-09, 6.404037e-09, 
    4.924009e-09, 3.466284e-09, 2.448327e-09, 1.638702e-09, 1.118257e-09,
  2.431663e-08, 2.426732e-08, 2.468715e-08, 2.424973e-08, 2.230307e-08, 
    1.937212e-08, 1.461972e-08, 1.011133e-08, 7.875457e-09, 6.241315e-09, 
    4.739647e-09, 3.276934e-09, 2.290471e-09, 1.518665e-09, 1.035326e-09,
  2.403045e-08, 2.404476e-08, 2.465994e-08, 2.424376e-08, 2.266931e-08, 
    1.93403e-08, 1.443371e-08, 9.819711e-09, 7.565314e-09, 6.034711e-09, 
    4.525928e-09, 3.09563e-09, 2.139149e-09, 1.407653e-09, 9.621365e-10,
  2.422199e-08, 2.418387e-08, 2.449463e-08, 2.367333e-08, 2.235314e-08, 
    1.953992e-08, 1.432332e-08, 9.725584e-09, 7.515367e-09, 5.877459e-09, 
    4.304241e-09, 2.93201e-09, 1.997736e-09, 1.302581e-09, 9.013329e-10,
  2.434291e-08, 2.408197e-08, 2.424587e-08, 2.354287e-08, 2.28323e-08, 
    1.976215e-08, 1.402417e-08, 9.481887e-09, 7.317956e-09, 5.677779e-09, 
    4.10668e-09, 2.787607e-09, 1.865142e-09, 1.202647e-09, 8.525115e-10,
  2.496491e-08, 2.653528e-08, 2.505048e-08, 2.057403e-08, 1.638548e-08, 
    1.296708e-08, 1.143076e-08, 1.037506e-08, 8.691939e-09, 7.213458e-09, 
    6.310703e-09, 5.402886e-09, 4.544568e-09, 3.856026e-09, 3.303885e-09,
  2.403061e-08, 2.614e-08, 2.717806e-08, 2.365865e-08, 1.867049e-08, 
    1.462286e-08, 1.210541e-08, 1.086969e-08, 9.063915e-09, 7.446145e-09, 
    6.42921e-09, 5.492022e-09, 4.614557e-09, 3.895507e-09, 3.322889e-09,
  2.302641e-08, 2.478873e-08, 2.731862e-08, 2.656368e-08, 2.179912e-08, 
    1.644943e-08, 1.307249e-08, 1.149306e-08, 9.56293e-09, 7.698001e-09, 
    6.538562e-09, 5.563884e-09, 4.645254e-09, 3.901971e-09, 3.312609e-09,
  2.259045e-08, 2.313921e-08, 2.549801e-08, 2.784993e-08, 2.495102e-08, 
    1.918049e-08, 1.435668e-08, 1.201072e-08, 9.915906e-09, 7.982612e-09, 
    6.668434e-09, 5.61357e-09, 4.659165e-09, 3.89195e-09, 3.280197e-09,
  2.279745e-08, 2.268726e-08, 2.378598e-08, 2.719703e-08, 2.691273e-08, 
    2.221423e-08, 1.614827e-08, 1.292516e-08, 1.036396e-08, 8.271352e-09, 
    6.806207e-09, 5.66305e-09, 4.659032e-09, 3.865416e-09, 3.232859e-09,
  2.245434e-08, 2.239186e-08, 2.257745e-08, 2.524324e-08, 2.740177e-08, 
    2.499974e-08, 1.829252e-08, 1.364264e-08, 1.06804e-08, 8.546526e-09, 
    6.96132e-09, 5.690901e-09, 4.649855e-09, 3.839764e-09, 3.191117e-09,
  2.273575e-08, 2.252746e-08, 2.20966e-08, 2.375564e-08, 2.639151e-08, 
    2.593035e-08, 2.152672e-08, 1.523503e-08, 1.118579e-08, 8.760952e-09, 
    7.08206e-09, 5.717189e-09, 4.637702e-09, 3.811816e-09, 3.142385e-09,
  2.248892e-08, 2.233298e-08, 2.166827e-08, 2.248555e-08, 2.548088e-08, 
    2.633602e-08, 2.287501e-08, 1.650886e-08, 1.146236e-08, 8.871536e-09, 
    7.179201e-09, 5.734045e-09, 4.632344e-09, 3.788119e-09, 3.089083e-09,
  2.231508e-08, 2.206269e-08, 2.154336e-08, 2.199961e-08, 2.452065e-08, 
    2.576475e-08, 2.395962e-08, 1.773126e-08, 1.202254e-08, 9.056356e-09, 
    7.264334e-09, 5.758737e-09, 4.63656e-09, 3.754756e-09, 3.022774e-09,
  2.27078e-08, 2.221653e-08, 2.158772e-08, 2.178331e-08, 2.362065e-08, 
    2.523432e-08, 2.465448e-08, 1.937838e-08, 1.268539e-08, 9.170297e-09, 
    7.313406e-09, 5.781547e-09, 4.628661e-09, 3.706066e-09, 2.938633e-09,
  1.347016e-08, 1.324567e-08, 1.359958e-08, 1.424377e-08, 1.377809e-08, 
    1.287465e-08, 1.154136e-08, 1.009484e-08, 9.383479e-09, 8.707511e-09, 
    7.685466e-09, 6.438408e-09, 5.351009e-09, 4.320738e-09, 3.38693e-09,
  1.394912e-08, 1.332016e-08, 1.332848e-08, 1.420537e-08, 1.419202e-08, 
    1.27651e-08, 1.144229e-08, 1.006462e-08, 9.307756e-09, 8.668774e-09, 
    7.726248e-09, 6.464138e-09, 5.341035e-09, 4.323519e-09, 3.412929e-09,
  1.470226e-08, 1.372925e-08, 1.307334e-08, 1.418374e-08, 1.463516e-08, 
    1.303109e-08, 1.132023e-08, 1.007698e-08, 9.2252e-09, 8.603501e-09, 
    7.724711e-09, 6.492397e-09, 5.339456e-09, 4.334014e-09, 3.412674e-09,
  1.527712e-08, 1.422786e-08, 1.329933e-08, 1.396384e-08, 1.528909e-08, 
    1.37355e-08, 1.152562e-08, 1.021144e-08, 9.130672e-09, 8.513706e-09, 
    7.717061e-09, 6.533909e-09, 5.351701e-09, 4.317607e-09, 3.41841e-09,
  1.594257e-08, 1.526849e-08, 1.408358e-08, 1.381732e-08, 1.552236e-08, 
    1.476079e-08, 1.192694e-08, 1.041355e-08, 9.16174e-09, 8.461753e-09, 
    7.696594e-09, 6.560017e-09, 5.377554e-09, 4.297223e-09, 3.409147e-09,
  1.631619e-08, 1.626681e-08, 1.524542e-08, 1.423188e-08, 1.544188e-08, 
    1.584687e-08, 1.290644e-08, 1.059115e-08, 9.256646e-09, 8.442997e-09, 
    7.682734e-09, 6.563317e-09, 5.416199e-09, 4.280049e-09, 3.399746e-09,
  1.670683e-08, 1.697025e-08, 1.596839e-08, 1.456886e-08, 1.497158e-08, 
    1.634984e-08, 1.402799e-08, 1.12033e-08, 9.459918e-09, 8.46487e-09, 
    7.694909e-09, 6.576726e-09, 5.44516e-09, 4.281204e-09, 3.380466e-09,
  1.77828e-08, 1.712614e-08, 1.652168e-08, 1.521619e-08, 1.503738e-08, 
    1.655268e-08, 1.467865e-08, 1.150785e-08, 9.438044e-09, 8.372941e-09, 
    7.7027e-09, 6.622879e-09, 5.473698e-09, 4.298766e-09, 3.36589e-09,
  1.871998e-08, 1.770757e-08, 1.701343e-08, 1.652072e-08, 1.564511e-08, 
    1.597239e-08, 1.486243e-08, 1.178746e-08, 9.736588e-09, 8.602991e-09, 
    7.796237e-09, 6.68794e-09, 5.529185e-09, 4.34509e-09, 3.364603e-09,
  2.009341e-08, 1.861753e-08, 1.794183e-08, 1.759011e-08, 1.653977e-08, 
    1.606565e-08, 1.565475e-08, 1.299975e-08, 1.026343e-08, 8.768465e-09, 
    7.82028e-09, 6.767343e-09, 5.6064e-09, 4.406218e-09, 3.380838e-09,
  1.611129e-08, 1.542586e-08, 1.51785e-08, 1.37676e-08, 1.362363e-08, 
    1.264896e-08, 1.162036e-08, 1.062405e-08, 9.812711e-09, 8.712726e-09, 
    7.260569e-09, 5.81671e-09, 4.705742e-09, 3.495953e-09, 2.693855e-09,
  1.592415e-08, 1.553228e-08, 1.48419e-08, 1.428555e-08, 1.445904e-08, 
    1.356416e-08, 1.221614e-08, 1.107266e-08, 1.023497e-08, 9.280521e-09, 
    8.014724e-09, 6.399439e-09, 5.127418e-09, 3.883103e-09, 2.940492e-09,
  1.619863e-08, 1.575856e-08, 1.510187e-08, 1.526839e-08, 1.477525e-08, 
    1.425864e-08, 1.284265e-08, 1.151903e-08, 1.069802e-08, 9.772244e-09, 
    8.656488e-09, 7.027163e-09, 5.556103e-09, 4.263669e-09, 3.188971e-09,
  1.650413e-08, 1.623026e-08, 1.542031e-08, 1.531332e-08, 1.488793e-08, 
    1.475785e-08, 1.337528e-08, 1.195868e-08, 1.117028e-08, 1.022474e-08, 
    9.173153e-09, 7.605069e-09, 6.002496e-09, 4.646405e-09, 3.441881e-09,
  1.68718e-08, 1.654114e-08, 1.573632e-08, 1.547648e-08, 1.482693e-08, 
    1.504657e-08, 1.394851e-08, 1.247137e-08, 1.166009e-08, 1.065305e-08, 
    9.642029e-09, 8.12951e-09, 6.386871e-09, 4.986141e-09, 3.700722e-09,
  1.735802e-08, 1.691039e-08, 1.60596e-08, 1.571501e-08, 1.520623e-08, 
    1.501218e-08, 1.432701e-08, 1.269571e-08, 1.198572e-08, 1.102505e-08, 
    1.003608e-08, 8.633467e-09, 6.793581e-09, 5.310004e-09, 3.943204e-09,
  1.673351e-08, 1.648575e-08, 1.612855e-08, 1.595601e-08, 1.546175e-08, 
    1.517013e-08, 1.471922e-08, 1.311578e-08, 1.22245e-08, 1.134084e-08, 
    1.036023e-08, 9.129458e-09, 7.205624e-09, 5.621056e-09, 4.174501e-09,
  1.618321e-08, 1.628464e-08, 1.620413e-08, 1.625614e-08, 1.598227e-08, 
    1.588367e-08, 1.524934e-08, 1.350195e-08, 1.222964e-08, 1.149005e-08, 
    1.062642e-08, 9.494558e-09, 7.597131e-09, 5.920052e-09, 4.409862e-09,
  1.667134e-08, 1.62164e-08, 1.623165e-08, 1.65125e-08, 1.617621e-08, 
    1.600029e-08, 1.528315e-08, 1.389014e-08, 1.275141e-08, 1.20618e-08, 
    1.089727e-08, 9.788537e-09, 7.954434e-09, 6.20541e-09, 4.641021e-09,
  1.709467e-08, 1.626513e-08, 1.613249e-08, 1.652402e-08, 1.649622e-08, 
    1.605089e-08, 1.527491e-08, 1.41483e-08, 1.30736e-08, 1.241391e-08, 
    1.118365e-08, 1.008724e-08, 8.317122e-09, 6.478837e-09, 4.853658e-09,
  1.441506e-08, 1.307382e-08, 1.18775e-08, 1.063903e-08, 9.480372e-09, 
    8.293994e-09, 6.89377e-09, 5.39638e-09, 4.100366e-09, 3.151718e-09, 
    2.469583e-09, 1.911429e-09, 1.528074e-09, 1.230364e-09, 9.994828e-10,
  1.47413e-08, 1.367293e-08, 1.253939e-08, 1.1372e-08, 1.018188e-08, 
    9.076468e-09, 7.799845e-09, 6.264534e-09, 4.790997e-09, 3.665484e-09, 
    2.84442e-09, 2.223692e-09, 1.699231e-09, 1.360809e-09, 1.092232e-09,
  1.490137e-08, 1.417298e-08, 1.325757e-08, 1.205403e-08, 1.088506e-08, 
    9.718755e-09, 8.64587e-09, 7.19315e-09, 5.615197e-09, 4.268841e-09, 
    3.314885e-09, 2.609814e-09, 1.99996e-09, 1.550191e-09, 1.234825e-09,
  1.513807e-08, 1.430564e-08, 1.373162e-08, 1.286688e-08, 1.160052e-08, 
    1.044907e-08, 9.312905e-09, 8.055576e-09, 6.417745e-09, 4.986065e-09, 
    3.8541e-09, 3.057539e-09, 2.399875e-09, 1.827317e-09, 1.411194e-09,
  1.556909e-08, 1.480831e-08, 1.411635e-08, 1.342993e-08, 1.235179e-08, 
    1.110291e-08, 1.000493e-08, 8.958644e-09, 7.414268e-09, 5.812579e-09, 
    4.521223e-09, 3.537769e-09, 2.813366e-09, 2.18493e-09, 1.666797e-09,
  1.549634e-08, 1.495983e-08, 1.452955e-08, 1.383378e-08, 1.303791e-08, 
    1.193875e-08, 1.061997e-08, 9.521115e-09, 8.184806e-09, 6.690393e-09, 
    5.305954e-09, 4.121246e-09, 3.249045e-09, 2.57313e-09, 1.982869e-09,
  1.559902e-08, 1.521458e-08, 1.486984e-08, 1.434792e-08, 1.351284e-08, 
    1.251393e-08, 1.148862e-08, 1.044268e-08, 9.142507e-09, 7.53636e-09, 
    6.136011e-09, 4.78902e-09, 3.734726e-09, 2.970473e-09, 2.336535e-09,
  1.551904e-08, 1.508695e-08, 1.50345e-08, 1.454008e-08, 1.424096e-08, 
    1.325532e-08, 1.225335e-08, 1.118147e-08, 9.889271e-09, 8.457187e-09, 
    6.966693e-09, 5.499178e-09, 4.274632e-09, 3.370977e-09, 2.688537e-09,
  1.557305e-08, 1.525944e-08, 1.511583e-08, 1.504196e-08, 1.445637e-08, 
    1.33132e-08, 1.233189e-08, 1.156237e-08, 1.072137e-08, 9.474691e-09, 
    7.889922e-09, 6.309022e-09, 4.900199e-09, 3.803451e-09, 3.021661e-09,
  1.554776e-08, 1.530209e-08, 1.518037e-08, 1.526761e-08, 1.502431e-08, 
    1.384952e-08, 1.259836e-08, 1.194897e-08, 1.143056e-08, 1.041017e-08, 
    8.809231e-09, 7.217215e-09, 5.64173e-09, 4.322586e-09, 3.379679e-09,
  1.264999e-08, 1.073296e-08, 9.112397e-09, 7.313664e-09, 5.465311e-09, 
    3.510098e-09, 2.222719e-09, 1.684763e-09, 1.273835e-09, 9.943979e-10, 
    6.670345e-10, 3.78873e-10, 2.856969e-10, 3.09102e-10, 4.427989e-10,
  1.342272e-08, 1.16714e-08, 9.972673e-09, 8.207299e-09, 6.406211e-09, 
    4.410281e-09, 2.767683e-09, 1.912795e-09, 1.454359e-09, 1.127463e-09, 
    8.343712e-10, 4.692476e-10, 3.044783e-10, 2.608092e-10, 3.699707e-10,
  1.40526e-08, 1.24845e-08, 1.084271e-08, 9.125119e-09, 7.367836e-09, 
    5.313193e-09, 3.46414e-09, 2.234011e-09, 1.680822e-09, 1.287698e-09, 
    9.968087e-10, 6.315707e-10, 3.607418e-10, 2.405894e-10, 3.032768e-10,
  1.483084e-08, 1.318237e-08, 1.173561e-08, 1.015482e-08, 8.362705e-09, 
    6.399381e-09, 4.336367e-09, 2.734381e-09, 1.928132e-09, 1.464008e-09, 
    1.14875e-09, 8.248675e-10, 4.872583e-10, 2.707128e-10, 2.410622e-10,
  1.564211e-08, 1.405557e-08, 1.268761e-08, 1.113988e-08, 9.315894e-09, 
    7.396399e-09, 5.274674e-09, 3.473105e-09, 2.256461e-09, 1.675319e-09, 
    1.304646e-09, 1.008762e-09, 6.654136e-10, 3.677801e-10, 2.323671e-10,
  1.622362e-08, 1.474653e-08, 1.353718e-08, 1.208217e-08, 1.044149e-08, 
    8.560189e-09, 6.327513e-09, 4.272493e-09, 2.754533e-09, 1.904471e-09, 
    1.46804e-09, 1.164586e-09, 8.663362e-10, 5.312217e-10, 2.856129e-10,
  1.656057e-08, 1.572075e-08, 1.460395e-08, 1.319756e-08, 1.132415e-08, 
    9.60718e-09, 7.523477e-09, 5.346379e-09, 3.501574e-09, 2.282737e-09, 
    1.67763e-09, 1.324506e-09, 1.042814e-09, 7.315007e-10, 4.175892e-10,
  1.673375e-08, 1.599402e-08, 1.538882e-08, 1.421807e-08, 1.281632e-08, 
    1.084794e-08, 8.703847e-09, 6.432441e-09, 4.355496e-09, 2.7909e-09, 
    1.945862e-09, 1.514669e-09, 1.198734e-09, 9.229427e-10, 6.053561e-10,
  1.712726e-08, 1.64499e-08, 1.599286e-08, 1.558729e-08, 1.415246e-08, 
    1.162087e-08, 9.599467e-09, 7.487809e-09, 5.379845e-09, 3.595673e-09, 
    2.328102e-09, 1.719257e-09, 1.366588e-09, 1.089202e-09, 7.992604e-10,
  1.763532e-08, 1.678172e-08, 1.654121e-08, 1.643538e-08, 1.511286e-08, 
    1.277894e-08, 1.065521e-08, 8.668171e-09, 6.625217e-09, 4.605533e-09, 
    2.94068e-09, 2.007029e-09, 1.551335e-09, 1.240536e-09, 9.792355e-10,
  1.573582e-08, 1.257273e-08, 9.669238e-09, 6.682316e-09, 4.096316e-09, 
    2.519269e-09, 1.646774e-09, 1.350108e-09, 1.10138e-09, 9.035087e-10, 
    7.186565e-10, 4.802535e-10, 3.479157e-10, 3.527888e-10, 4.294382e-10,
  1.651622e-08, 1.377313e-08, 1.083718e-08, 7.833572e-09, 5.056297e-09, 
    3.06279e-09, 1.927994e-09, 1.484882e-09, 1.221889e-09, 9.93537e-10, 
    7.966499e-10, 5.55445e-10, 3.85685e-10, 3.647304e-10, 4.630556e-10,
  1.767262e-08, 1.495372e-08, 1.201798e-08, 9.012784e-09, 6.070208e-09, 
    3.788748e-09, 2.300482e-09, 1.661812e-09, 1.369199e-09, 1.102694e-09, 
    8.772167e-10, 6.385215e-10, 4.006663e-10, 3.558863e-10, 4.589277e-10,
  1.815897e-08, 1.560602e-08, 1.3149e-08, 1.028039e-08, 7.115477e-09, 
    4.633602e-09, 2.814848e-09, 1.894493e-09, 1.518486e-09, 1.223488e-09, 
    9.711724e-10, 7.371208e-10, 4.515801e-10, 3.36481e-10, 4.035217e-10,
  1.856192e-08, 1.639214e-08, 1.421194e-08, 1.15384e-08, 8.310942e-09, 
    5.509974e-09, 3.420475e-09, 2.177565e-09, 1.67638e-09, 1.370749e-09, 
    1.082404e-09, 8.333965e-10, 5.498544e-10, 3.489844e-10, 3.454506e-10,
  1.927632e-08, 1.699268e-08, 1.508243e-08, 1.275083e-08, 9.592263e-09, 
    6.610126e-09, 4.227564e-09, 2.568925e-09, 1.834285e-09, 1.486308e-09, 
    1.199231e-09, 9.282025e-10, 6.738349e-10, 4.020064e-10, 3.275472e-10,
  2.035526e-08, 1.811575e-08, 1.608625e-08, 1.391092e-08, 1.078812e-08, 
    7.744967e-09, 5.164645e-09, 3.29092e-09, 2.178291e-09, 1.654075e-09, 
    1.335885e-09, 1.034997e-09, 7.804299e-10, 4.947322e-10, 3.535191e-10,
  2.122388e-08, 1.866721e-08, 1.680194e-08, 1.48343e-08, 1.228574e-08, 
    9.007239e-09, 6.046124e-09, 3.79699e-09, 2.481889e-09, 1.854435e-09, 
    1.487165e-09, 1.165664e-09, 8.98523e-10, 5.911073e-10, 4.002637e-10,
  2.251608e-08, 1.960837e-08, 1.749491e-08, 1.59239e-08, 1.346514e-08, 
    1.01597e-08, 7.171022e-09, 4.519972e-09, 2.724866e-09, 1.959936e-09, 
    1.616046e-09, 1.308413e-09, 1.025953e-09, 7.004211e-10, 4.584725e-10,
  2.323213e-08, 2.066443e-08, 1.825772e-08, 1.666704e-08, 1.454748e-08, 
    1.139347e-08, 8.387955e-09, 5.557298e-09, 3.400296e-09, 2.194428e-09, 
    1.729286e-09, 1.430509e-09, 1.158671e-09, 8.298339e-10, 5.391951e-10,
  2.123591e-08, 1.696635e-08, 1.261825e-08, 9.168039e-09, 6.025056e-09, 
    3.655204e-09, 2.530784e-09, 2.053765e-09, 1.695313e-09, 1.304909e-09, 
    1.018244e-09, 7.392277e-10, 5.518935e-10, 6.397952e-10, 8.142126e-10,
  2.261084e-08, 1.851904e-08, 1.406242e-08, 1.01386e-08, 6.947729e-09, 
    4.273052e-09, 2.747891e-09, 2.167123e-09, 1.774096e-09, 1.382759e-09, 
    1.061253e-09, 8.038599e-10, 6.201476e-10, 6.119263e-10, 7.925119e-10,
  2.433767e-08, 2.006347e-08, 1.549221e-08, 1.13431e-08, 7.86703e-09, 
    5.100311e-09, 3.131485e-09, 2.301588e-09, 1.872148e-09, 1.470293e-09, 
    1.116782e-09, 8.62263e-10, 6.716439e-10, 6.610947e-10, 7.717434e-10,
  2.630702e-08, 2.16283e-08, 1.705366e-08, 1.273708e-08, 8.968878e-09, 
    6.037135e-09, 3.744838e-09, 2.517426e-09, 1.990812e-09, 1.562729e-09, 
    1.175759e-09, 8.93605e-10, 7.214231e-10, 7.08031e-10, 7.872022e-10,
  2.83409e-08, 2.384026e-08, 1.896696e-08, 1.424947e-08, 1.021319e-08, 
    6.988199e-09, 4.510428e-09, 2.875701e-09, 2.12025e-09, 1.669755e-09, 
    1.268355e-09, 9.421582e-10, 7.224346e-10, 7.171143e-10, 7.911982e-10,
  2.904339e-08, 2.561126e-08, 2.099012e-08, 1.600868e-08, 1.158743e-08, 
    8.127544e-09, 5.451214e-09, 3.471433e-09, 2.37565e-09, 1.795158e-09, 
    1.379571e-09, 1.047105e-09, 7.518044e-10, 6.964405e-10, 7.586162e-10,
  2.914417e-08, 2.70813e-08, 2.296567e-08, 1.798305e-08, 1.322439e-08, 
    9.377518e-09, 6.527695e-09, 4.470224e-09, 2.910288e-09, 1.994193e-09, 
    1.498301e-09, 1.166106e-09, 8.283788e-10, 6.967196e-10, 7.287729e-10,
  2.846057e-08, 2.764006e-08, 2.458498e-08, 2.001793e-08, 1.527917e-08, 
    1.082438e-08, 7.354724e-09, 4.957431e-09, 3.320332e-09, 2.249406e-09, 
    1.62771e-09, 1.269131e-09, 9.328668e-10, 7.200812e-10, 7.052466e-10,
  2.838617e-08, 2.803859e-08, 2.583823e-08, 2.203062e-08, 1.725284e-08, 
    1.223371e-08, 8.293767e-09, 5.578859e-09, 3.754951e-09, 2.567749e-09, 
    1.774753e-09, 1.360007e-09, 1.036479e-09, 7.589384e-10, 6.847377e-10,
  2.835365e-08, 2.843963e-08, 2.683276e-08, 2.35735e-08, 1.958939e-08, 
    1.443733e-08, 9.773651e-09, 6.592572e-09, 4.590586e-09, 3.041343e-09, 
    1.981364e-09, 1.449357e-09, 1.133252e-09, 8.268413e-10, 6.646777e-10,
  2.44121e-08, 2.377345e-08, 2.293788e-08, 2.455037e-08, 2.423355e-08, 
    2.267921e-08, 1.859636e-08, 1.381809e-08, 9.674327e-09, 7.552275e-09, 
    6.165179e-09, 4.810977e-09, 3.826868e-09, 2.853071e-09, 2.040214e-09,
  2.479438e-08, 2.423538e-08, 2.361451e-08, 2.366074e-08, 2.354942e-08, 
    2.328893e-08, 1.949106e-08, 1.446096e-08, 1.00242e-08, 7.703812e-09, 
    6.231641e-09, 4.875179e-09, 3.869832e-09, 2.935728e-09, 2.088527e-09,
  2.5075e-08, 2.439309e-08, 2.356287e-08, 2.241155e-08, 2.310627e-08, 
    2.315381e-08, 2.023113e-08, 1.509202e-08, 1.044564e-08, 7.846983e-09, 
    6.29351e-09, 4.91762e-09, 3.911492e-09, 3.005762e-09, 2.155172e-09,
  2.535814e-08, 2.425854e-08, 2.372611e-08, 2.275544e-08, 2.254761e-08, 
    2.290955e-08, 2.091771e-08, 1.582456e-08, 1.081319e-08, 7.992973e-09, 
    6.333631e-09, 4.913137e-09, 3.903552e-09, 3.045359e-09, 2.19937e-09,
  2.540476e-08, 2.444358e-08, 2.383318e-08, 2.262246e-08, 2.198286e-08, 
    2.234055e-08, 2.13874e-08, 1.679807e-08, 1.145353e-08, 8.203558e-09, 
    6.404405e-09, 4.895496e-09, 3.882183e-09, 3.046258e-09, 2.218387e-09,
  2.646538e-08, 2.447816e-08, 2.383949e-08, 2.293053e-08, 2.179186e-08, 
    2.161821e-08, 2.144814e-08, 1.741148e-08, 1.190431e-08, 8.490815e-09, 
    6.456924e-09, 4.851952e-09, 3.829923e-09, 3.021055e-09, 2.20999e-09,
  2.750852e-08, 2.526954e-08, 2.424639e-08, 2.311859e-08, 2.159504e-08, 
    2.102429e-08, 2.123548e-08, 1.832145e-08, 1.264672e-08, 8.764104e-09, 
    6.479403e-09, 4.785027e-09, 3.783502e-09, 2.972243e-09, 2.191753e-09,
  2.848835e-08, 2.613063e-08, 2.464184e-08, 2.348551e-08, 2.173796e-08, 
    2.054788e-08, 2.063027e-08, 1.87727e-08, 1.351613e-08, 9.149518e-09, 
    6.591596e-09, 4.747933e-09, 3.725048e-09, 2.92671e-09, 2.159845e-09,
  2.891268e-08, 2.70689e-08, 2.522155e-08, 2.381235e-08, 2.18704e-08, 
    2.053156e-08, 2.055528e-08, 1.914505e-08, 1.412239e-08, 9.417581e-09, 
    6.712402e-09, 4.71846e-09, 3.650862e-09, 2.871625e-09, 2.125835e-09,
  2.854596e-08, 2.769717e-08, 2.61561e-08, 2.435895e-08, 2.256187e-08, 
    2.084439e-08, 2.030703e-08, 1.905181e-08, 1.451117e-08, 9.694059e-09, 
    6.865409e-09, 4.743654e-09, 3.586504e-09, 2.817724e-09, 2.091963e-09,
  2.660859e-08, 2.586202e-08, 2.511796e-08, 2.291843e-08, 1.880257e-08, 
    1.598538e-08, 1.385324e-08, 1.136832e-08, 1.04222e-08, 1.083943e-08, 
    9.825266e-09, 7.818924e-09, 6.139881e-09, 4.932548e-09, 3.964387e-09,
  2.810686e-08, 2.680088e-08, 2.59847e-08, 2.453228e-08, 2.178914e-08, 
    1.733973e-08, 1.484129e-08, 1.233806e-08, 1.064514e-08, 1.058104e-08, 
    1.033074e-08, 8.665268e-09, 6.609166e-09, 5.292793e-09, 4.193637e-09,
  3.045418e-08, 2.860719e-08, 2.722338e-08, 2.56401e-08, 2.34267e-08, 
    1.940719e-08, 1.593547e-08, 1.336379e-08, 1.154979e-08, 1.059481e-08, 
    1.050389e-08, 9.238543e-09, 7.140053e-09, 5.576417e-09, 4.416185e-09,
  3.053106e-08, 3.096689e-08, 2.854157e-08, 2.687667e-08, 2.478906e-08, 
    2.175669e-08, 1.765625e-08, 1.462606e-08, 1.24169e-08, 1.07864e-08, 
    1.065745e-08, 9.777375e-09, 7.668587e-09, 5.914222e-09, 4.660186e-09,
  2.89653e-08, 3.153103e-08, 2.992002e-08, 2.791407e-08, 2.600893e-08, 
    2.312732e-08, 1.932063e-08, 1.662944e-08, 1.385745e-08, 1.148095e-08, 
    1.063048e-08, 1.010459e-08, 8.15058e-09, 6.294485e-09, 4.926108e-09,
  2.685477e-08, 2.940503e-08, 3.037561e-08, 2.839411e-08, 2.702149e-08, 
    2.474361e-08, 2.106316e-08, 1.805404e-08, 1.533465e-08, 1.268824e-08, 
    1.082824e-08, 1.035661e-08, 8.579901e-09, 6.694912e-09, 5.196883e-09,
  2.553655e-08, 2.783272e-08, 2.920843e-08, 2.951113e-08, 2.753871e-08, 
    2.588849e-08, 2.250328e-08, 2.003275e-08, 1.720327e-08, 1.400141e-08, 
    1.143728e-08, 1.039077e-08, 8.933608e-09, 7.075435e-09, 5.467446e-09,
  2.511818e-08, 2.741243e-08, 2.84294e-08, 2.861837e-08, 2.851588e-08, 
    2.719172e-08, 2.416487e-08, 2.156872e-08, 1.99169e-08, 1.609885e-08, 
    1.235104e-08, 1.051604e-08, 9.20434e-09, 7.453246e-09, 5.731751e-09,
  2.497409e-08, 2.738377e-08, 2.72532e-08, 2.737609e-08, 2.820465e-08, 
    2.856276e-08, 2.705209e-08, 2.349591e-08, 2.116789e-08, 1.801403e-08, 
    1.355914e-08, 1.07037e-08, 9.422545e-09, 7.751964e-09, 5.975595e-09,
  2.4666e-08, 2.696433e-08, 2.706014e-08, 2.659232e-08, 2.750495e-08, 
    2.862496e-08, 2.85222e-08, 2.529587e-08, 2.230416e-08, 2.000663e-08, 
    1.516365e-08, 1.124891e-08, 9.597564e-09, 7.99936e-09, 6.197082e-09,
  1.820302e-08, 1.719683e-08, 1.586148e-08, 1.48014e-08, 1.468544e-08, 
    1.488073e-08, 1.489784e-08, 1.463782e-08, 1.373004e-08, 1.170687e-08, 
    9.554114e-09, 7.659147e-09, 5.708909e-09, 4.336433e-09, 3.628205e-09,
  1.818239e-08, 1.777332e-08, 1.662102e-08, 1.524688e-08, 1.456528e-08, 
    1.453893e-08, 1.477322e-08, 1.463809e-08, 1.418431e-08, 1.275073e-08, 
    1.04854e-08, 8.616469e-09, 6.640048e-09, 4.868561e-09, 3.897443e-09,
  1.795264e-08, 1.864191e-08, 1.782551e-08, 1.614067e-08, 1.493328e-08, 
    1.446736e-08, 1.451334e-08, 1.44906e-08, 1.433001e-08, 1.347733e-08, 
    1.159944e-08, 9.549479e-09, 7.473536e-09, 5.541437e-09, 4.257021e-09,
  1.806243e-08, 1.8891e-08, 1.888915e-08, 1.724246e-08, 1.564054e-08, 
    1.465802e-08, 1.440526e-08, 1.414509e-08, 1.39722e-08, 1.38726e-08, 
    1.271429e-08, 1.069932e-08, 8.455912e-09, 6.259904e-09, 4.652144e-09,
  1.981438e-08, 1.930499e-08, 1.960398e-08, 1.843532e-08, 1.653545e-08, 
    1.484463e-08, 1.43142e-08, 1.404153e-08, 1.375498e-08, 1.372007e-08, 
    1.316426e-08, 1.191269e-08, 9.479666e-09, 7.021681e-09, 5.059909e-09,
  2.085919e-08, 2.00996e-08, 1.996462e-08, 1.912723e-08, 1.758845e-08, 
    1.542656e-08, 1.412599e-08, 1.328768e-08, 1.304368e-08, 1.319182e-08, 
    1.297617e-08, 1.269276e-08, 1.064574e-08, 7.854974e-09, 5.570811e-09,
  2.141874e-08, 2.041166e-08, 2.009337e-08, 1.990989e-08, 1.839423e-08, 
    1.57563e-08, 1.414982e-08, 1.29457e-08, 1.263584e-08, 1.270099e-08, 
    1.238695e-08, 1.293341e-08, 1.160703e-08, 8.654551e-09, 6.169894e-09,
  2.255257e-08, 2.118236e-08, 2.041545e-08, 2.031757e-08, 1.955698e-08, 
    1.696703e-08, 1.515332e-08, 1.466288e-08, 1.400649e-08, 1.27484e-08, 
    1.222639e-08, 1.324313e-08, 1.224376e-08, 9.586598e-09, 6.874476e-09,
  2.425669e-08, 2.232639e-08, 2.079461e-08, 2.023036e-08, 2.047354e-08, 
    1.929865e-08, 1.739204e-08, 1.564976e-08, 1.406987e-08, 1.246617e-08, 
    1.208686e-08, 1.286351e-08, 1.283031e-08, 1.043864e-08, 7.572225e-09,
  2.476939e-08, 2.368177e-08, 2.151144e-08, 2.037346e-08, 2.111406e-08, 
    2.083123e-08, 1.897819e-08, 1.624751e-08, 1.369515e-08, 1.235484e-08, 
    1.205438e-08, 1.242354e-08, 1.299485e-08, 1.126578e-08, 8.210307e-09,
  2.13889e-08, 1.98865e-08, 1.910479e-08, 1.949268e-08, 1.963806e-08, 
    1.864421e-08, 1.762073e-08, 1.617328e-08, 1.439019e-08, 1.224058e-08, 
    1.00389e-08, 8.20067e-09, 6.477542e-09, 4.96901e-09, 4.041572e-09,
  2.289962e-08, 2.061603e-08, 1.95045e-08, 1.915079e-08, 1.967061e-08, 
    1.937063e-08, 1.829143e-08, 1.692245e-08, 1.532254e-08, 1.342132e-08, 
    1.113746e-08, 9.098549e-09, 7.310838e-09, 5.603584e-09, 4.459493e-09,
  2.477331e-08, 2.182529e-08, 2.007632e-08, 1.925289e-08, 1.935743e-08, 
    1.966333e-08, 1.883591e-08, 1.757772e-08, 1.62015e-08, 1.441911e-08, 
    1.223675e-08, 1.006672e-08, 8.142286e-09, 6.283353e-09, 4.878419e-09,
  2.630572e-08, 2.325017e-08, 2.106728e-08, 1.965315e-08, 1.924686e-08, 
    1.972401e-08, 1.940936e-08, 1.818138e-08, 1.681127e-08, 1.533362e-08, 
    1.327803e-08, 1.096256e-08, 8.999876e-09, 7.066409e-09, 5.357628e-09,
  2.853632e-08, 2.503185e-08, 2.248145e-08, 2.019162e-08, 1.941408e-08, 
    1.952106e-08, 1.976393e-08, 1.893334e-08, 1.749573e-08, 1.61163e-08, 
    1.41845e-08, 1.190751e-08, 9.788546e-09, 7.825784e-09, 5.925359e-09,
  2.842519e-08, 2.621431e-08, 2.367849e-08, 2.121401e-08, 1.980042e-08, 
    1.953088e-08, 1.977446e-08, 1.92388e-08, 1.803648e-08, 1.685101e-08, 
    1.522129e-08, 1.291683e-08, 1.06003e-08, 8.623699e-09, 6.563871e-09,
  2.730616e-08, 2.638082e-08, 2.431945e-08, 2.225505e-08, 2.014451e-08, 
    1.964097e-08, 1.969616e-08, 1.968248e-08, 1.864928e-08, 1.741488e-08, 
    1.597251e-08, 1.393386e-08, 1.152814e-08, 9.457236e-09, 7.268277e-09,
  2.636711e-08, 2.631849e-08, 2.500038e-08, 2.299949e-08, 2.098045e-08, 
    1.965533e-08, 1.946753e-08, 1.947587e-08, 1.860092e-08, 1.749568e-08, 
    1.631336e-08, 1.468866e-08, 1.230847e-08, 1.017387e-08, 7.992519e-09,
  2.585362e-08, 2.629508e-08, 2.537001e-08, 2.327211e-08, 2.137409e-08, 
    2.007426e-08, 1.935235e-08, 1.931527e-08, 1.890519e-08, 1.792992e-08, 
    1.658892e-08, 1.527482e-08, 1.327557e-08, 1.091547e-08, 8.628133e-09,
  2.555878e-08, 2.596561e-08, 2.543451e-08, 2.377731e-08, 2.221302e-08, 
    2.0575e-08, 1.921404e-08, 1.919861e-08, 1.898424e-08, 1.818029e-08, 
    1.678906e-08, 1.565312e-08, 1.395415e-08, 1.165933e-08, 9.169504e-09,
  2.328502e-08, 2.398401e-08, 2.433226e-08, 2.306829e-08, 2.186615e-08, 
    2.145866e-08, 2.044255e-08, 1.825954e-08, 1.57008e-08, 1.314702e-08, 
    1.100622e-08, 8.709944e-09, 6.469849e-09, 5.329732e-09, 4.354221e-09,
  2.341143e-08, 2.382565e-08, 2.419564e-08, 2.394995e-08, 2.254172e-08, 
    2.178389e-08, 2.128361e-08, 1.983301e-08, 1.747084e-08, 1.484125e-08, 
    1.256159e-08, 1.045599e-08, 8.145478e-09, 6.161109e-09, 4.826944e-09,
  2.380074e-08, 2.400903e-08, 2.434514e-08, 2.427412e-08, 2.342559e-08, 
    2.219203e-08, 2.157011e-08, 2.083193e-08, 1.91038e-08, 1.648224e-08, 
    1.402116e-08, 1.191598e-08, 9.685934e-09, 7.463989e-09, 5.507797e-09,
  2.455631e-08, 2.380622e-08, 2.389972e-08, 2.425046e-08, 2.395466e-08, 
    2.291048e-08, 2.190283e-08, 2.129385e-08, 2.030594e-08, 1.81117e-08, 
    1.561924e-08, 1.330921e-08, 1.122495e-08, 8.979857e-09, 6.717923e-09,
  2.531853e-08, 2.453206e-08, 2.368682e-08, 2.412608e-08, 2.410178e-08, 
    2.344396e-08, 2.239641e-08, 2.164369e-08, 2.106279e-08, 1.95173e-08, 
    1.711225e-08, 1.472461e-08, 1.254138e-08, 1.037102e-08, 8.067093e-09,
  2.486308e-08, 2.430269e-08, 2.345546e-08, 2.343407e-08, 2.406694e-08, 
    2.404165e-08, 2.299657e-08, 2.188891e-08, 2.143591e-08, 2.053961e-08, 
    1.851322e-08, 1.603687e-08, 1.368761e-08, 1.147651e-08, 9.269224e-09,
  2.51349e-08, 2.474959e-08, 2.366987e-08, 2.317533e-08, 2.340668e-08, 
    2.38391e-08, 2.37975e-08, 2.273827e-08, 2.181962e-08, 2.107954e-08, 
    1.962514e-08, 1.712843e-08, 1.479049e-08, 1.249485e-08, 1.02558e-08,
  2.552992e-08, 2.539547e-08, 2.439041e-08, 2.297444e-08, 2.371131e-08, 
    2.373356e-08, 2.382212e-08, 2.323154e-08, 2.235564e-08, 2.145112e-08, 
    2.038314e-08, 1.810803e-08, 1.573497e-08, 1.350799e-08, 1.122536e-08,
  2.562438e-08, 2.563462e-08, 2.503647e-08, 2.310498e-08, 2.329172e-08, 
    2.369903e-08, 2.366656e-08, 2.308161e-08, 2.236906e-08, 2.159855e-08, 
    2.083575e-08, 1.898296e-08, 1.668088e-08, 1.453233e-08, 1.230668e-08,
  2.518362e-08, 2.565117e-08, 2.580084e-08, 2.371078e-08, 2.277905e-08, 
    2.333539e-08, 2.44448e-08, 2.340617e-08, 2.26505e-08, 2.177734e-08, 
    2.105932e-08, 1.963496e-08, 1.754475e-08, 1.548339e-08, 1.329508e-08,
  2.215906e-08, 2.13376e-08, 2.131901e-08, 2.259941e-08, 2.302009e-08, 
    2.303131e-08, 2.200641e-08, 1.930485e-08, 1.545383e-08, 1.158768e-08, 
    7.987027e-09, 5.531999e-09, 4.018191e-09, 3.236687e-09, 2.214414e-09,
  2.316925e-08, 2.198493e-08, 2.133769e-08, 2.183512e-08, 2.283432e-08, 
    2.313745e-08, 2.295963e-08, 2.129781e-08, 1.805417e-08, 1.421474e-08, 
    1.034549e-08, 7.27494e-09, 4.777866e-09, 3.510196e-09, 2.494e-09,
  2.402055e-08, 2.316306e-08, 2.173521e-08, 2.151809e-08, 2.209028e-08, 
    2.284717e-08, 2.331365e-08, 2.242104e-08, 2.025492e-08, 1.673231e-08, 
    1.272174e-08, 9.188943e-09, 6.073913e-09, 3.949813e-09, 2.806772e-09,
  2.319854e-08, 2.369334e-08, 2.252761e-08, 2.166646e-08, 2.177591e-08, 
    2.2397e-08, 2.304919e-08, 2.323492e-08, 2.163512e-08, 1.90405e-08, 
    1.512027e-08, 1.144027e-08, 7.913367e-09, 4.890376e-09, 3.328624e-09,
  2.255e-08, 2.374771e-08, 2.342472e-08, 2.205047e-08, 2.167843e-08, 
    2.206358e-08, 2.259601e-08, 2.350433e-08, 2.257232e-08, 2.070278e-08, 
    1.729473e-08, 1.370246e-08, 9.944365e-09, 6.558944e-09, 4.17154e-09,
  2.124192e-08, 2.26569e-08, 2.333172e-08, 2.278078e-08, 2.187116e-08, 
    2.193125e-08, 2.231534e-08, 2.298719e-08, 2.324997e-08, 2.198713e-08, 
    1.92511e-08, 1.586288e-08, 1.208148e-08, 8.596332e-09, 5.429266e-09,
  2.149863e-08, 2.200557e-08, 2.298111e-08, 2.310458e-08, 2.222322e-08, 
    2.185843e-08, 2.224174e-08, 2.270646e-08, 2.307659e-08, 2.266184e-08, 
    2.074513e-08, 1.780324e-08, 1.419317e-08, 1.059647e-08, 7.153712e-09,
  2.229218e-08, 2.202996e-08, 2.252673e-08, 2.305359e-08, 2.288624e-08, 
    2.208604e-08, 2.211495e-08, 2.288131e-08, 2.360203e-08, 2.31876e-08, 
    2.177607e-08, 1.940366e-08, 1.614614e-08, 1.244896e-08, 8.886402e-09,
  2.314032e-08, 2.210792e-08, 2.2211e-08, 2.285971e-08, 2.319327e-08, 
    2.276889e-08, 2.238472e-08, 2.256364e-08, 2.310736e-08, 2.331104e-08, 
    2.249967e-08, 2.070484e-08, 1.771486e-08, 1.429271e-08, 1.053909e-08,
  2.429238e-08, 2.249076e-08, 2.213029e-08, 2.249037e-08, 2.334852e-08, 
    2.303856e-08, 2.28893e-08, 2.254453e-08, 2.263644e-08, 2.314208e-08, 
    2.290093e-08, 2.167504e-08, 1.904411e-08, 1.590713e-08, 1.203199e-08,
  2.254005e-08, 2.341998e-08, 2.342813e-08, 2.306427e-08, 2.324285e-08, 
    2.310905e-08, 2.152856e-08, 1.856496e-08, 1.533703e-08, 1.218621e-08, 
    8.490326e-09, 5.429742e-09, 3.844245e-09, 2.115641e-09, 1.018208e-09,
  2.135363e-08, 2.298719e-08, 2.367356e-08, 2.342247e-08, 2.313905e-08, 
    2.351631e-08, 2.287323e-08, 2.072652e-08, 1.764651e-08, 1.430677e-08, 
    1.086241e-08, 7.02258e-09, 4.653413e-09, 2.66351e-09, 1.208171e-09,
  2.102627e-08, 2.206182e-08, 2.335157e-08, 2.37093e-08, 2.326711e-08, 
    2.314983e-08, 2.347604e-08, 2.22895e-08, 1.966397e-08, 1.638212e-08, 
    1.304288e-08, 8.96973e-09, 5.654478e-09, 3.268513e-09, 1.498922e-09,
  2.092704e-08, 2.16086e-08, 2.258168e-08, 2.369662e-08, 2.38281e-08, 
    2.332229e-08, 2.335654e-08, 2.324168e-08, 2.151747e-08, 1.847898e-08, 
    1.523894e-08, 1.119067e-08, 7.157999e-09, 4.077418e-09, 1.941688e-09,
  2.095068e-08, 2.108719e-08, 2.188707e-08, 2.282543e-08, 2.371216e-08, 
    2.368248e-08, 2.332903e-08, 2.358909e-08, 2.266468e-08, 2.018901e-08, 
    1.730588e-08, 1.345313e-08, 8.971154e-09, 5.116903e-09, 2.483367e-09,
  2.084641e-08, 2.069609e-08, 2.121174e-08, 2.225342e-08, 2.332196e-08, 
    2.413896e-08, 2.366328e-08, 2.348779e-08, 2.368662e-08, 2.181688e-08, 
    1.907748e-08, 1.5648e-08, 1.105621e-08, 6.463138e-09, 3.139361e-09,
  2.154945e-08, 2.111937e-08, 2.100705e-08, 2.187874e-08, 2.266968e-08, 
    2.3663e-08, 2.420316e-08, 2.382578e-08, 2.383659e-08, 2.296265e-08, 
    2.06982e-08, 1.761775e-08, 1.32182e-08, 8.149279e-09, 4.057011e-09,
  2.219604e-08, 2.179099e-08, 2.122642e-08, 2.129917e-08, 2.260565e-08, 
    2.330993e-08, 2.396987e-08, 2.369752e-08, 2.398168e-08, 2.367124e-08, 
    2.20088e-08, 1.938692e-08, 1.524234e-08, 1.006287e-08, 5.242235e-09,
  2.266984e-08, 2.208536e-08, 2.157517e-08, 2.151358e-08, 2.189318e-08, 
    2.225426e-08, 2.352791e-08, 2.349834e-08, 2.385518e-08, 2.402618e-08, 
    2.293206e-08, 2.06321e-08, 1.707639e-08, 1.199427e-08, 6.608018e-09,
  2.379136e-08, 2.23826e-08, 2.183317e-08, 2.181581e-08, 2.128167e-08, 
    2.186816e-08, 2.304485e-08, 2.372201e-08, 2.390562e-08, 2.418007e-08, 
    2.358176e-08, 2.171539e-08, 1.842954e-08, 1.37251e-08, 8.182059e-09,
  2.349361e-08, 2.315629e-08, 2.263979e-08, 2.382002e-08, 2.535508e-08, 
    2.364507e-08, 2.010024e-08, 1.62298e-08, 1.142967e-08, 6.715184e-09, 
    3.567636e-09, 2.42038e-09, 1.790148e-09, 9.534479e-10, 5.273003e-10,
  2.276761e-08, 2.352068e-08, 2.307521e-08, 2.315962e-08, 2.450577e-08, 
    2.48715e-08, 2.231382e-08, 1.895179e-08, 1.447981e-08, 9.238976e-09, 
    4.9399e-09, 2.910628e-09, 2.171743e-09, 1.314066e-09, 6.471773e-10,
  2.108916e-08, 2.307917e-08, 2.322654e-08, 2.303828e-08, 2.348944e-08, 
    2.457271e-08, 2.396929e-08, 2.099507e-08, 1.724187e-08, 1.225861e-08, 
    6.962529e-09, 3.772763e-09, 2.569356e-09, 1.718519e-09, 8.764962e-10,
  1.972116e-08, 2.208363e-08, 2.312794e-08, 2.32035e-08, 2.332629e-08, 
    2.380003e-08, 2.445458e-08, 2.278239e-08, 1.951805e-08, 1.518612e-08, 
    9.478137e-09, 5.109828e-09, 3.125969e-09, 2.169722e-09, 1.207496e-09,
  1.921473e-08, 2.036922e-08, 2.239981e-08, 2.291265e-08, 2.337107e-08, 
    2.340817e-08, 2.387819e-08, 2.376652e-08, 2.134384e-08, 1.777212e-08, 
    1.256239e-08, 6.989795e-09, 3.898282e-09, 2.646751e-09, 1.594195e-09,
  1.968897e-08, 1.938027e-08, 2.133889e-08, 2.229528e-08, 2.319769e-08, 
    2.360402e-08, 2.361258e-08, 2.411552e-08, 2.276854e-08, 1.971497e-08, 
    1.533617e-08, 9.416363e-09, 5.113264e-09, 3.180212e-09, 2.019524e-09,
  2.114443e-08, 1.95802e-08, 2.004293e-08, 2.167746e-08, 2.262772e-08, 
    2.35131e-08, 2.379221e-08, 2.405047e-08, 2.367752e-08, 2.155112e-08, 
    1.779501e-08, 1.221806e-08, 6.806205e-09, 3.898637e-09, 2.47618e-09,
  2.272131e-08, 2.067426e-08, 1.970846e-08, 2.074916e-08, 2.214733e-08, 
    2.3212e-08, 2.377764e-08, 2.373457e-08, 2.393371e-08, 2.254497e-08, 
    1.962887e-08, 1.493359e-08, 8.984688e-09, 4.960222e-09, 2.978291e-09,
  2.345022e-08, 2.161275e-08, 2.006824e-08, 2.025593e-08, 2.142047e-08, 
    2.27473e-08, 2.356824e-08, 2.321204e-08, 2.362976e-08, 2.32968e-08, 
    2.128172e-08, 1.723951e-08, 1.145789e-08, 6.411735e-09, 3.634221e-09,
  2.363749e-08, 2.254574e-08, 2.063902e-08, 2.015408e-08, 2.070363e-08, 
    2.187537e-08, 2.329773e-08, 2.338311e-08, 2.356481e-08, 2.361644e-08, 
    2.259607e-08, 1.922142e-08, 1.390948e-08, 8.210159e-09, 4.517044e-09,
  2.343225e-08, 2.370188e-08, 2.408551e-08, 2.321572e-08, 2.111164e-08, 
    1.780246e-08, 1.424632e-08, 1.031931e-08, 6.855942e-09, 3.654033e-09, 
    1.821043e-09, 9.608138e-10, 1.126328e-09, 9.295715e-10, 7.073737e-10,
  2.313e-08, 2.388305e-08, 2.413663e-08, 2.374649e-08, 2.216787e-08, 
    1.93169e-08, 1.580979e-08, 1.19095e-08, 8.354654e-09, 5.070447e-09, 
    2.487073e-09, 1.147057e-09, 1.122582e-09, 1.306001e-09, 7.808617e-10,
  2.276217e-08, 2.437805e-08, 2.454336e-08, 2.405181e-08, 2.302706e-08, 
    2.086096e-08, 1.737972e-08, 1.357341e-08, 9.904718e-09, 6.729429e-09, 
    3.61521e-09, 1.575199e-09, 1.105673e-09, 1.468963e-09, 9.762682e-10,
  2.186244e-08, 2.469319e-08, 2.532544e-08, 2.454328e-08, 2.381191e-08, 
    2.210991e-08, 1.934536e-08, 1.535582e-08, 1.150608e-08, 8.291745e-09, 
    5.036573e-09, 2.192651e-09, 1.273054e-09, 1.690617e-09, 1.352658e-09,
  2.212921e-08, 2.444455e-08, 2.606092e-08, 2.562025e-08, 2.467709e-08, 
    2.294327e-08, 2.085211e-08, 1.758761e-08, 1.340988e-08, 1.000366e-08, 
    6.647154e-09, 3.247377e-09, 1.406883e-09, 1.745593e-09, 1.708598e-09,
  2.253288e-08, 2.340392e-08, 2.57094e-08, 2.572254e-08, 2.530106e-08, 
    2.39728e-08, 2.201559e-08, 1.9099e-08, 1.514551e-08, 1.153822e-08, 
    8.38036e-09, 4.833524e-09, 2.052866e-09, 1.701735e-09, 1.918598e-09,
  2.250553e-08, 2.238617e-08, 2.429463e-08, 2.578488e-08, 2.51564e-08, 
    2.427703e-08, 2.244054e-08, 2.058677e-08, 1.75788e-08, 1.338197e-08, 
    1.019022e-08, 6.648173e-09, 3.284721e-09, 1.671413e-09, 1.807091e-09,
  2.327644e-08, 2.247655e-08, 2.332165e-08, 2.495974e-08, 2.510562e-08, 
    2.454211e-08, 2.323353e-08, 2.160895e-08, 1.984846e-08, 1.575815e-08, 
    1.210567e-08, 8.66536e-09, 4.930788e-09, 2.279923e-09, 1.554973e-09,
  2.37628e-08, 2.278736e-08, 2.258696e-08, 2.361468e-08, 2.505874e-08, 
    2.599601e-08, 2.520775e-08, 2.27486e-08, 2.021617e-08, 1.698979e-08, 
    1.395551e-08, 1.056362e-08, 6.727899e-09, 3.365971e-09, 1.689305e-09,
  2.399902e-08, 2.317627e-08, 2.248114e-08, 2.278794e-08, 2.450425e-08, 
    2.589802e-08, 2.584466e-08, 2.358939e-08, 2.088445e-08, 1.843185e-08, 
    1.569756e-08, 1.220523e-08, 8.628007e-09, 4.831203e-09, 2.183873e-09,
  2.664916e-08, 2.754799e-08, 2.673706e-08, 2.380721e-08, 1.933846e-08, 
    1.443127e-08, 9.60567e-09, 5.587617e-09, 3.171233e-09, 1.734569e-09, 
    1.030078e-09, 8.042607e-10, 8.024942e-10, 7.68161e-10, 5.394382e-10,
  2.609715e-08, 2.734972e-08, 2.727942e-08, 2.487976e-08, 2.060255e-08, 
    1.56695e-08, 1.074073e-08, 6.46203e-09, 3.626801e-09, 2.019483e-09, 
    1.121966e-09, 8.073788e-10, 7.732295e-10, 7.222791e-10, 5.106091e-10,
  2.572769e-08, 2.723954e-08, 2.757736e-08, 2.573475e-08, 2.184034e-08, 
    1.689124e-08, 1.194495e-08, 7.438704e-09, 4.204868e-09, 2.347713e-09, 
    1.247893e-09, 8.280446e-10, 7.401765e-10, 6.85331e-10, 4.920211e-10,
  2.502635e-08, 2.678997e-08, 2.781917e-08, 2.632528e-08, 2.301728e-08, 
    1.814656e-08, 1.307755e-08, 8.404565e-09, 4.847035e-09, 2.666203e-09, 
    1.400909e-09, 8.576503e-10, 7.09598e-10, 6.552234e-10, 5.013671e-10,
  2.509054e-08, 2.646526e-08, 2.773253e-08, 2.697736e-08, 2.396827e-08, 
    1.940656e-08, 1.424628e-08, 9.50226e-09, 5.624408e-09, 3.015145e-09, 
    1.594176e-09, 9.020671e-10, 6.98651e-10, 6.518894e-10, 5.274704e-10,
  2.448965e-08, 2.576348e-08, 2.733947e-08, 2.721908e-08, 2.488727e-08, 
    2.060411e-08, 1.53702e-08, 1.042548e-08, 6.359583e-09, 3.423561e-09, 
    1.820481e-09, 9.804757e-10, 7.102018e-10, 6.606298e-10, 5.559496e-10,
  2.402745e-08, 2.499944e-08, 2.668579e-08, 2.73757e-08, 2.547499e-08, 
    2.168327e-08, 1.654091e-08, 1.153069e-08, 7.259942e-09, 4.057052e-09, 
    2.088443e-09, 1.100495e-09, 7.487644e-10, 6.583619e-10, 5.712616e-10,
  2.40045e-08, 2.47101e-08, 2.613833e-08, 2.719311e-08, 2.598807e-08, 
    2.256833e-08, 1.764747e-08, 1.256205e-08, 8.242868e-09, 4.769556e-09, 
    2.388259e-09, 1.26917e-09, 8.052129e-10, 6.684752e-10, 5.765126e-10,
  2.415461e-08, 2.445825e-08, 2.576988e-08, 2.682823e-08, 2.635872e-08, 
    2.372337e-08, 1.916342e-08, 1.393998e-08, 9.282365e-09, 5.439682e-09, 
    2.745041e-09, 1.465573e-09, 8.724592e-10, 6.760625e-10, 5.638343e-10,
  2.420157e-08, 2.428283e-08, 2.524601e-08, 2.654678e-08, 2.659015e-08, 
    2.445777e-08, 2.023221e-08, 1.496923e-08, 1.021444e-08, 6.181029e-09, 
    3.221525e-09, 1.697921e-09, 9.544295e-10, 6.960959e-10, 5.46852e-10,
  2.280635e-08, 2.178086e-08, 2.18427e-08, 2.326549e-08, 2.07079e-08, 
    1.538367e-08, 1.008931e-08, 5.361775e-09, 2.895192e-09, 2.165158e-09, 
    1.618855e-09, 1.079371e-09, 6.882033e-10, 5.69992e-10, 4.656917e-10,
  2.329551e-08, 2.203699e-08, 2.168459e-08, 2.323997e-08, 2.185161e-08, 
    1.663862e-08, 1.137623e-08, 6.249575e-09, 3.217667e-09, 2.340478e-09, 
    1.774e-09, 1.188431e-09, 7.558646e-10, 6.262313e-10, 4.788571e-10,
  2.374657e-08, 2.244916e-08, 2.167875e-08, 2.286945e-08, 2.272766e-08, 
    1.802528e-08, 1.260485e-08, 7.309986e-09, 3.630869e-09, 2.514255e-09, 
    1.928624e-09, 1.275821e-09, 7.893641e-10, 6.236173e-10, 5.031293e-10,
  2.444135e-08, 2.304029e-08, 2.182777e-08, 2.256116e-08, 2.335238e-08, 
    1.952025e-08, 1.384292e-08, 8.384686e-09, 4.095217e-09, 2.721898e-09, 
    2.066481e-09, 1.34928e-09, 7.928118e-10, 6.036125e-10, 5.22446e-10,
  2.509247e-08, 2.378911e-08, 2.230517e-08, 2.215175e-08, 2.365343e-08, 
    2.063963e-08, 1.526847e-08, 9.605315e-09, 4.736227e-09, 2.944479e-09, 
    2.216918e-09, 1.445554e-09, 8.049568e-10, 5.80768e-10, 5.23619e-10,
  2.529308e-08, 2.415618e-08, 2.27512e-08, 2.200468e-08, 2.362441e-08, 
    2.167647e-08, 1.657306e-08, 1.065888e-08, 5.42993e-09, 3.158749e-09, 
    2.366644e-09, 1.542428e-09, 8.190451e-10, 5.726262e-10, 5.406894e-10,
  2.512366e-08, 2.461185e-08, 2.319835e-08, 2.217249e-08, 2.322187e-08, 
    2.236523e-08, 1.786272e-08, 1.194494e-08, 6.263458e-09, 3.472725e-09, 
    2.534469e-09, 1.639849e-09, 8.50417e-10, 5.796958e-10, 5.791985e-10,
  2.512147e-08, 2.503869e-08, 2.3857e-08, 2.256259e-08, 2.29561e-08, 
    2.277926e-08, 1.912757e-08, 1.349241e-08, 7.386991e-09, 3.846379e-09, 
    2.72598e-09, 1.772051e-09, 9.212377e-10, 5.942227e-10, 5.948685e-10,
  2.471316e-08, 2.518876e-08, 2.437648e-08, 2.290466e-08, 2.296067e-08, 
    2.358135e-08, 2.065192e-08, 1.509806e-08, 8.396039e-09, 4.073467e-09, 
    2.87407e-09, 1.911592e-09, 1.007758e-09, 6.238871e-10, 5.967858e-10,
  2.415178e-08, 2.505224e-08, 2.481407e-08, 2.364176e-08, 2.278018e-08, 
    2.381559e-08, 2.164277e-08, 1.643624e-08, 9.417584e-09, 4.487995e-09, 
    3.024686e-09, 2.06153e-09, 1.091577e-09, 6.748448e-10, 6.116539e-10,
  2.486714e-08, 2.470898e-08, 2.459292e-08, 2.43784e-08, 2.408729e-08, 
    2.325891e-08, 2.167287e-08, 1.87389e-08, 1.524239e-08, 1.172412e-08, 
    7.984863e-09, 5.281465e-09, 3.222177e-09, 1.970264e-09, 1.4453e-09,
  2.507297e-08, 2.502798e-08, 2.468803e-08, 2.453981e-08, 2.426937e-08, 
    2.344933e-08, 2.19178e-08, 1.887647e-08, 1.553065e-08, 1.209067e-08, 
    8.42183e-09, 5.569363e-09, 3.389292e-09, 2.100168e-09, 1.505963e-09,
  2.5036e-08, 2.506467e-08, 2.490001e-08, 2.475253e-08, 2.453191e-08, 
    2.364568e-08, 2.208184e-08, 1.905456e-08, 1.56062e-08, 1.228536e-08, 
    8.644484e-09, 5.71486e-09, 3.482768e-09, 2.196234e-09, 1.583922e-09,
  2.528337e-08, 2.479133e-08, 2.480213e-08, 2.486796e-08, 2.44781e-08, 
    2.354389e-08, 2.206005e-08, 1.905241e-08, 1.562769e-08, 1.232269e-08, 
    8.747103e-09, 5.787609e-09, 3.583365e-09, 2.216578e-09, 1.638162e-09,
  2.534234e-08, 2.519318e-08, 2.478928e-08, 2.452633e-08, 2.427432e-08, 
    2.339197e-08, 2.190435e-08, 1.907307e-08, 1.562226e-08, 1.226963e-08, 
    8.750484e-09, 5.848283e-09, 3.649257e-09, 2.187644e-09, 1.637542e-09,
  2.515795e-08, 2.503042e-08, 2.433522e-08, 2.412142e-08, 2.381363e-08, 
    2.261753e-08, 2.129464e-08, 1.875224e-08, 1.54841e-08, 1.212328e-08, 
    8.690237e-09, 5.822709e-09, 3.668701e-09, 2.157225e-09, 1.615524e-09,
  2.495238e-08, 2.457401e-08, 2.396916e-08, 2.335793e-08, 2.313911e-08, 
    2.224371e-08, 2.096686e-08, 1.867346e-08, 1.524781e-08, 1.193949e-08, 
    8.523735e-09, 5.67699e-09, 3.653755e-09, 2.154934e-09, 1.583232e-09,
  2.457015e-08, 2.411e-08, 2.363715e-08, 2.294725e-08, 2.21269e-08, 
    2.202104e-08, 2.177366e-08, 1.945199e-08, 1.545199e-08, 1.174055e-08, 
    8.25978e-09, 5.476355e-09, 3.634043e-09, 2.198804e-09, 1.575064e-09,
  2.4747e-08, 2.414942e-08, 2.345669e-08, 2.238559e-08, 2.226477e-08, 
    2.294728e-08, 2.262002e-08, 2.026572e-08, 1.531739e-08, 1.150784e-08, 
    7.836384e-09, 5.245363e-09, 3.621611e-09, 2.269926e-09, 1.591063e-09,
  2.479123e-08, 2.422776e-08, 2.333073e-08, 2.220784e-08, 2.288996e-08, 
    2.314562e-08, 2.262566e-08, 2.014768e-08, 1.496604e-08, 1.112651e-08, 
    7.367953e-09, 5.021957e-09, 3.599111e-09, 2.342296e-09, 1.600483e-09,
  2.286865e-08, 2.364675e-08, 2.509753e-08, 2.390268e-08, 2.064251e-08, 
    1.819776e-08, 1.674201e-08, 1.438321e-08, 1.181407e-08, 8.384541e-09, 
    4.779766e-09, 2.721347e-09, 1.674764e-09, 1.260582e-09, 1.094773e-09,
  2.357659e-08, 2.322859e-08, 2.435722e-08, 2.470898e-08, 2.262067e-08, 
    1.949538e-08, 1.756203e-08, 1.554004e-08, 1.329539e-08, 1.006448e-08, 
    6.238944e-09, 3.38063e-09, 1.979874e-09, 1.364985e-09, 1.181652e-09,
  2.490689e-08, 2.349798e-08, 2.380811e-08, 2.467741e-08, 2.383458e-08, 
    2.09717e-08, 1.862649e-08, 1.655884e-08, 1.460557e-08, 1.165218e-08, 
    7.809613e-09, 4.281175e-09, 2.369881e-09, 1.503032e-09, 1.265761e-09,
  2.600259e-08, 2.411246e-08, 2.370679e-08, 2.448745e-08, 2.449877e-08, 
    2.242781e-08, 1.981402e-08, 1.740196e-08, 1.558742e-08, 1.314081e-08, 
    9.361722e-09, 5.420739e-09, 2.857515e-09, 1.691612e-09, 1.34486e-09,
  2.640648e-08, 2.497716e-08, 2.373464e-08, 2.405825e-08, 2.470363e-08, 
    2.335467e-08, 2.095498e-08, 1.852621e-08, 1.647333e-08, 1.447677e-08, 
    1.08718e-08, 6.665513e-09, 3.435157e-09, 1.89052e-09, 1.39292e-09,
  2.611792e-08, 2.507479e-08, 2.386023e-08, 2.3746e-08, 2.450679e-08, 
    2.409409e-08, 2.194058e-08, 1.935085e-08, 1.719319e-08, 1.544864e-08, 
    1.227875e-08, 7.928154e-09, 4.172332e-09, 2.105723e-09, 1.435313e-09,
  2.56924e-08, 2.559664e-08, 2.41696e-08, 2.373693e-08, 2.430814e-08, 
    2.436956e-08, 2.306156e-08, 2.080339e-08, 1.811186e-08, 1.637534e-08, 
    1.361783e-08, 9.173478e-09, 5.02453e-09, 2.328114e-09, 1.500876e-09,
  2.555733e-08, 2.575673e-08, 2.449095e-08, 2.380896e-08, 2.473917e-08, 
    2.486843e-08, 2.359711e-08, 2.134232e-08, 1.880308e-08, 1.694585e-08, 
    1.473466e-08, 1.034535e-08, 5.900768e-09, 2.588247e-09, 1.577843e-09,
  2.518498e-08, 2.569094e-08, 2.469965e-08, 2.41507e-08, 2.501138e-08, 
    2.507977e-08, 2.414925e-08, 2.180517e-08, 1.94426e-08, 1.749884e-08, 
    1.565457e-08, 1.140987e-08, 6.795821e-09, 2.88737e-09, 1.660903e-09,
  2.509148e-08, 2.55064e-08, 2.478229e-08, 2.4353e-08, 2.465437e-08, 
    2.517817e-08, 2.521154e-08, 2.267977e-08, 2.01436e-08, 1.794252e-08, 
    1.625461e-08, 1.231043e-08, 7.579324e-09, 3.247203e-09, 1.724041e-09,
  2.752415e-08, 2.678666e-08, 2.480331e-08, 2.24514e-08, 2.106641e-08, 
    2.025309e-08, 1.88013e-08, 1.502654e-08, 1.103427e-08, 6.224156e-09, 
    4.050532e-09, 2.887999e-09, 2.014362e-09, 1.318834e-09, 9.585972e-10,
  2.6673e-08, 2.757453e-08, 2.666984e-08, 2.468285e-08, 2.236707e-08, 
    2.102869e-08, 2.009956e-08, 1.74681e-08, 1.338656e-08, 8.625152e-09, 
    4.986529e-09, 3.343974e-09, 2.408611e-09, 1.551056e-09, 1.078286e-09,
  2.636999e-08, 2.691988e-08, 2.720025e-08, 2.634441e-08, 2.418746e-08, 
    2.195726e-08, 2.09557e-08, 1.931433e-08, 1.56313e-08, 1.123153e-08, 
    6.576285e-09, 3.934988e-09, 2.769705e-09, 1.876574e-09, 1.245504e-09,
  2.599319e-08, 2.563277e-08, 2.645856e-08, 2.739457e-08, 2.615507e-08, 
    2.360861e-08, 2.176987e-08, 2.063715e-08, 1.777087e-08, 1.344404e-08, 
    8.630497e-09, 4.875733e-09, 3.14673e-09, 2.20378e-09, 1.454967e-09,
  2.715764e-08, 2.563639e-08, 2.553861e-08, 2.676672e-08, 2.751942e-08, 
    2.553809e-08, 2.306223e-08, 2.159482e-08, 1.960571e-08, 1.575747e-08, 
    1.096513e-08, 6.140446e-09, 3.572226e-09, 2.454045e-09, 1.669738e-09,
  2.870266e-08, 2.633173e-08, 2.533689e-08, 2.544118e-08, 2.723434e-08, 
    2.712592e-08, 2.476435e-08, 2.250297e-08, 2.068657e-08, 1.757213e-08, 
    1.310794e-08, 7.929603e-09, 4.249256e-09, 2.664841e-09, 1.860329e-09,
  2.90023e-08, 2.858673e-08, 2.686201e-08, 2.478354e-08, 2.603172e-08, 
    2.743574e-08, 2.657134e-08, 2.444793e-08, 2.215493e-08, 1.941865e-08, 
    1.514199e-08, 1.005853e-08, 5.218762e-09, 2.97567e-09, 2.004037e-09,
  2.907222e-08, 2.956608e-08, 2.818582e-08, 2.556111e-08, 2.512349e-08, 
    2.689915e-08, 2.711124e-08, 2.547917e-08, 2.33171e-08, 2.092156e-08, 
    1.706634e-08, 1.208121e-08, 6.630575e-09, 3.484163e-09, 2.145561e-09,
  2.782888e-08, 2.896239e-08, 2.873447e-08, 2.678462e-08, 2.4946e-08, 
    2.549289e-08, 2.696863e-08, 2.632907e-08, 2.445741e-08, 2.191562e-08, 
    1.878169e-08, 1.375886e-08, 8.310935e-09, 4.199518e-09, 2.365806e-09,
  2.663896e-08, 2.826587e-08, 2.893835e-08, 2.752001e-08, 2.489982e-08, 
    2.473635e-08, 2.642907e-08, 2.699786e-08, 2.568703e-08, 2.319969e-08, 
    2.03525e-08, 1.531641e-08, 9.838082e-09, 4.992143e-09, 2.690267e-09,
  2.57889e-08, 2.644026e-08, 2.618198e-08, 2.35634e-08, 2.12487e-08, 
    1.788033e-08, 1.412105e-08, 1.056677e-08, 7.073898e-09, 4.345925e-09, 
    3.316984e-09, 2.628769e-09, 2.092792e-09, 1.527677e-09, 1.03193e-09,
  2.540196e-08, 2.594153e-08, 2.666564e-08, 2.5223e-08, 2.254412e-08, 
    2.001736e-08, 1.634968e-08, 1.261449e-08, 8.830613e-09, 5.454081e-09, 
    3.721558e-09, 2.846067e-09, 2.213186e-09, 1.64563e-09, 1.094293e-09,
  2.528153e-08, 2.562217e-08, 2.611719e-08, 2.598534e-08, 2.395462e-08, 
    2.135247e-08, 1.8254e-08, 1.477022e-08, 1.076072e-08, 6.974024e-09, 
    4.368408e-09, 3.146787e-09, 2.415118e-09, 1.822409e-09, 1.240906e-09,
  2.550575e-08, 2.532828e-08, 2.53178e-08, 2.589354e-08, 2.509824e-08, 
    2.262391e-08, 2.006021e-08, 1.670811e-08, 1.285269e-08, 8.646138e-09, 
    5.350625e-09, 3.625559e-09, 2.690394e-09, 2.007106e-09, 1.408139e-09,
  2.553284e-08, 2.541117e-08, 2.498818e-08, 2.534924e-08, 2.565163e-08, 
    2.387723e-08, 2.116296e-08, 1.856527e-08, 1.505833e-08, 1.065901e-08, 
    6.677455e-09, 4.187919e-09, 3.02131e-09, 2.20678e-09, 1.586985e-09,
  2.606657e-08, 2.533295e-08, 2.500492e-08, 2.494235e-08, 2.574747e-08, 
    2.501199e-08, 2.250852e-08, 1.986895e-08, 1.679761e-08, 1.283622e-08, 
    8.482934e-09, 5.046791e-09, 3.441003e-09, 2.464033e-09, 1.750715e-09,
  2.589657e-08, 2.571926e-08, 2.550428e-08, 2.494751e-08, 2.518965e-08, 
    2.557498e-08, 2.393605e-08, 2.147116e-08, 1.873665e-08, 1.484022e-08, 
    1.05663e-08, 6.403107e-09, 4.017002e-09, 2.794662e-09, 1.926527e-09,
  2.471625e-08, 2.590128e-08, 2.60611e-08, 2.54549e-08, 2.499851e-08, 
    2.541314e-08, 2.470002e-08, 2.24347e-08, 2.006438e-08, 1.678834e-08, 
    1.266907e-08, 8.267498e-09, 4.813566e-09, 3.248969e-09, 2.131715e-09,
  2.41269e-08, 2.603842e-08, 2.655419e-08, 2.605118e-08, 2.557329e-08, 
    2.526432e-08, 2.508612e-08, 2.314821e-08, 2.102195e-08, 1.825829e-08, 
    1.44628e-08, 1.030274e-08, 5.965094e-09, 3.784842e-09, 2.405104e-09,
  2.331533e-08, 2.505348e-08, 2.599316e-08, 2.613268e-08, 2.588172e-08, 
    2.577815e-08, 2.559344e-08, 2.388691e-08, 2.196334e-08, 1.957969e-08, 
    1.6113e-08, 1.204383e-08, 7.592134e-09, 4.470659e-09, 2.761525e-09,
  2.283962e-08, 2.407923e-08, 2.429216e-08, 2.372814e-08, 2.220815e-08, 
    2.08905e-08, 1.873381e-08, 1.533913e-08, 1.153829e-08, 8.461391e-09, 
    5.937154e-09, 4.014176e-09, 2.317105e-09, 1.410221e-09, 9.316802e-10,
  2.215291e-08, 2.374303e-08, 2.446676e-08, 2.401337e-08, 2.262249e-08, 
    2.134042e-08, 1.940887e-08, 1.63504e-08, 1.241684e-08, 9.179264e-09, 
    6.360051e-09, 4.267094e-09, 2.520839e-09, 1.487635e-09, 9.867827e-10,
  2.194503e-08, 2.313166e-08, 2.427616e-08, 2.402164e-08, 2.318334e-08, 
    2.190716e-08, 2.007524e-08, 1.731597e-08, 1.347342e-08, 9.817588e-09, 
    6.841854e-09, 4.561797e-09, 2.723729e-09, 1.595791e-09, 1.064194e-09,
  2.185491e-08, 2.266306e-08, 2.387499e-08, 2.415176e-08, 2.3575e-08, 
    2.250739e-08, 2.07642e-08, 1.811161e-08, 1.443507e-08, 1.051061e-08, 
    7.340117e-09, 4.882078e-09, 2.931413e-09, 1.707018e-09, 1.121108e-09,
  2.264935e-08, 2.262072e-08, 2.347966e-08, 2.42781e-08, 2.391501e-08, 
    2.30114e-08, 2.153314e-08, 1.908736e-08, 1.550279e-08, 1.124243e-08, 
    7.74944e-09, 5.189124e-09, 3.135123e-09, 1.812822e-09, 1.172439e-09,
  2.290088e-08, 2.256003e-08, 2.3232e-08, 2.430429e-08, 2.431951e-08, 
    2.354715e-08, 2.217188e-08, 1.971823e-08, 1.643985e-08, 1.222202e-08, 
    8.171195e-09, 5.433036e-09, 3.323689e-09, 1.881325e-09, 1.233868e-09,
  2.32899e-08, 2.277075e-08, 2.31082e-08, 2.446059e-08, 2.453877e-08, 
    2.369839e-08, 2.293786e-08, 2.076852e-08, 1.749615e-08, 1.326137e-08, 
    8.785865e-09, 5.635703e-09, 3.468352e-09, 1.996191e-09, 1.301417e-09,
  2.411549e-08, 2.314185e-08, 2.319549e-08, 2.42798e-08, 2.458858e-08, 
    2.392667e-08, 2.339313e-08, 2.171731e-08, 1.860351e-08, 1.433446e-08, 
    9.602415e-09, 5.932907e-09, 3.571035e-09, 2.095678e-09, 1.382453e-09,
  2.534384e-08, 2.37333e-08, 2.314816e-08, 2.356892e-08, 2.424131e-08, 
    2.461498e-08, 2.429392e-08, 2.267509e-08, 1.947278e-08, 1.538328e-08, 
    1.054724e-08, 6.310878e-09, 3.694432e-09, 2.181253e-09, 1.461835e-09,
  2.576715e-08, 2.411527e-08, 2.300506e-08, 2.333986e-08, 2.469782e-08, 
    2.506781e-08, 2.440898e-08, 2.315562e-08, 2.016029e-08, 1.637418e-08, 
    1.15344e-08, 6.839408e-09, 3.866766e-09, 2.2496e-09, 1.554239e-09,
  2.264971e-08, 2.287414e-08, 2.291807e-08, 2.210146e-08, 1.914296e-08, 
    1.8615e-08, 1.896067e-08, 1.723854e-08, 1.636752e-08, 1.562553e-08, 
    1.433615e-08, 1.060253e-08, 6.511821e-09, 4.107098e-09, 2.365298e-09,
  2.383559e-08, 2.370118e-08, 2.324407e-08, 2.321495e-08, 2.163267e-08, 
    1.937267e-08, 1.936064e-08, 1.846607e-08, 1.721829e-08, 1.615802e-08, 
    1.559859e-08, 1.254307e-08, 8.228278e-09, 5.024873e-09, 2.861823e-09,
  2.420404e-08, 2.37454e-08, 2.373808e-08, 2.388994e-08, 2.361603e-08, 
    2.105139e-08, 1.997574e-08, 1.922956e-08, 1.825895e-08, 1.672887e-08, 
    1.632364e-08, 1.414553e-08, 1.005797e-08, 6.097711e-09, 3.470007e-09,
  2.483653e-08, 2.392244e-08, 2.31264e-08, 2.404162e-08, 2.468892e-08, 
    2.321501e-08, 2.111755e-08, 2.015916e-08, 1.904255e-08, 1.758456e-08, 
    1.665339e-08, 1.58103e-08, 1.165745e-08, 7.358084e-09, 4.186135e-09,
  2.430483e-08, 2.481008e-08, 2.438356e-08, 2.378657e-08, 2.479833e-08, 
    2.493284e-08, 2.286588e-08, 2.12098e-08, 2.032583e-08, 1.869949e-08, 
    1.719267e-08, 1.672245e-08, 1.317412e-08, 8.688237e-09, 4.92923e-09,
  2.459717e-08, 2.367554e-08, 2.446636e-08, 2.421602e-08, 2.418928e-08, 
    2.542317e-08, 2.465243e-08, 2.244087e-08, 2.092456e-08, 1.985226e-08, 
    1.79152e-08, 1.735257e-08, 1.48408e-08, 9.928164e-09, 5.760606e-09,
  2.515992e-08, 2.460516e-08, 2.414655e-08, 2.432001e-08, 2.390277e-08, 
    2.463225e-08, 2.553302e-08, 2.440922e-08, 2.257914e-08, 2.111735e-08, 
    1.886767e-08, 1.766092e-08, 1.627883e-08, 1.105969e-08, 6.595382e-09,
  2.627389e-08, 2.548467e-08, 2.474403e-08, 2.386451e-08, 2.397912e-08, 
    2.399676e-08, 2.509523e-08, 2.516424e-08, 2.401399e-08, 2.219999e-08, 
    2.014396e-08, 1.809696e-08, 1.723603e-08, 1.227908e-08, 7.434015e-09,
  2.626615e-08, 2.53589e-08, 2.462964e-08, 2.454508e-08, 2.366906e-08, 
    2.358783e-08, 2.406912e-08, 2.493831e-08, 2.466367e-08, 2.306131e-08, 
    2.124387e-08, 1.868896e-08, 1.774997e-08, 1.351757e-08, 8.211602e-09,
  2.641937e-08, 2.590099e-08, 2.473762e-08, 2.479541e-08, 2.402226e-08, 
    2.364519e-08, 2.373624e-08, 2.424433e-08, 2.43031e-08, 2.418043e-08, 
    2.258888e-08, 1.955972e-08, 1.778394e-08, 1.45296e-08, 8.916481e-09,
  1.896836e-08, 1.80153e-08, 1.645341e-08, 1.617535e-08, 1.637248e-08, 
    1.566346e-08, 1.489261e-08, 1.34026e-08, 1.116749e-08, 8.836007e-09, 
    7.18428e-09, 5.335007e-09, 4.168204e-09, 3.61651e-09, 2.621327e-09,
  2.000973e-08, 1.927725e-08, 1.779514e-08, 1.608575e-08, 1.63084e-08, 
    1.619321e-08, 1.574153e-08, 1.462844e-08, 1.271136e-08, 1.022023e-08, 
    8.235194e-09, 6.432268e-09, 4.753872e-09, 4.048272e-09, 3.005462e-09,
  1.964083e-08, 2.04068e-08, 1.938589e-08, 1.719862e-08, 1.615484e-08, 
    1.624795e-08, 1.605713e-08, 1.552439e-08, 1.414102e-08, 1.170834e-08, 
    9.435581e-09, 7.552368e-09, 5.632048e-09, 4.579129e-09, 3.436746e-09,
  1.930894e-08, 2.098924e-08, 2.061178e-08, 1.890999e-08, 1.67253e-08, 
    1.628925e-08, 1.611884e-08, 1.60492e-08, 1.517752e-08, 1.314915e-08, 
    1.070631e-08, 8.712185e-09, 6.625882e-09, 5.259863e-09, 4.01445e-09,
  2.143722e-08, 2.140387e-08, 2.135785e-08, 2.058494e-08, 1.866964e-08, 
    1.664359e-08, 1.60798e-08, 1.594143e-08, 1.600713e-08, 1.460721e-08, 
    1.219762e-08, 9.975814e-09, 7.708079e-09, 6.088229e-09, 4.695708e-09,
  2.365945e-08, 2.186633e-08, 2.118434e-08, 2.101089e-08, 2.009754e-08, 
    1.866176e-08, 1.696137e-08, 1.589618e-08, 1.588004e-08, 1.5452e-08, 
    1.371523e-08, 1.137543e-08, 8.906122e-09, 6.965064e-09, 5.508579e-09,
  2.454251e-08, 2.311955e-08, 2.153054e-08, 2.109197e-08, 2.102394e-08, 
    1.974617e-08, 1.84599e-08, 1.714139e-08, 1.626828e-08, 1.595271e-08, 
    1.474132e-08, 1.290009e-08, 1.026166e-08, 7.880599e-09, 6.362077e-09,
  2.726304e-08, 2.56637e-08, 2.346048e-08, 2.162681e-08, 2.172323e-08, 
    2.113612e-08, 1.936419e-08, 1.754215e-08, 1.657079e-08, 1.639901e-08, 
    1.561786e-08, 1.41699e-08, 1.175241e-08, 8.917807e-09, 7.162135e-09,
  2.856352e-08, 2.761706e-08, 2.544071e-08, 2.337104e-08, 2.215412e-08, 
    2.203373e-08, 2.073502e-08, 1.864089e-08, 1.706951e-08, 1.656669e-08, 
    1.612358e-08, 1.508727e-08, 1.327563e-08, 1.00952e-08, 7.94478e-09,
  2.829985e-08, 2.863946e-08, 2.711885e-08, 2.518195e-08, 2.364812e-08, 
    2.279326e-08, 2.198158e-08, 2.018393e-08, 1.838207e-08, 1.728171e-08, 
    1.666897e-08, 1.574563e-08, 1.45695e-08, 1.153605e-08, 8.812983e-09,
  1.828208e-08, 1.627403e-08, 1.539486e-08, 1.363342e-08, 1.292754e-08, 
    1.215156e-08, 1.116671e-08, 1.056908e-08, 9.724519e-09, 8.307651e-09, 
    6.169198e-09, 4.048105e-09, 3.038714e-09, 2.399272e-09, 1.915927e-09,
  1.864588e-08, 1.778641e-08, 1.593922e-08, 1.451065e-08, 1.345089e-08, 
    1.2906e-08, 1.169231e-08, 1.065214e-08, 1.007096e-08, 8.946892e-09, 
    7.087677e-09, 4.697383e-09, 3.347218e-09, 2.590959e-09, 2.012518e-09,
  1.840217e-08, 1.895651e-08, 1.730472e-08, 1.513408e-08, 1.38871e-08, 
    1.362928e-08, 1.230738e-08, 1.093005e-08, 1.022429e-08, 9.49085e-09, 
    7.93542e-09, 5.546905e-09, 3.783995e-09, 2.812496e-09, 2.116735e-09,
  1.791732e-08, 1.897326e-08, 1.852024e-08, 1.615165e-08, 1.44952e-08, 
    1.418031e-08, 1.324133e-08, 1.145643e-08, 1.029257e-08, 9.894615e-09, 
    8.602516e-09, 6.42966e-09, 4.337503e-09, 3.079807e-09, 2.283052e-09,
  2.085621e-08, 1.902992e-08, 1.868538e-08, 1.722442e-08, 1.518269e-08, 
    1.433066e-08, 1.415048e-08, 1.237982e-08, 1.063549e-08, 1.00717e-08, 
    9.191007e-09, 7.301697e-09, 5.073217e-09, 3.442127e-09, 2.532342e-09,
  2.323966e-08, 1.90161e-08, 1.83893e-08, 1.791374e-08, 1.621759e-08, 
    1.500694e-08, 1.465751e-08, 1.340595e-08, 1.125793e-08, 1.021384e-08, 
    9.675881e-09, 8.05051e-09, 5.903093e-09, 3.899889e-09, 2.812502e-09,
  2.373083e-08, 1.857117e-08, 1.714924e-08, 1.770485e-08, 1.764266e-08, 
    1.588429e-08, 1.521499e-08, 1.472027e-08, 1.22957e-08, 1.049468e-08, 
    1.007368e-08, 8.739603e-09, 6.737781e-09, 4.539784e-09, 3.128343e-09,
  2.550295e-08, 1.947545e-08, 1.607505e-08, 1.628127e-08, 1.902381e-08, 
    1.748495e-08, 1.583542e-08, 1.524802e-08, 1.351894e-08, 1.118299e-08, 
    1.02774e-08, 9.363476e-09, 7.507963e-09, 5.285244e-09, 3.528839e-09,
  2.941659e-08, 2.231839e-08, 1.685198e-08, 1.51498e-08, 1.853933e-08, 
    1.943994e-08, 1.647653e-08, 1.525451e-08, 1.449226e-08, 1.247983e-08, 
    1.077518e-08, 9.82751e-09, 8.220412e-09, 6.114826e-09, 4.023991e-09,
  3.271598e-08, 2.401225e-08, 1.87123e-08, 1.495735e-08, 1.677697e-08, 
    1.999505e-08, 1.867154e-08, 1.607628e-08, 1.555778e-08, 1.370115e-08, 
    1.139653e-08, 1.024267e-08, 8.822274e-09, 6.948224e-09, 4.662411e-09,
  2.288401e-08, 1.982525e-08, 1.73326e-08, 1.490253e-08, 1.313382e-08, 
    1.177109e-08, 1.075266e-08, 9.360418e-09, 7.569765e-09, 5.898762e-09, 
    4.863481e-09, 3.736456e-09, 2.691846e-09, 2.041725e-09, 1.513301e-09,
  2.40831e-08, 2.158725e-08, 1.864895e-08, 1.602035e-08, 1.369442e-08, 
    1.216404e-08, 1.102398e-08, 9.951259e-09, 8.293022e-09, 6.480358e-09, 
    5.262955e-09, 4.282488e-09, 3.02885e-09, 2.286944e-09, 1.671167e-09,
  2.462446e-08, 2.310888e-08, 2.005214e-08, 1.703098e-08, 1.425623e-08, 
    1.2487e-08, 1.130176e-08, 1.038622e-08, 9.035748e-09, 7.15719e-09, 
    5.703459e-09, 4.711916e-09, 3.413095e-09, 2.551198e-09, 1.855352e-09,
  2.497285e-08, 2.345015e-08, 2.146426e-08, 1.833337e-08, 1.528553e-08, 
    1.305198e-08, 1.160097e-08, 1.067843e-08, 9.575641e-09, 7.849857e-09, 
    6.215287e-09, 5.099635e-09, 3.863464e-09, 2.830162e-09, 2.067405e-09,
  2.594137e-08, 2.447733e-08, 2.222092e-08, 1.992482e-08, 1.662973e-08, 
    1.367791e-08, 1.206821e-08, 1.109358e-08, 1.020634e-08, 8.545606e-09, 
    6.810304e-09, 5.437797e-09, 4.339486e-09, 3.134708e-09, 2.306933e-09,
  2.576918e-08, 2.442916e-08, 2.269541e-08, 2.100434e-08, 1.814439e-08, 
    1.47741e-08, 1.251872e-08, 1.133356e-08, 1.052489e-08, 9.17658e-09, 
    7.516346e-09, 5.860428e-09, 4.756435e-09, 3.473471e-09, 2.576034e-09,
  2.604849e-08, 2.426306e-08, 2.295015e-08, 2.179562e-08, 1.924723e-08, 
    1.582771e-08, 1.328677e-08, 1.185421e-08, 1.095472e-08, 9.760029e-09, 
    8.154229e-09, 6.406647e-09, 5.132904e-09, 3.858753e-09, 2.863808e-09,
  2.667947e-08, 2.464446e-08, 2.329783e-08, 2.21264e-08, 2.063483e-08, 
    1.725347e-08, 1.43663e-08, 1.260992e-08, 1.134216e-08, 1.017256e-08, 
    8.745916e-09, 7.013166e-09, 5.533832e-09, 4.255379e-09, 3.174716e-09,
  2.713437e-08, 2.510359e-08, 2.350631e-08, 2.215099e-08, 2.118696e-08, 
    1.842798e-08, 1.512104e-08, 1.282377e-08, 1.162647e-08, 1.062689e-08, 
    9.166889e-09, 7.590732e-09, 6.024286e-09, 4.661211e-09, 3.495116e-09,
  2.733651e-08, 2.56917e-08, 2.349212e-08, 2.233305e-08, 2.174137e-08, 
    1.933645e-08, 1.555911e-08, 1.267732e-08, 1.166248e-08, 1.088511e-08, 
    9.506466e-09, 8.110221e-09, 6.534895e-09, 5.088893e-09, 3.832696e-09,
  2.504034e-08, 2.569193e-08, 2.526292e-08, 2.34775e-08, 2.094271e-08, 
    1.874277e-08, 1.579463e-08, 1.201943e-08, 8.960947e-09, 6.447945e-09, 
    4.156682e-09, 2.35882e-09, 1.422255e-09, 1.094397e-09, 9.359704e-10,
  2.46375e-08, 2.606759e-08, 2.625282e-08, 2.510274e-08, 2.263756e-08, 
    2.005597e-08, 1.716023e-08, 1.348076e-08, 1.007423e-08, 7.269274e-09, 
    4.930816e-09, 2.873682e-09, 1.696549e-09, 1.18355e-09, 9.111601e-10,
  2.421432e-08, 2.501231e-08, 2.644945e-08, 2.593022e-08, 2.436952e-08, 
    2.133076e-08, 1.852106e-08, 1.500342e-08, 1.120218e-08, 8.070675e-09, 
    5.640399e-09, 3.411598e-09, 1.996801e-09, 1.3086e-09, 9.027821e-10,
  2.479912e-08, 2.421273e-08, 2.572158e-08, 2.665896e-08, 2.550354e-08, 
    2.320867e-08, 1.99875e-08, 1.648383e-08, 1.250552e-08, 8.993095e-09, 
    6.333039e-09, 3.992512e-09, 2.35411e-09, 1.489585e-09, 9.385415e-10,
  2.530332e-08, 2.44755e-08, 2.493048e-08, 2.657412e-08, 2.627486e-08, 
    2.448765e-08, 2.156588e-08, 1.814243e-08, 1.390318e-08, 9.979042e-09, 
    7.041987e-09, 4.589126e-09, 2.747129e-09, 1.728116e-09, 1.019811e-09,
  2.505518e-08, 2.437329e-08, 2.407173e-08, 2.587759e-08, 2.654481e-08, 
    2.576442e-08, 2.299314e-08, 1.948064e-08, 1.53924e-08, 1.106821e-08, 
    7.768187e-09, 5.192198e-09, 3.16167e-09, 2.006546e-09, 1.152484e-09,
  2.699005e-08, 2.540865e-08, 2.397886e-08, 2.5205e-08, 2.639857e-08, 
    2.626336e-08, 2.481879e-08, 2.137769e-08, 1.681487e-08, 1.223387e-08, 
    8.561585e-09, 5.775626e-09, 3.576069e-09, 2.307327e-09, 1.340079e-09,
  2.828711e-08, 2.670763e-08, 2.470643e-08, 2.432908e-08, 2.63602e-08, 
    2.687653e-08, 2.563565e-08, 2.310146e-08, 1.845841e-08, 1.344204e-08, 
    9.381128e-09, 6.392767e-09, 3.991719e-09, 2.59729e-09, 1.571098e-09,
  2.81559e-08, 2.78e-08, 2.571887e-08, 2.410768e-08, 2.579183e-08, 
    2.691752e-08, 2.600306e-08, 2.344348e-08, 1.99911e-08, 1.496934e-08, 
    1.030021e-08, 7.029395e-09, 4.411078e-09, 2.872034e-09, 1.815512e-09,
  2.805197e-08, 2.820691e-08, 2.704428e-08, 2.462962e-08, 2.503879e-08, 
    2.668738e-08, 2.680433e-08, 2.442057e-08, 2.109568e-08, 1.627278e-08, 
    1.127652e-08, 7.720582e-09, 4.852387e-09, 3.142167e-09, 2.050598e-09,
  2.499217e-08, 2.416035e-08, 2.418621e-08, 2.460801e-08, 2.583127e-08, 
    2.617937e-08, 2.531813e-08, 2.37874e-08, 2.212558e-08, 1.851383e-08, 
    1.468121e-08, 1.000421e-08, 5.908817e-09, 3.036095e-09, 1.099832e-09,
  2.580451e-08, 2.500453e-08, 2.422323e-08, 2.400004e-08, 2.495773e-08, 
    2.642894e-08, 2.601076e-08, 2.460065e-08, 2.313161e-08, 1.997565e-08, 
    1.620603e-08, 1.139467e-08, 6.823725e-09, 3.651382e-09, 1.39388e-09,
  2.582067e-08, 2.495819e-08, 2.439221e-08, 2.387505e-08, 2.431469e-08, 
    2.578182e-08, 2.643043e-08, 2.5159e-08, 2.40442e-08, 2.129286e-08, 
    1.742442e-08, 1.276205e-08, 7.770601e-09, 4.285806e-09, 1.710488e-09,
  2.646927e-08, 2.50744e-08, 2.487191e-08, 2.388811e-08, 2.367798e-08, 
    2.510555e-08, 2.681699e-08, 2.564093e-08, 2.445888e-08, 2.247621e-08, 
    1.854751e-08, 1.403097e-08, 8.707199e-09, 4.877773e-09, 2.047548e-09,
  2.712338e-08, 2.575945e-08, 2.498853e-08, 2.4459e-08, 2.374094e-08, 
    2.40176e-08, 2.629837e-08, 2.673876e-08, 2.506291e-08, 2.335238e-08, 
    1.957487e-08, 1.512457e-08, 9.592466e-09, 5.429115e-09, 2.375437e-09,
  2.608247e-08, 2.504269e-08, 2.508324e-08, 2.459125e-08, 2.382086e-08, 
    2.395293e-08, 2.554928e-08, 2.637106e-08, 2.534963e-08, 2.387881e-08, 
    2.047169e-08, 1.605905e-08, 1.03996e-08, 5.90917e-09, 2.654959e-09,
  2.729508e-08, 2.605934e-08, 2.553365e-08, 2.523548e-08, 2.401125e-08, 
    2.340789e-08, 2.550957e-08, 2.76351e-08, 2.617834e-08, 2.441992e-08, 
    2.112189e-08, 1.677874e-08, 1.109697e-08, 6.32829e-09, 2.898392e-09,
  2.784809e-08, 2.667717e-08, 2.57412e-08, 2.528933e-08, 2.491418e-08, 
    2.367391e-08, 2.425562e-08, 2.674249e-08, 2.658381e-08, 2.476036e-08, 
    2.170054e-08, 1.739599e-08, 1.170142e-08, 6.652137e-09, 3.086666e-09,
  2.760945e-08, 2.718683e-08, 2.612665e-08, 2.608769e-08, 2.511663e-08, 
    2.339758e-08, 2.383066e-08, 2.603698e-08, 2.660864e-08, 2.516109e-08, 
    2.219724e-08, 1.785001e-08, 1.21315e-08, 6.895396e-09, 3.213151e-09,
  2.722133e-08, 2.741215e-08, 2.636903e-08, 2.63636e-08, 2.560815e-08, 
    2.380554e-08, 2.352374e-08, 2.566768e-08, 2.677769e-08, 2.552228e-08, 
    2.257559e-08, 1.819119e-08, 1.2439e-08, 7.06422e-09, 3.269822e-09,
  2.529622e-08, 2.413966e-08, 2.408707e-08, 2.479674e-08, 2.547051e-08, 
    2.609851e-08, 2.597129e-08, 2.566839e-08, 2.402873e-08, 2.043365e-08, 
    1.559416e-08, 1.097128e-08, 7.433137e-09, 4.695872e-09, 2.611411e-09,
  2.633916e-08, 2.562555e-08, 2.436354e-08, 2.432632e-08, 2.515907e-08, 
    2.597631e-08, 2.64687e-08, 2.608941e-08, 2.50621e-08, 2.237358e-08, 
    1.783715e-08, 1.279388e-08, 8.657303e-09, 5.538575e-09, 3.18401e-09,
  2.71022e-08, 2.616703e-08, 2.50006e-08, 2.387993e-08, 2.457306e-08, 
    2.564564e-08, 2.624346e-08, 2.630346e-08, 2.552967e-08, 2.376944e-08, 
    1.974011e-08, 1.461724e-08, 9.915154e-09, 6.390303e-09, 3.735341e-09,
  2.776257e-08, 2.670721e-08, 2.568609e-08, 2.434993e-08, 2.404814e-08, 
    2.53124e-08, 2.619748e-08, 2.637158e-08, 2.584607e-08, 2.478395e-08, 
    2.138383e-08, 1.637217e-08, 1.114328e-08, 7.223406e-09, 4.236932e-09,
  2.650565e-08, 2.734866e-08, 2.660749e-08, 2.495912e-08, 2.390403e-08, 
    2.447022e-08, 2.590896e-08, 2.652016e-08, 2.60623e-08, 2.536624e-08, 
    2.258613e-08, 1.790068e-08, 1.234386e-08, 7.994885e-09, 4.69905e-09,
  2.542057e-08, 2.614929e-08, 2.685383e-08, 2.593016e-08, 2.429005e-08, 
    2.431272e-08, 2.553626e-08, 2.634531e-08, 2.610751e-08, 2.568206e-08, 
    2.365509e-08, 1.914658e-08, 1.342523e-08, 8.657266e-09, 5.089857e-09,
  2.61151e-08, 2.618003e-08, 2.688333e-08, 2.681364e-08, 2.474082e-08, 
    2.377153e-08, 2.573474e-08, 2.685771e-08, 2.617054e-08, 2.568543e-08, 
    2.424022e-08, 2.00395e-08, 1.436288e-08, 9.242612e-09, 5.411068e-09,
  2.63491e-08, 2.612823e-08, 2.672314e-08, 2.682383e-08, 2.616193e-08, 
    2.395671e-08, 2.494659e-08, 2.719201e-08, 2.638234e-08, 2.562585e-08, 
    2.474611e-08, 2.073464e-08, 1.503738e-08, 9.65441e-09, 5.605835e-09,
  2.632424e-08, 2.607717e-08, 2.643371e-08, 2.736693e-08, 2.634856e-08, 
    2.4302e-08, 2.438894e-08, 2.60636e-08, 2.658897e-08, 2.569106e-08, 
    2.495846e-08, 2.117294e-08, 1.550458e-08, 9.952872e-09, 5.688981e-09,
  2.660479e-08, 2.620506e-08, 2.613226e-08, 2.738719e-08, 2.645597e-08, 
    2.477079e-08, 2.422755e-08, 2.61356e-08, 2.662471e-08, 2.565284e-08, 
    2.510948e-08, 2.145969e-08, 1.573343e-08, 1.000429e-08, 5.642977e-09,
  2.667729e-08, 2.611027e-08, 2.587194e-08, 2.486059e-08, 2.494026e-08, 
    2.524924e-08, 2.409802e-08, 2.18922e-08, 1.861743e-08, 1.601311e-08, 
    1.344693e-08, 9.993092e-09, 6.789015e-09, 4.661982e-09, 3.598057e-09,
  2.634876e-08, 2.631745e-08, 2.622294e-08, 2.551249e-08, 2.495932e-08, 
    2.513562e-08, 2.490876e-08, 2.357399e-08, 2.071293e-08, 1.765693e-08, 
    1.498617e-08, 1.155009e-08, 8.139351e-09, 5.29372e-09, 3.943578e-09,
  2.703542e-08, 2.603494e-08, 2.609062e-08, 2.605355e-08, 2.532795e-08, 
    2.494273e-08, 2.510222e-08, 2.468467e-08, 2.265647e-08, 1.941876e-08, 
    1.661986e-08, 1.313389e-08, 9.468899e-09, 6.206861e-09, 4.296858e-09,
  2.899849e-08, 2.605573e-08, 2.581174e-08, 2.62569e-08, 2.580482e-08, 
    2.524928e-08, 2.50773e-08, 2.511191e-08, 2.40259e-08, 2.11299e-08, 
    1.798115e-08, 1.465099e-08, 1.082045e-08, 7.207347e-09, 4.712276e-09,
  2.763733e-08, 2.749897e-08, 2.672772e-08, 2.631908e-08, 2.63067e-08, 
    2.546134e-08, 2.51165e-08, 2.534496e-08, 2.521563e-08, 2.28466e-08, 
    1.943373e-08, 1.592237e-08, 1.201965e-08, 8.194054e-09, 5.220825e-09,
  2.684343e-08, 2.662131e-08, 2.676057e-08, 2.696586e-08, 2.641591e-08, 
    2.625695e-08, 2.528516e-08, 2.514352e-08, 2.549524e-08, 2.413851e-08, 
    2.093283e-08, 1.7141e-08, 1.315192e-08, 9.138266e-09, 5.790808e-09,
  2.78117e-08, 2.844777e-08, 2.811126e-08, 2.767059e-08, 2.748113e-08, 
    2.624765e-08, 2.624876e-08, 2.578567e-08, 2.61062e-08, 2.52503e-08, 
    2.22215e-08, 1.83239e-08, 1.4103e-08, 9.965364e-09, 6.335164e-09,
  2.78165e-08, 2.866989e-08, 2.871604e-08, 2.797806e-08, 2.883969e-08, 
    2.735111e-08, 2.636322e-08, 2.529768e-08, 2.555187e-08, 2.568335e-08, 
    2.337135e-08, 1.943125e-08, 1.495469e-08, 1.065944e-08, 6.825059e-09,
  2.696146e-08, 2.796967e-08, 2.840873e-08, 2.922655e-08, 2.984991e-08, 
    2.745747e-08, 2.617293e-08, 2.53122e-08, 2.577628e-08, 2.62205e-08, 
    2.433094e-08, 2.03951e-08, 1.572697e-08, 1.12025e-08, 7.174247e-09,
  2.674638e-08, 2.780786e-08, 2.779779e-08, 2.929129e-08, 2.951485e-08, 
    2.897443e-08, 2.687241e-08, 2.553439e-08, 2.595741e-08, 2.641126e-08, 
    2.500981e-08, 2.118543e-08, 1.637547e-08, 1.159794e-08, 7.421233e-09,
  2.554235e-08, 2.449118e-08, 2.386509e-08, 2.313514e-08, 2.291033e-08, 
    2.240166e-08, 2.125357e-08, 1.963026e-08, 1.765047e-08, 1.537361e-08, 
    1.320389e-08, 1.055486e-08, 8.144428e-09, 6.080105e-09, 4.466189e-09,
  2.587672e-08, 2.56509e-08, 2.439741e-08, 2.374125e-08, 2.30163e-08, 
    2.274258e-08, 2.214656e-08, 2.085901e-08, 1.899888e-08, 1.680979e-08, 
    1.476175e-08, 1.216231e-08, 9.369671e-09, 7.024836e-09, 5.224663e-09,
  2.526222e-08, 2.585105e-08, 2.513642e-08, 2.412792e-08, 2.356209e-08, 
    2.280682e-08, 2.232306e-08, 2.157312e-08, 2.017929e-08, 1.810205e-08, 
    1.609094e-08, 1.364297e-08, 1.079156e-08, 8.004942e-09, 5.98392e-09,
  2.51306e-08, 2.529798e-08, 2.571203e-08, 2.50745e-08, 2.409962e-08, 
    2.377774e-08, 2.284135e-08, 2.198016e-08, 2.076043e-08, 1.90155e-08, 
    1.721707e-08, 1.491562e-08, 1.225472e-08, 9.0878e-09, 6.764649e-09,
  2.423239e-08, 2.565183e-08, 2.586381e-08, 2.563302e-08, 2.466349e-08, 
    2.35813e-08, 2.337763e-08, 2.275846e-08, 2.177429e-08, 1.996269e-08, 
    1.816253e-08, 1.606826e-08, 1.357544e-08, 1.027131e-08, 7.553047e-09,
  2.332172e-08, 2.417592e-08, 2.591221e-08, 2.613271e-08, 2.549376e-08, 
    2.455053e-08, 2.360701e-08, 2.272229e-08, 2.187871e-08, 2.067752e-08, 
    1.89542e-08, 1.706646e-08, 1.468584e-08, 1.147965e-08, 8.37925e-09,
  2.52293e-08, 2.419653e-08, 2.515296e-08, 2.629699e-08, 2.563699e-08, 
    2.4712e-08, 2.414129e-08, 2.392544e-08, 2.293962e-08, 2.147274e-08, 
    1.963734e-08, 1.790679e-08, 1.562783e-08, 1.258354e-08, 9.193223e-09,
  2.527504e-08, 2.467531e-08, 2.456115e-08, 2.57198e-08, 2.68788e-08, 
    2.584685e-08, 2.476441e-08, 2.429405e-08, 2.311269e-08, 2.186769e-08, 
    2.023577e-08, 1.849432e-08, 1.650903e-08, 1.352647e-08, 1.003028e-08,
  2.427536e-08, 2.478023e-08, 2.4426e-08, 2.577172e-08, 2.698013e-08, 
    2.538566e-08, 2.47162e-08, 2.39717e-08, 2.366771e-08, 2.252547e-08, 
    2.083652e-08, 1.898206e-08, 1.71045e-08, 1.433242e-08, 1.079993e-08,
  2.411769e-08, 2.413007e-08, 2.477933e-08, 2.515091e-08, 2.678138e-08, 
    2.648796e-08, 2.459369e-08, 2.38781e-08, 2.39712e-08, 2.302644e-08, 
    2.135934e-08, 1.934185e-08, 1.75909e-08, 1.500362e-08, 1.147543e-08,
  1.500704e-08, 1.343327e-08, 1.21959e-08, 1.10216e-08, 1.009835e-08, 
    9.061839e-09, 7.844134e-09, 6.478428e-09, 5.048936e-09, 4.350735e-09, 
    4.177098e-09, 4.232391e-09, 4.044074e-09, 3.883232e-09, 3.314435e-09,
  1.540375e-08, 1.408874e-08, 1.292718e-08, 1.167076e-08, 1.066254e-08, 
    9.797942e-09, 8.835094e-09, 7.639468e-09, 6.188978e-09, 4.810891e-09, 
    4.461883e-09, 4.564941e-09, 4.41556e-09, 4.141633e-09, 3.772715e-09,
  1.601436e-08, 1.483275e-08, 1.3849e-08, 1.258106e-08, 1.14456e-08, 
    1.050824e-08, 9.690122e-09, 8.657468e-09, 7.371834e-09, 5.889528e-09, 
    5.006531e-09, 4.906429e-09, 4.667261e-09, 4.429445e-09, 4.176171e-09,
  1.710558e-08, 1.569257e-08, 1.451664e-08, 1.339577e-08, 1.233996e-08, 
    1.128632e-08, 1.042119e-08, 9.548787e-09, 8.448681e-09, 7.092751e-09, 
    6.001161e-09, 5.380247e-09, 5.033736e-09, 4.774941e-09, 4.429459e-09,
  1.855777e-08, 1.694241e-08, 1.550518e-08, 1.4245e-08, 1.320152e-08, 
    1.216425e-08, 1.12217e-08, 1.032039e-08, 9.445203e-09, 8.270748e-09, 
    7.168456e-09, 6.267539e-09, 5.461211e-09, 5.080997e-09, 4.790242e-09,
  1.993106e-08, 1.808787e-08, 1.632381e-08, 1.495168e-08, 1.400892e-08, 
    1.318592e-08, 1.223586e-08, 1.107569e-08, 1.016142e-08, 9.34144e-09, 
    8.208058e-09, 7.497748e-09, 6.2736e-09, 5.469005e-09, 5.312744e-09,
  2.051294e-08, 1.93101e-08, 1.72835e-08, 1.584158e-08, 1.467168e-08, 
    1.397329e-08, 1.311657e-08, 1.216216e-08, 1.124458e-08, 1.04042e-08, 
    9.311924e-09, 8.479738e-09, 7.422015e-09, 6.12602e-09, 5.872446e-09,
  2.078962e-08, 2.020762e-08, 1.867528e-08, 1.691116e-08, 1.566216e-08, 
    1.49001e-08, 1.422345e-08, 1.338573e-08, 1.265137e-08, 1.165366e-08, 
    1.047182e-08, 9.558418e-09, 8.546897e-09, 7.080631e-09, 6.492573e-09,
  2.143967e-08, 2.097288e-08, 1.981434e-08, 1.802454e-08, 1.672982e-08, 
    1.628811e-08, 1.56938e-08, 1.465999e-08, 1.345886e-08, 1.249368e-08, 
    1.172394e-08, 1.063388e-08, 9.710281e-09, 8.246633e-09, 7.052211e-09,
  2.200244e-08, 2.147198e-08, 2.068709e-08, 1.92372e-08, 1.802941e-08, 
    1.766311e-08, 1.668296e-08, 1.567627e-08, 1.437135e-08, 1.347666e-08, 
    1.282834e-08, 1.188167e-08, 1.088068e-08, 9.514296e-09, 7.918292e-09,
  2.38817e-08, 2.335647e-08, 2.331692e-08, 2.222882e-08, 1.945498e-08, 
    1.787456e-08, 1.682168e-08, 1.534505e-08, 1.340284e-08, 1.087848e-08, 
    7.917362e-09, 5.366765e-09, 3.436579e-09, 2.084585e-09, 1.634715e-09,
  2.351106e-08, 2.30319e-08, 2.295933e-08, 2.206252e-08, 2.027311e-08, 
    1.788719e-08, 1.689606e-08, 1.564514e-08, 1.374687e-08, 1.131289e-08, 
    8.382581e-09, 5.761894e-09, 3.770743e-09, 2.312496e-09, 1.761673e-09,
  2.288304e-08, 2.21531e-08, 2.263453e-08, 2.164386e-08, 2.056397e-08, 
    1.824931e-08, 1.689126e-08, 1.570772e-08, 1.402629e-08, 1.163133e-08, 
    8.700014e-09, 6.073603e-09, 4.059999e-09, 2.515699e-09, 1.875192e-09,
  2.227905e-08, 2.178067e-08, 2.238091e-08, 2.143094e-08, 2.059892e-08, 
    1.857589e-08, 1.699036e-08, 1.58181e-08, 1.410255e-08, 1.182389e-08, 
    8.936271e-09, 6.31728e-09, 4.295082e-09, 2.720044e-09, 2.021769e-09,
  2.266946e-08, 2.2372e-08, 2.276392e-08, 2.127763e-08, 2.039043e-08, 
    1.865276e-08, 1.696854e-08, 1.579171e-08, 1.424852e-08, 1.187427e-08, 
    9.07044e-09, 6.466424e-09, 4.482933e-09, 2.916977e-09, 2.155589e-09,
  2.41692e-08, 2.317674e-08, 2.280166e-08, 2.13889e-08, 1.983437e-08, 
    1.870053e-08, 1.711869e-08, 1.561404e-08, 1.411008e-08, 1.190538e-08, 
    9.087742e-09, 6.518877e-09, 4.614471e-09, 3.081461e-09, 2.281589e-09,
  2.350035e-08, 2.251369e-08, 2.198794e-08, 2.129155e-08, 1.898301e-08, 
    1.806863e-08, 1.712997e-08, 1.59011e-08, 1.420786e-08, 1.191058e-08, 
    9.117862e-09, 6.507793e-09, 4.685035e-09, 3.239711e-09, 2.404981e-09,
  2.27439e-08, 2.177783e-08, 2.156662e-08, 2.108487e-08, 1.829375e-08, 
    1.777858e-08, 1.694164e-08, 1.535609e-08, 1.400329e-08, 1.17891e-08, 
    8.98379e-09, 6.427814e-09, 4.719165e-09, 3.346185e-09, 2.498258e-09,
  2.371679e-08, 2.175422e-08, 2.13568e-08, 2.084668e-08, 1.760772e-08, 
    1.674074e-08, 1.62296e-08, 1.497633e-08, 1.381568e-08, 1.167676e-08, 
    8.894327e-09, 6.328602e-09, 4.661062e-09, 3.367294e-09, 2.556671e-09,
  2.2911e-08, 2.14662e-08, 2.113649e-08, 2.057979e-08, 1.833448e-08, 
    1.637607e-08, 1.539988e-08, 1.454143e-08, 1.348398e-08, 1.148037e-08, 
    8.785417e-09, 6.208201e-09, 4.536172e-09, 3.329625e-09, 2.566915e-09,
  2.64141e-08, 2.647152e-08, 2.743233e-08, 2.760633e-08, 2.352126e-08, 
    2.06414e-08, 1.915407e-08, 1.686308e-08, 1.453853e-08, 1.11158e-08, 
    7.476199e-09, 4.685781e-09, 2.911845e-09, 1.870045e-09, 1.21305e-09,
  2.679964e-08, 2.663868e-08, 2.608802e-08, 2.735947e-08, 2.597668e-08, 
    2.265002e-08, 2.039228e-08, 1.829797e-08, 1.596231e-08, 1.300337e-08, 
    9.179838e-09, 5.869746e-09, 3.455717e-09, 2.168594e-09, 1.383559e-09,
  2.730795e-08, 2.687444e-08, 2.640766e-08, 2.626747e-08, 2.672443e-08, 
    2.445922e-08, 2.194392e-08, 1.97737e-08, 1.747809e-08, 1.473878e-08, 
    1.107637e-08, 7.237415e-09, 4.185183e-09, 2.513468e-09, 1.59724e-09,
  2.777557e-08, 2.632216e-08, 2.629417e-08, 2.651101e-08, 2.638233e-08, 
    2.573505e-08, 2.385378e-08, 2.131639e-08, 1.888554e-08, 1.610331e-08, 
    1.287601e-08, 8.836753e-09, 5.194936e-09, 2.935224e-09, 1.836761e-09,
  2.680176e-08, 2.663386e-08, 2.59382e-08, 2.667011e-08, 2.684779e-08, 
    2.611726e-08, 2.528439e-08, 2.382965e-08, 2.091319e-08, 1.766064e-08, 
    1.444694e-08, 1.051183e-08, 6.451487e-09, 3.515413e-09, 2.120223e-09,
  2.549388e-08, 2.567957e-08, 2.612149e-08, 2.634437e-08, 2.699429e-08, 
    2.676472e-08, 2.589595e-08, 2.499119e-08, 2.26593e-08, 1.935755e-08, 
    1.588595e-08, 1.218601e-08, 7.884744e-09, 4.23551e-09, 2.498985e-09,
  2.540049e-08, 2.544987e-08, 2.584372e-08, 2.606e-08, 2.672297e-08, 
    2.704152e-08, 2.729145e-08, 2.729211e-08, 2.498781e-08, 2.118149e-08, 
    1.734358e-08, 1.359189e-08, 9.454943e-09, 5.161712e-09, 2.978058e-09,
  2.522927e-08, 2.560052e-08, 2.560009e-08, 2.552102e-08, 2.627622e-08, 
    2.697759e-08, 2.680792e-08, 2.761825e-08, 2.758832e-08, 2.366918e-08, 
    1.906717e-08, 1.494887e-08, 1.090504e-08, 6.271168e-09, 3.535037e-09,
  2.464365e-08, 2.496357e-08, 2.534726e-08, 2.565698e-08, 2.588681e-08, 
    2.61862e-08, 2.708157e-08, 2.635461e-08, 2.706137e-08, 2.504502e-08, 
    2.08529e-08, 1.635499e-08, 1.227963e-08, 7.480343e-09, 4.180533e-09,
  2.447696e-08, 2.461669e-08, 2.526845e-08, 2.565865e-08, 2.528317e-08, 
    2.501695e-08, 2.716818e-08, 2.693073e-08, 2.65253e-08, 2.632881e-08, 
    2.335349e-08, 1.786872e-08, 1.35063e-08, 8.711833e-09, 4.903106e-09,
  2.214114e-08, 2.145165e-08, 1.980004e-08, 1.725267e-08, 1.400895e-08, 
    1.147113e-08, 9.418029e-09, 9.052917e-09, 8.712237e-09, 8.589731e-09, 
    7.99416e-09, 6.49128e-09, 4.140188e-09, 2.289902e-09, 1.467833e-09,
  2.224218e-08, 2.253223e-08, 2.120002e-08, 1.861422e-08, 1.576318e-08, 
    1.29632e-08, 1.058702e-08, 9.526997e-09, 8.857897e-09, 8.602837e-09, 
    8.572022e-09, 7.139346e-09, 4.916385e-09, 2.843894e-09, 1.632252e-09,
  2.261974e-08, 2.348401e-08, 2.261157e-08, 2.023361e-08, 1.763532e-08, 
    1.477267e-08, 1.180462e-08, 1.018464e-08, 9.240559e-09, 8.795199e-09, 
    8.864915e-09, 7.900175e-09, 5.713732e-09, 3.455368e-09, 1.939255e-09,
  2.416082e-08, 2.490177e-08, 2.423966e-08, 2.172464e-08, 1.943269e-08, 
    1.684403e-08, 1.356477e-08, 1.103465e-08, 9.70658e-09, 8.76231e-09, 
    8.756138e-09, 8.675949e-09, 6.434964e-09, 4.110376e-09, 2.38033e-09,
  2.852863e-08, 2.630634e-08, 2.538595e-08, 2.332869e-08, 2.082494e-08, 
    1.878016e-08, 1.553376e-08, 1.238882e-08, 1.046243e-08, 9.029569e-09, 
    8.418369e-09, 9.089267e-09, 7.238002e-09, 4.917089e-09, 2.916978e-09,
  3.02182e-08, 2.848592e-08, 2.622354e-08, 2.429529e-08, 2.249784e-08, 
    2.064372e-08, 1.790922e-08, 1.387838e-08, 1.122585e-08, 9.718547e-09, 
    8.481863e-09, 9.07547e-09, 8.056817e-09, 5.777103e-09, 3.530424e-09,
  2.822595e-08, 2.831271e-08, 2.742482e-08, 2.535172e-08, 2.312312e-08, 
    2.170678e-08, 1.960323e-08, 1.61535e-08, 1.27839e-08, 1.061607e-08, 
    9.057573e-09, 9.075769e-09, 8.872182e-09, 6.620953e-09, 4.222511e-09,
  2.897184e-08, 2.908366e-08, 2.772875e-08, 2.708138e-08, 2.425806e-08, 
    2.277985e-08, 2.122171e-08, 1.851691e-08, 1.538947e-08, 1.225519e-08, 
    9.985757e-09, 9.267049e-09, 9.436379e-09, 7.4201e-09, 4.99278e-09,
  2.931519e-08, 3.005643e-08, 2.866608e-08, 2.665397e-08, 2.576004e-08, 
    2.532793e-08, 2.403945e-08, 2.071013e-08, 1.698093e-08, 1.39811e-08, 
    1.142943e-08, 9.794393e-09, 9.800235e-09, 8.129972e-09, 5.731967e-09,
  2.935039e-08, 3.013439e-08, 2.969443e-08, 2.784561e-08, 2.631025e-08, 
    2.673276e-08, 2.605599e-08, 2.253743e-08, 1.88506e-08, 1.586235e-08, 
    1.328259e-08, 1.083468e-08, 1.002276e-08, 8.819748e-09, 6.507631e-09,
  1.969035e-08, 1.770539e-08, 1.572467e-08, 1.735148e-08, 1.921659e-08, 
    2.034226e-08, 2.04018e-08, 1.891953e-08, 1.718556e-08, 1.570839e-08, 
    1.338178e-08, 9.740151e-09, 5.315408e-09, 2.394384e-09, 1.287291e-09,
  1.896214e-08, 1.709118e-08, 1.572365e-08, 1.540383e-08, 1.797572e-08, 
    1.963289e-08, 2.004569e-08, 1.856199e-08, 1.688832e-08, 1.536526e-08, 
    1.332073e-08, 1.019318e-08, 5.828898e-09, 2.709587e-09, 1.422678e-09,
  1.886253e-08, 1.700591e-08, 1.521008e-08, 1.424468e-08, 1.669352e-08, 
    1.865788e-08, 1.98835e-08, 1.792914e-08, 1.674225e-08, 1.52855e-08, 
    1.307643e-08, 1.018015e-08, 6.145801e-09, 2.899539e-09, 1.473442e-09,
  1.916827e-08, 1.727729e-08, 1.495338e-08, 1.434297e-08, 1.543046e-08, 
    1.752322e-08, 1.910684e-08, 1.770204e-08, 1.607805e-08, 1.53447e-08, 
    1.305536e-08, 1.007973e-08, 6.196991e-09, 3.034563e-09, 1.526729e-09,
  2.075051e-08, 1.902725e-08, 1.519722e-08, 1.445273e-08, 1.398242e-08, 
    1.62413e-08, 1.819416e-08, 1.746699e-08, 1.58339e-08, 1.516525e-08, 
    1.313718e-08, 9.94539e-09, 6.138578e-09, 3.086065e-09, 1.592071e-09,
  2.254659e-08, 2.110462e-08, 1.569588e-08, 1.418627e-08, 1.279005e-08, 
    1.491274e-08, 1.734456e-08, 1.754307e-08, 1.532528e-08, 1.465759e-08, 
    1.305473e-08, 9.81958e-09, 6.074539e-09, 3.138122e-09, 1.669547e-09,
  2.163579e-08, 2.04105e-08, 1.611165e-08, 1.381885e-08, 1.227431e-08, 
    1.338335e-08, 1.589552e-08, 1.692413e-08, 1.56351e-08, 1.408243e-08, 
    1.255863e-08, 9.623574e-09, 6.035235e-09, 3.232721e-09, 1.757383e-09,
  2.25104e-08, 2.056271e-08, 1.70409e-08, 1.344968e-08, 1.230006e-08, 
    1.256598e-08, 1.491987e-08, 1.687593e-08, 1.595586e-08, 1.385303e-08, 
    1.182586e-08, 9.104916e-09, 5.950633e-09, 3.358842e-09, 1.915917e-09,
  2.477295e-08, 2.204241e-08, 1.853466e-08, 1.345402e-08, 1.195642e-08, 
    1.306527e-08, 1.423696e-08, 1.577116e-08, 1.532546e-08, 1.377087e-08, 
    1.128619e-08, 8.530313e-09, 5.900074e-09, 3.604849e-09, 2.12683e-09,
  2.734848e-08, 2.244132e-08, 1.950212e-08, 1.442234e-08, 1.32058e-08, 
    1.432513e-08, 1.346225e-08, 1.494851e-08, 1.474219e-08, 1.359791e-08, 
    1.093994e-08, 8.187538e-09, 5.86901e-09, 3.939221e-09, 2.436483e-09,
  2.162593e-08, 2.17356e-08, 2.10066e-08, 2.063556e-08, 2.165204e-08, 
    2.215488e-08, 2.174836e-08, 2.049838e-08, 1.93222e-08, 1.87132e-08, 
    1.691902e-08, 1.51694e-08, 1.210902e-08, 8.355007e-09, 4.074574e-09,
  2.222528e-08, 2.217615e-08, 2.213885e-08, 2.121735e-08, 2.079728e-08, 
    2.142884e-08, 2.219596e-08, 2.200394e-08, 2.095805e-08, 1.980551e-08, 
    1.858227e-08, 1.751724e-08, 1.466341e-08, 1.116463e-08, 6.353238e-09,
  2.50413e-08, 2.382542e-08, 2.294299e-08, 2.173768e-08, 2.140481e-08, 
    2.131476e-08, 2.202636e-08, 2.236852e-08, 2.210158e-08, 2.127091e-08, 
    1.969802e-08, 1.915111e-08, 1.710499e-08, 1.359428e-08, 8.790791e-09,
  2.712391e-08, 2.596066e-08, 2.49771e-08, 2.319646e-08, 2.225209e-08, 
    2.216444e-08, 2.22735e-08, 2.297699e-08, 2.230783e-08, 2.238908e-08, 
    2.12361e-08, 2.062698e-08, 1.888479e-08, 1.599273e-08, 1.126528e-08,
  2.723558e-08, 2.782376e-08, 2.782176e-08, 2.574073e-08, 2.421115e-08, 
    2.311404e-08, 2.276112e-08, 2.280563e-08, 2.296315e-08, 2.249467e-08, 
    2.243879e-08, 2.205529e-08, 2.058132e-08, 1.795201e-08, 1.354908e-08,
  2.555375e-08, 2.562749e-08, 2.749697e-08, 2.829602e-08, 2.688515e-08, 
    2.575703e-08, 2.411657e-08, 2.301288e-08, 2.301185e-08, 2.383357e-08, 
    2.343379e-08, 2.36596e-08, 2.206269e-08, 1.945357e-08, 1.562716e-08,
  2.451463e-08, 2.509621e-08, 2.619391e-08, 2.73841e-08, 2.814032e-08, 
    2.773348e-08, 2.665721e-08, 2.654645e-08, 2.497218e-08, 2.475799e-08, 
    2.443829e-08, 2.51823e-08, 2.331109e-08, 2.065857e-08, 1.716701e-08,
  2.593791e-08, 2.570823e-08, 2.608272e-08, 2.639581e-08, 2.732385e-08, 
    2.747201e-08, 2.701984e-08, 2.585377e-08, 2.47851e-08, 2.48546e-08, 
    2.558424e-08, 2.613103e-08, 2.504498e-08, 2.153616e-08, 1.860526e-08,
  2.46134e-08, 2.545494e-08, 2.575887e-08, 2.666194e-08, 2.742967e-08, 
    2.705685e-08, 2.632817e-08, 2.555346e-08, 2.536114e-08, 2.562132e-08, 
    2.584591e-08, 2.672996e-08, 2.599256e-08, 2.280239e-08, 1.950364e-08,
  2.298316e-08, 2.364662e-08, 2.435874e-08, 2.582039e-08, 2.607021e-08, 
    2.640716e-08, 2.66381e-08, 2.635204e-08, 2.705008e-08, 2.681302e-08, 
    2.567632e-08, 2.610315e-08, 2.585359e-08, 2.367157e-08, 2.039121e-08,
  1.910246e-08, 1.803106e-08, 1.759973e-08, 1.645888e-08, 1.507983e-08, 
    1.392178e-08, 1.236226e-08, 1.015653e-08, 7.971289e-09, 5.951566e-09, 
    3.86712e-09, 3.020328e-09, 3.307946e-09, 4.129174e-09, 3.344849e-09,
  1.954296e-08, 1.854761e-08, 1.804223e-08, 1.699707e-08, 1.55688e-08, 
    1.450783e-08, 1.338844e-08, 1.175333e-08, 9.532805e-09, 7.551643e-09, 
    5.346609e-09, 3.971449e-09, 3.340067e-09, 3.344863e-09, 3.880609e-09,
  1.972727e-08, 1.970715e-08, 1.897253e-08, 1.757209e-08, 1.608903e-08, 
    1.493263e-08, 1.397866e-08, 1.289173e-08, 1.109366e-08, 9.153399e-09, 
    7.010232e-09, 5.095499e-09, 4.084074e-09, 3.597996e-09, 3.601034e-09,
  1.914111e-08, 2.009692e-08, 1.979482e-08, 1.865749e-08, 1.704008e-08, 
    1.556959e-08, 1.442997e-08, 1.361827e-08, 1.22815e-08, 1.059726e-08, 
    8.761619e-09, 6.658881e-09, 5.000301e-09, 4.179497e-09, 3.735046e-09,
  1.933183e-08, 1.960344e-08, 1.951214e-08, 1.90144e-08, 1.804001e-08, 
    1.659653e-08, 1.516021e-08, 1.413106e-08, 1.328644e-08, 1.193717e-08, 
    1.028577e-08, 8.449533e-09, 6.469859e-09, 4.981565e-09, 4.124322e-09,
  1.93404e-08, 1.951797e-08, 1.90984e-08, 1.890904e-08, 1.850292e-08, 
    1.77511e-08, 1.648201e-08, 1.507214e-08, 1.385318e-08, 1.316624e-08, 
    1.168892e-08, 9.985984e-09, 8.201262e-09, 6.3288e-09, 4.928077e-09,
  1.816697e-08, 1.879655e-08, 1.915643e-08, 1.923825e-08, 1.909464e-08, 
    1.8826e-08, 1.779249e-08, 1.677168e-08, 1.537454e-08, 1.405234e-08, 
    1.274729e-08, 1.148735e-08, 9.831871e-09, 7.98612e-09, 6.162471e-09,
  1.903224e-08, 1.891425e-08, 1.917974e-08, 1.95757e-08, 2.021744e-08, 
    1.985087e-08, 1.862877e-08, 1.761572e-08, 1.624803e-08, 1.452705e-08, 
    1.358414e-08, 1.250738e-08, 1.12255e-08, 9.706311e-09, 7.740249e-09,
  1.99265e-08, 1.969618e-08, 1.968723e-08, 2.009868e-08, 2.088917e-08, 
    2.053268e-08, 1.977459e-08, 1.826166e-08, 1.717056e-08, 1.589355e-08, 
    1.451382e-08, 1.331216e-08, 1.218381e-08, 1.103812e-08, 9.441804e-09,
  2.144214e-08, 2.114161e-08, 2.087565e-08, 2.107567e-08, 2.140191e-08, 
    2.170635e-08, 2.106532e-08, 1.994567e-08, 1.887245e-08, 1.761202e-08, 
    1.587666e-08, 1.441451e-08, 1.304889e-08, 1.200681e-08, 1.085011e-08,
  2.431512e-08, 2.503455e-08, 2.453015e-08, 2.297579e-08, 2.15432e-08, 
    1.902548e-08, 1.608048e-08, 1.315847e-08, 1.010096e-08, 6.270918e-09, 
    3.305176e-09, 1.842386e-09, 1.225957e-09, 8.673314e-10, 5.295147e-10,
  2.392876e-08, 2.494565e-08, 2.494571e-08, 2.374238e-08, 2.220301e-08, 
    2.019639e-08, 1.710028e-08, 1.425289e-08, 1.164539e-08, 8.037589e-09, 
    4.505092e-09, 2.304825e-09, 1.196569e-09, 9.161095e-10, 6.884952e-10,
  2.357984e-08, 2.458671e-08, 2.506607e-08, 2.428824e-08, 2.27511e-08, 
    2.113503e-08, 1.809732e-08, 1.518121e-08, 1.281125e-08, 9.885567e-09, 
    6.22297e-09, 3.242175e-09, 1.211797e-09, 8.161917e-10, 7.401584e-10,
  2.342078e-08, 2.397763e-08, 2.499367e-08, 2.470292e-08, 2.334949e-08, 
    2.194805e-08, 1.921806e-08, 1.608725e-08, 1.370487e-08, 1.146178e-08, 
    8.107361e-09, 4.698804e-09, 1.779659e-09, 7.807235e-10, 6.309313e-10,
  2.354514e-08, 2.370367e-08, 2.450609e-08, 2.500293e-08, 2.37748e-08, 
    2.228609e-08, 2.028507e-08, 1.723707e-08, 1.470142e-08, 1.276568e-08, 
    9.703453e-09, 6.481287e-09, 2.873782e-09, 9.771463e-10, 4.409217e-10,
  2.360363e-08, 2.354366e-08, 2.405775e-08, 2.476314e-08, 2.449231e-08, 
    2.314718e-08, 2.133255e-08, 1.839771e-08, 1.573095e-08, 1.365675e-08, 
    1.114593e-08, 7.921692e-09, 4.65259e-09, 1.684385e-09, 3.451772e-10,
  2.360973e-08, 2.34469e-08, 2.359122e-08, 2.446457e-08, 2.426962e-08, 
    2.34584e-08, 2.223723e-08, 1.992604e-08, 1.732838e-08, 1.480073e-08, 
    1.238102e-08, 9.285338e-09, 6.402197e-09, 2.969514e-09, 6.286253e-10,
  2.344933e-08, 2.332399e-08, 2.324658e-08, 2.382898e-08, 2.456323e-08, 
    2.400614e-08, 2.27737e-08, 2.117119e-08, 1.859079e-08, 1.579686e-08, 
    1.334357e-08, 1.081675e-08, 8.030979e-09, 4.882556e-09, 1.418974e-09,
  2.378357e-08, 2.351774e-08, 2.330793e-08, 2.340698e-08, 2.411737e-08, 
    2.430999e-08, 2.349773e-08, 2.20791e-08, 1.903734e-08, 1.627111e-08, 
    1.385443e-08, 1.201223e-08, 9.549007e-09, 6.793777e-09, 2.949938e-09,
  2.373062e-08, 2.357317e-08, 2.332221e-08, 2.343416e-08, 2.390583e-08, 
    2.434037e-08, 2.373103e-08, 2.256281e-08, 2.017335e-08, 1.714611e-08, 
    1.458709e-08, 1.284053e-08, 1.080238e-08, 8.294093e-09, 4.980108e-09,
  2.513044e-08, 2.626442e-08, 2.651292e-08, 2.566889e-08, 2.398697e-08, 
    2.088805e-08, 1.844326e-08, 1.596718e-08, 1.426525e-08, 1.225924e-08, 
    9.432362e-09, 7.25888e-09, 4.798545e-09, 3.121118e-09, 1.985928e-09,
  2.508018e-08, 2.601335e-08, 2.66046e-08, 2.592263e-08, 2.457634e-08, 
    2.190532e-08, 1.935816e-08, 1.665476e-08, 1.464908e-08, 1.310345e-08, 
    1.022641e-08, 7.808656e-09, 5.444766e-09, 3.536411e-09, 2.142585e-09,
  2.525238e-08, 2.600616e-08, 2.676324e-08, 2.60996e-08, 2.476408e-08, 
    2.256535e-08, 2.011713e-08, 1.751052e-08, 1.52026e-08, 1.377938e-08, 
    1.125763e-08, 8.442935e-09, 6.034585e-09, 3.9412e-09, 2.329409e-09,
  2.546374e-08, 2.621588e-08, 2.657511e-08, 2.624484e-08, 2.50676e-08, 
    2.315376e-08, 2.086082e-08, 1.832991e-08, 1.58273e-08, 1.429619e-08, 
    1.222449e-08, 9.224232e-09, 6.610085e-09, 4.36666e-09, 2.613468e-09,
  2.66977e-08, 2.644674e-08, 2.622979e-08, 2.627423e-08, 2.537472e-08, 
    2.360519e-08, 2.149813e-08, 1.929757e-08, 1.663201e-08, 1.478451e-08, 
    1.305777e-08, 1.001148e-08, 7.106421e-09, 4.775305e-09, 2.906162e-09,
  2.760891e-08, 2.659161e-08, 2.593312e-08, 2.564363e-08, 2.567777e-08, 
    2.441832e-08, 2.208575e-08, 2.001368e-08, 1.733612e-08, 1.517293e-08, 
    1.375822e-08, 1.095132e-08, 7.720272e-09, 5.248788e-09, 3.236009e-09,
  2.682446e-08, 2.617814e-08, 2.557353e-08, 2.540313e-08, 2.524824e-08, 
    2.459202e-08, 2.25104e-08, 2.10162e-08, 1.860737e-08, 1.590445e-08, 
    1.444434e-08, 1.172639e-08, 8.412978e-09, 5.703185e-09, 3.582856e-09,
  2.669929e-08, 2.612431e-08, 2.56024e-08, 2.490965e-08, 2.51535e-08, 
    2.466043e-08, 2.241013e-08, 2.148938e-08, 1.980529e-08, 1.665191e-08, 
    1.488623e-08, 1.23561e-08, 9.225079e-09, 6.213737e-09, 3.931186e-09,
  2.733512e-08, 2.695799e-08, 2.591135e-08, 2.419846e-08, 2.442837e-08, 
    2.524858e-08, 2.360021e-08, 2.214271e-08, 2.057714e-08, 1.728587e-08, 
    1.52919e-08, 1.292866e-08, 9.970673e-09, 6.816397e-09, 4.330762e-09,
  2.769799e-08, 2.74973e-08, 2.647611e-08, 2.410655e-08, 2.397328e-08, 
    2.49589e-08, 2.428582e-08, 2.300582e-08, 2.131664e-08, 1.801395e-08, 
    1.58589e-08, 1.351537e-08, 1.066356e-08, 7.548307e-09, 4.846819e-09,
  2.822324e-08, 2.986584e-08, 3.204457e-08, 3.231858e-08, 2.807509e-08, 
    2.585736e-08, 2.571478e-08, 2.185304e-08, 1.831172e-08, 1.635204e-08, 
    1.454935e-08, 1.204406e-08, 1.007461e-08, 7.794449e-09, 5.666863e-09,
  2.754952e-08, 3.075723e-08, 3.277364e-08, 3.417841e-08, 2.985131e-08, 
    2.58995e-08, 2.546773e-08, 2.288758e-08, 1.908565e-08, 1.663947e-08, 
    1.472541e-08, 1.24688e-08, 1.07096e-08, 8.54415e-09, 6.085675e-09,
  2.726564e-08, 3.080024e-08, 3.331208e-08, 3.441188e-08, 3.081428e-08, 
    2.580781e-08, 2.487294e-08, 2.382344e-08, 2.028991e-08, 1.700611e-08, 
    1.476249e-08, 1.313826e-08, 1.142307e-08, 9.200671e-09, 6.589783e-09,
  2.680976e-08, 3.070682e-08, 3.335207e-08, 3.394301e-08, 3.240991e-08, 
    2.685484e-08, 2.4804e-08, 2.46272e-08, 2.157646e-08, 1.735862e-08, 
    1.485657e-08, 1.375003e-08, 1.217528e-08, 9.839606e-09, 7.063234e-09,
  2.712518e-08, 3.022796e-08, 3.344789e-08, 3.425124e-08, 3.373927e-08, 
    2.790639e-08, 2.475144e-08, 2.482127e-08, 2.240779e-08, 1.803632e-08, 
    1.502313e-08, 1.446954e-08, 1.294549e-08, 1.053597e-08, 7.563816e-09,
  2.724401e-08, 2.954786e-08, 3.299266e-08, 3.401092e-08, 3.457185e-08, 
    2.945053e-08, 2.496494e-08, 2.381829e-08, 2.176126e-08, 1.832386e-08, 
    1.570786e-08, 1.520903e-08, 1.35012e-08, 1.119172e-08, 8.038587e-09,
  2.708946e-08, 2.857455e-08, 3.228204e-08, 3.345377e-08, 3.46841e-08, 
    3.028323e-08, 2.507713e-08, 2.306952e-08, 2.11791e-08, 1.894973e-08, 
    1.673499e-08, 1.603568e-08, 1.401737e-08, 1.175576e-08, 8.554861e-09,
  2.696396e-08, 2.794573e-08, 3.195248e-08, 3.306497e-08, 3.390752e-08, 
    3.130338e-08, 2.578294e-08, 2.298149e-08, 2.094902e-08, 1.971503e-08, 
    1.764398e-08, 1.669782e-08, 1.441866e-08, 1.219043e-08, 9.074448e-09,
  2.691787e-08, 2.781145e-08, 3.119229e-08, 3.194813e-08, 3.234456e-08, 
    3.434443e-08, 2.716195e-08, 2.290562e-08, 1.996193e-08, 1.918862e-08, 
    1.789053e-08, 1.712298e-08, 1.47273e-08, 1.261186e-08, 9.542971e-09,
  2.703637e-08, 2.770349e-08, 3.063496e-08, 3.141926e-08, 3.137913e-08, 
    3.404464e-08, 2.782998e-08, 2.291172e-08, 1.989323e-08, 1.859663e-08, 
    1.812664e-08, 1.683145e-08, 1.484327e-08, 1.289734e-08, 9.96798e-09,
  2.666822e-08, 2.643164e-08, 2.6094e-08, 2.607372e-08, 2.599234e-08, 
    2.437722e-08, 2.38e-08, 2.372911e-08, 2.301425e-08, 2.168622e-08, 
    1.962071e-08, 1.563684e-08, 1.221271e-08, 9.62318e-09, 7.367719e-09,
  2.731278e-08, 2.69766e-08, 2.629824e-08, 2.628629e-08, 2.668271e-08, 
    2.597375e-08, 2.451499e-08, 2.383141e-08, 2.347138e-08, 2.219211e-08, 
    2.038497e-08, 1.690429e-08, 1.304929e-08, 1.022783e-08, 7.804281e-09,
  2.730649e-08, 2.734999e-08, 2.67976e-08, 2.641957e-08, 2.685938e-08, 
    2.67079e-08, 2.53691e-08, 2.425979e-08, 2.369861e-08, 2.272767e-08, 
    2.104242e-08, 1.809394e-08, 1.403075e-08, 1.084694e-08, 8.287404e-09,
  2.724229e-08, 2.702846e-08, 2.707858e-08, 2.679212e-08, 2.685942e-08, 
    2.69895e-08, 2.621284e-08, 2.492362e-08, 2.384489e-08, 2.319856e-08, 
    2.159015e-08, 1.907958e-08, 1.512317e-08, 1.152431e-08, 8.808883e-09,
  2.668395e-08, 2.705143e-08, 2.726809e-08, 2.728213e-08, 2.721064e-08, 
    2.692157e-08, 2.660366e-08, 2.562192e-08, 2.456206e-08, 2.360977e-08, 
    2.249488e-08, 1.983913e-08, 1.627472e-08, 1.227975e-08, 9.382627e-09,
  2.530481e-08, 2.600149e-08, 2.72187e-08, 2.749646e-08, 2.767497e-08, 
    2.696524e-08, 2.68354e-08, 2.632353e-08, 2.51438e-08, 2.368787e-08, 
    2.28372e-08, 2.054854e-08, 1.72745e-08, 1.305094e-08, 9.900119e-09,
  2.56408e-08, 2.610924e-08, 2.700635e-08, 2.762271e-08, 2.791783e-08, 
    2.70599e-08, 2.699564e-08, 2.728228e-08, 2.605927e-08, 2.385935e-08, 
    2.31165e-08, 2.128038e-08, 1.811063e-08, 1.388014e-08, 1.042183e-08,
  2.678663e-08, 2.671757e-08, 2.742046e-08, 2.742625e-08, 2.849052e-08, 
    2.799909e-08, 2.774926e-08, 2.814041e-08, 2.644685e-08, 2.383277e-08, 
    2.296888e-08, 2.187393e-08, 1.887831e-08, 1.488089e-08, 1.096214e-08,
  2.734241e-08, 2.730784e-08, 2.7577e-08, 2.737053e-08, 2.873252e-08, 
    2.972083e-08, 2.834543e-08, 2.840334e-08, 2.643239e-08, 2.327239e-08, 
    2.284367e-08, 2.293242e-08, 1.960809e-08, 1.597803e-08, 1.167188e-08,
  2.767915e-08, 2.803475e-08, 2.815449e-08, 2.674825e-08, 2.830143e-08, 
    3.181478e-08, 2.788552e-08, 2.757777e-08, 2.595465e-08, 2.296254e-08, 
    2.266681e-08, 2.395228e-08, 2.054672e-08, 1.685028e-08, 1.247683e-08,
  2.412443e-08, 2.120132e-08, 2.021196e-08, 1.802506e-08, 1.71692e-08, 
    1.631932e-08, 1.603685e-08, 1.615641e-08, 1.716518e-08, 1.699217e-08, 
    1.548651e-08, 1.331217e-08, 1.117696e-08, 9.325277e-09, 7.593913e-09,
  2.784038e-08, 2.329082e-08, 2.113195e-08, 1.907034e-08, 1.754922e-08, 
    1.672074e-08, 1.633255e-08, 1.639642e-08, 1.713658e-08, 1.758198e-08, 
    1.656121e-08, 1.458593e-08, 1.218293e-08, 1.006954e-08, 8.383415e-09,
  2.972873e-08, 2.556287e-08, 2.275444e-08, 2.065408e-08, 1.83485e-08, 
    1.708998e-08, 1.669414e-08, 1.660419e-08, 1.703623e-08, 1.78061e-08, 
    1.744885e-08, 1.582257e-08, 1.344835e-08, 1.093282e-08, 9.074687e-09,
  2.835581e-08, 2.781515e-08, 2.473837e-08, 2.150992e-08, 1.925796e-08, 
    1.778662e-08, 1.712683e-08, 1.678505e-08, 1.704739e-08, 1.761877e-08, 
    1.792498e-08, 1.697532e-08, 1.468597e-08, 1.203732e-08, 9.771499e-09,
  2.887564e-08, 2.85792e-08, 2.56649e-08, 2.213712e-08, 1.950389e-08, 
    1.85225e-08, 1.753404e-08, 1.712106e-08, 1.717398e-08, 1.76226e-08, 
    1.797242e-08, 1.783156e-08, 1.602012e-08, 1.339267e-08, 1.064175e-08,
  2.811921e-08, 2.766741e-08, 2.552091e-08, 2.258771e-08, 1.972571e-08, 
    1.893249e-08, 1.850389e-08, 1.773489e-08, 1.729535e-08, 1.744424e-08, 
    1.796289e-08, 1.807445e-08, 1.713888e-08, 1.485214e-08, 1.169588e-08,
  2.683512e-08, 2.687119e-08, 2.548498e-08, 2.329401e-08, 2.030279e-08, 
    1.892602e-08, 1.894398e-08, 1.873902e-08, 1.796055e-08, 1.75981e-08, 
    1.802598e-08, 1.810553e-08, 1.790836e-08, 1.624951e-08, 1.303797e-08,
  2.647011e-08, 2.789007e-08, 2.690405e-08, 2.425944e-08, 2.128022e-08, 
    1.957264e-08, 1.935645e-08, 1.893141e-08, 1.847451e-08, 1.811333e-08, 
    1.812438e-08, 1.815797e-08, 1.813494e-08, 1.731416e-08, 1.457669e-08,
  2.829684e-08, 2.866742e-08, 2.824325e-08, 2.544558e-08, 2.230056e-08, 
    2.061783e-08, 1.987377e-08, 1.919663e-08, 1.873352e-08, 1.848532e-08, 
    1.829009e-08, 1.828937e-08, 1.818025e-08, 1.791729e-08, 1.594776e-08,
  2.688378e-08, 2.846503e-08, 2.875778e-08, 2.637785e-08, 2.335624e-08, 
    2.149976e-08, 2.082136e-08, 2.029526e-08, 1.954407e-08, 1.897545e-08, 
    1.84317e-08, 1.835775e-08, 1.833216e-08, 1.812588e-08, 1.707238e-08,
  2.493863e-08, 2.162491e-08, 1.828145e-08, 1.51304e-08, 1.240631e-08, 
    1.056162e-08, 7.440388e-09, 5.499909e-09, 5.832717e-09, 7.14597e-09, 
    8.281566e-09, 1.050196e-08, 9.570464e-09, 9.409916e-09, 8.017849e-09,
  2.74604e-08, 2.390298e-08, 1.969049e-08, 1.537021e-08, 1.265865e-08, 
    1.132896e-08, 8.476739e-09, 5.944158e-09, 4.790473e-09, 6.397257e-09, 
    8.037191e-09, 9.564933e-09, 9.440733e-09, 9.573201e-09, 8.790567e-09,
  3.024718e-08, 2.556848e-08, 2.188249e-08, 1.569273e-08, 1.307439e-08, 
    1.184113e-08, 9.726907e-09, 6.587431e-09, 4.407798e-09, 5.237593e-09, 
    7.720642e-09, 8.989393e-09, 9.584589e-09, 9.51975e-09, 9.350582e-09,
  3.213545e-08, 2.783179e-08, 2.383401e-08, 1.709501e-08, 1.387687e-08, 
    1.269686e-08, 1.062251e-08, 7.603282e-09, 5.151495e-09, 4.407786e-09, 
    6.706777e-09, 8.680521e-09, 9.395994e-09, 9.624799e-09, 9.588733e-09,
  3.471395e-08, 3.241889e-08, 2.426252e-08, 1.982207e-08, 1.465649e-08, 
    1.341143e-08, 1.14814e-08, 8.79681e-09, 6.133464e-09, 4.591531e-09, 
    6.094939e-09, 8.234393e-09, 9.369473e-09, 9.581012e-09, 9.56978e-09,
  3.373152e-08, 3.339239e-08, 2.453424e-08, 2.092336e-08, 1.657426e-08, 
    1.453576e-08, 1.263736e-08, 9.744811e-09, 7.125163e-09, 4.908769e-09, 
    5.269838e-09, 7.768967e-09, 9.05157e-09, 9.585837e-09, 9.693037e-09,
  3.1808e-08, 3.092926e-08, 2.539471e-08, 2.11837e-08, 1.839707e-08, 
    1.515316e-08, 1.253116e-08, 1.012349e-08, 7.445624e-09, 5.662847e-09, 
    5.234111e-09, 7.148692e-09, 8.816814e-09, 9.324958e-09, 9.565351e-09,
  3.082273e-08, 3.089755e-08, 2.621477e-08, 2.231103e-08, 1.969238e-08, 
    1.597921e-08, 1.392539e-08, 1.286291e-08, 9.502471e-09, 6.938772e-09, 
    5.515293e-09, 6.718766e-09, 8.53399e-09, 9.148916e-09, 9.664604e-09,
  3.351099e-08, 3.215322e-08, 2.831591e-08, 2.423527e-08, 2.079688e-08, 
    1.884947e-08, 1.586726e-08, 1.323968e-08, 9.918224e-09, 7.137539e-09, 
    6.25325e-09, 6.943073e-09, 8.169547e-09, 8.930386e-09, 9.682019e-09,
  3.587262e-08, 3.240596e-08, 3.057382e-08, 2.429691e-08, 2.203307e-08, 
    2.066843e-08, 1.733802e-08, 1.424652e-08, 1.062588e-08, 8.134504e-09, 
    7.232796e-09, 7.507451e-09, 8.316997e-09, 8.943085e-09, 9.546252e-09,
  1.050807e-08, 1.019088e-08, 9.78105e-09, 8.936952e-09, 8.536527e-09, 
    9.351491e-09, 9.611103e-09, 9.674717e-09, 8.669214e-09, 7.226675e-09, 
    6.640727e-09, 5.988633e-09, 5.653757e-09, 6.184805e-09, 6.420293e-09,
  1.116699e-08, 1.050595e-08, 1.049915e-08, 9.825693e-09, 8.72479e-09, 
    9.053312e-09, 9.455319e-09, 9.561151e-09, 8.967707e-09, 7.656338e-09, 
    6.862523e-09, 6.442499e-09, 6.041219e-09, 6.087712e-09, 6.489339e-09,
  1.29051e-08, 1.155057e-08, 1.086994e-08, 1.056832e-08, 9.454726e-09, 
    9.168057e-09, 9.477164e-09, 9.567581e-09, 9.319134e-09, 7.876743e-09, 
    7.112502e-09, 6.823484e-09, 6.597511e-09, 6.077117e-09, 6.59648e-09,
  1.417836e-08, 1.286607e-08, 1.185568e-08, 1.126721e-08, 1.041942e-08, 
    9.586386e-09, 9.71402e-09, 9.726051e-09, 9.45831e-09, 8.067363e-09, 
    7.126146e-09, 6.903752e-09, 7.142817e-09, 6.471788e-09, 6.636821e-09,
  1.621265e-08, 1.460169e-08, 1.288162e-08, 1.216575e-08, 1.149454e-08, 
    1.037864e-08, 1.004123e-08, 1.002477e-08, 9.790094e-09, 8.643504e-09, 
    7.013657e-09, 6.758095e-09, 7.349221e-09, 6.981799e-09, 6.591491e-09,
  1.947072e-08, 1.644218e-08, 1.443688e-08, 1.310819e-08, 1.244813e-08, 
    1.154372e-08, 1.052079e-08, 1.029863e-08, 9.941997e-09, 9.09507e-09, 
    7.197889e-09, 6.682212e-09, 7.031158e-09, 7.441486e-09, 6.657754e-09,
  2.369992e-08, 1.974021e-08, 1.636753e-08, 1.464377e-08, 1.375884e-08, 
    1.280436e-08, 1.164717e-08, 1.095751e-08, 1.021792e-08, 9.383689e-09, 
    7.815281e-09, 6.448505e-09, 6.799739e-09, 7.874969e-09, 6.791661e-09,
  2.582995e-08, 2.395565e-08, 2.002803e-08, 1.633824e-08, 1.457496e-08, 
    1.417718e-08, 1.308006e-08, 1.181588e-08, 1.050245e-08, 9.032091e-09, 
    8.252964e-09, 6.680537e-09, 6.586672e-09, 8.063153e-09, 7.338835e-09,
  2.642096e-08, 2.649793e-08, 2.31489e-08, 1.975243e-08, 1.634187e-08, 
    1.4539e-08, 1.407709e-08, 1.25784e-08, 1.131471e-08, 9.460126e-09, 
    8.073774e-09, 7.211462e-09, 6.542596e-09, 7.373979e-09, 7.953735e-09,
  2.827233e-08, 2.824008e-08, 2.571111e-08, 2.2327e-08, 1.869314e-08, 
    1.636335e-08, 1.677266e-08, 1.337679e-08, 1.227076e-08, 1.029654e-08, 
    7.923037e-09, 7.111332e-09, 6.939978e-09, 7.002769e-09, 8.309891e-09,
  8.215027e-09, 7.891654e-09, 7.984005e-09, 7.999507e-09, 7.318405e-09, 
    6.390259e-09, 5.972991e-09, 5.763913e-09, 5.597723e-09, 5.821652e-09, 
    5.836925e-09, 5.413006e-09, 4.876511e-09, 4.404407e-09, 4.184925e-09,
  8.670267e-09, 8.044409e-09, 8.132216e-09, 8.175166e-09, 7.564125e-09, 
    6.592927e-09, 5.813358e-09, 5.415105e-09, 5.53233e-09, 5.753705e-09, 
    5.850163e-09, 5.619771e-09, 5.209223e-09, 4.657819e-09, 4.269332e-09,
  9.058302e-09, 8.187347e-09, 8.337845e-09, 8.400794e-09, 7.934944e-09, 
    6.814374e-09, 5.842674e-09, 5.509857e-09, 5.126845e-09, 5.565689e-09, 
    5.862284e-09, 5.732003e-09, 5.473074e-09, 4.952077e-09, 4.588364e-09,
  9.741344e-09, 8.603121e-09, 8.658972e-09, 8.60673e-09, 8.329795e-09, 
    7.159226e-09, 6.219274e-09, 5.482959e-09, 5.063573e-09, 5.460318e-09, 
    5.783982e-09, 5.798533e-09, 5.613527e-09, 5.175224e-09, 5.057228e-09,
  1.108501e-08, 9.556427e-09, 9.041642e-09, 8.779057e-09, 8.523384e-09, 
    7.391807e-09, 6.36404e-09, 5.506718e-09, 5.120514e-09, 5.313989e-09, 
    5.624045e-09, 5.755063e-09, 5.75695e-09, 5.34964e-09, 5.344053e-09,
  1.253212e-08, 1.039259e-08, 9.335943e-09, 8.84677e-09, 8.639562e-09, 
    7.651913e-09, 6.386845e-09, 5.213106e-09, 4.706727e-09, 4.996731e-09, 
    5.356432e-09, 5.501243e-09, 5.786545e-09, 5.625706e-09, 5.559688e-09,
  1.313091e-08, 1.11606e-08, 9.652848e-09, 8.919812e-09, 8.39063e-09, 
    7.489666e-09, 6.214047e-09, 4.902154e-09, 4.351376e-09, 4.63435e-09, 
    5.271545e-09, 5.410519e-09, 5.638028e-09, 5.773205e-09, 5.554136e-09,
  1.292578e-08, 1.17802e-08, 1.005117e-08, 8.965805e-09, 7.967966e-09, 
    7.423576e-09, 6.660093e-09, 5.383165e-09, 4.39556e-09, 4.269344e-09, 
    5.165854e-09, 5.332962e-09, 5.561501e-09, 5.882825e-09, 5.782161e-09,
  1.32016e-08, 1.225628e-08, 1.074531e-08, 9.06823e-09, 7.97348e-09, 
    7.943057e-09, 7.776701e-09, 6.911169e-09, 5.297305e-09, 4.260008e-09, 
    5.025409e-09, 5.444437e-09, 5.519558e-09, 5.881737e-09, 5.99753e-09,
  1.380528e-08, 1.241734e-08, 1.155353e-08, 9.610702e-09, 8.560056e-09, 
    8.683576e-09, 8.50042e-09, 7.609562e-09, 5.595867e-09, 4.277042e-09, 
    4.708954e-09, 5.419622e-09, 5.764198e-09, 5.800824e-09, 6.152085e-09,
  2.014455e-08, 1.797232e-08, 1.466991e-08, 1.332006e-08, 1.225323e-08, 
    1.07637e-08, 9.085302e-09, 7.333932e-09, 5.658844e-09, 4.364895e-09, 
    3.649773e-09, 3.404725e-09, 3.126003e-09, 2.60645e-09, 2.240455e-09,
  2.073845e-08, 1.952696e-08, 1.69959e-08, 1.417151e-08, 1.28269e-08, 
    1.146718e-08, 9.868902e-09, 8.085608e-09, 6.51171e-09, 4.922303e-09, 
    3.92167e-09, 3.506243e-09, 3.398391e-09, 2.920872e-09, 2.433219e-09,
  2.330565e-08, 2.093402e-08, 1.912045e-08, 1.584402e-08, 1.36636e-08, 
    1.204552e-08, 1.066681e-08, 8.882385e-09, 7.229519e-09, 5.649624e-09, 
    4.34813e-09, 3.683841e-09, 3.572007e-09, 3.215726e-09, 2.560068e-09,
  2.453796e-08, 2.278505e-08, 2.057665e-08, 1.816445e-08, 1.456921e-08, 
    1.320032e-08, 1.116849e-08, 9.67823e-09, 7.826941e-09, 6.381156e-09, 
    4.847635e-09, 3.974046e-09, 3.738013e-09, 3.486701e-09, 2.808486e-09,
  2.673696e-08, 2.383118e-08, 2.186477e-08, 2.002765e-08, 1.692736e-08, 
    1.3747e-08, 1.226232e-08, 1.041223e-08, 8.693886e-09, 7.047626e-09, 
    5.492226e-09, 4.331175e-09, 3.912321e-09, 3.734697e-09, 3.051831e-09,
  2.681953e-08, 2.495818e-08, 2.229454e-08, 2.096622e-08, 1.914066e-08, 
    1.580823e-08, 1.29775e-08, 1.12561e-08, 9.28215e-09, 7.69936e-09, 
    6.252201e-09, 4.797684e-09, 4.175412e-09, 3.973301e-09, 3.302991e-09,
  2.790751e-08, 2.566746e-08, 2.349405e-08, 2.195192e-08, 2.003438e-08, 
    1.756856e-08, 1.424099e-08, 1.229721e-08, 1.021928e-08, 8.327298e-09, 
    6.921834e-09, 5.387477e-09, 4.562711e-09, 4.17182e-09, 3.578855e-09,
  2.831743e-08, 2.636492e-08, 2.441552e-08, 2.283043e-08, 2.071469e-08, 
    1.926379e-08, 1.583635e-08, 1.299524e-08, 1.127685e-08, 9.173895e-09, 
    7.505186e-09, 6.016888e-09, 4.956919e-09, 4.393829e-09, 3.85675e-09,
  2.788945e-08, 2.741152e-08, 2.492072e-08, 2.294794e-08, 2.140744e-08, 
    1.948268e-08, 1.777583e-08, 1.411609e-08, 1.187725e-08, 9.848486e-09, 
    8.070305e-09, 6.624274e-09, 5.386018e-09, 4.580497e-09, 4.050525e-09,
  2.76182e-08, 2.746257e-08, 2.578833e-08, 2.30306e-08, 2.201467e-08, 
    2.017163e-08, 1.845059e-08, 1.534348e-08, 1.238995e-08, 1.046566e-08, 
    8.681595e-09, 7.127028e-09, 5.791757e-09, 4.83491e-09, 4.252347e-09,
  2.217528e-08, 2.166746e-08, 1.95502e-08, 1.857207e-08, 1.842648e-08, 
    1.689698e-08, 1.445441e-08, 1.196179e-08, 9.113429e-09, 6.071883e-09, 
    4.360487e-09, 4.670413e-09, 5.353501e-09, 5.037041e-09, 5.003691e-09,
  2.004833e-08, 2.205756e-08, 2.091546e-08, 1.92666e-08, 1.837212e-08, 
    1.778567e-08, 1.557912e-08, 1.306738e-08, 1.060524e-08, 7.457463e-09, 
    5.093928e-09, 4.211102e-09, 4.968208e-09, 4.979661e-09, 5.067448e-09,
  1.95561e-08, 2.077163e-08, 2.169689e-08, 2.034132e-08, 1.882811e-08, 
    1.821519e-08, 1.671701e-08, 1.418917e-08, 1.159963e-08, 8.768088e-09, 
    6.062596e-09, 4.412967e-09, 4.667109e-09, 4.812257e-09, 5.034744e-09,
  2.162728e-08, 2.016422e-08, 2.089318e-08, 2.110008e-08, 1.98725e-08, 
    1.85119e-08, 1.757627e-08, 1.528243e-08, 1.272872e-08, 9.825385e-09, 
    7.155819e-09, 4.93102e-09, 4.583827e-09, 4.74373e-09, 4.905127e-09,
  2.526959e-08, 2.192746e-08, 2.107472e-08, 2.064054e-08, 2.075889e-08, 
    1.942122e-08, 1.811916e-08, 1.638836e-08, 1.40203e-08, 1.110902e-08, 
    8.491095e-09, 5.538152e-09, 4.745426e-09, 4.962488e-09, 5.039902e-09,
  2.887476e-08, 2.522791e-08, 2.254934e-08, 2.163232e-08, 2.034812e-08, 
    2.03703e-08, 1.909493e-08, 1.71706e-08, 1.496454e-08, 1.222826e-08, 
    9.652961e-09, 6.550491e-09, 4.883562e-09, 4.946363e-09, 5.166711e-09,
  3.142654e-08, 3.016909e-08, 2.624041e-08, 2.279748e-08, 2.188318e-08, 
    2.013502e-08, 1.977866e-08, 1.836598e-08, 1.609331e-08, 1.338981e-08, 
    1.067024e-08, 7.971297e-09, 5.300504e-09, 4.883527e-09, 5.402268e-09,
  3.323107e-08, 3.355809e-08, 3.124742e-08, 2.685041e-08, 2.30029e-08, 
    2.179931e-08, 2.020023e-08, 1.910773e-08, 1.752713e-08, 1.488096e-08, 
    1.192159e-08, 9.411669e-09, 6.13542e-09, 4.981467e-09, 5.420947e-09,
  3.221925e-08, 3.403919e-08, 3.46064e-08, 3.197603e-08, 2.716144e-08, 
    2.286357e-08, 2.189509e-08, 1.95474e-08, 1.800009e-08, 1.58465e-08, 
    1.345168e-08, 1.078444e-08, 7.370949e-09, 5.218586e-09, 5.151619e-09,
  3.038294e-08, 3.22398e-08, 3.51254e-08, 3.554636e-08, 3.273811e-08, 
    2.696554e-08, 2.33185e-08, 2.127748e-08, 1.860476e-08, 1.725258e-08, 
    1.517702e-08, 1.220986e-08, 8.939946e-09, 5.719945e-09, 4.951149e-09,
  2.242478e-08, 2.03752e-08, 1.884208e-08, 1.707668e-08, 1.386554e-08, 
    1.384652e-08, 1.356878e-08, 1.061918e-08, 8.089779e-09, 7.596549e-09, 
    8.56455e-09, 8.296241e-09, 8.070434e-09, 9.086999e-09, 9.731609e-09,
  2.187109e-08, 2.123905e-08, 2.02772e-08, 1.948351e-08, 1.579003e-08, 
    1.401322e-08, 1.418093e-08, 1.284559e-08, 9.747655e-09, 8.10417e-09, 
    8.039527e-09, 8.271692e-09, 7.968073e-09, 8.712366e-09, 9.293542e-09,
  2.192526e-08, 2.169697e-08, 2.125175e-08, 2.074746e-08, 1.85572e-08, 
    1.534153e-08, 1.409425e-08, 1.410995e-08, 1.209751e-08, 9.435107e-09, 
    8.149168e-09, 7.884204e-09, 7.970191e-09, 8.37778e-09, 8.947681e-09,
  2.129135e-08, 2.199041e-08, 2.162715e-08, 2.097864e-08, 2.093584e-08, 
    1.793124e-08, 1.535448e-08, 1.437276e-08, 1.386284e-08, 1.15669e-08, 
    8.906452e-09, 7.820665e-09, 7.445847e-09, 8.051671e-09, 8.892302e-09,
  2.095656e-08, 2.206112e-08, 2.193291e-08, 2.09946e-08, 2.083948e-08, 
    2.037764e-08, 1.748461e-08, 1.522059e-08, 1.437463e-08, 1.357268e-08, 
    1.122995e-08, 8.721117e-09, 7.261451e-09, 7.594354e-09, 8.608206e-09,
  1.78073e-08, 2.10276e-08, 2.234039e-08, 2.185732e-08, 2.058855e-08, 
    2.058544e-08, 2.003995e-08, 1.714236e-08, 1.485708e-08, 1.425549e-08, 
    1.317083e-08, 1.069942e-08, 8.043719e-09, 7.133268e-09, 8.183241e-09,
  1.802366e-08, 1.822012e-08, 2.0374e-08, 2.20116e-08, 2.129735e-08, 
    2.011141e-08, 2.051536e-08, 2.005235e-08, 1.741623e-08, 1.520927e-08, 
    1.449322e-08, 1.285337e-08, 9.97662e-09, 7.785665e-09, 7.629736e-09,
  2.019754e-08, 1.87499e-08, 1.852076e-08, 2.030207e-08, 2.176158e-08, 
    2.111773e-08, 2.027366e-08, 2.06608e-08, 1.965699e-08, 1.720834e-08, 
    1.528577e-08, 1.450868e-08, 1.18101e-08, 9.454268e-09, 7.870875e-09,
  2.330001e-08, 2.065487e-08, 1.907907e-08, 1.853481e-08, 2.011235e-08, 
    2.15875e-08, 2.095512e-08, 2.047615e-08, 2.041426e-08, 1.929655e-08, 
    1.694485e-08, 1.537518e-08, 1.404034e-08, 1.076678e-08, 8.977434e-09,
  2.651617e-08, 2.443887e-08, 2.197256e-08, 1.965009e-08, 1.902606e-08, 
    2.060705e-08, 2.1658e-08, 2.062733e-08, 2.075725e-08, 2.090252e-08, 
    1.924923e-08, 1.714435e-08, 1.54093e-08, 1.305684e-08, 9.961262e-09,
  1.811523e-08, 1.899734e-08, 1.875215e-08, 1.782809e-08, 1.728537e-08, 
    1.684524e-08, 1.654088e-08, 1.512638e-08, 1.493501e-08, 1.493836e-08, 
    1.193022e-08, 9.826589e-09, 7.343913e-09, 6.888988e-09, 6.819005e-09,
  1.639871e-08, 1.853996e-08, 1.938495e-08, 1.903109e-08, 1.806862e-08, 
    1.777183e-08, 1.71564e-08, 1.439644e-08, 1.371845e-08, 1.341287e-08, 
    1.153685e-08, 1.087121e-08, 9.921783e-09, 8.767567e-09, 7.823552e-09,
  1.52592e-08, 1.669802e-08, 1.88751e-08, 1.908853e-08, 1.908993e-08, 
    1.806264e-08, 1.812177e-08, 1.533452e-08, 1.343734e-08, 1.267299e-08, 
    1.067293e-08, 1.066604e-08, 1.055245e-08, 1.055158e-08, 9.585072e-09,
  1.624472e-08, 1.642196e-08, 1.767302e-08, 1.858217e-08, 1.908112e-08, 
    1.894485e-08, 1.859939e-08, 1.696624e-08, 1.400313e-08, 1.284326e-08, 
    1.151648e-08, 9.649143e-09, 1.022354e-08, 1.0577e-08, 1.086921e-08,
  1.657603e-08, 1.676771e-08, 1.748687e-08, 1.82834e-08, 1.881241e-08, 
    1.899193e-08, 1.88426e-08, 1.874776e-08, 1.501328e-08, 1.336723e-08, 
    1.220138e-08, 1.076756e-08, 9.519588e-09, 9.153385e-09, 1.04593e-08,
  1.684842e-08, 1.712797e-08, 1.692708e-08, 1.804067e-08, 1.848929e-08, 
    1.879867e-08, 1.891601e-08, 1.900597e-08, 1.683586e-08, 1.392725e-08, 
    1.251069e-08, 1.138372e-08, 9.96859e-09, 8.845013e-09, 9.10757e-09,
  1.928747e-08, 1.827782e-08, 1.799479e-08, 1.775898e-08, 1.841146e-08, 
    1.837392e-08, 1.820714e-08, 1.9059e-08, 1.906194e-08, 1.545898e-08, 
    1.291272e-08, 1.169746e-08, 1.067336e-08, 9.650262e-09, 8.562326e-09,
  2.288436e-08, 2.097764e-08, 1.960283e-08, 1.901568e-08, 1.892139e-08, 
    1.890628e-08, 1.861126e-08, 1.934031e-08, 1.968741e-08, 1.788533e-08, 
    1.398427e-08, 1.171446e-08, 1.09906e-08, 1.007927e-08, 8.893689e-09,
  2.696176e-08, 2.412721e-08, 2.188453e-08, 2.027719e-08, 1.981685e-08, 
    2.005591e-08, 2.007546e-08, 1.959056e-08, 1.958211e-08, 1.784234e-08, 
    1.513651e-08, 1.195945e-08, 1.097755e-08, 1.045525e-08, 9.362543e-09,
  3.22222e-08, 3.098638e-08, 2.701295e-08, 2.26189e-08, 2.11285e-08, 
    2.180096e-08, 2.157609e-08, 1.969635e-08, 1.960164e-08, 1.846097e-08, 
    1.662119e-08, 1.294955e-08, 1.098731e-08, 1.041687e-08, 9.727245e-09,
  9.126961e-09, 8.895383e-09, 8.67941e-09, 8.292546e-09, 8.009331e-09, 
    7.5182e-09, 7.22856e-09, 7.175011e-09, 7.222591e-09, 8.64233e-09, 
    7.482482e-09, 5.247231e-09, 4.488375e-09, 5.355094e-09, 5.793264e-09,
  1.077817e-08, 1.036753e-08, 1.012068e-08, 9.7755e-09, 9.434635e-09, 
    9.20063e-09, 8.830005e-09, 8.301726e-09, 8.162649e-09, 8.649611e-09, 
    7.581202e-09, 6.306915e-09, 4.837315e-09, 4.489824e-09, 4.518472e-09,
  1.301456e-08, 1.264087e-08, 1.232181e-08, 1.194948e-08, 1.162512e-08, 
    1.113825e-08, 1.090577e-08, 1.045211e-08, 9.767835e-09, 9.497447e-09, 
    9.090882e-09, 7.198484e-09, 5.997273e-09, 4.722336e-09, 4.430787e-09,
  1.419652e-08, 1.400836e-08, 1.409815e-08, 1.381349e-08, 1.351199e-08, 
    1.317451e-08, 1.28177e-08, 1.281389e-08, 1.238102e-08, 1.156473e-08, 
    1.176863e-08, 9.09273e-09, 7.345283e-09, 6.032726e-09, 5.07906e-09,
  1.375391e-08, 1.402273e-08, 1.448534e-08, 1.49292e-08, 1.498761e-08, 
    1.484193e-08, 1.43706e-08, 1.419782e-08, 1.426834e-08, 1.383626e-08, 
    1.351151e-08, 1.211795e-08, 9.330925e-09, 7.76841e-09, 6.412465e-09,
  1.430647e-08, 1.426903e-08, 1.404296e-08, 1.454398e-08, 1.478407e-08, 
    1.495424e-08, 1.494759e-08, 1.45946e-08, 1.471836e-08, 1.490897e-08, 
    1.474696e-08, 1.463211e-08, 1.146523e-08, 9.45564e-09, 7.905712e-09,
  1.712157e-08, 1.644349e-08, 1.595443e-08, 1.545357e-08, 1.567321e-08, 
    1.551405e-08, 1.536292e-08, 1.516635e-08, 1.480296e-08, 1.511934e-08, 
    1.541623e-08, 1.511723e-08, 1.368677e-08, 1.117382e-08, 9.56151e-09,
  2.061289e-08, 2.005737e-08, 1.91611e-08, 1.810561e-08, 1.754028e-08, 
    1.723691e-08, 1.671413e-08, 1.611543e-08, 1.543283e-08, 1.515914e-08, 
    1.522431e-08, 1.534313e-08, 1.471822e-08, 1.225938e-08, 1.07935e-08,
  2.328666e-08, 2.304492e-08, 2.20934e-08, 2.163931e-08, 2.046571e-08, 
    1.906065e-08, 1.861883e-08, 1.771276e-08, 1.702488e-08, 1.622082e-08, 
    1.584687e-08, 1.578589e-08, 1.508364e-08, 1.37238e-08, 1.13831e-08,
  2.512001e-08, 2.5347e-08, 2.495479e-08, 2.468226e-08, 2.360777e-08, 
    2.195755e-08, 2.066056e-08, 1.987399e-08, 1.902652e-08, 1.789362e-08, 
    1.705368e-08, 1.656523e-08, 1.574007e-08, 1.465867e-08, 1.251181e-08,
  3.996579e-09, 4.034214e-09, 3.858974e-09, 3.679501e-09, 3.534682e-09, 
    3.534532e-09, 3.691776e-09, 3.926408e-09, 4.040929e-09, 4.308599e-09, 
    4.805817e-09, 4.80131e-09, 4.283526e-09, 3.948425e-09, 3.981949e-09,
  4.218716e-09, 4.291032e-09, 4.3333e-09, 4.184862e-09, 4.055695e-09, 
    3.923128e-09, 3.864268e-09, 3.997371e-09, 4.14805e-09, 4.207257e-09, 
    4.421691e-09, 5.145438e-09, 5.351954e-09, 4.520838e-09, 4.04397e-09,
  4.364594e-09, 4.495023e-09, 4.618352e-09, 4.603075e-09, 4.451488e-09, 
    4.246817e-09, 4.141651e-09, 4.161427e-09, 4.292909e-09, 4.389837e-09, 
    4.462281e-09, 4.613417e-09, 5.330887e-09, 5.508354e-09, 4.805706e-09,
  4.462579e-09, 4.675564e-09, 4.780477e-09, 4.852892e-09, 4.811913e-09, 
    4.659123e-09, 4.429726e-09, 4.326112e-09, 4.333945e-09, 4.448356e-09, 
    4.598419e-09, 4.801117e-09, 5.019689e-09, 5.562593e-09, 5.739622e-09,
  4.643836e-09, 4.687283e-09, 4.674185e-09, 4.764014e-09, 4.969597e-09, 
    4.920453e-09, 4.704543e-09, 4.518166e-09, 4.484431e-09, 4.551137e-09, 
    4.75218e-09, 4.948768e-09, 5.21735e-09, 5.485066e-09, 5.905621e-09,
  5.388734e-09, 5.250339e-09, 5.049414e-09, 4.924039e-09, 4.913133e-09, 
    4.987181e-09, 4.922468e-09, 4.772332e-09, 4.71191e-09, 4.743871e-09, 
    4.922438e-09, 5.210617e-09, 5.453509e-09, 5.68294e-09, 6.103213e-09,
  5.771275e-09, 5.567858e-09, 5.406013e-09, 5.275735e-09, 5.153465e-09, 
    5.097948e-09, 5.091953e-09, 5.11551e-09, 5.129918e-09, 5.133897e-09, 
    5.157465e-09, 5.307528e-09, 5.577325e-09, 5.813461e-09, 6.038252e-09,
  6.128208e-09, 6.10085e-09, 6.056103e-09, 5.91741e-09, 5.779774e-09, 
    5.824311e-09, 5.919542e-09, 5.984968e-09, 6.082817e-09, 5.967214e-09, 
    5.857857e-09, 5.843035e-09, 5.920648e-09, 6.080196e-09, 6.175933e-09,
  6.690727e-09, 6.716205e-09, 6.714485e-09, 6.763649e-09, 6.802999e-09, 
    6.927991e-09, 7.081793e-09, 7.176283e-09, 7.137269e-09, 7.072789e-09, 
    6.990704e-09, 6.901126e-09, 6.895638e-09, 6.890144e-09, 6.876137e-09,
  7.522432e-09, 7.537729e-09, 7.543486e-09, 7.725993e-09, 7.978441e-09, 
    8.187894e-09, 8.316017e-09, 8.527643e-09, 8.597705e-09, 8.623302e-09, 
    8.59353e-09, 8.487488e-09, 8.337854e-09, 8.144406e-09, 8.038286e-09,
  1.270988e-09, 1.258117e-09, 1.197224e-09, 1.196752e-09, 1.224022e-09, 
    1.289125e-09, 1.30816e-09, 1.248359e-09, 1.162385e-09, 1.074869e-09, 
    1.102771e-09, 1.194559e-09, 1.406034e-09, 1.742679e-09, 1.946987e-09,
  1.311416e-09, 1.243475e-09, 1.151671e-09, 1.13646e-09, 1.189698e-09, 
    1.267061e-09, 1.290078e-09, 1.263623e-09, 1.172971e-09, 1.141744e-09, 
    1.170922e-09, 1.24572e-09, 1.38178e-09, 1.611897e-09, 1.856771e-09,
  1.356443e-09, 1.306541e-09, 1.169947e-09, 1.111533e-09, 1.200301e-09, 
    1.35174e-09, 1.42863e-09, 1.411945e-09, 1.30476e-09, 1.276889e-09, 
    1.287653e-09, 1.31437e-09, 1.411763e-09, 1.591485e-09, 1.8689e-09,
  1.35173e-09, 1.369477e-09, 1.271475e-09, 1.161267e-09, 1.191313e-09, 
    1.421567e-09, 1.67664e-09, 1.826754e-09, 1.876192e-09, 1.753462e-09, 
    1.659873e-09, 1.621375e-09, 1.695801e-09, 1.83417e-09, 2.102549e-09,
  1.441248e-09, 1.541988e-09, 1.364496e-09, 1.214819e-09, 1.140673e-09, 
    1.347372e-09, 1.759002e-09, 2.153035e-09, 2.395142e-09, 2.529816e-09, 
    2.406111e-09, 2.23693e-09, 2.171049e-09, 2.223842e-09, 2.438963e-09,
  1.543907e-09, 1.555263e-09, 1.451835e-09, 1.279306e-09, 1.197868e-09, 
    1.309383e-09, 1.705829e-09, 2.132911e-09, 2.535321e-09, 2.778945e-09, 
    2.830315e-09, 2.877107e-09, 2.812939e-09, 2.796721e-09, 2.972035e-09,
  1.460769e-09, 1.528985e-09, 1.489349e-09, 1.433896e-09, 1.395855e-09, 
    1.395678e-09, 1.578431e-09, 1.827256e-09, 2.274402e-09, 2.675123e-09, 
    2.915692e-09, 2.929946e-09, 3.075639e-09, 3.274967e-09, 3.470208e-09,
  1.47882e-09, 1.512483e-09, 1.558985e-09, 1.579956e-09, 1.512173e-09, 
    1.55685e-09, 1.669858e-09, 1.980642e-09, 2.263836e-09, 2.567371e-09, 
    2.802959e-09, 3.012113e-09, 3.201293e-09, 3.467854e-09, 3.753448e-09,
  1.647296e-09, 1.605527e-09, 1.648529e-09, 1.680695e-09, 1.620072e-09, 
    1.691306e-09, 1.809886e-09, 2.143003e-09, 2.403964e-09, 2.614212e-09, 
    2.895915e-09, 3.116384e-09, 3.246995e-09, 3.535183e-09, 3.841051e-09,
  1.903767e-09, 1.769324e-09, 1.717968e-09, 1.71334e-09, 1.75836e-09, 
    1.820079e-09, 1.79774e-09, 1.972115e-09, 2.237252e-09, 2.520609e-09, 
    2.764227e-09, 2.957357e-09, 3.218756e-09, 3.552749e-09, 3.921527e-09,
  1.922267e-09, 2.053052e-09, 2.330203e-09, 2.497895e-09, 2.572206e-09, 
    2.551698e-09, 2.5529e-09, 2.560949e-09, 2.536096e-09, 2.503521e-09, 
    2.354005e-09, 2.024221e-09, 1.540847e-09, 1.142176e-09, 9.560562e-10,
  1.741539e-09, 1.966662e-09, 2.285164e-09, 2.485338e-09, 2.559161e-09, 
    2.55451e-09, 2.558611e-09, 2.574633e-09, 2.551271e-09, 2.548409e-09, 
    2.396656e-09, 2.021648e-09, 1.483012e-09, 1.051167e-09, 8.657544e-10,
  1.597981e-09, 1.917599e-09, 2.22523e-09, 2.421758e-09, 2.537447e-09, 
    2.548479e-09, 2.55917e-09, 2.599668e-09, 2.582049e-09, 2.596505e-09, 
    2.46762e-09, 2.059769e-09, 1.542594e-09, 1.05024e-09, 8.615585e-10,
  1.647296e-09, 1.880281e-09, 2.152089e-09, 2.371254e-09, 2.520444e-09, 
    2.581682e-09, 2.572122e-09, 2.569561e-09, 2.575543e-09, 2.619364e-09, 
    2.518328e-09, 2.165146e-09, 1.643037e-09, 1.115073e-09, 8.996757e-10,
  1.885649e-09, 1.891905e-09, 2.033798e-09, 2.294703e-09, 2.468864e-09, 
    2.529034e-09, 2.551278e-09, 2.589782e-09, 2.586926e-09, 2.59546e-09, 
    2.557834e-09, 2.266106e-09, 1.780918e-09, 1.309362e-09, 1.10058e-09,
  2.093001e-09, 1.874658e-09, 1.879717e-09, 2.105441e-09, 2.382e-09, 
    2.521478e-09, 2.53144e-09, 2.518518e-09, 2.539651e-09, 2.575561e-09, 
    2.530741e-09, 2.366689e-09, 1.831009e-09, 1.397725e-09, 1.195222e-09,
  2.330188e-09, 1.787917e-09, 1.699129e-09, 1.921114e-09, 2.21645e-09, 
    2.356442e-09, 2.496739e-09, 2.52506e-09, 2.503055e-09, 2.515904e-09, 
    2.526215e-09, 2.211006e-09, 1.950748e-09, 1.424688e-09, 1.222438e-09,
  2.710374e-09, 1.928864e-09, 1.687799e-09, 1.733867e-09, 2.115277e-09, 
    2.301982e-09, 2.423292e-09, 2.531001e-09, 2.592574e-09, 2.581636e-09, 
    2.458806e-09, 2.232995e-09, 1.961187e-09, 1.685544e-09, 1.37276e-09,
  3.128127e-09, 2.175945e-09, 1.819692e-09, 1.652519e-09, 1.900352e-09, 
    2.272418e-09, 2.476737e-09, 2.54122e-09, 2.502365e-09, 2.520764e-09, 
    2.467329e-09, 2.357539e-09, 2.00703e-09, 1.729622e-09, 1.508237e-09,
  3.631899e-09, 2.577451e-09, 1.978637e-09, 1.714772e-09, 1.779654e-09, 
    2.18585e-09, 2.461457e-09, 2.535312e-09, 2.421248e-09, 2.463489e-09, 
    2.488707e-09, 2.315601e-09, 2.098493e-09, 1.719095e-09, 1.448153e-09,
  7.013481e-09, 5.573901e-09, 4.411722e-09, 3.435191e-09, 2.776961e-09, 
    2.218264e-09, 1.812875e-09, 1.5363e-09, 1.429867e-09, 1.423888e-09, 
    1.604096e-09, 1.986867e-09, 2.744658e-09, 3.282164e-09, 3.254952e-09,
  7.267344e-09, 5.921045e-09, 4.655171e-09, 3.634115e-09, 2.960079e-09, 
    2.369141e-09, 1.930931e-09, 1.593583e-09, 1.515398e-09, 1.460535e-09, 
    1.544139e-09, 1.864255e-09, 2.492272e-09, 3.118755e-09, 3.169282e-09,
  7.45996e-09, 6.22892e-09, 4.971709e-09, 3.862943e-09, 3.134167e-09, 
    2.504005e-09, 2.036169e-09, 1.647217e-09, 1.562695e-09, 1.515444e-09, 
    1.556674e-09, 1.820531e-09, 2.290751e-09, 2.859393e-09, 2.973146e-09,
  7.855547e-09, 6.495989e-09, 5.302895e-09, 4.047858e-09, 3.332134e-09, 
    2.67443e-09, 2.198816e-09, 1.717631e-09, 1.614567e-09, 1.569703e-09, 
    1.563468e-09, 1.7792e-09, 2.164755e-09, 2.698332e-09, 2.787577e-09,
  8.336952e-09, 6.798217e-09, 5.605103e-09, 4.354747e-09, 3.554389e-09, 
    2.802695e-09, 2.300435e-09, 1.778953e-09, 1.635909e-09, 1.623195e-09, 
    1.601693e-09, 1.769967e-09, 2.117048e-09, 2.557606e-09, 2.637339e-09,
  8.745985e-09, 7.23468e-09, 5.959611e-09, 4.646847e-09, 3.782606e-09, 
    2.982418e-09, 2.443961e-09, 1.849859e-09, 1.622794e-09, 1.559781e-09, 
    1.620195e-09, 1.697521e-09, 2.040791e-09, 2.487409e-09, 2.578724e-09,
  9.134987e-09, 7.597738e-09, 6.305095e-09, 5.035085e-09, 3.971466e-09, 
    3.076112e-09, 2.600568e-09, 2.068739e-09, 1.720778e-09, 1.511504e-09, 
    1.595612e-09, 1.6738e-09, 1.957192e-09, 2.371582e-09, 2.549773e-09,
  9.594864e-09, 8.066897e-09, 6.661586e-09, 5.34088e-09, 4.324507e-09, 
    3.309802e-09, 2.638722e-09, 2.122424e-09, 1.788317e-09, 1.610421e-09, 
    1.619447e-09, 1.685573e-09, 1.91429e-09, 2.304737e-09, 2.508261e-09,
  9.772402e-09, 8.359745e-09, 7.041654e-09, 5.655679e-09, 4.658999e-09, 
    3.73268e-09, 2.951293e-09, 2.286516e-09, 1.843525e-09, 1.768167e-09, 
    1.722797e-09, 1.749727e-09, 1.84886e-09, 2.224808e-09, 2.444964e-09,
  1.01066e-08, 8.617923e-09, 7.403583e-09, 6.121363e-09, 4.981007e-09, 
    4.118891e-09, 3.213147e-09, 2.532223e-09, 2.006306e-09, 1.87354e-09, 
    1.779633e-09, 1.829846e-09, 1.83067e-09, 2.129374e-09, 2.378433e-09,
  8.539391e-09, 6.847142e-09, 5.740885e-09, 4.589539e-09, 3.469102e-09, 
    2.632347e-09, 2.084457e-09, 1.918657e-09, 2.230729e-09, 2.250291e-09, 
    2.068733e-09, 2.059781e-09, 2.271183e-09, 2.344061e-09, 2.280855e-09,
  9.256756e-09, 7.467584e-09, 6.233905e-09, 5.089658e-09, 3.960154e-09, 
    2.949417e-09, 2.231759e-09, 1.813142e-09, 2.139689e-09, 2.236817e-09, 
    2.0525e-09, 1.981099e-09, 2.147424e-09, 2.203574e-09, 2.218407e-09,
  1.013652e-08, 8.231831e-09, 6.808281e-09, 5.546078e-09, 4.464328e-09, 
    3.305385e-09, 2.453602e-09, 1.849981e-09, 2.038333e-09, 2.24103e-09, 
    2.073295e-09, 1.948517e-09, 2.043325e-09, 2.069384e-09, 2.149679e-09,
  1.101695e-08, 9.05723e-09, 7.511191e-09, 6.040621e-09, 5.017532e-09, 
    3.742465e-09, 2.753577e-09, 1.979343e-09, 1.94691e-09, 2.182526e-09, 
    2.046721e-09, 1.910073e-09, 1.97505e-09, 2.008224e-09, 2.094303e-09,
  1.250846e-08, 9.921014e-09, 8.274421e-09, 6.699428e-09, 5.565511e-09, 
    4.227587e-09, 3.074187e-09, 2.18343e-09, 1.934291e-09, 2.122725e-09, 
    2.038359e-09, 1.888842e-09, 1.949383e-09, 1.982807e-09, 2.028507e-09,
  1.395529e-08, 1.082194e-08, 9.097671e-09, 7.443608e-09, 6.203657e-09, 
    4.801241e-09, 3.516514e-09, 2.456193e-09, 2.025994e-09, 2.044998e-09, 
    1.979897e-09, 1.853846e-09, 1.922245e-09, 1.964914e-09, 1.95674e-09,
  1.504093e-08, 1.171442e-08, 9.86908e-09, 8.229631e-09, 6.722119e-09, 
    5.278632e-09, 3.995152e-09, 2.927956e-09, 2.313249e-09, 2.067888e-09, 
    1.942966e-09, 1.759401e-09, 1.87817e-09, 1.881368e-09, 1.886252e-09,
  1.665191e-08, 1.304054e-08, 1.092084e-08, 8.975253e-09, 7.307813e-09, 
    5.912635e-09, 4.3731e-09, 3.054659e-09, 2.329739e-09, 2.18825e-09, 
    1.988041e-09, 1.722736e-09, 1.766972e-09, 1.77148e-09, 1.820487e-09,
  1.842982e-08, 1.477602e-08, 1.18913e-08, 9.466963e-09, 7.810041e-09, 
    6.675686e-09, 4.931264e-09, 3.420066e-09, 2.54236e-09, 2.453532e-09, 
    2.122757e-09, 1.744459e-09, 1.613905e-09, 1.656125e-09, 1.765668e-09,
  1.970379e-08, 1.642749e-08, 1.308589e-08, 1.017991e-08, 8.398829e-09, 
    7.240622e-09, 5.335974e-09, 3.826592e-09, 3.06213e-09, 2.725077e-09, 
    2.271719e-09, 1.776431e-09, 1.467013e-09, 1.548173e-09, 1.710425e-09,
  9.308747e-09, 7.202391e-09, 5.444159e-09, 4.17528e-09, 3.435892e-09, 
    3.413302e-09, 3.132056e-09, 2.993664e-09, 3.160489e-09, 3.392248e-09, 
    3.658984e-09, 3.967832e-09, 4.150039e-09, 4.062831e-09, 3.80773e-09,
  1.032914e-08, 7.965158e-09, 5.96524e-09, 4.473649e-09, 3.389554e-09, 
    3.143291e-09, 3.127159e-09, 2.922189e-09, 3.053238e-09, 3.26203e-09, 
    3.524961e-09, 3.852719e-09, 4.144235e-09, 4.200685e-09, 4.009932e-09,
  1.148686e-08, 8.750055e-09, 6.523402e-09, 4.806527e-09, 3.600132e-09, 
    3.016724e-09, 3.072233e-09, 2.967097e-09, 3.08394e-09, 3.227777e-09, 
    3.410105e-09, 3.712434e-09, 4.047605e-09, 4.174848e-09, 4.035745e-09,
  1.231019e-08, 9.59382e-09, 7.143597e-09, 5.268163e-09, 3.938667e-09, 
    3.057231e-09, 3.037701e-09, 3.053862e-09, 3.119799e-09, 3.169169e-09, 
    3.311656e-09, 3.538711e-09, 3.882954e-09, 4.04314e-09, 3.93131e-09,
  1.302849e-08, 1.046046e-08, 7.895668e-09, 5.731974e-09, 4.291773e-09, 
    3.133553e-09, 3.047514e-09, 3.072161e-09, 3.042692e-09, 3.101591e-09, 
    3.275309e-09, 3.312816e-09, 3.586268e-09, 3.808306e-09, 3.717032e-09,
  1.398275e-08, 1.103159e-08, 8.433135e-09, 6.138159e-09, 4.622287e-09, 
    3.291092e-09, 2.942287e-09, 2.934795e-09, 2.97797e-09, 3.038829e-09, 
    3.08485e-09, 3.111202e-09, 3.232443e-09, 3.535993e-09, 3.5701e-09,
  1.486011e-08, 1.134793e-08, 8.78588e-09, 6.685813e-09, 4.812655e-09, 
    3.31904e-09, 2.697603e-09, 2.664491e-09, 2.752e-09, 2.939878e-09, 
    2.985299e-09, 2.991591e-09, 2.937655e-09, 3.274923e-09, 3.467046e-09,
  1.608642e-08, 1.192528e-08, 9.188331e-09, 7.18568e-09, 5.095368e-09, 
    3.510842e-09, 2.779078e-09, 2.894377e-09, 2.878842e-09, 2.923422e-09, 
    2.965391e-09, 2.875273e-09, 2.789018e-09, 3.102801e-09, 3.453039e-09,
  1.772506e-08, 1.276986e-08, 9.578951e-09, 7.584283e-09, 5.593434e-09, 
    4.117394e-09, 3.240884e-09, 3.216214e-09, 2.897436e-09, 2.764625e-09, 
    2.948676e-09, 2.78882e-09, 2.777185e-09, 3.004652e-09, 3.394891e-09,
  1.940474e-08, 1.39487e-08, 1.00079e-08, 8.056773e-09, 6.193871e-09, 
    4.432053e-09, 3.318726e-09, 2.973122e-09, 2.677202e-09, 2.592342e-09, 
    2.930109e-09, 2.81469e-09, 2.773239e-09, 3.042083e-09, 3.3099e-09,
  8.123167e-09, 6.52563e-09, 5.223638e-09, 4.377969e-09, 4.168469e-09, 
    4.102803e-09, 3.89886e-09, 3.473356e-09, 3.769955e-09, 3.913545e-09, 
    3.496493e-09, 3.142687e-09, 3.058715e-09, 2.884828e-09, 2.536165e-09,
  8.532664e-09, 7.116138e-09, 5.793764e-09, 4.712898e-09, 4.390512e-09, 
    4.197812e-09, 4.175227e-09, 3.746375e-09, 3.724835e-09, 4.039041e-09, 
    3.727974e-09, 3.294657e-09, 3.224357e-09, 3.23811e-09, 2.966332e-09,
  8.968042e-09, 7.645148e-09, 6.35586e-09, 5.077748e-09, 4.570631e-09, 
    4.304646e-09, 4.166911e-09, 4.078424e-09, 3.848769e-09, 4.067257e-09, 
    3.929292e-09, 3.513064e-09, 3.336201e-09, 3.432214e-09, 3.383426e-09,
  9.760593e-09, 8.420974e-09, 7.039914e-09, 5.516398e-09, 4.845796e-09, 
    4.471098e-09, 4.133885e-09, 4.036882e-09, 3.880988e-09, 4.015285e-09, 
    4.077197e-09, 3.797437e-09, 3.525499e-09, 3.580786e-09, 3.693243e-09,
  1.118801e-08, 9.419018e-09, 7.729735e-09, 5.970823e-09, 5.109455e-09, 
    4.619951e-09, 4.150276e-09, 3.939882e-09, 3.850253e-09, 3.959706e-09, 
    4.184012e-09, 3.957003e-09, 3.805747e-09, 3.747989e-09, 3.873159e-09,
  1.262258e-08, 1.05493e-08, 8.39362e-09, 6.363792e-09, 5.425056e-09, 
    4.861596e-09, 4.230155e-09, 3.747442e-09, 3.667693e-09, 3.871787e-09, 
    4.356137e-09, 4.006952e-09, 4.011579e-09, 3.962349e-09, 4.065697e-09,
  1.354281e-08, 1.131428e-08, 8.900704e-09, 6.775196e-09, 5.573445e-09, 
    4.982268e-09, 4.46155e-09, 3.967427e-09, 3.675223e-09, 3.936949e-09, 
    4.556417e-09, 4.085563e-09, 4.142349e-09, 4.148831e-09, 4.244875e-09,
  1.453011e-08, 1.225851e-08, 9.675373e-09, 7.223789e-09, 5.797076e-09, 
    5.037186e-09, 4.45125e-09, 3.99253e-09, 3.935885e-09, 4.10476e-09, 
    4.737009e-09, 4.172946e-09, 4.243886e-09, 4.270673e-09, 4.299533e-09,
  1.548619e-08, 1.299649e-08, 1.041311e-08, 7.61433e-09, 6.104119e-09, 
    5.598676e-09, 5.063947e-09, 4.313329e-09, 3.849972e-09, 3.980756e-09, 
    4.780549e-09, 4.271226e-09, 4.294331e-09, 4.331153e-09, 4.310917e-09,
  1.659499e-08, 1.391707e-08, 1.120695e-08, 8.385951e-09, 6.532924e-09, 
    5.91031e-09, 5.528137e-09, 4.742319e-09, 4.071875e-09, 3.958927e-09, 
    4.76034e-09, 4.27944e-09, 4.219517e-09, 4.278054e-09, 4.295906e-09,
  1.007379e-08, 7.35205e-09, 5.377621e-09, 3.991105e-09, 3.347615e-09, 
    3.085744e-09, 2.930564e-09, 3.054538e-09, 3.260569e-09, 3.051718e-09, 
    2.862266e-09, 2.696563e-09, 2.539279e-09, 2.387657e-09, 2.164217e-09,
  1.114006e-08, 8.680204e-09, 6.442278e-09, 4.716139e-09, 3.786248e-09, 
    3.272967e-09, 3.088492e-09, 3.178029e-09, 3.348431e-09, 3.314828e-09, 
    2.990761e-09, 2.761255e-09, 2.638043e-09, 2.5283e-09, 2.357021e-09,
  1.224742e-08, 9.816851e-09, 7.575137e-09, 5.602937e-09, 4.294247e-09, 
    3.595406e-09, 3.252661e-09, 3.254986e-09, 3.375055e-09, 3.46108e-09, 
    3.119249e-09, 2.756776e-09, 2.683745e-09, 2.640814e-09, 2.461867e-09,
  1.33769e-08, 1.090546e-08, 8.624628e-09, 6.552802e-09, 4.986519e-09, 
    4.036163e-09, 3.451022e-09, 3.286863e-09, 3.321989e-09, 3.393734e-09, 
    3.223768e-09, 2.75093e-09, 2.710965e-09, 2.720461e-09, 2.523329e-09,
  1.472235e-08, 1.179228e-08, 9.549506e-09, 7.491137e-09, 5.695807e-09, 
    4.529862e-09, 3.685226e-09, 3.393059e-09, 3.347808e-09, 3.35171e-09, 
    3.268517e-09, 2.869356e-09, 2.696704e-09, 2.746373e-09, 2.584316e-09,
  1.559738e-08, 1.276223e-08, 1.033412e-08, 8.240365e-09, 6.466572e-09, 
    5.16534e-09, 4.070388e-09, 3.546421e-09, 3.369381e-09, 3.320301e-09, 
    3.246688e-09, 3.02281e-09, 2.771541e-09, 2.732973e-09, 2.61012e-09,
  1.670908e-08, 1.392573e-08, 1.131523e-08, 9.03328e-09, 7.040982e-09, 
    5.634706e-09, 4.575635e-09, 3.873974e-09, 3.563636e-09, 3.408594e-09, 
    3.219106e-09, 3.121592e-09, 2.886609e-09, 2.781048e-09, 2.644842e-09,
  1.724964e-08, 1.487156e-08, 1.224181e-08, 9.773614e-09, 7.810375e-09, 
    6.107854e-09, 4.805127e-09, 3.990644e-09, 3.693184e-09, 3.51742e-09, 
    3.257944e-09, 3.197411e-09, 2.981824e-09, 2.814423e-09, 2.650661e-09,
  1.762102e-08, 1.571561e-08, 1.322168e-08, 1.057881e-08, 8.420251e-09, 
    6.848814e-09, 5.418031e-09, 4.26614e-09, 3.778478e-09, 3.555019e-09, 
    3.299079e-09, 3.248219e-09, 3.070515e-09, 2.859105e-09, 2.642798e-09,
  1.803746e-08, 1.63601e-08, 1.407783e-08, 1.148289e-08, 9.021962e-09, 
    7.259724e-09, 5.9378e-09, 4.71479e-09, 3.964514e-09, 3.650651e-09, 
    3.367176e-09, 3.271087e-09, 3.132062e-09, 2.968663e-09, 2.714837e-09,
  1.200303e-08, 8.717308e-09, 6.46096e-09, 4.715556e-09, 3.443043e-09, 
    2.698336e-09, 2.206198e-09, 1.918027e-09, 1.592208e-09, 1.466712e-09, 
    1.524639e-09, 1.546422e-09, 1.119503e-09, 7.457981e-10, 5.264711e-10,
  1.230664e-08, 9.214836e-09, 6.7646e-09, 4.90539e-09, 3.612967e-09, 
    2.843595e-09, 2.287897e-09, 2.148809e-09, 1.858111e-09, 1.451214e-09, 
    1.34418e-09, 1.265513e-09, 1.3665e-09, 1.184208e-09, 9.37927e-10,
  1.241899e-08, 9.519376e-09, 7.03093e-09, 5.005724e-09, 3.705089e-09, 
    2.859304e-09, 2.315197e-09, 2.272179e-09, 2.150374e-09, 1.557881e-09, 
    1.2953e-09, 1.180759e-09, 1.204239e-09, 1.345959e-09, 1.250541e-09,
  1.256116e-08, 9.835775e-09, 7.320874e-09, 5.07502e-09, 3.69239e-09, 
    2.869769e-09, 2.412172e-09, 2.436837e-09, 2.496984e-09, 1.881672e-09, 
    1.39179e-09, 1.19128e-09, 1.197074e-09, 1.277594e-09, 1.349411e-09,
  1.255544e-08, 9.964888e-09, 7.526368e-09, 5.192659e-09, 3.745166e-09, 
    2.841348e-09, 2.437061e-09, 2.589757e-09, 2.685036e-09, 2.216711e-09, 
    1.603164e-09, 1.289786e-09, 1.216455e-09, 1.287505e-09, 1.333555e-09,
  1.274032e-08, 1.005529e-08, 7.625708e-09, 5.31606e-09, 3.77863e-09, 
    2.925143e-09, 2.46949e-09, 2.67884e-09, 2.841624e-09, 2.425787e-09, 
    1.775694e-09, 1.460619e-09, 1.354539e-09, 1.349733e-09, 1.369768e-09,
  1.25809e-08, 9.729617e-09, 7.45809e-09, 5.371918e-09, 3.687742e-09, 
    2.880096e-09, 2.593977e-09, 2.825967e-09, 3.088009e-09, 2.669752e-09, 
    2.038208e-09, 1.730063e-09, 1.532178e-09, 1.485173e-09, 1.478807e-09,
  1.224438e-08, 9.513273e-09, 7.407441e-09, 5.421489e-09, 3.578176e-09, 
    2.870529e-09, 2.795161e-09, 3.096889e-09, 3.485853e-09, 2.963511e-09, 
    2.280053e-09, 1.994798e-09, 1.740422e-09, 1.635607e-09, 1.617388e-09,
  1.229113e-08, 9.634664e-09, 7.529155e-09, 5.423062e-09, 3.576181e-09, 
    3.249727e-09, 3.297123e-09, 3.262348e-09, 3.533647e-09, 3.071767e-09, 
    2.487833e-09, 2.278101e-09, 2.003616e-09, 1.858744e-09, 1.800754e-09,
  1.234256e-08, 9.858096e-09, 7.724997e-09, 5.636036e-09, 3.808582e-09, 
    3.373468e-09, 3.611133e-09, 3.457967e-09, 3.574195e-09, 3.208362e-09, 
    2.660819e-09, 2.462207e-09, 2.234345e-09, 2.065095e-09, 1.956913e-09,
  2.63908e-08, 2.221625e-08, 1.932457e-08, 1.586763e-08, 1.125937e-08, 
    7.45261e-09, 4.93636e-09, 3.138904e-09, 2.099854e-09, 1.421327e-09, 
    1.04944e-09, 8.638095e-10, 5.659157e-10, 4.293096e-10, 3.466095e-10,
  2.670307e-08, 2.359389e-08, 1.988687e-08, 1.684093e-08, 1.239964e-08, 
    8.370952e-09, 5.675134e-09, 3.719237e-09, 2.521104e-09, 1.731292e-09, 
    1.233512e-09, 1.037477e-09, 7.225802e-10, 5.62088e-10, 4.111442e-10,
  2.685413e-08, 2.436665e-08, 2.047027e-08, 1.760132e-08, 1.339457e-08, 
    9.118593e-09, 6.247999e-09, 4.284945e-09, 2.986885e-09, 2.110753e-09, 
    1.466472e-09, 1.207782e-09, 9.262646e-10, 6.893617e-10, 5.215188e-10,
  2.662639e-08, 2.47992e-08, 2.081517e-08, 1.799176e-08, 1.414184e-08, 
    9.754562e-09, 6.702658e-09, 4.724475e-09, 3.378305e-09, 2.467822e-09, 
    1.769943e-09, 1.399607e-09, 1.096842e-09, 8.758773e-10, 6.618395e-10,
  2.77104e-08, 2.481511e-08, 2.083858e-08, 1.809236e-08, 1.455418e-08, 
    1.019103e-08, 7.132339e-09, 5.162959e-09, 3.762925e-09, 2.778437e-09, 
    2.061778e-09, 1.584812e-09, 1.274387e-09, 1.075458e-09, 8.57706e-10,
  2.823483e-08, 2.455788e-08, 2.068924e-08, 1.795935e-08, 1.478973e-08, 
    1.050721e-08, 7.391955e-09, 5.437578e-09, 4.097461e-09, 2.99896e-09, 
    2.281148e-09, 1.771282e-09, 1.466027e-09, 1.288338e-09, 1.097838e-09,
  2.743407e-08, 2.406344e-08, 2.04043e-08, 1.774495e-08, 1.462215e-08, 
    1.062701e-08, 7.614218e-09, 5.703383e-09, 4.316595e-09, 3.108027e-09, 
    2.39592e-09, 1.931665e-09, 1.581782e-09, 1.507295e-09, 1.314557e-09,
  2.64521e-08, 2.383227e-08, 2.028474e-08, 1.741268e-08, 1.450604e-08, 
    1.064295e-08, 7.830768e-09, 5.949514e-09, 4.460879e-09, 3.06175e-09, 
    2.36711e-09, 2.046215e-09, 1.656145e-09, 1.60819e-09, 1.484649e-09,
  2.702133e-08, 2.386771e-08, 2.004843e-08, 1.697315e-08, 1.403635e-08, 
    1.042837e-08, 7.702778e-09, 5.852858e-09, 4.296129e-09, 2.917387e-09, 
    2.313581e-09, 2.097843e-09, 1.795499e-09, 1.673657e-09, 1.607269e-09,
  2.773828e-08, 2.34874e-08, 1.956674e-08, 1.640976e-08, 1.371521e-08, 
    1.007359e-08, 7.097825e-09, 5.341977e-09, 4.01654e-09, 2.854029e-09, 
    2.268703e-09, 2.05487e-09, 1.931636e-09, 1.751319e-09, 1.690555e-09,
  2.679755e-08, 2.761335e-08, 2.671065e-08, 2.512756e-08, 2.182126e-08, 
    1.510501e-08, 1.054536e-08, 7.468532e-09, 5.732069e-09, 3.840424e-09, 
    2.471807e-09, 1.765724e-09, 1.278905e-09, 1.022437e-09, 8.700244e-10,
  2.641975e-08, 2.769169e-08, 2.799576e-08, 2.619036e-08, 2.426243e-08, 
    1.938891e-08, 1.371078e-08, 9.770424e-09, 6.971547e-09, 5.168725e-09, 
    3.356685e-09, 2.370363e-09, 1.680266e-09, 1.236605e-09, 1.013375e-09,
  2.688494e-08, 2.640024e-08, 2.827035e-08, 2.763776e-08, 2.561446e-08, 
    2.255293e-08, 1.667587e-08, 1.2288e-08, 8.729205e-09, 6.495761e-09, 
    4.526339e-09, 3.052121e-09, 2.212339e-09, 1.581621e-09, 1.217364e-09,
  2.770629e-08, 2.646712e-08, 2.820133e-08, 2.798551e-08, 2.722324e-08, 
    2.440641e-08, 1.951891e-08, 1.442754e-08, 1.064503e-08, 7.786967e-09, 
    5.750472e-09, 3.912317e-09, 2.805992e-09, 2.038336e-09, 1.540979e-09,
  2.878249e-08, 2.701606e-08, 2.7214e-08, 2.838956e-08, 2.839105e-08, 
    2.555791e-08, 2.172229e-08, 1.651068e-08, 1.235996e-08, 9.440622e-09, 
    7.0191e-09, 4.92799e-09, 3.470906e-09, 2.507532e-09, 1.921501e-09,
  2.996481e-08, 2.853293e-08, 2.732783e-08, 2.849723e-08, 2.90128e-08, 
    2.74031e-08, 2.321753e-08, 1.794394e-08, 1.34735e-08, 1.067133e-08, 
    8.256611e-09, 6.035874e-09, 4.270909e-09, 3.039222e-09, 2.296162e-09,
  2.809309e-08, 2.855225e-08, 2.739951e-08, 2.807433e-08, 2.912519e-08, 
    2.859804e-08, 2.478123e-08, 1.996217e-08, 1.487634e-08, 1.172762e-08, 
    9.372678e-09, 7.027432e-09, 5.109801e-09, 3.647274e-09, 2.690972e-09,
  2.750961e-08, 2.869742e-08, 2.748057e-08, 2.74267e-08, 2.94747e-08, 
    2.894234e-08, 2.583924e-08, 2.07037e-08, 1.560119e-08, 1.221253e-08, 
    1.013247e-08, 7.872376e-09, 5.825895e-09, 4.22528e-09, 3.113152e-09,
  2.711326e-08, 2.89263e-08, 2.804951e-08, 2.717416e-08, 2.880302e-08, 
    2.9422e-08, 2.681035e-08, 2.112393e-08, 1.630908e-08, 1.255408e-08, 
    1.052216e-08, 8.394084e-09, 6.360379e-09, 4.739614e-09, 3.490909e-09,
  2.918865e-08, 2.90029e-08, 2.817399e-08, 2.690953e-08, 2.845809e-08, 
    2.978613e-08, 2.713637e-08, 2.104378e-08, 1.667389e-08, 1.270341e-08, 
    1.062302e-08, 8.729138e-09, 6.713815e-09, 5.139016e-09, 3.801248e-09,
  2.582724e-08, 2.353584e-08, 1.975566e-08, 1.493724e-08, 9.748935e-09, 
    6.034891e-09, 3.852781e-09, 2.791197e-09, 1.94279e-09, 1.106958e-09, 
    7.651808e-10, 6.595275e-10, 6.646255e-10, 6.268827e-10, 5.392403e-10,
  2.510065e-08, 2.533454e-08, 2.280936e-08, 1.92937e-08, 1.450809e-08, 
    9.660448e-09, 5.94526e-09, 3.977454e-09, 2.852836e-09, 1.939076e-09, 
    1.129344e-09, 8.575654e-10, 7.243662e-10, 7.095636e-10, 6.455671e-10,
  2.367241e-08, 2.545796e-08, 2.502809e-08, 2.22118e-08, 1.8666e-08, 
    1.406042e-08, 9.271004e-09, 5.907635e-09, 4.041633e-09, 2.980368e-09, 
    1.958018e-09, 1.200502e-09, 9.385053e-10, 8.310462e-10, 7.772356e-10,
  2.31853e-08, 2.411653e-08, 2.543238e-08, 2.438145e-08, 2.158604e-08, 
    1.795781e-08, 1.336003e-08, 8.98079e-09, 5.746049e-09, 3.920097e-09, 
    2.92218e-09, 1.88744e-09, 1.313407e-09, 1.060219e-09, 9.34325e-10,
  2.335216e-08, 2.365768e-08, 2.420921e-08, 2.517191e-08, 2.388516e-08, 
    2.101851e-08, 1.710491e-08, 1.275213e-08, 8.920185e-09, 5.93001e-09, 
    4.015617e-09, 2.870278e-09, 1.82191e-09, 1.423563e-09, 1.197666e-09,
  2.418633e-08, 2.381254e-08, 2.390215e-08, 2.442328e-08, 2.502136e-08, 
    2.344158e-08, 2.030335e-08, 1.614531e-08, 1.181243e-08, 8.325343e-09, 
    5.701849e-09, 4.086605e-09, 2.729659e-09, 1.92619e-09, 1.568226e-09,
  2.455164e-08, 2.384389e-08, 2.406317e-08, 2.399074e-08, 2.48614e-08, 
    2.460425e-08, 2.292017e-08, 1.974641e-08, 1.570938e-08, 1.138876e-08, 
    7.942618e-09, 5.502339e-09, 3.982848e-09, 2.613306e-09, 2.055595e-09,
  2.597212e-08, 2.481662e-08, 2.455515e-08, 2.392263e-08, 2.434856e-08, 
    2.491261e-08, 2.425852e-08, 2.215413e-08, 1.891294e-08, 1.48993e-08, 
    1.081886e-08, 7.487535e-09, 5.417351e-09, 3.632312e-09, 2.728419e-09,
  2.768706e-08, 2.60245e-08, 2.486049e-08, 2.433407e-08, 2.402528e-08, 
    2.487843e-08, 2.534559e-08, 2.379207e-08, 2.103292e-08, 1.776651e-08, 
    1.392882e-08, 9.947177e-09, 6.995084e-09, 4.969091e-09, 3.485545e-09,
  2.886238e-08, 2.745145e-08, 2.593131e-08, 2.481467e-08, 2.441037e-08, 
    2.4728e-08, 2.555184e-08, 2.519468e-08, 2.296341e-08, 2.007268e-08, 
    1.668797e-08, 1.27247e-08, 8.883041e-09, 6.443241e-09, 4.376392e-09,
  1.290474e-08, 1.040775e-08, 6.422978e-09, 4.001923e-09, 2.506175e-09, 
    1.740967e-09, 1.311235e-09, 1.141055e-09, 9.759117e-10, 7.556999e-10, 
    3.640876e-10, 1.522944e-10, 1.045941e-10, 1.088489e-10, 2.194875e-10,
  1.51689e-08, 1.197961e-08, 9.068096e-09, 5.956959e-09, 3.634226e-09, 
    2.499838e-09, 1.788291e-09, 1.321885e-09, 1.190504e-09, 9.884426e-10, 
    6.988053e-10, 3.699428e-10, 1.556924e-10, 8.974439e-11, 1.085268e-10,
  1.774771e-08, 1.452164e-08, 1.113643e-08, 8.009351e-09, 5.442528e-09, 
    3.519343e-09, 2.498545e-09, 1.74574e-09, 1.36425e-09, 1.233827e-09, 
    1.013928e-09, 7.279056e-10, 3.926016e-10, 1.638846e-10, 9.771448e-11,
  1.903269e-08, 1.668526e-08, 1.319978e-08, 9.78461e-09, 7.300631e-09, 
    5.109305e-09, 3.580867e-09, 2.471116e-09, 1.704716e-09, 1.390255e-09, 
    1.242285e-09, 1.035792e-09, 7.5816e-10, 4.397549e-10, 2.087428e-10,
  2.104397e-08, 1.750051e-08, 1.511784e-08, 1.190646e-08, 9.001853e-09, 
    6.738313e-09, 4.944265e-09, 3.436064e-09, 2.369415e-09, 1.739571e-09, 
    1.450711e-09, 1.276623e-09, 1.093499e-09, 7.819748e-10, 4.728323e-10,
  2.227911e-08, 1.874337e-08, 1.594755e-08, 1.391092e-08, 1.100446e-08, 
    8.448342e-09, 6.581344e-09, 4.635604e-09, 3.074288e-09, 2.165235e-09, 
    1.708709e-09, 1.476774e-09, 1.391861e-09, 1.159639e-09, 7.549251e-10,
  2.3434e-08, 2.018236e-08, 1.709462e-08, 1.559072e-08, 1.321278e-08, 
    1.033418e-08, 8.182035e-09, 6.538445e-09, 4.38357e-09, 2.874549e-09, 
    2.094792e-09, 1.714169e-09, 1.612284e-09, 1.446874e-09, 1.099279e-09,
  2.498378e-08, 2.177433e-08, 1.877213e-08, 1.656812e-08, 1.508385e-08, 
    1.291421e-08, 1.009715e-08, 7.87911e-09, 5.806871e-09, 3.790942e-09, 
    2.655036e-09, 2.040805e-09, 1.795812e-09, 1.678281e-09, 1.415878e-09,
  2.656314e-08, 2.352329e-08, 2.025988e-08, 1.779445e-08, 1.639033e-08, 
    1.486561e-08, 1.247079e-08, 9.632557e-09, 7.404307e-09, 5.005361e-09, 
    3.403213e-09, 2.514804e-09, 2.081896e-09, 1.881911e-09, 1.763732e-09,
  2.822862e-08, 2.484254e-08, 2.190339e-08, 1.91138e-08, 1.729363e-08, 
    1.616686e-08, 1.457476e-08, 1.173378e-08, 9.382054e-09, 6.593693e-09, 
    4.507727e-09, 3.193847e-09, 2.544834e-09, 2.163517e-09, 2.068652e-09,
  2.234651e-08, 1.857321e-08, 1.29083e-08, 7.705e-09, 4.577825e-09, 
    2.60064e-09, 1.552473e-09, 8.317406e-10, 5.213479e-10, 3.952935e-10, 
    3.15702e-10, 2.379879e-10, 2.790338e-10, 2.870252e-10, 2.861089e-10,
  2.371907e-08, 2.062703e-08, 1.578016e-08, 1.032711e-08, 5.939898e-09, 
    3.235069e-09, 1.86901e-09, 9.947725e-10, 5.693601e-10, 4.115064e-10, 
    3.42526e-10, 2.748847e-10, 2.65087e-10, 2.853252e-10, 2.481376e-10,
  2.462519e-08, 2.251396e-08, 1.819683e-08, 1.294173e-08, 7.846366e-09, 
    4.151677e-09, 2.264217e-09, 1.207623e-09, 6.293945e-10, 4.178128e-10, 
    3.558301e-10, 3.064568e-10, 2.737239e-10, 2.758632e-10, 2.133029e-10,
  2.470508e-08, 2.312775e-08, 1.997257e-08, 1.523819e-08, 9.959454e-09, 
    5.452041e-09, 2.812854e-09, 1.431043e-09, 7.273994e-10, 4.180885e-10, 
    3.559163e-10, 3.130381e-10, 2.802682e-10, 2.616221e-10, 1.934981e-10,
  2.522172e-08, 2.365149e-08, 2.10834e-08, 1.694047e-08, 1.207407e-08, 
    7.053135e-09, 3.575203e-09, 1.836469e-09, 8.704256e-10, 4.387803e-10, 
    3.448223e-10, 3.116577e-10, 2.631008e-10, 2.252365e-10, 1.898249e-10,
  2.59178e-08, 2.393671e-08, 2.180434e-08, 1.805318e-08, 1.368797e-08, 
    8.763116e-09, 4.51086e-09, 2.222817e-09, 1.054766e-09, 5.045104e-10, 
    3.307582e-10, 3.038155e-10, 2.483947e-10, 2.21047e-10, 2.286567e-10,
  2.63224e-08, 2.468601e-08, 2.250937e-08, 1.902419e-08, 1.479832e-08, 
    1.019562e-08, 5.812399e-09, 2.738886e-09, 1.273011e-09, 5.720863e-10, 
    3.27652e-10, 2.828978e-10, 2.498326e-10, 2.214453e-10, 2.751839e-10,
  2.625054e-08, 2.516081e-08, 2.330749e-08, 2.01212e-08, 1.561555e-08, 
    1.138667e-08, 6.935514e-09, 3.527199e-09, 1.692475e-09, 6.912354e-10, 
    3.360746e-10, 2.559487e-10, 2.450496e-10, 2.124808e-10, 2.366837e-10,
  2.625298e-08, 2.528502e-08, 2.369067e-08, 2.116933e-08, 1.655787e-08, 
    1.219769e-08, 7.947771e-09, 4.427036e-09, 2.09085e-09, 8.187103e-10, 
    3.609119e-10, 2.477843e-10, 2.501452e-10, 2.19013e-10, 2.023831e-10,
  2.620714e-08, 2.517503e-08, 2.396042e-08, 2.188516e-08, 1.739514e-08, 
    1.279689e-08, 8.487796e-09, 5.035499e-09, 2.42083e-09, 9.771687e-10, 
    4.220645e-10, 2.520162e-10, 2.566068e-10, 2.373077e-10, 1.97128e-10,
  1.320634e-08, 1.130323e-08, 9.980114e-09, 8.572673e-09, 7.133821e-09, 
    5.436197e-09, 3.827958e-09, 2.68884e-09, 2.195908e-09, 1.459908e-09, 
    8.921787e-10, 5.321129e-10, 3.372105e-10, 1.684772e-10, 1.5219e-10,
  1.468988e-08, 1.27329e-08, 1.100582e-08, 9.630618e-09, 8.27168e-09, 
    6.653835e-09, 4.858793e-09, 3.279316e-09, 2.451196e-09, 1.827867e-09, 
    1.060434e-09, 6.499831e-10, 4.194364e-10, 2.538581e-10, 1.951501e-10,
  1.662877e-08, 1.461846e-08, 1.244101e-08, 1.06977e-08, 9.316981e-09, 
    7.813101e-09, 6.031397e-09, 4.151188e-09, 2.884968e-09, 2.233194e-09, 
    1.381279e-09, 7.861034e-10, 4.988971e-10, 3.307446e-10, 2.293559e-10,
  1.814597e-08, 1.636026e-08, 1.424189e-08, 1.203634e-08, 1.034284e-08, 
    8.844729e-09, 7.273489e-09, 5.213157e-09, 3.554966e-09, 2.569545e-09, 
    1.81863e-09, 1.034025e-09, 6.086599e-10, 3.917957e-10, 2.706357e-10,
  1.998727e-08, 1.807701e-08, 1.609319e-08, 1.353267e-08, 1.15542e-08, 
    9.814268e-09, 8.301166e-09, 6.454634e-09, 4.511352e-09, 3.05323e-09, 
    2.20785e-09, 1.400948e-09, 7.589641e-10, 4.69212e-10, 3.144074e-10,
  2.100968e-08, 1.90079e-08, 1.764891e-08, 1.538315e-08, 1.302597e-08, 
    1.103459e-08, 9.319566e-09, 7.428628e-09, 5.480012e-09, 3.722616e-09, 
    2.578534e-09, 1.763559e-09, 1.024573e-09, 5.683432e-10, 3.696929e-10,
  2.26102e-08, 2.005081e-08, 1.873697e-08, 1.719398e-08, 1.493203e-08, 
    1.238887e-08, 1.037273e-08, 8.724594e-09, 6.588733e-09, 4.597644e-09, 
    3.058385e-09, 2.075457e-09, 1.321624e-09, 7.37322e-10, 4.351671e-10,
  2.427036e-08, 2.209777e-08, 2.00902e-08, 1.868762e-08, 1.703012e-08, 
    1.441136e-08, 1.163454e-08, 9.746257e-09, 7.656532e-09, 5.528127e-09, 
    3.675126e-09, 2.459662e-09, 1.557913e-09, 9.273141e-10, 5.122329e-10,
  2.626416e-08, 2.422177e-08, 2.20141e-08, 2.006423e-08, 1.854567e-08, 
    1.633343e-08, 1.331414e-08, 1.085926e-08, 8.854729e-09, 6.636849e-09, 
    4.473591e-09, 2.918734e-09, 1.844998e-09, 1.141593e-09, 6.136553e-10,
  2.718534e-08, 2.584884e-08, 2.359654e-08, 2.128574e-08, 1.992155e-08, 
    1.842455e-08, 1.520712e-08, 1.214937e-08, 9.732294e-09, 7.608564e-09, 
    5.394158e-09, 3.471287e-09, 2.188808e-09, 1.358345e-09, 7.595432e-10,
  1.265991e-08, 9.18336e-09, 6.882043e-09, 5.158708e-09, 3.504286e-09, 
    2.579152e-09, 1.983486e-09, 1.623835e-09, 1.339117e-09, 1.067719e-09, 
    8.172689e-10, 6.051983e-10, 3.937931e-10, 3.528019e-10, 2.286266e-10,
  1.442838e-08, 1.090835e-08, 8.024727e-09, 6.020529e-09, 4.284068e-09, 
    3.00636e-09, 2.271828e-09, 1.761025e-09, 1.469388e-09, 1.211196e-09, 
    1.018222e-09, 7.939513e-10, 5.051263e-10, 3.58805e-10, 2.600676e-10,
  1.562032e-08, 1.267576e-08, 9.505564e-09, 7.035568e-09, 5.063217e-09, 
    3.541435e-09, 2.623093e-09, 1.98673e-09, 1.593715e-09, 1.360962e-09, 
    1.159246e-09, 9.531421e-10, 6.694468e-10, 4.099266e-10, 2.831126e-10,
  1.6466e-08, 1.398514e-08, 1.096782e-08, 8.252737e-09, 5.9922e-09, 
    4.220209e-09, 3.052317e-09, 2.285156e-09, 1.742968e-09, 1.481438e-09, 
    1.255911e-09, 1.079899e-09, 8.444541e-10, 5.24397e-10, 3.225596e-10,
  1.758084e-08, 1.48675e-08, 1.200035e-08, 9.425489e-09, 7.053487e-09, 
    4.98149e-09, 3.523628e-09, 2.673654e-09, 2.003386e-09, 1.607044e-09, 
    1.352167e-09, 1.131429e-09, 9.72539e-10, 6.909562e-10, 3.990585e-10,
  1.813356e-08, 1.520874e-08, 1.254505e-08, 1.020118e-08, 8.138551e-09, 
    5.9256e-09, 4.106565e-09, 3.003471e-09, 2.242409e-09, 1.745572e-09, 
    1.44948e-09, 1.176336e-09, 1.042149e-09, 8.612078e-10, 5.564319e-10,
  1.828308e-08, 1.592639e-08, 1.329137e-08, 1.088314e-08, 8.856161e-09, 
    6.761587e-09, 4.834216e-09, 3.505933e-09, 2.593557e-09, 1.932342e-09, 
    1.569348e-09, 1.306292e-09, 1.096624e-09, 1.056178e-09, 7.486124e-10,
  1.859345e-08, 1.665738e-08, 1.416541e-08, 1.167179e-08, 9.540224e-09, 
    7.624971e-09, 5.669991e-09, 4.045829e-09, 2.951854e-09, 2.156941e-09, 
    1.67462e-09, 1.38009e-09, 1.188358e-09, 1.024295e-09, 8.188404e-10,
  1.942944e-08, 1.765364e-08, 1.511004e-08, 1.248094e-08, 1.017367e-08, 
    8.308e-09, 6.3352e-09, 4.663115e-09, 3.381597e-09, 2.447595e-09, 
    1.829717e-09, 1.456303e-09, 1.313132e-09, 1.092062e-09, 9.493457e-10,
  1.965959e-08, 1.817763e-08, 1.607284e-08, 1.322561e-08, 1.073569e-08, 
    8.992822e-09, 6.92639e-09, 5.1874e-09, 3.919367e-09, 2.804543e-09, 
    2.000506e-09, 1.555182e-09, 1.392635e-09, 1.160396e-09, 1.108916e-09,
  1.855759e-08, 1.248862e-08, 8.062214e-09, 5.823479e-09, 3.495638e-09, 
    2.426359e-09, 1.991185e-09, 1.925289e-09, 1.782994e-09, 1.642941e-09, 
    1.275375e-09, 8.319697e-10, 6.122251e-10, 6.248986e-10, 5.962927e-10,
  2.216399e-08, 1.626097e-08, 1.074148e-08, 7.32491e-09, 4.698511e-09, 
    3.055302e-09, 2.206374e-09, 1.958051e-09, 1.831752e-09, 1.7474e-09, 
    1.414836e-09, 9.857497e-10, 6.621428e-10, 6.337462e-10, 6.107407e-10,
  2.530047e-08, 2.01513e-08, 1.404762e-08, 9.363673e-09, 6.087101e-09, 
    3.93285e-09, 2.609918e-09, 2.074794e-09, 1.934559e-09, 1.860946e-09, 
    1.51518e-09, 1.127163e-09, 7.86026e-10, 6.68976e-10, 6.458644e-10,
  2.743819e-08, 2.208768e-08, 1.723458e-08, 1.224836e-08, 7.904656e-09, 
    5.068594e-09, 3.328614e-09, 2.321836e-09, 2.010365e-09, 1.899677e-09, 
    1.666492e-09, 1.256624e-09, 9.397434e-10, 7.244794e-10, 6.888852e-10,
  2.946505e-08, 2.409086e-08, 1.91262e-08, 1.506178e-08, 1.038266e-08, 
    6.563452e-09, 4.267852e-09, 2.832832e-09, 2.198696e-09, 2.000252e-09, 
    1.827786e-09, 1.440793e-09, 1.121656e-09, 8.329478e-10, 7.185498e-10,
  3.092205e-08, 2.622737e-08, 2.109937e-08, 1.675681e-08, 1.276804e-08, 
    8.533667e-09, 5.510095e-09, 3.433486e-09, 2.368066e-09, 2.077291e-09, 
    1.921841e-09, 1.666653e-09, 1.296065e-09, 9.730493e-10, 7.60577e-10,
  3.054368e-08, 2.780022e-08, 2.27998e-08, 1.821645e-08, 1.424013e-08, 
    1.029987e-08, 6.913546e-09, 4.514562e-09, 2.829206e-09, 2.19097e-09, 
    1.930043e-09, 1.856837e-09, 1.511892e-09, 1.144575e-09, 8.606737e-10,
  2.95295e-08, 2.828697e-08, 2.429991e-08, 1.951433e-08, 1.535988e-08, 
    1.186453e-08, 8.251454e-09, 5.472625e-09, 3.534855e-09, 2.350675e-09, 
    1.922267e-09, 1.955381e-09, 1.790705e-09, 1.331137e-09, 9.96118e-10,
  2.910749e-08, 2.849353e-08, 2.585696e-08, 2.079314e-08, 1.617818e-08, 
    1.24867e-08, 9.455232e-09, 6.48328e-09, 4.104022e-09, 2.361122e-09, 
    1.901472e-09, 2.025715e-09, 1.990507e-09, 1.526249e-09, 1.134864e-09,
  2.937876e-08, 2.794951e-08, 2.608351e-08, 2.176005e-08, 1.722313e-08, 
    1.310003e-08, 9.998926e-09, 7.337979e-09, 4.807031e-09, 2.779898e-09, 
    2.122324e-09, 2.051908e-09, 2.067284e-09, 1.704186e-09, 1.273236e-09,
  5.423514e-09, 4.718796e-09, 4.605285e-09, 4.339961e-09, 3.268162e-09, 
    2.647513e-09, 2.422391e-09, 2.499695e-09, 2.443111e-09, 2.226619e-09, 
    2.047012e-09, 1.861031e-09, 1.839635e-09, 1.701624e-09, 1.322968e-09,
  6.406133e-09, 5.66219e-09, 4.912439e-09, 4.458784e-09, 4.041257e-09, 
    3.172666e-09, 2.552635e-09, 2.442385e-09, 2.533624e-09, 2.43142e-09, 
    2.142512e-09, 1.94381e-09, 1.833662e-09, 1.846236e-09, 1.595191e-09,
  7.876208e-09, 6.864359e-09, 5.840445e-09, 4.98843e-09, 4.486733e-09, 
    3.817472e-09, 3.048722e-09, 2.494996e-09, 2.464606e-09, 2.541568e-09, 
    2.375854e-09, 2.084349e-09, 1.86648e-09, 1.832389e-09, 1.793397e-09,
  1.03623e-08, 8.492573e-09, 6.785179e-09, 5.668662e-09, 5.035836e-09, 
    4.549837e-09, 3.654111e-09, 2.946419e-09, 2.509991e-09, 2.450947e-09, 
    2.529073e-09, 2.317218e-09, 2.034242e-09, 1.854011e-09, 1.825057e-09,
  1.394794e-08, 1.106013e-08, 8.818274e-09, 6.710305e-09, 5.680381e-09, 
    5.223374e-09, 4.500938e-09, 3.515346e-09, 2.843599e-09, 2.543218e-09, 
    2.501453e-09, 2.483726e-09, 2.213272e-09, 1.951938e-09, 1.826148e-09,
  1.710069e-08, 1.358714e-08, 1.07589e-08, 8.741118e-09, 6.971225e-09, 
    6.026529e-09, 5.449786e-09, 4.335162e-09, 3.285868e-09, 2.704818e-09, 
    2.53601e-09, 2.492963e-09, 2.370992e-09, 2.101227e-09, 1.892593e-09,
  2.000906e-08, 1.655665e-08, 1.260293e-08, 1.039657e-08, 8.961988e-09, 
    7.21818e-09, 6.245601e-09, 5.487284e-09, 4.210943e-09, 3.141043e-09, 
    2.573054e-09, 2.569624e-09, 2.420429e-09, 2.217429e-09, 1.977925e-09,
  2.501785e-08, 2.194379e-08, 1.783897e-08, 1.324804e-08, 1.10311e-08, 
    9.377914e-09, 7.431936e-09, 6.24052e-09, 5.037438e-09, 3.789923e-09, 
    2.795421e-09, 2.441212e-09, 2.420464e-09, 2.321455e-09, 2.09827e-09,
  2.779538e-08, 2.623871e-08, 2.275122e-08, 1.814698e-08, 1.418478e-08, 
    1.164068e-08, 9.509038e-09, 7.221982e-09, 5.989282e-09, 4.529639e-09, 
    3.293118e-09, 2.505457e-09, 2.275106e-09, 2.315671e-09, 2.222202e-09,
  3.162701e-08, 2.879876e-08, 2.708894e-08, 2.378257e-08, 1.968498e-08, 
    1.566544e-08, 1.210302e-08, 9.095524e-09, 7.240575e-09, 5.850758e-09, 
    3.936437e-09, 2.873392e-09, 2.261497e-09, 2.162415e-09, 2.200879e-09,
  6.229779e-09, 4.672016e-09, 3.99486e-09, 3.552862e-09, 3.429659e-09, 
    3.440205e-09, 3.199103e-09, 2.768704e-09, 2.146868e-09, 1.887154e-09, 
    2.12742e-09, 2.11296e-09, 1.834444e-09, 1.602349e-09, 1.409006e-09,
  7.500461e-09, 5.631855e-09, 4.405924e-09, 3.732651e-09, 3.345644e-09, 
    3.31956e-09, 3.355893e-09, 3.138332e-09, 2.674334e-09, 2.084405e-09, 
    1.916839e-09, 2.029801e-09, 2.088371e-09, 1.863062e-09, 1.65419e-09,
  9.103064e-09, 6.893345e-09, 5.260018e-09, 4.157429e-09, 3.558774e-09, 
    3.22539e-09, 3.247622e-09, 3.270548e-09, 3.111504e-09, 2.600639e-09, 
    2.121203e-09, 1.918444e-09, 2.034893e-09, 2.079671e-09, 1.895443e-09,
  1.106341e-08, 8.453304e-09, 6.45905e-09, 4.903536e-09, 3.941495e-09, 
    3.432342e-09, 3.212561e-09, 3.158386e-09, 3.223121e-09, 3.052999e-09, 
    2.55968e-09, 2.133669e-09, 1.965114e-09, 2.074199e-09, 2.074486e-09,
  1.428518e-08, 1.052567e-08, 8.05621e-09, 6.057844e-09, 4.681191e-09, 
    3.772584e-09, 3.380298e-09, 3.154241e-09, 3.171448e-09, 3.307971e-09, 
    3.00769e-09, 2.543293e-09, 2.16454e-09, 2.02293e-09, 2.078151e-09,
  1.679696e-08, 1.264676e-08, 9.767652e-09, 7.430098e-09, 5.761112e-09, 
    4.52932e-09, 3.769843e-09, 3.372358e-09, 3.082307e-09, 3.269197e-09, 
    3.384492e-09, 3.003356e-09, 2.576321e-09, 2.223881e-09, 2.032811e-09,
  1.87665e-08, 1.542356e-08, 1.185948e-08, 9.057457e-09, 6.863937e-09, 
    5.480906e-09, 4.44043e-09, 3.910932e-09, 3.491852e-09, 3.215597e-09, 
    3.456381e-09, 3.436849e-09, 3.055532e-09, 2.652526e-09, 2.290551e-09,
  2.010138e-08, 1.745489e-08, 1.444386e-08, 1.111084e-08, 8.426554e-09, 
    6.566946e-09, 5.303817e-09, 4.453979e-09, 4.084048e-09, 3.611314e-09, 
    3.439642e-09, 3.640442e-09, 3.434094e-09, 3.004705e-09, 2.65639e-09,
  2.162826e-08, 1.923157e-08, 1.635414e-08, 1.327363e-08, 1.034177e-08, 
    8.235615e-09, 6.637509e-09, 5.294655e-09, 4.543474e-09, 4.121066e-09, 
    3.731883e-09, 3.70656e-09, 3.758458e-09, 3.292657e-09, 2.957508e-09,
  2.291615e-08, 2.065852e-08, 1.847581e-08, 1.542979e-08, 1.252702e-08, 
    9.869335e-09, 8.232496e-09, 6.606179e-09, 5.371139e-09, 4.744082e-09, 
    4.170287e-09, 3.931819e-09, 3.891631e-09, 3.583696e-09, 3.121392e-09,
  1.092603e-08, 8.70168e-09, 7.313486e-09, 5.962068e-09, 5.016708e-09, 
    3.938018e-09, 2.579679e-09, 1.916867e-09, 2.014556e-09, 2.588157e-09, 
    2.838902e-09, 2.415362e-09, 1.887749e-09, 1.445664e-09, 1.187198e-09,
  1.284225e-08, 1.017775e-08, 8.273078e-09, 6.959123e-09, 5.85551e-09, 
    4.944037e-09, 3.85559e-09, 2.49781e-09, 1.993637e-09, 1.863236e-09, 
    2.365856e-09, 2.466051e-09, 2.372869e-09, 2.057797e-09, 1.711105e-09,
  1.686911e-08, 1.256995e-08, 9.763714e-09, 7.965108e-09, 6.593653e-09, 
    5.67541e-09, 4.915507e-09, 3.637178e-09, 2.369291e-09, 1.858955e-09, 
    1.807676e-09, 2.259013e-09, 2.401727e-09, 2.401488e-09, 2.200737e-09,
  1.951841e-08, 1.563528e-08, 1.194611e-08, 9.42075e-09, 7.761757e-09, 
    6.282036e-09, 5.698454e-09, 5.011275e-09, 3.536868e-09, 2.357711e-09, 
    1.751919e-09, 1.69365e-09, 2.045084e-09, 2.348442e-09, 2.471952e-09,
  2.217579e-08, 1.871406e-08, 1.488219e-08, 1.135056e-08, 9.162442e-09, 
    7.328133e-09, 6.251148e-09, 5.608832e-09, 4.927641e-09, 3.563358e-09, 
    2.482547e-09, 1.843945e-09, 1.658094e-09, 1.932289e-09, 2.27992e-09,
  2.755608e-08, 2.16103e-08, 1.791286e-08, 1.369939e-08, 1.094178e-08, 
    8.741462e-09, 6.8646e-09, 5.839556e-09, 5.096124e-09, 4.560087e-09, 
    3.431087e-09, 2.620393e-09, 2.066793e-09, 1.761093e-09, 1.834142e-09,
  2.935906e-08, 2.634196e-08, 2.120939e-08, 1.667e-08, 1.2872e-08, 
    1.01064e-08, 7.922478e-09, 6.330152e-09, 5.55052e-09, 4.488629e-09, 
    4.35755e-09, 3.389723e-09, 2.802069e-09, 2.236107e-09, 1.861159e-09,
  2.907099e-08, 2.837874e-08, 2.523007e-08, 1.978422e-08, 1.59749e-08, 
    1.216922e-08, 9.312197e-09, 7.086105e-09, 6.149599e-09, 4.879988e-09, 
    4.168192e-09, 4.081463e-09, 3.433726e-09, 2.923118e-09, 2.324198e-09,
  2.812796e-08, 2.856928e-08, 2.818649e-08, 2.336061e-08, 1.832626e-08, 
    1.516709e-08, 1.155606e-08, 8.370377e-09, 6.504083e-09, 5.326768e-09, 
    4.542918e-09, 4.144717e-09, 4.069498e-09, 3.477582e-09, 2.993013e-09,
  2.663817e-08, 2.76036e-08, 2.754241e-08, 2.67733e-08, 2.106983e-08, 
    1.73267e-08, 1.403973e-08, 9.856024e-09, 7.027933e-09, 5.664805e-09, 
    4.933681e-09, 4.32733e-09, 4.123261e-09, 3.946002e-09, 3.389804e-09,
  1.651959e-08, 1.578972e-08, 1.537162e-08, 1.50669e-08, 1.390237e-08, 
    1.148975e-08, 9.055083e-09, 6.464382e-09, 5.302781e-09, 4.772632e-09, 
    4.115255e-09, 3.22372e-09, 2.600884e-09, 2.288469e-09, 1.915974e-09,
  1.706783e-08, 1.662307e-08, 1.591905e-08, 1.534928e-08, 1.503272e-08, 
    1.341636e-08, 1.194453e-08, 9.313134e-09, 6.650833e-09, 5.381997e-09, 
    4.701295e-09, 4.211431e-09, 3.466442e-09, 2.743227e-09, 2.301239e-09,
  1.692523e-08, 1.692431e-08, 1.663085e-08, 1.598374e-08, 1.555225e-08, 
    1.459244e-08, 1.342182e-08, 1.193943e-08, 9.250161e-09, 6.689515e-09, 
    5.453836e-09, 4.656704e-09, 4.07616e-09, 3.453489e-09, 2.871012e-09,
  1.622102e-08, 1.646033e-08, 1.684085e-08, 1.65845e-08, 1.614094e-08, 
    1.543386e-08, 1.435309e-08, 1.335282e-08, 1.15621e-08, 8.975966e-09, 
    6.64423e-09, 5.470401e-09, 4.67969e-09, 3.88342e-09, 3.209387e-09,
  1.543437e-08, 1.590666e-08, 1.651624e-08, 1.681835e-08, 1.663028e-08, 
    1.616877e-08, 1.506578e-08, 1.425637e-08, 1.315359e-08, 1.11536e-08, 
    8.563568e-09, 6.521196e-09, 5.215218e-09, 4.425978e-09, 3.69928e-09,
  1.568093e-08, 1.567741e-08, 1.570038e-08, 1.6347e-08, 1.647904e-08, 
    1.630672e-08, 1.559916e-08, 1.455378e-08, 1.352608e-08, 1.245717e-08, 
    1.037128e-08, 8.186934e-09, 6.304132e-09, 4.980948e-09, 4.25032e-09,
  1.739561e-08, 1.761949e-08, 1.692933e-08, 1.652211e-08, 1.673684e-08, 
    1.665248e-08, 1.616421e-08, 1.514791e-08, 1.440263e-08, 1.322277e-08, 
    1.159542e-08, 9.42777e-09, 7.775207e-09, 6.003085e-09, 4.711168e-09,
  1.797093e-08, 1.848476e-08, 1.850054e-08, 1.771941e-08, 1.727466e-08, 
    1.708629e-08, 1.70409e-08, 1.618027e-08, 1.470148e-08, 1.371194e-08, 
    1.269102e-08, 1.071672e-08, 8.727816e-09, 7.103224e-09, 5.595198e-09,
  1.875951e-08, 1.870547e-08, 1.92661e-08, 1.994112e-08, 1.914665e-08, 
    1.786205e-08, 1.765286e-08, 1.744217e-08, 1.62766e-08, 1.449639e-08, 
    1.314427e-08, 1.182919e-08, 9.907557e-09, 8.104144e-09, 6.514984e-09,
  2.052692e-08, 2.048709e-08, 2.03426e-08, 2.146822e-08, 2.109612e-08, 
    1.992913e-08, 1.894724e-08, 1.857775e-08, 1.83883e-08, 1.622364e-08, 
    1.412472e-08, 1.246087e-08, 1.072415e-08, 9.02751e-09, 7.400242e-09,
  4.224474e-09, 4.012255e-09, 3.768378e-09, 3.476066e-09, 3.164231e-09, 
    2.955623e-09, 2.750767e-09, 2.553933e-09, 2.388093e-09, 2.151149e-09, 
    1.922236e-09, 1.676838e-09, 1.4618e-09, 1.193038e-09, 1.087628e-09,
  4.690549e-09, 4.558584e-09, 4.471936e-09, 4.212153e-09, 3.945522e-09, 
    3.614872e-09, 3.364025e-09, 3.204102e-09, 3.062125e-09, 2.894106e-09, 
    2.713792e-09, 2.467796e-09, 2.285549e-09, 1.99881e-09, 1.797908e-09,
  5.349948e-09, 5.250145e-09, 5.238602e-09, 5.06003e-09, 4.810779e-09, 
    4.546552e-09, 4.202782e-09, 3.927746e-09, 3.722678e-09, 3.653757e-09, 
    3.50531e-09, 3.280915e-09, 3.128409e-09, 2.855189e-09, 2.535884e-09,
  6.188294e-09, 6.062335e-09, 5.975642e-09, 5.899838e-09, 5.679226e-09, 
    5.518279e-09, 5.297236e-09, 4.949753e-09, 4.682102e-09, 4.437987e-09, 
    4.422585e-09, 4.39729e-09, 4.3823e-09, 3.927555e-09, 3.399206e-09,
  6.937164e-09, 6.810029e-09, 6.735414e-09, 6.734991e-09, 6.699681e-09, 
    6.549484e-09, 6.459393e-09, 6.319865e-09, 6.031113e-09, 5.78834e-09, 
    5.58799e-09, 5.592302e-09, 5.507251e-09, 4.248287e-09, 3.908056e-09,
  7.976934e-09, 7.956621e-09, 7.631984e-09, 7.474886e-09, 7.57885e-09, 
    7.596373e-09, 7.677047e-09, 7.650915e-09, 7.421002e-09, 7.061612e-09, 
    6.949431e-09, 7.083822e-09, 6.025612e-09, 3.799859e-09, 4.138425e-09,
  7.636119e-09, 8.124312e-09, 8.302965e-09, 8.284228e-09, 8.522904e-09, 
    8.530918e-09, 8.535514e-09, 8.558612e-09, 8.886063e-09, 8.727148e-09, 
    8.411821e-09, 8.02104e-09, 6.863572e-09, 5.609679e-09, 5.12384e-09,
  6.841515e-09, 7.529079e-09, 8.362468e-09, 8.618005e-09, 8.755469e-09, 
    9.359479e-09, 9.700848e-09, 9.567299e-09, 9.597414e-09, 9.516383e-09, 
    9.738485e-09, 9.263323e-09, 8.695169e-09, 8.496871e-09, 7.575305e-09,
  7.380043e-09, 7.669176e-09, 8.020758e-09, 8.68018e-09, 9.017215e-09, 
    9.474137e-09, 1.026855e-08, 1.082998e-08, 1.077406e-08, 1.063721e-08, 
    1.030265e-08, 1.054422e-08, 1.040264e-08, 1.008608e-08, 1.001329e-08,
  8.146682e-09, 7.969838e-09, 7.958346e-09, 8.353347e-09, 8.850177e-09, 
    9.533576e-09, 9.839003e-09, 1.049439e-08, 1.123898e-08, 1.151785e-08, 
    1.153258e-08, 1.123497e-08, 1.13194e-08, 1.142974e-08, 1.160771e-08,
  4.426776e-09, 3.179184e-09, 2.073287e-09, 1.246035e-09, 7.56031e-10, 
    4.288008e-10, 2.832438e-10, 2.12369e-10, 1.598889e-10, 1.469742e-10, 
    1.46123e-10, 1.36072e-10, 1.111624e-10, 1.200397e-10, 1.171099e-10,
  5.124122e-09, 3.805735e-09, 2.642687e-09, 1.671957e-09, 1.061286e-09, 
    6.489106e-10, 4.020205e-10, 2.918655e-10, 2.331702e-10, 1.906404e-10, 
    1.847248e-10, 1.780404e-10, 1.560256e-10, 1.492323e-10, 1.378744e-10,
  5.677033e-09, 4.347334e-09, 3.247392e-09, 2.225806e-09, 1.494433e-09, 
    9.57503e-10, 6.037595e-10, 4.050347e-10, 3.243672e-10, 2.68604e-10, 
    2.383735e-10, 2.257922e-10, 2.151784e-10, 2.125265e-10, 2.110652e-10,
  6.230007e-09, 4.793293e-09, 3.706623e-09, 2.856861e-09, 2.005814e-09, 
    1.377827e-09, 9.212735e-10, 6.054405e-10, 4.504399e-10, 3.712268e-10, 
    3.170684e-10, 2.863326e-10, 2.729016e-10, 2.80125e-10, 2.927735e-10,
  6.66807e-09, 5.125966e-09, 4.100414e-09, 3.31171e-09, 2.562308e-09, 
    1.87273e-09, 1.300237e-09, 8.893367e-10, 6.398781e-10, 5.065945e-10, 
    4.406349e-10, 3.922236e-10, 3.668154e-10, 3.627538e-10, 3.73521e-10,
  7.442424e-09, 5.483018e-09, 4.379867e-09, 3.632107e-09, 2.899567e-09, 
    2.362031e-09, 1.848899e-09, 1.305583e-09, 9.245776e-10, 7.092067e-10, 
    5.981651e-10, 5.310987e-10, 4.882527e-10, 4.781444e-10, 5.014461e-10,
  7.78465e-09, 5.913603e-09, 4.756379e-09, 3.784713e-09, 3.088212e-09, 
    2.500577e-09, 2.209813e-09, 1.880688e-09, 1.423389e-09, 1.074202e-09, 
    8.740775e-10, 7.471113e-10, 6.760138e-10, 6.590564e-10, 6.958158e-10,
  7.678627e-09, 5.863455e-09, 4.748851e-09, 3.99425e-09, 3.178809e-09, 
    2.523947e-09, 2.218532e-09, 2.121294e-09, 1.87647e-09, 1.554139e-09, 
    1.283387e-09, 1.094293e-09, 9.826658e-10, 9.434383e-10, 9.720681e-10,
  7.484882e-09, 5.607852e-09, 4.393149e-09, 3.930524e-09, 3.350541e-09, 
    2.558741e-09, 2.172314e-09, 2.021344e-09, 2.031345e-09, 1.911227e-09, 
    1.741481e-09, 1.581376e-09, 1.44966e-09, 1.371848e-09, 1.356313e-09,
  7.516971e-09, 5.810395e-09, 4.438867e-09, 3.678573e-09, 3.358199e-09, 
    2.841574e-09, 2.179059e-09, 1.950889e-09, 1.929334e-09, 1.992067e-09, 
    1.962246e-09, 1.954218e-09, 1.902322e-09, 1.8919e-09, 1.927697e-09,
  8.222112e-09, 5.161726e-09, 3.101368e-09, 1.721233e-09, 9.65411e-10, 
    5.347133e-10, 2.928598e-10, 2.074362e-10, 1.729266e-10, 2.120596e-10, 
    2.913682e-10, 3.351202e-10, 3.602178e-10, 3.919636e-10, 4.581902e-10,
  1.056682e-08, 7.200704e-09, 4.661302e-09, 2.708555e-09, 1.527447e-09, 
    9.024335e-10, 5.032896e-10, 3.068817e-10, 2.106473e-10, 1.928222e-10, 
    2.335579e-10, 2.964033e-10, 3.293111e-10, 3.588307e-10, 4.195393e-10,
  1.420848e-08, 9.476917e-09, 6.324025e-09, 4.056353e-09, 2.345753e-09, 
    1.337273e-09, 8.2604e-10, 4.950662e-10, 3.051533e-10, 2.305717e-10, 
    2.210109e-10, 2.61143e-10, 2.694551e-10, 3.059991e-10, 3.598145e-10,
  1.795592e-08, 1.252487e-08, 8.410348e-09, 5.640636e-09, 3.528385e-09, 
    2.033849e-09, 1.193677e-09, 7.802368e-10, 4.806872e-10, 3.123845e-10, 
    2.403064e-10, 2.265566e-10, 2.307801e-10, 2.606653e-10, 2.977409e-10,
  2.079151e-08, 1.578672e-08, 1.098851e-08, 7.463264e-09, 4.907605e-09, 
    3.048895e-09, 1.743946e-09, 1.076064e-09, 7.377326e-10, 4.973786e-10, 
    3.282737e-10, 2.406129e-10, 2.040978e-10, 2.204498e-10, 2.495472e-10,
  2.259603e-08, 1.898144e-08, 1.394066e-08, 9.727696e-09, 6.522662e-09, 
    4.292724e-09, 2.645577e-09, 1.53983e-09, 9.548773e-10, 6.562335e-10, 
    4.705956e-10, 3.3158e-10, 2.32073e-10, 2.036314e-10, 2.128573e-10,
  2.453398e-08, 2.089211e-08, 1.680006e-08, 1.216708e-08, 8.440946e-09, 
    5.525282e-09, 3.666734e-09, 2.300459e-09, 1.452654e-09, 9.351393e-10, 
    6.295342e-10, 4.564341e-10, 3.2534e-10, 2.486242e-10, 2.108412e-10,
  2.608235e-08, 2.237067e-08, 1.909897e-08, 1.454969e-08, 1.06914e-08, 
    7.301316e-09, 4.813539e-09, 3.151911e-09, 1.988832e-09, 1.308296e-09, 
    8.680798e-10, 6.158807e-10, 4.630899e-10, 3.43463e-10, 2.629786e-10,
  2.661213e-08, 2.443793e-08, 2.07678e-08, 1.687416e-08, 1.266e-08, 
    8.963915e-09, 6.132922e-09, 4.136397e-09, 2.703164e-09, 1.752678e-09, 
    1.182428e-09, 8.079807e-10, 6.014788e-10, 4.51959e-10, 3.427884e-10,
  2.587276e-08, 2.487246e-08, 2.243346e-08, 1.854874e-08, 1.477598e-08, 
    1.089211e-08, 7.588843e-09, 5.195646e-09, 3.532023e-09, 2.371916e-09, 
    1.59821e-09, 1.058697e-09, 7.558443e-10, 5.619168e-10, 4.181924e-10,
  1.931896e-09, 1.197647e-09, 7.567424e-10, 5.802587e-10, 4.768628e-10, 
    4.748263e-10, 3.933193e-10, 2.421168e-10, 1.43956e-10, 1.022098e-10, 
    4.955929e-11, -2.881093e-11, -1.003646e-10, -1.520051e-10, -1.370085e-10,
  2.833654e-09, 1.776769e-09, 1.081942e-09, 7.205252e-10, 5.602818e-10, 
    4.979384e-10, 4.775068e-10, 3.595272e-10, 2.451852e-10, 1.358439e-10, 
    5.252748e-11, -1.807517e-11, -4.532272e-11, -1.033824e-10, -1.310308e-10,
  4.143695e-09, 2.646116e-09, 1.667469e-09, 1.016302e-09, 7.054958e-10, 
    5.883261e-10, 5.501261e-10, 4.589767e-10, 3.616382e-10, 2.454963e-10, 
    1.201108e-10, 6.799011e-11, 2.632647e-11, -2.501769e-11, -6.729453e-11,
  5.469094e-09, 3.825948e-09, 2.512223e-09, 1.576961e-09, 9.880197e-10, 
    7.154964e-10, 6.246925e-10, 5.837786e-10, 4.511174e-10, 3.376764e-10, 
    2.4059e-10, 1.725804e-10, 1.058085e-10, 2.578384e-11, -3.617978e-11,
  7.140406e-09, 5.296229e-09, 3.732894e-09, 2.456818e-09, 1.552267e-09, 
    9.845085e-10, 7.185472e-10, 6.70258e-10, 5.869696e-10, 4.245605e-10, 
    3.084499e-10, 2.762085e-10, 2.041117e-10, 1.060027e-10, 2.538345e-11,
  9.493379e-09, 6.980901e-09, 5.083871e-09, 3.582847e-09, 2.390582e-09, 
    1.556509e-09, 1.027416e-09, 7.618789e-10, 7.017639e-10, 5.733927e-10, 
    3.846235e-10, 3.500166e-10, 3.080243e-10, 2.202841e-10, 1.29857e-10,
  1.212898e-08, 9.442425e-09, 6.804923e-09, 4.945361e-09, 3.462267e-09, 
    2.338022e-09, 1.572727e-09, 1.087824e-09, 8.433471e-10, 7.381832e-10, 
    5.510019e-10, 4.384227e-10, 3.888822e-10, 3.11941e-10, 2.427182e-10,
  1.549888e-08, 1.162469e-08, 9.109081e-09, 6.563132e-09, 4.709843e-09, 
    3.450087e-09, 2.436962e-09, 1.674474e-09, 1.184989e-09, 9.172647e-10, 
    7.175596e-10, 5.577862e-10, 4.962571e-10, 4.007265e-10, 3.316582e-10,
  2.086417e-08, 1.613802e-08, 1.224253e-08, 8.930392e-09, 6.325569e-09, 
    4.593651e-09, 3.44796e-09, 2.514582e-09, 1.778873e-09, 1.365667e-09, 
    1.028187e-09, 7.227643e-10, 6.107604e-10, 5.249671e-10, 4.497436e-10,
  2.423363e-08, 2.096263e-08, 1.651923e-08, 1.243123e-08, 8.923398e-09, 
    6.270312e-09, 4.555867e-09, 3.477996e-09, 2.538681e-09, 1.912785e-09, 
    1.585234e-09, 1.142028e-09, 7.813112e-10, 6.472437e-10, 5.943665e-10,
  6.003923e-09, 3.33592e-09, 1.97435e-09, 1.084407e-09, 5.49166e-10, 
    3.816388e-10, 2.546784e-10, 1.28911e-10, 9.637583e-11, 1.098305e-10, 
    7.777254e-11, 2.049559e-10, 3.145603e-10, 3.018652e-10, 5.774685e-10,
  7.848541e-09, 4.637808e-09, 2.589848e-09, 1.441463e-09, 7.278271e-10, 
    4.042085e-10, 2.953899e-10, 1.918208e-10, 1.196999e-10, 1.132197e-10, 
    4.556709e-11, 1.072489e-10, 2.270214e-10, 3.238501e-10, 3.768892e-10,
  1.001783e-08, 6.067622e-09, 3.524631e-09, 1.93493e-09, 1.036885e-09, 
    5.360797e-10, 3.731763e-10, 2.582104e-10, 1.707324e-10, 1.402923e-10, 
    6.23399e-11, 4.125666e-11, 1.688347e-10, 2.85987e-10, 3.370033e-10,
  1.258374e-08, 7.54576e-09, 4.731644e-09, 2.715281e-09, 1.460531e-09, 
    7.85266e-10, 4.970274e-10, 3.767465e-10, 2.434647e-10, 1.844226e-10, 
    9.776023e-11, 3.591401e-11, 1.103063e-10, 1.900131e-10, 2.776341e-10,
  1.530918e-08, 9.826521e-09, 6.012714e-09, 3.678832e-09, 2.094082e-09, 
    1.132553e-09, 6.592691e-10, 4.942278e-10, 3.600606e-10, 2.458022e-10, 
    1.605092e-10, 6.448821e-11, 5.565643e-11, 9.796793e-11, 1.902967e-10,
  1.701383e-08, 1.248514e-08, 8.036366e-09, 4.749216e-09, 2.866753e-09, 
    1.616486e-09, 8.499188e-10, 5.547792e-10, 3.814672e-10, 2.635621e-10, 
    2.157683e-10, 1.172823e-10, 5.564797e-11, 6.59644e-11, 7.681138e-11,
  1.890692e-08, 1.477122e-08, 1.04301e-08, 6.514971e-09, 3.69468e-09, 
    2.228361e-09, 1.12787e-09, 6.278012e-10, 4.572164e-10, 2.957944e-10, 
    2.183391e-10, 1.986729e-10, 1.00524e-10, 8.064502e-11, 6.542909e-11,
  2.075137e-08, 1.698308e-08, 1.275694e-08, 8.532947e-09, 5.125252e-09, 
    3.035314e-09, 1.608771e-09, 8.811375e-10, 7.031791e-10, 4.649741e-10, 
    2.659107e-10, 2.522536e-10, 1.995933e-10, 1.411509e-10, 1.225728e-10,
  2.244125e-08, 1.921569e-08, 1.502468e-08, 1.083689e-08, 7.016969e-09, 
    4.019029e-09, 2.435168e-09, 1.248042e-09, 8.802357e-10, 5.728697e-10, 
    3.634719e-10, 2.596753e-10, 2.902829e-10, 2.306627e-10, 1.67795e-10,
  2.340642e-08, 2.126496e-08, 1.758171e-08, 1.312942e-08, 9.134214e-09, 
    5.451e-09, 3.252517e-09, 1.743077e-09, 9.935629e-10, 6.718829e-10, 
    4.617398e-10, 2.875891e-10, 3.505407e-10, 3.248389e-10, 2.660494e-10,
  1.302766e-08, 8.982263e-09, 5.536155e-09, 2.581074e-09, 1.059966e-09, 
    5.177309e-10, 1.279333e-10, -1.291562e-10, -1.931235e-11, 1.75589e-10, 
    2.56368e-10, 2.735093e-10, 3.245276e-10, 3.505027e-10, 3.679266e-10,
  1.50648e-08, 1.088658e-08, 7.125825e-09, 4.04314e-09, 1.656908e-09, 
    7.034505e-10, 3.726143e-10, -7.220206e-11, -7.824218e-11, 1.062595e-10, 
    2.756467e-10, 2.751719e-10, 3.266234e-10, 3.582371e-10, 3.62975e-10,
  1.706077e-08, 1.257998e-08, 8.654941e-09, 5.515429e-09, 2.676188e-09, 
    1.027117e-09, 5.484703e-10, 6.206558e-11, -1.108824e-10, 2.326488e-11, 
    2.37183e-10, 3.082832e-10, 3.104702e-10, 3.430528e-10, 3.506826e-10,
  1.847165e-08, 1.434439e-08, 1.029388e-08, 7.06067e-09, 4.112865e-09, 
    1.676773e-09, 7.272957e-10, 2.840786e-10, -1.230603e-10, -4.547752e-11, 
    1.629125e-10, 2.676593e-10, 2.643039e-10, 3.243555e-10, 3.276957e-10,
  1.946556e-08, 1.601311e-08, 1.213044e-08, 8.541017e-09, 5.611047e-09, 
    2.861388e-09, 1.02118e-09, 5.518274e-10, -4.733062e-11, -1.02265e-10, 
    1.139424e-10, 1.997404e-10, 1.905775e-10, 2.650698e-10, 3.023998e-10,
  2.020068e-08, 1.753638e-08, 1.417135e-08, 1.02817e-08, 7.142303e-09, 
    4.35454e-09, 1.784526e-09, 8.570271e-10, 1.675617e-10, -1.54044e-10, 
    4.428926e-12, 1.545428e-10, 1.269702e-10, 1.804476e-10, 2.451173e-10,
  2.104513e-08, 1.884121e-08, 1.619756e-08, 1.236396e-08, 8.713703e-09, 
    5.868766e-09, 3.016611e-09, 1.181181e-09, 5.353299e-10, -4.692201e-11, 
    -1.026203e-10, 1.13309e-10, 1.059751e-10, 1.385402e-10, 2.28981e-10,
  2.189573e-08, 1.99571e-08, 1.77558e-08, 1.441115e-08, 1.070262e-08, 
    7.55908e-09, 4.613864e-09, 1.981345e-09, 8.118765e-10, 9.142145e-11, 
    -1.664272e-10, 3.376187e-11, 8.629047e-11, 1.40897e-10, 2.20175e-10,
  2.275013e-08, 2.099661e-08, 1.904055e-08, 1.668927e-08, 1.267903e-08, 
    8.929179e-09, 6.063923e-09, 3.409271e-09, 1.359459e-09, 4.413631e-10, 
    -7.210781e-11, -8.317341e-11, 7.731711e-11, 1.653706e-10, 2.615274e-10,
  2.476526e-08, 2.20919e-08, 2.014799e-08, 1.841274e-08, 1.495749e-08, 
    1.092899e-08, 7.538571e-09, 4.899478e-09, 2.527897e-09, 8.971973e-10, 
    1.22567e-10, -1.101395e-10, 2.512316e-11, 1.774213e-10, 2.623325e-10,
  2.560038e-08, 2.099905e-08, 1.536467e-08, 1.10575e-08, 7.99888e-09, 
    4.811255e-09, 2.678612e-09, 1.805145e-09, 1.414827e-09, 1.151608e-09, 
    8.854405e-10, 5.725586e-10, 2.767712e-10, 2.905324e-10, 3.730304e-10,
  2.730875e-08, 2.437249e-08, 1.879116e-08, 1.332504e-08, 9.339836e-09, 
    6.271219e-09, 3.58144e-09, 2.135635e-09, 1.522924e-09, 1.200863e-09, 
    9.946476e-10, 7.35019e-10, 4.25448e-10, 2.839433e-10, 3.409333e-10,
  2.931617e-08, 2.733046e-08, 2.156587e-08, 1.593079e-08, 1.124926e-08, 
    7.565689e-09, 4.705654e-09, 2.738876e-09, 1.756298e-09, 1.307043e-09, 
    1.059153e-09, 8.57191e-10, 5.94584e-10, 3.262369e-10, 3.277958e-10,
  2.884861e-08, 2.918325e-08, 2.551279e-08, 1.878463e-08, 1.338992e-08, 
    9.061226e-09, 5.937432e-09, 3.4404e-09, 2.088911e-09, 1.447786e-09, 
    1.139801e-09, 9.69175e-10, 7.276846e-10, 4.515467e-10, 3.177919e-10,
  2.687791e-08, 2.839485e-08, 2.789527e-08, 2.292312e-08, 1.573846e-08, 
    1.079875e-08, 7.177154e-09, 4.44155e-09, 2.619012e-09, 1.690173e-09, 
    1.250831e-09, 1.005296e-09, 8.078997e-10, 5.614744e-10, 3.461163e-10,
  2.69272e-08, 2.65749e-08, 2.741196e-08, 2.568047e-08, 1.921456e-08, 
    1.276501e-08, 8.601194e-09, 5.373334e-09, 3.177716e-09, 1.99491e-09, 
    1.34919e-09, 1.047136e-09, 8.347953e-10, 6.369815e-10, 4.205543e-10,
  2.763167e-08, 2.675947e-08, 2.621582e-08, 2.613151e-08, 2.204811e-08, 
    1.534072e-08, 1.027281e-08, 6.615268e-09, 3.899782e-09, 2.323668e-09, 
    1.490091e-09, 1.112528e-09, 8.838845e-10, 6.985753e-10, 4.81554e-10,
  2.819246e-08, 2.723963e-08, 2.56384e-08, 2.47129e-08, 2.280823e-08, 
    1.7696e-08, 1.209764e-08, 7.851683e-09, 4.717859e-09, 2.747434e-09, 
    1.653535e-09, 1.230255e-09, 9.36527e-10, 7.33961e-10, 5.290122e-10,
  2.768101e-08, 2.743695e-08, 2.570395e-08, 2.389658e-08, 2.191441e-08, 
    1.815072e-08, 1.354061e-08, 9.211766e-09, 5.706407e-09, 3.333328e-09, 
    1.897315e-09, 1.329713e-09, 9.876678e-10, 7.227843e-10, 5.527691e-10,
  2.740577e-08, 2.775805e-08, 2.648559e-08, 2.403676e-08, 2.088927e-08, 
    1.771468e-08, 1.401654e-08, 1.016102e-08, 6.635334e-09, 3.896673e-09, 
    2.274602e-09, 1.479679e-09, 1.040307e-09, 7.092919e-10, 5.334623e-10,
  1.683746e-08, 1.475629e-08, 1.260153e-08, 1.050195e-08, 8.695741e-09, 
    6.535864e-09, 4.549511e-09, 3.114216e-09, 1.81056e-09, 1.22404e-09, 
    1.048281e-09, 8.417946e-10, 5.120446e-10, 1.982367e-10, 4.707014e-13,
  1.760717e-08, 1.590823e-08, 1.357053e-08, 1.139561e-08, 9.367864e-09, 
    7.472775e-09, 5.28498e-09, 3.664645e-09, 2.30943e-09, 1.441368e-09, 
    1.172931e-09, 1.002167e-09, 6.727254e-10, 3.524564e-10, 1.690526e-11,
  1.815808e-08, 1.671619e-08, 1.468156e-08, 1.258121e-08, 1.027274e-08, 
    8.369503e-09, 6.147357e-09, 4.27529e-09, 2.801091e-09, 1.759982e-09, 
    1.335383e-09, 1.145615e-09, 8.438586e-10, 5.302276e-10, 1.151572e-10,
  1.856228e-08, 1.684164e-08, 1.568239e-08, 1.395294e-08, 1.146394e-08, 
    9.337207e-09, 7.139175e-09, 4.972251e-09, 3.347958e-09, 2.111828e-09, 
    1.518917e-09, 1.304708e-09, 1.029909e-09, 7.052828e-10, 3.031613e-10,
  1.899729e-08, 1.775183e-08, 1.61493e-08, 1.511512e-08, 1.296738e-08, 
    1.043545e-08, 8.277057e-09, 5.971694e-09, 4.079425e-09, 2.591407e-09, 
    1.754119e-09, 1.443148e-09, 1.23109e-09, 9.000374e-10, 5.409241e-10,
  1.876531e-08, 1.839821e-08, 1.708145e-08, 1.584937e-08, 1.432509e-08, 
    1.18781e-08, 9.314547e-09, 7.008866e-09, 4.815022e-09, 3.149287e-09, 
    2.043681e-09, 1.614361e-09, 1.393295e-09, 1.123396e-09, 7.774336e-10,
  1.859498e-08, 1.886383e-08, 1.845065e-08, 1.689747e-08, 1.539432e-08, 
    1.312059e-08, 1.060554e-08, 8.33023e-09, 6.006692e-09, 3.973045e-09, 
    2.486304e-09, 1.812105e-09, 1.572991e-09, 1.354341e-09, 1.037669e-09,
  1.898806e-08, 1.920603e-08, 1.960319e-08, 1.872923e-08, 1.716698e-08, 
    1.479129e-08, 1.21053e-08, 9.614368e-09, 7.20008e-09, 4.950737e-09, 
    3.094119e-09, 2.09805e-09, 1.740704e-09, 1.567092e-09, 1.298228e-09,
  1.964582e-08, 1.950762e-08, 1.976067e-08, 2.062726e-08, 1.887033e-08, 
    1.655975e-08, 1.370983e-08, 1.124873e-08, 8.718649e-09, 6.218582e-09, 
    3.976451e-09, 2.526422e-09, 1.931337e-09, 1.74286e-09, 1.549628e-09,
  2.059665e-08, 1.992345e-08, 1.992573e-08, 2.105523e-08, 2.072993e-08, 
    1.846651e-08, 1.59211e-08, 1.310966e-08, 1.045364e-08, 7.636729e-09, 
    5.02246e-09, 3.141748e-09, 2.204853e-09, 1.879169e-09, 1.731819e-09,
  2.059696e-08, 1.89327e-08, 1.781986e-08, 1.552847e-08, 1.232598e-08, 
    8.656231e-09, 5.815125e-09, 3.179961e-09, 1.765047e-09, 1.21269e-09, 
    7.571744e-10, 4.347685e-10, 3.384448e-10, 5.578311e-10, 5.26729e-10,
  1.953785e-08, 1.704872e-08, 1.54934e-08, 1.511235e-08, 1.592935e-08, 
    1.043388e-08, 6.031149e-09, 3.42447e-09, 1.828394e-09, 1.269854e-09, 
    8.073428e-10, 3.220557e-10, 2.252039e-10, 4.920532e-10, 6.150589e-10,
  1.909307e-08, 1.667869e-08, 1.363822e-08, 1.256882e-08, 1.397586e-08, 
    1.361234e-08, 7.692503e-09, 4.007287e-09, 2.053748e-09, 1.302906e-09, 
    8.769114e-10, 3.532097e-10, 7.521326e-11, 5.664323e-10, 6.702008e-10,
  1.935368e-08, 1.691077e-08, 1.323191e-08, 1.081338e-08, 1.18443e-08, 
    1.275228e-08, 9.872923e-09, 5.564933e-09, 2.436885e-09, 1.306447e-09, 
    9.059351e-10, 4.169341e-10, 3.238008e-11, 4.638106e-10, 6.793424e-10,
  2.05395e-08, 1.748833e-08, 1.400521e-08, 1.02521e-08, 8.780832e-09, 
    1.06554e-08, 9.890492e-09, 6.976385e-09, 3.29349e-09, 1.437159e-09, 
    9.878455e-10, 5.3693e-10, 1.431388e-10, 2.441312e-10, 5.736652e-10,
  2.173131e-08, 1.863235e-08, 1.46753e-08, 1.045511e-08, 8.074442e-09, 
    8.003142e-09, 9.169296e-09, 7.605784e-09, 4.249318e-09, 1.674159e-09, 
    1.030831e-09, 6.734875e-10, 2.476871e-10, 1.500083e-10, 3.132547e-10,
  2.257992e-08, 1.956079e-08, 1.521113e-08, 1.163316e-08, 9.177868e-09, 
    7.825236e-09, 8.730439e-09, 8.336778e-09, 5.014617e-09, 2.138271e-09, 
    1.133312e-09, 7.693506e-10, 3.33541e-10, 2.251406e-10, 2.585477e-10,
  2.283763e-08, 2.029779e-08, 1.63099e-08, 1.267777e-08, 1.053854e-08, 
    9.051613e-09, 8.655738e-09, 8.362052e-09, 5.420095e-09, 2.593864e-09, 
    1.299095e-09, 8.432383e-10, 4.023044e-10, 2.572967e-10, 3.02294e-10,
  2.330994e-08, 2.086006e-08, 1.743943e-08, 1.397202e-08, 1.165194e-08, 
    9.788078e-09, 8.440577e-09, 8.230204e-09, 6.082728e-09, 3.235831e-09, 
    1.597668e-09, 1.019011e-09, 5.078599e-10, 2.887083e-10, 2.89527e-10,
  2.350011e-08, 2.134458e-08, 1.80528e-08, 1.502665e-08, 1.277682e-08, 
    1.08482e-08, 9.033627e-09, 8.330615e-09, 6.895475e-09, 3.94715e-09, 
    2.104264e-09, 1.241938e-09, 6.894501e-10, 3.282124e-10, 2.640898e-10,
  2.481781e-08, 2.365902e-08, 2.307065e-08, 2.337951e-08, 2.285282e-08, 
    2.194098e-08, 2.014085e-08, 1.726688e-08, 1.426803e-08, 1.101187e-08, 
    7.895239e-09, 5.859597e-09, 4.298093e-09, 3.256057e-09, 2.308381e-09,
  2.180415e-08, 2.140388e-08, 2.290006e-08, 2.322175e-08, 2.285287e-08, 
    2.144204e-08, 1.996588e-08, 1.843575e-08, 1.548806e-08, 1.244884e-08, 
    9.217817e-09, 6.569354e-09, 4.698788e-09, 3.694465e-09, 2.487403e-09,
  1.854215e-08, 1.987148e-08, 2.196562e-08, 2.268314e-08, 2.281991e-08, 
    2.278979e-08, 2.021327e-08, 1.809881e-08, 1.584356e-08, 1.31809e-08, 
    1.018998e-08, 7.21439e-09, 5.103618e-09, 3.724284e-09, 2.526438e-09,
  1.699915e-08, 1.840558e-08, 1.908472e-08, 2.000334e-08, 2.020451e-08, 
    1.985517e-08, 1.963878e-08, 1.806888e-08, 1.544269e-08, 1.283395e-08, 
    1.01657e-08, 7.149373e-09, 5.123597e-09, 3.548731e-09, 2.315593e-09,
  1.645746e-08, 1.701458e-08, 1.727274e-08, 1.739309e-08, 1.708385e-08, 
    1.73954e-08, 1.664467e-08, 1.695217e-08, 1.416732e-08, 1.180762e-08, 
    9.36859e-09, 6.573963e-09, 4.865951e-09, 3.301839e-09, 2.000225e-09,
  1.653576e-08, 1.641786e-08, 1.577399e-08, 1.329232e-08, 1.349717e-08, 
    1.371067e-08, 1.336329e-08, 1.364385e-08, 1.239932e-08, 1.029238e-08, 
    8.032069e-09, 5.382283e-09, 3.420561e-09, 2.413491e-09, 1.558763e-09,
  1.67439e-08, 1.415934e-08, 1.189685e-08, 1.080608e-08, 1.008033e-08, 
    9.360668e-09, 1.018872e-08, 1.041341e-08, 1.009861e-08, 8.322103e-09, 
    5.841968e-09, 3.660579e-09, 2.53688e-09, 1.61223e-09, 8.01571e-10,
  1.564073e-08, 1.079334e-08, 7.969318e-09, 8.273008e-09, 7.713703e-09, 
    6.616915e-09, 7.258679e-09, 7.116451e-09, 6.874322e-09, 5.630067e-09, 
    3.585987e-09, 2.551756e-09, 1.990178e-09, 1.314043e-09, 7.737764e-10,
  1.290085e-08, 7.826968e-09, 5.596536e-09, 6.472024e-09, 5.588367e-09, 
    4.63668e-09, 4.459892e-09, 4.231951e-09, 4.365464e-09, 3.824337e-09, 
    2.490686e-09, 1.956659e-09, 1.557183e-09, 1.072045e-09, 7.608832e-10,
  1.090494e-08, 6.456839e-09, 4.596815e-09, 4.428615e-09, 4.117884e-09, 
    3.068303e-09, 2.7994e-09, 2.835973e-09, 2.908028e-09, 2.636715e-09, 
    1.843277e-09, 1.541534e-09, 1.308522e-09, 9.42097e-10, 7.376445e-10,
  3.792928e-09, 3.540559e-09, 3.367796e-09, 3.279457e-09, 3.078442e-09, 
    2.783924e-09, 2.532482e-09, 2.293392e-09, 2.062537e-09, 1.97117e-09, 
    2.006835e-09, 2.02636e-09, 2.071461e-09, 2.143859e-09, 2.249807e-09,
  4.772184e-09, 4.502414e-09, 4.414606e-09, 4.318996e-09, 4.1657e-09, 
    3.919031e-09, 3.70378e-09, 3.397651e-09, 3.050222e-09, 2.889332e-09, 
    2.89384e-09, 2.875715e-09, 2.735735e-09, 2.703433e-09, 2.824834e-09,
  6.479048e-09, 6.283237e-09, 6.054028e-09, 5.61867e-09, 5.259503e-09, 
    5.05702e-09, 4.874244e-09, 4.755254e-09, 4.479604e-09, 4.280214e-09, 
    4.178365e-09, 4.128481e-09, 3.978305e-09, 3.81137e-09, 3.756074e-09,
  8.215109e-09, 7.938297e-09, 7.444165e-09, 6.718872e-09, 6.276166e-09, 
    6.160319e-09, 6.133428e-09, 6.238216e-09, 6.101707e-09, 5.986152e-09, 
    5.991478e-09, 6.014719e-09, 5.961831e-09, 5.561811e-09, 5.05729e-09,
  9.612356e-09, 8.988899e-09, 8.348852e-09, 7.806793e-09, 7.468888e-09, 
    7.639961e-09, 7.99409e-09, 8.261315e-09, 8.269655e-09, 8.223808e-09, 
    8.271496e-09, 8.515666e-09, 8.486449e-09, 8.117187e-09, 7.201993e-09,
  1.070595e-08, 1.065711e-08, 9.715877e-09, 9.072814e-09, 8.952663e-09, 
    9.55133e-09, 9.974438e-09, 1.028095e-08, 1.010464e-08, 1.029489e-08, 
    1.026591e-08, 1.056228e-08, 1.052197e-08, 1.001321e-08, 9.153179e-09,
  1.268322e-08, 1.174502e-08, 1.075774e-08, 1.055008e-08, 1.050633e-08, 
    1.095573e-08, 1.155061e-08, 1.275897e-08, 1.304093e-08, 1.284664e-08, 
    1.28994e-08, 1.287893e-08, 1.251068e-08, 1.15757e-08, 1.015652e-08,
  1.420711e-08, 1.262863e-08, 1.17911e-08, 1.130369e-08, 1.193257e-08, 
    1.255627e-08, 1.298377e-08, 1.337977e-08, 1.439376e-08, 1.470314e-08, 
    1.49485e-08, 1.467182e-08, 1.381505e-08, 1.245191e-08, 1.098581e-08,
  1.395201e-08, 1.261559e-08, 1.226029e-08, 1.242945e-08, 1.339241e-08, 
    1.383733e-08, 1.339146e-08, 1.33311e-08, 1.498624e-08, 1.59163e-08, 
    1.607301e-08, 1.506355e-08, 1.423338e-08, 1.296396e-08, 1.111589e-08,
  1.354094e-08, 1.266194e-08, 1.246363e-08, 1.320589e-08, 1.444958e-08, 
    1.409723e-08, 1.484963e-08, 1.505003e-08, 1.586735e-08, 1.597986e-08, 
    1.54637e-08, 1.484774e-08, 1.407839e-08, 1.241803e-08, 1.025534e-08,
  1.599987e-09, 1.06999e-09, 8.21855e-10, 6.477095e-10, 5.846957e-10, 
    5.25094e-10, 4.066555e-10, 2.780557e-10, 2.782362e-10, 2.368671e-10, 
    2.301761e-10, 3.212633e-10, 4.31728e-10, 4.917572e-10, 3.668967e-10,
  1.732089e-09, 1.197873e-09, 9.004336e-10, 7.305008e-10, 6.078503e-10, 
    5.897401e-10, 5.040469e-10, 3.196841e-10, 2.685092e-10, 2.591878e-10, 
    2.357996e-10, 2.739926e-10, 2.72562e-10, 2.827903e-10, 2.991217e-10,
  2.176212e-09, 1.453581e-09, 1.13415e-09, 8.595215e-10, 6.53063e-10, 
    6.054143e-10, 5.682439e-10, 4.101367e-10, 3.222546e-10, 3.298296e-10, 
    3.46808e-10, 2.972595e-10, 2.214793e-10, 1.729866e-10, 1.606876e-10,
  2.693067e-09, 1.920301e-09, 1.413112e-09, 1.010606e-09, 7.307127e-10, 
    6.001922e-10, 5.871809e-10, 5.15775e-10, 3.633429e-10, 4.074113e-10, 
    4.480193e-10, 3.991557e-10, 2.562094e-10, 1.656455e-10, 1.342793e-10,
  3.411882e-09, 2.335542e-09, 1.705464e-09, 1.214542e-09, 8.334508e-10, 
    6.302285e-10, 5.591719e-10, 5.807528e-10, 4.472779e-10, 4.339558e-10, 
    5.344343e-10, 4.863365e-10, 3.646975e-10, 2.165507e-10, 1.428061e-10,
  3.899568e-09, 2.607064e-09, 1.796992e-09, 1.344044e-09, 9.891908e-10, 
    7.137255e-10, 6.339951e-10, 6.419894e-10, 5.819748e-10, 4.6424e-10, 
    4.976718e-10, 4.872485e-10, 4.553471e-10, 3.128983e-10, 2.255388e-10,
  4.12998e-09, 2.626994e-09, 1.857263e-09, 1.423291e-09, 1.116897e-09, 
    8.784249e-10, 7.604937e-10, 6.682649e-10, 6.138491e-10, 4.837663e-10, 
    5.136582e-10, 4.996339e-10, 4.544093e-10, 4.073437e-10, 3.184912e-10,
  4.768767e-09, 3.010218e-09, 2.057235e-09, 1.576641e-09, 1.244438e-09, 
    1.114031e-09, 9.389128e-10, 7.827241e-10, 6.910322e-10, 5.741292e-10, 
    4.821372e-10, 5.046243e-10, 5.154162e-10, 5.116184e-10, 4.579954e-10,
  5.588551e-09, 3.642317e-09, 2.406978e-09, 1.71847e-09, 1.439106e-09, 
    1.387226e-09, 1.156839e-09, 8.727641e-10, 5.957828e-10, 5.37263e-10, 
    4.6858e-10, 4.664327e-10, 5.132405e-10, 5.360961e-10, 5.545584e-10,
  6.167149e-09, 4.159764e-09, 2.794428e-09, 1.981605e-09, 1.673133e-09, 
    1.515879e-09, 1.30364e-09, 9.325737e-10, 6.162e-10, 5.670807e-10, 
    5.488906e-10, 4.423265e-10, 4.839467e-10, 5.506635e-10, 6.393331e-10,
  1.124003e-08, 6.269889e-09, 3.005501e-09, 1.305877e-09, 6.760809e-10, 
    4.427108e-10, 3.464709e-10, 3.923864e-10, 4.011187e-10, 3.88888e-10, 
    4.219235e-10, 5.07661e-10, 5.646497e-10, 5.538264e-10, 6.466511e-10,
  1.223863e-08, 7.661655e-09, 3.765651e-09, 1.745772e-09, 8.327949e-10, 
    4.945801e-10, 3.509552e-10, 3.686315e-10, 3.77333e-10, 3.665776e-10, 
    4.054103e-10, 4.716358e-10, 5.063022e-10, 4.865537e-10, 5.978166e-10,
  1.325242e-08, 9.067162e-09, 4.621295e-09, 2.202663e-09, 1.022882e-09, 
    5.514185e-10, 3.646187e-10, 3.494104e-10, 3.676871e-10, 3.443487e-10, 
    3.711377e-10, 4.205707e-10, 4.821215e-10, 4.511589e-10, 4.700262e-10,
  1.415114e-08, 1.0166e-08, 5.484248e-09, 2.654619e-09, 1.267978e-09, 
    6.598878e-10, 3.925106e-10, 3.434256e-10, 3.545413e-10, 3.324673e-10, 
    3.465425e-10, 3.826389e-10, 4.845357e-10, 4.315201e-10, 4.184542e-10,
  1.498785e-08, 1.091404e-08, 6.125234e-09, 3.126259e-09, 1.525781e-09, 
    7.732603e-10, 4.432879e-10, 3.505822e-10, 3.524284e-10, 3.21292e-10, 
    3.256091e-10, 3.598758e-10, 4.548107e-10, 4.515177e-10, 4.444344e-10,
  1.547609e-08, 1.131473e-08, 6.591434e-09, 3.527946e-09, 1.792469e-09, 
    9.088328e-10, 5.095971e-10, 3.64175e-10, 3.364574e-10, 3.179852e-10, 
    3.142725e-10, 3.456232e-10, 4.302532e-10, 4.281346e-10, 4.449692e-10,
  1.544031e-08, 1.130343e-08, 6.91628e-09, 3.920642e-09, 2.054238e-09, 
    1.041998e-09, 6.289309e-10, 4.254242e-10, 3.438451e-10, 3.042696e-10, 
    3.113657e-10, 3.416636e-10, 3.955896e-10, 4.157247e-10, 4.097505e-10,
  1.512703e-08, 1.121837e-08, 7.005007e-09, 4.231762e-09, 2.30123e-09, 
    1.215695e-09, 7.210501e-10, 4.749693e-10, 3.188655e-10, 2.853442e-10, 
    2.935254e-10, 3.294873e-10, 3.956155e-10, 3.821851e-10, 3.798726e-10,
  1.492558e-08, 1.123754e-08, 6.95995e-09, 4.144698e-09, 2.401953e-09, 
    1.416085e-09, 8.678124e-10, 5.086914e-10, 3.101616e-10, 2.801979e-10, 
    2.887111e-10, 3.167541e-10, 3.839783e-10, 3.613361e-10, 3.530309e-10,
  1.443233e-08, 1.086437e-08, 6.757221e-09, 3.938772e-09, 2.328916e-09, 
    1.456383e-09, 1.043079e-09, 5.873985e-10, 3.209854e-10, 2.731905e-10, 
    2.662593e-10, 3.024294e-10, 3.73019e-10, 3.612871e-10, 3.417253e-10,
  2.589939e-08, 2.302173e-08, 2.038544e-08, 1.618796e-08, 1.087693e-08, 
    5.713016e-09, 3.155879e-09, 2.025178e-09, 7.907548e-10, 1.106547e-10, 
    -2.950929e-11, 1.452889e-10, 3.877896e-10, 4.357253e-10, 4.591145e-10,
  2.648629e-08, 2.377622e-08, 2.094932e-08, 1.730569e-08, 1.273674e-08, 
    7.339932e-09, 3.855203e-09, 2.54194e-09, 1.393977e-09, 3.244121e-10, 
    -1.309222e-11, 7.105334e-11, 2.995164e-10, 3.842391e-10, 4.20015e-10,
  2.695944e-08, 2.423941e-08, 2.133972e-08, 1.78978e-08, 1.39036e-08, 
    8.811138e-09, 4.65771e-09, 2.959473e-09, 1.941096e-09, 6.919648e-10, 
    8.052568e-11, 6.732571e-11, 2.46726e-10, 3.271042e-10, 3.787582e-10,
  2.702214e-08, 2.439647e-08, 2.159764e-08, 1.815496e-08, 1.447995e-08, 
    9.862543e-09, 5.464162e-09, 3.332259e-09, 2.212946e-09, 1.077957e-09, 
    2.39696e-10, 1.081463e-10, 2.544518e-10, 3.279061e-10, 3.314743e-10,
  2.724213e-08, 2.455467e-08, 2.161263e-08, 1.81166e-08, 1.470514e-08, 
    1.036071e-08, 6.133726e-09, 3.805707e-09, 2.480401e-09, 1.411282e-09, 
    5.091591e-10, 2.196061e-10, 2.848882e-10, 3.651552e-10, 2.57178e-10,
  2.633034e-08, 2.43819e-08, 2.153135e-08, 1.791103e-08, 1.461359e-08, 
    1.053134e-08, 6.510898e-09, 4.111954e-09, 2.732171e-09, 1.745667e-09, 
    8.529255e-10, 3.254105e-10, 2.471802e-10, 2.948815e-10, 2.180591e-10,
  2.628528e-08, 2.423709e-08, 2.12153e-08, 1.756818e-08, 1.428145e-08, 
    1.040705e-08, 6.658644e-09, 4.29586e-09, 2.869489e-09, 2.016668e-09, 
    1.21303e-09, 5.587883e-10, 2.630048e-10, 2.326057e-10, 2.343911e-10,
  2.632843e-08, 2.410019e-08, 2.087892e-08, 1.712249e-08, 1.391701e-08, 
    9.96837e-09, 6.632206e-09, 4.497562e-09, 2.930399e-09, 2.019428e-09, 
    1.270495e-09, 6.077151e-10, 2.616539e-10, 2.053126e-10, 2.952613e-10,
  2.605807e-08, 2.374901e-08, 2.026714e-08, 1.643788e-08, 1.332913e-08, 
    9.548612e-09, 6.450992e-09, 4.241578e-09, 2.468216e-09, 1.625827e-09, 
    1.081908e-09, 6.095529e-10, 2.930301e-10, 1.8783e-10, 3.139616e-10,
  2.589473e-08, 2.333102e-08, 1.94759e-08, 1.56201e-08, 1.257042e-08, 
    8.736306e-09, 5.918825e-09, 3.570422e-09, 1.975e-09, 1.410678e-09, 
    9.812144e-10, 5.376249e-10, 3.176732e-10, 2.405221e-10, 3.1359e-10,
  2.277505e-08, 2.111159e-08, 2.021505e-08, 1.730232e-08, 1.244977e-08, 
    8.886957e-09, 6.280866e-09, 4.17532e-09, 2.775856e-09, 1.886503e-09, 
    1.08843e-09, 5.709012e-10, 3.826421e-10, 2.723241e-10, 1.677553e-10,
  2.489825e-08, 2.353226e-08, 2.218768e-08, 2.057984e-08, 1.615289e-08, 
    1.116934e-08, 7.912409e-09, 5.471203e-09, 3.568128e-09, 2.390392e-09, 
    1.559595e-09, 9.849119e-10, 4.595802e-10, 2.854725e-10, 2.16534e-10,
  2.661921e-08, 2.527455e-08, 2.330116e-08, 2.304686e-08, 1.960184e-08, 
    1.436158e-08, 9.756356e-09, 7.025681e-09, 4.766902e-09, 3.13335e-09, 
    2.044964e-09, 1.397609e-09, 7.849218e-10, 4.686539e-10, 2.778369e-10,
  2.690169e-08, 2.645633e-08, 2.488952e-08, 2.382719e-08, 2.289441e-08, 
    1.769885e-08, 1.206729e-08, 8.425959e-09, 5.845073e-09, 3.901726e-09, 
    2.553842e-09, 1.846688e-09, 1.136051e-09, 6.98562e-10, 4.62607e-10,
  2.654648e-08, 2.757049e-08, 2.667648e-08, 2.483823e-08, 2.472787e-08, 
    2.102736e-08, 1.470842e-08, 1.005316e-08, 7.239914e-09, 4.924424e-09, 
    3.212439e-09, 2.226548e-09, 1.55387e-09, 9.997377e-10, 6.592304e-10,
  2.605657e-08, 2.692803e-08, 2.791593e-08, 2.64732e-08, 2.554091e-08, 
    2.330099e-08, 1.747878e-08, 1.15495e-08, 8.025517e-09, 5.638329e-09, 
    3.80829e-09, 2.619329e-09, 1.908587e-09, 1.320012e-09, 7.916214e-10,
  2.64613e-08, 2.715136e-08, 2.849075e-08, 2.787601e-08, 2.682151e-08, 
    2.502799e-08, 1.999505e-08, 1.367126e-08, 9.27075e-09, 6.270084e-09, 
    4.269947e-09, 2.942154e-09, 2.205488e-09, 1.545843e-09, 8.486634e-10,
  2.765263e-08, 2.814438e-08, 2.880317e-08, 2.888862e-08, 2.825683e-08, 
    2.697247e-08, 2.159252e-08, 1.53135e-08, 1.036112e-08, 6.974615e-09, 
    4.721799e-09, 3.245022e-09, 2.350129e-09, 1.72402e-09, 9.254315e-10,
  2.745961e-08, 2.843066e-08, 2.92073e-08, 2.976474e-08, 2.910002e-08, 
    2.747408e-08, 2.344244e-08, 1.678531e-08, 1.130159e-08, 7.481398e-09, 
    5.036755e-09, 3.338452e-09, 2.452901e-09, 1.795733e-09, 1.016316e-09,
  2.775805e-08, 2.845348e-08, 2.920456e-08, 2.985182e-08, 2.923189e-08, 
    2.760227e-08, 2.514893e-08, 1.830444e-08, 1.206439e-08, 7.950392e-09, 
    5.162168e-09, 3.357669e-09, 2.483478e-09, 1.865587e-09, 1.055592e-09,
  1.010396e-08, 8.485152e-09, 7.274485e-09, 6.016869e-09, 4.149672e-09, 
    2.877151e-09, 1.940188e-09, 1.521175e-09, 1.063087e-09, 6.637848e-10, 
    4.515752e-10, 5.329392e-10, 4.278383e-10, 2.665045e-10, 8.736328e-11,
  1.108403e-08, 9.549534e-09, 8.134102e-09, 6.941644e-09, 5.386476e-09, 
    3.665712e-09, 2.522887e-09, 2.087285e-09, 1.444072e-09, 1.005496e-09, 
    6.512986e-10, 4.623185e-10, 4.270444e-10, 2.924447e-10, 1.855013e-10,
  1.201048e-08, 1.05743e-08, 9.152104e-09, 7.924744e-09, 6.551998e-09, 
    4.865881e-09, 3.235845e-09, 2.607289e-09, 2.028883e-09, 1.466783e-09, 
    9.671709e-10, 6.692057e-10, 3.970893e-10, 3.950442e-10, 3.167825e-10,
  1.317234e-08, 1.168516e-08, 1.030801e-08, 8.961077e-09, 7.885684e-09, 
    6.27535e-09, 4.235495e-09, 3.08037e-09, 2.593898e-09, 1.861997e-09, 
    1.205232e-09, 9.110382e-10, 5.7508e-10, 4.378773e-10, 3.500917e-10,
  1.457124e-08, 1.278798e-08, 1.140222e-08, 1.015482e-08, 9.286465e-09, 
    7.81545e-09, 5.206453e-09, 3.534397e-09, 3.018979e-09, 2.299259e-09, 
    1.530518e-09, 1.24004e-09, 8.272239e-10, 5.475408e-10, 3.137896e-10,
  1.579916e-08, 1.376726e-08, 1.246853e-08, 1.148386e-08, 1.054186e-08, 
    9.23436e-09, 6.725584e-09, 4.685929e-09, 3.77545e-09, 2.837109e-09, 
    2.081625e-09, 1.472325e-09, 1.208231e-09, 7.402764e-10, 3.563153e-10,
  1.666652e-08, 1.441146e-08, 1.292233e-08, 1.210958e-08, 1.168733e-08, 
    1.070886e-08, 8.102099e-09, 5.754567e-09, 4.441934e-09, 3.449074e-09, 
    2.748077e-09, 1.915822e-09, 1.534848e-09, 1.125191e-09, 7.33931e-10,
  1.779882e-08, 1.513809e-08, 1.325326e-08, 1.23256e-08, 1.212641e-08, 
    1.162226e-08, 9.527968e-09, 6.351275e-09, 5.01887e-09, 4.265145e-09, 
    3.341547e-09, 2.357278e-09, 1.895076e-09, 1.533137e-09, 1.15176e-09,
  1.930689e-08, 1.648108e-08, 1.374482e-08, 1.240805e-08, 1.20585e-08, 
    1.119044e-08, 1.007645e-08, 7.760204e-09, 6.434368e-09, 5.12496e-09, 
    3.924992e-09, 2.920954e-09, 2.334036e-09, 2.005614e-09, 1.637173e-09,
  2.03848e-08, 1.763195e-08, 1.459116e-08, 1.272927e-08, 1.199999e-08, 
    1.056744e-08, 9.778073e-09, 8.415863e-09, 7.451772e-09, 5.896845e-09, 
    4.528901e-09, 3.433572e-09, 2.720717e-09, 2.36071e-09, 1.998639e-09,
  1.267115e-08, 8.783401e-09, 4.816642e-09, 2.177639e-09, 9.763147e-10, 
    5.283682e-10, 6.943445e-10, 7.649755e-10, 7.729099e-10, 7.770748e-10, 
    7.84621e-10, 7.083212e-10, 6.928199e-10, 5.968555e-10, 5.835233e-10,
  1.321321e-08, 9.61481e-09, 5.675176e-09, 2.695291e-09, 1.235093e-09, 
    5.967865e-10, 7.204227e-10, 7.579869e-10, 6.214334e-10, 5.151415e-10, 
    7.134952e-10, 7.378743e-10, 5.607069e-10, 5.50804e-10, 7.390271e-10,
  1.348698e-08, 1.004983e-08, 6.343121e-09, 3.250577e-09, 1.558764e-09, 
    7.519984e-10, 7.107876e-10, 7.804357e-10, 5.167898e-10, 3.088085e-10, 
    5.827958e-10, 5.985313e-10, 4.303002e-10, 4.614523e-10, 6.912791e-10,
  1.335057e-08, 1.017193e-08, 6.883005e-09, 3.833788e-09, 1.924431e-09, 
    1.080514e-09, 8.000364e-10, 7.421946e-10, 4.880632e-10, 1.632632e-10, 
    2.826861e-10, 5.249395e-10, 4.59651e-10, 4.68265e-10, 6.25849e-10,
  1.317573e-08, 1.01678e-08, 7.171622e-09, 4.320319e-09, 2.324493e-09, 
    1.423371e-09, 9.549173e-10, 7.758917e-10, 4.863329e-10, 1.284938e-10, 
    1.757499e-10, 3.221401e-10, 3.804598e-10, 3.882233e-10, 5.848321e-10,
  1.280236e-08, 9.949932e-09, 7.215598e-09, 4.694026e-09, 2.716938e-09, 
    1.705629e-09, 1.097113e-09, 9.177796e-10, 5.538238e-10, 1.584356e-10, 
    1.76754e-10, 1.958023e-10, 2.05319e-10, 2.557605e-10, 3.652052e-10,
  1.250679e-08, 9.731133e-09, 7.141832e-09, 4.914623e-09, 2.812078e-09, 
    1.951741e-09, 1.453941e-09, 1.272029e-09, 9.899681e-10, 3.904248e-10, 
    3.321078e-10, 1.93604e-10, 1.852736e-10, 1.551978e-10, 1.680287e-10,
  1.199552e-08, 9.386182e-09, 7.086948e-09, 5.038612e-09, 3.150022e-09, 
    2.60386e-09, 1.896095e-09, 1.996861e-09, 1.560044e-09, 9.669884e-10, 
    6.033077e-10, 3.760988e-10, 2.115282e-10, 1.676276e-10, 2.049483e-10,
  1.163683e-08, 9.190035e-09, 7.240111e-09, 5.535761e-09, 3.674727e-09, 
    2.777568e-09, 2.374662e-09, 2.289581e-09, 2.106446e-09, 1.617951e-09, 
    1.176095e-09, 7.95192e-10, 5.929287e-10, 4.382469e-10, 2.817347e-10,
  1.128858e-08, 9.027688e-09, 7.088441e-09, 4.735976e-09, 2.603411e-09, 
    1.635542e-09, 1.438531e-09, 2.172979e-09, 2.162537e-09, 1.911971e-09, 
    1.638447e-09, 1.202174e-09, 9.762401e-10, 9.737261e-10, 6.320711e-10,
  1.394005e-08, 9.404836e-09, 6.106539e-09, 3.750401e-09, 2.360995e-09, 
    1.73665e-09, 1.415804e-09, 1.299267e-09, 1.491372e-09, 1.256207e-09, 
    5.24738e-10, 2.502782e-10, 3.808499e-10, 5.136062e-10, 4.644413e-10,
  1.470073e-08, 9.869219e-09, 6.368932e-09, 3.801085e-09, 2.34692e-09, 
    1.701328e-09, 1.379897e-09, 1.294904e-09, 1.462362e-09, 1.231425e-09, 
    3.999369e-10, 2.351681e-10, 2.747757e-10, 5.039396e-10, 3.373047e-10,
  1.551087e-08, 1.033774e-08, 6.606494e-09, 3.864908e-09, 2.309036e-09, 
    1.670332e-09, 1.379366e-09, 1.403544e-09, 1.437729e-09, 1.254014e-09, 
    3.927809e-10, 3.077795e-10, 4.313235e-10, 5.331615e-10, 3.120283e-10,
  1.623121e-08, 1.085512e-08, 6.890733e-09, 3.908256e-09, 2.367873e-09, 
    1.625643e-09, 1.419015e-09, 1.480532e-09, 1.49535e-09, 1.126135e-09, 
    5.161023e-10, 3.280742e-10, 4.155039e-10, 5.557984e-10, 3.766495e-10,
  1.689609e-08, 1.151121e-08, 7.277911e-09, 4.094741e-09, 2.466331e-09, 
    1.615913e-09, 1.432627e-09, 1.558077e-09, 1.594736e-09, 1.001715e-09, 
    4.576592e-10, 4.627624e-10, 4.797653e-10, 6.217357e-10, 4.176252e-10,
  1.733268e-08, 1.183294e-08, 7.570297e-09, 4.271409e-09, 2.624345e-09, 
    1.648469e-09, 1.36908e-09, 1.482245e-09, 1.54444e-09, 8.527786e-10, 
    4.129931e-10, 4.434222e-10, 5.416396e-10, 6.488758e-10, 3.336199e-10,
  1.818586e-08, 1.239986e-08, 7.818087e-09, 4.471788e-09, 2.75471e-09, 
    1.545309e-09, 1.220217e-09, 1.424893e-09, 1.490949e-09, 6.578657e-10, 
    3.911069e-10, 5.410083e-10, 6.338732e-10, 5.927353e-10, 3.424132e-10,
  1.910981e-08, 1.280362e-08, 7.98898e-09, 4.59859e-09, 2.66412e-09, 
    1.415547e-09, 1.206469e-09, 1.447169e-09, 1.373434e-09, 5.728269e-10, 
    3.583467e-10, 4.756435e-10, 6.357955e-10, 4.368556e-10, 3.472253e-10,
  1.973535e-08, 1.313141e-08, 8.125381e-09, 4.584503e-09, 2.437526e-09, 
    1.289129e-09, 9.935831e-10, 1.525156e-09, 1.377242e-09, 5.457254e-10, 
    3.537939e-10, 4.213221e-10, 4.628052e-10, 3.57295e-10, 4.958463e-10,
  2.028331e-08, 1.342677e-08, 8.131081e-09, 4.451006e-09, 2.277831e-09, 
    1.030201e-09, 7.853996e-10, 1.43905e-09, 1.265491e-09, 5.5729e-10, 
    3.726002e-10, 3.24838e-10, 2.455382e-10, 2.963193e-10, 7.06178e-10,
  2.370052e-08, 2.072339e-08, 1.694461e-08, 1.29875e-08, 9.3764e-09, 
    6.791125e-09, 4.904551e-09, 3.671111e-09, 2.558753e-09, 1.823254e-09, 
    1.236904e-09, 9.029775e-10, 6.887573e-10, 6.586127e-10, 8.268999e-10,
  2.449105e-08, 2.131393e-08, 1.742238e-08, 1.333073e-08, 9.5231e-09, 
    6.94223e-09, 4.928334e-09, 3.641052e-09, 2.45462e-09, 1.644903e-09, 
    1.065254e-09, 7.520215e-10, 5.663296e-10, 5.587227e-10, 8.520409e-10,
  2.493519e-08, 2.130166e-08, 1.729376e-08, 1.341467e-08, 9.413029e-09, 
    6.852462e-09, 4.854226e-09, 3.481506e-09, 2.273055e-09, 1.426882e-09, 
    9.518802e-10, 7.277779e-10, 4.95895e-10, 7.978429e-10, 8.841873e-10,
  2.501628e-08, 2.116471e-08, 1.705101e-08, 1.29793e-08, 9.008974e-09, 
    6.391663e-09, 4.531708e-09, 3.183918e-09, 2.003693e-09, 1.163093e-09, 
    8.232091e-10, 3.981745e-10, 5.824753e-10, 5.2456e-10, 9.431848e-10,
  2.522793e-08, 2.112026e-08, 1.646684e-08, 1.234387e-08, 8.305784e-09, 
    5.675787e-09, 4.061533e-09, 2.815133e-09, 1.841412e-09, 1.022001e-09, 
    4.975125e-10, 1.36752e-10, -1.890717e-10, 1.086824e-10, 1.139747e-09,
  2.484392e-08, 2.047513e-08, 1.583428e-08, 1.14539e-08, 7.460404e-09, 
    4.86838e-09, 3.356699e-09, 2.413631e-09, 1.61432e-09, 7.587995e-10, 
    1.746637e-10, -1.507933e-10, -1.978117e-10, -1.891666e-10, 9.521453e-10,
  2.50594e-08, 2.017723e-08, 1.502706e-08, 1.043877e-08, 6.435384e-09, 
    4.005142e-09, 2.757703e-09, 2.028118e-09, 1.394276e-09, 5.524456e-10, 
    -4.144757e-11, 5.375095e-12, -6.343575e-10, -2.648037e-10, 7.944673e-10,
  2.48385e-08, 1.949185e-08, 1.402892e-08, 9.31919e-09, 5.440448e-09, 
    3.468831e-09, 2.633188e-09, 1.888748e-09, 1.261788e-09, 3.933579e-10, 
    -9.431683e-12, -1.026945e-10, -7.961823e-10, -3.185242e-10, 6.580713e-10,
  2.43951e-08, 1.870798e-08, 1.301944e-08, 8.156365e-09, 4.659281e-09, 
    3.080622e-09, 2.240755e-09, 1.717865e-09, 1.092633e-09, 3.486003e-10, 
    2.19006e-11, -3.746764e-10, -8.914254e-10, 3.675846e-11, 7.11932e-10,
  2.391738e-08, 1.790994e-08, 1.20116e-08, 7.163784e-09, 4.242105e-09, 
    2.816792e-09, 1.973117e-09, 1.480474e-09, 9.079364e-10, 2.316843e-10, 
    -1.358049e-10, -8.333781e-10, -2.357976e-10, 2.487259e-10, 7.54368e-10,
  2.364967e-08, 2.165975e-08, 1.925741e-08, 1.651584e-08, 1.358812e-08, 
    1.088773e-08, 8.378389e-09, 6.618952e-09, 5.633972e-09, 5.066033e-09, 
    4.311392e-09, 3.921315e-09, 3.369092e-09, 2.930867e-09, 2.580338e-09,
  2.47065e-08, 2.330541e-08, 2.093175e-08, 1.868077e-08, 1.581476e-08, 
    1.298979e-08, 1.067602e-08, 8.365404e-09, 6.718863e-09, 5.386589e-09, 
    4.536157e-09, 4.219308e-09, 3.646444e-09, 3.309449e-09, 2.86339e-09,
  2.588657e-08, 2.432262e-08, 2.211319e-08, 2.000835e-08, 1.744549e-08, 
    1.427613e-08, 1.243338e-08, 1.010903e-08, 8.033367e-09, 5.975143e-09, 
    4.882625e-09, 4.393442e-09, 4.105021e-09, 3.597391e-09, 2.794691e-09,
  2.695668e-08, 2.507179e-08, 2.308173e-08, 2.107155e-08, 1.885512e-08, 
    1.540435e-08, 1.331769e-08, 1.154841e-08, 9.162959e-09, 6.637585e-09, 
    5.431997e-09, 4.82237e-09, 4.169988e-09, 3.513182e-09, 2.400089e-09,
  2.839374e-08, 2.609698e-08, 2.366843e-08, 2.14773e-08, 1.944912e-08, 
    1.628467e-08, 1.38254e-08, 1.227656e-08, 9.938089e-09, 7.341678e-09, 
    6.005789e-09, 5.040284e-09, 4.016762e-09, 3.110422e-09, 2.106624e-09,
  2.786198e-08, 2.661365e-08, 2.408581e-08, 2.164729e-08, 1.968439e-08, 
    1.676767e-08, 1.386726e-08, 1.209506e-08, 9.964888e-09, 7.766199e-09, 
    6.120407e-09, 5.007876e-09, 3.790154e-09, 2.817333e-09, 2.165511e-09,
  3.040043e-08, 2.76777e-08, 2.458127e-08, 2.151601e-08, 1.92083e-08, 
    1.654419e-08, 1.394063e-08, 1.204287e-08, 9.661122e-09, 7.478857e-09, 
    6.045366e-09, 4.959502e-09, 3.544609e-09, 2.537047e-09, 2.017766e-09,
  3.12394e-08, 2.784014e-08, 2.411807e-08, 2.092476e-08, 1.853916e-08, 
    1.574202e-08, 1.336125e-08, 1.091817e-08, 8.582166e-09, 6.859358e-09, 
    5.89106e-09, 4.811348e-09, 3.218407e-09, 2.114177e-09, 1.998994e-09,
  3.068552e-08, 2.703257e-08, 2.311982e-08, 1.997454e-08, 1.718304e-08, 
    1.459326e-08, 1.201014e-08, 9.130042e-09, 7.559875e-09, 6.063458e-09, 
    5.378692e-09, 4.09219e-09, 2.557443e-09, 1.765926e-09, 1.804265e-09,
  2.955743e-08, 2.560829e-08, 2.16225e-08, 1.818406e-08, 1.553821e-08, 
    1.281776e-08, 9.92747e-09, 7.724487e-09, 6.336776e-09, 5.244309e-09, 
    4.377924e-09, 3.112715e-09, 1.834713e-09, 1.675733e-09, 1.746979e-09,
  1.76833e-08, 1.292789e-08, 8.28914e-09, 6.41998e-09, 5.14369e-09, 
    4.016273e-09, 2.980985e-09, 2.570591e-09, 2.277852e-09, 3.304816e-09, 
    3.483395e-09, 2.719263e-09, 1.832134e-09, 1.488205e-09, 9.770091e-10,
  2.096735e-08, 1.57127e-08, 1.111278e-08, 7.965636e-09, 6.202356e-09, 
    5.060984e-09, 3.801425e-09, 2.768652e-09, 2.440209e-09, 2.518494e-09, 
    3.619096e-09, 3.461577e-09, 2.547014e-09, 2.028817e-09, 1.416401e-09,
  2.384719e-08, 1.898843e-08, 1.428397e-08, 1.017371e-08, 7.698035e-09, 
    6.1823e-09, 4.826388e-09, 3.467571e-09, 2.713524e-09, 2.689456e-09, 
    3.136712e-09, 4.183213e-09, 3.415633e-09, 2.688691e-09, 1.943212e-09,
  2.484836e-08, 2.144919e-08, 1.709021e-08, 1.292296e-08, 9.792376e-09, 
    7.602228e-09, 6.133388e-09, 4.663543e-09, 3.161155e-09, 2.553847e-09, 
    2.73959e-09, 4.210986e-09, 4.368986e-09, 3.598424e-09, 2.617738e-09,
  2.519521e-08, 2.345463e-08, 1.982995e-08, 1.539586e-08, 1.236461e-08, 
    9.545763e-09, 7.470427e-09, 6.149792e-09, 4.472037e-09, 2.950776e-09, 
    2.642321e-09, 3.632891e-09, 4.773757e-09, 4.509028e-09, 3.55171e-09,
  2.346366e-08, 2.410043e-08, 2.180308e-08, 1.787232e-08, 1.438121e-08, 
    1.184591e-08, 9.323427e-09, 7.328542e-09, 5.752914e-09, 3.858636e-09, 
    2.862852e-09, 3.351442e-09, 4.059191e-09, 4.960363e-09, 4.411745e-09,
  2.410099e-08, 2.407231e-08, 2.307717e-08, 2.010576e-08, 1.630919e-08, 
    1.350504e-08, 1.123168e-08, 9.250365e-09, 7.627733e-09, 5.073138e-09, 
    3.333369e-09, 3.41602e-09, 3.651399e-09, 4.630496e-09, 4.551741e-09,
  2.487781e-08, 2.395488e-08, 2.375081e-08, 2.168174e-08, 1.852194e-08, 
    1.5658e-08, 1.285261e-08, 1.061326e-08, 8.91017e-09, 6.189703e-09, 
    4.22824e-09, 4.047747e-09, 3.850332e-09, 4.422708e-09, 4.564788e-09,
  2.566827e-08, 2.430564e-08, 2.394445e-08, 2.286778e-08, 2.018508e-08, 
    1.766606e-08, 1.489347e-08, 1.21727e-08, 9.910735e-09, 7.344984e-09, 
    5.435123e-09, 5.070893e-09, 4.494348e-09, 4.468976e-09, 4.600351e-09,
  2.63646e-08, 2.501139e-08, 2.408832e-08, 2.366367e-08, 2.15456e-08, 
    1.915186e-08, 1.668997e-08, 1.394528e-08, 1.132269e-08, 8.750259e-09, 
    6.691398e-09, 6.129669e-09, 5.265668e-09, 4.533852e-09, 4.678811e-09,
  1.959937e-08, 1.72058e-08, 1.475093e-08, 1.180552e-08, 8.358273e-09, 
    5.560168e-09, 3.994486e-09, 2.572699e-09, 1.416361e-09, 9.45564e-10, 
    7.637084e-10, 6.424006e-10, 6.805853e-10, 5.925754e-10, 6.143633e-10,
  2.023782e-08, 1.759379e-08, 1.520065e-08, 1.247658e-08, 9.213707e-09, 
    6.298267e-09, 4.343968e-09, 2.868018e-09, 1.643004e-09, 1.105659e-09, 
    7.960643e-10, 6.30434e-10, 5.286703e-10, 6.016286e-10, 5.610655e-10,
  2.119992e-08, 1.794439e-08, 1.549911e-08, 1.28809e-08, 9.894154e-09, 
    7.150844e-09, 4.851993e-09, 3.245117e-09, 1.836913e-09, 1.24435e-09, 
    8.690274e-10, 6.504867e-10, 5.634387e-10, 6.169684e-10, 6.689532e-10,
  2.231935e-08, 1.847195e-08, 1.603137e-08, 1.326854e-08, 1.029267e-08, 
    7.922223e-09, 5.418358e-09, 3.624268e-09, 2.005419e-09, 1.368447e-09, 
    9.776789e-10, 6.719326e-10, 5.369269e-10, 5.737366e-10, 6.703377e-10,
  2.348671e-08, 1.940491e-08, 1.615457e-08, 1.351039e-08, 1.091995e-08, 
    8.714474e-09, 6.074439e-09, 4.073692e-09, 2.22158e-09, 1.45536e-09, 
    1.095039e-09, 7.720775e-10, 5.453463e-10, 5.606393e-10, 6.267822e-10,
  2.34719e-08, 2.005361e-08, 1.667567e-08, 1.410656e-08, 1.11802e-08, 
    8.87825e-09, 6.56506e-09, 4.359646e-09, 2.470562e-09, 1.517848e-09, 
    1.187781e-09, 9.790595e-10, 7.241839e-10, 6.321426e-10, 6.331453e-10,
  2.400221e-08, 2.091593e-08, 1.72727e-08, 1.401447e-08, 1.127079e-08, 
    8.919592e-09, 6.929921e-09, 4.767683e-09, 2.783935e-09, 1.77316e-09, 
    1.437213e-09, 1.210405e-09, 9.014864e-10, 7.504318e-10, 7.262152e-10,
  2.464367e-08, 2.156196e-08, 1.776075e-08, 1.447591e-08, 1.116096e-08, 
    9.338544e-09, 7.166925e-09, 5.144851e-09, 3.240111e-09, 2.322589e-09, 
    1.794937e-09, 1.390798e-09, 9.861285e-10, 8.20901e-10, 7.012965e-10,
  2.529049e-08, 2.240053e-08, 1.85233e-08, 1.432341e-08, 1.082057e-08, 
    9.352936e-09, 7.32296e-09, 5.612597e-09, 3.902235e-09, 2.915317e-09, 
    2.116616e-09, 1.545636e-09, 1.109559e-09, 9.469986e-10, 6.680221e-10,
  2.659096e-08, 2.327162e-08, 1.904487e-08, 1.45443e-08, 1.135741e-08, 
    9.275815e-09, 7.335954e-09, 5.804579e-09, 4.17278e-09, 3.136445e-09, 
    2.245873e-09, 1.657985e-09, 1.209085e-09, 9.978345e-10, 7.050668e-10,
  2.750831e-08, 2.473818e-08, 2.311446e-08, 2.104967e-08, 1.773792e-08, 
    1.358134e-08, 8.354862e-09, 4.507896e-09, 2.037599e-09, 1.124657e-09, 
    1.049277e-09, 8.803072e-10, 6.60476e-10, 4.515337e-10, 3.6175e-10,
  2.594918e-08, 2.596429e-08, 2.455707e-08, 2.202911e-08, 1.903476e-08, 
    1.535004e-08, 1.041861e-08, 5.445845e-09, 2.718119e-09, 1.414866e-09, 
    1.159376e-09, 8.225419e-10, 5.761845e-10, 3.329296e-10, 2.388104e-10,
  2.556122e-08, 2.452647e-08, 2.472629e-08, 2.306399e-08, 2.027756e-08, 
    1.675615e-08, 1.202976e-08, 6.62119e-09, 3.453311e-09, 1.80044e-09, 
    1.201111e-09, 7.426009e-10, 4.585373e-10, 4.129247e-10, 2.234395e-10,
  2.553372e-08, 2.367347e-08, 2.360663e-08, 2.279686e-08, 2.093254e-08, 
    1.785351e-08, 1.350038e-08, 8.152905e-09, 4.029304e-09, 2.342723e-09, 
    1.307952e-09, 7.736209e-10, 4.445792e-10, 3.947389e-10, 2.543497e-10,
  2.421926e-08, 2.342194e-08, 2.260195e-08, 2.175326e-08, 2.070894e-08, 
    1.799294e-08, 1.423231e-08, 9.338409e-09, 4.810692e-09, 2.918191e-09, 
    1.546791e-09, 9.261423e-10, 5.583787e-10, 3.80149e-10, 3.093644e-10,
  2.327757e-08, 2.264045e-08, 2.174854e-08, 2.061626e-08, 1.982951e-08, 
    1.813159e-08, 1.467568e-08, 1.011958e-08, 5.793375e-09, 3.416796e-09, 
    2.039674e-09, 1.183482e-09, 5.734664e-10, 3.988503e-10, 3.457148e-10,
  2.322491e-08, 2.22617e-08, 2.132587e-08, 2.002003e-08, 1.935427e-08, 
    1.747327e-08, 1.442209e-08, 1.003567e-08, 6.346401e-09, 3.850585e-09, 
    2.430149e-09, 1.362865e-09, 6.119441e-10, 3.738919e-10, 3.524205e-10,
  2.336574e-08, 2.228329e-08, 2.110305e-08, 2.005999e-08, 1.922359e-08, 
    1.787802e-08, 1.436721e-08, 1.026501e-08, 6.814822e-09, 4.286982e-09, 
    2.795082e-09, 1.632755e-09, 6.640426e-10, 3.992649e-10, 3.506439e-10,
  2.388596e-08, 2.283073e-08, 2.1804e-08, 2.086475e-08, 1.964836e-08, 
    1.716467e-08, 1.335656e-08, 9.987533e-09, 7.222767e-09, 4.461398e-09, 
    3.018503e-09, 1.854727e-09, 7.285469e-10, 3.89341e-10, 3.514745e-10,
  2.47433e-08, 2.366675e-08, 2.155836e-08, 1.937478e-08, 1.784173e-08, 
    1.594174e-08, 1.22657e-08, 9.895891e-09, 7.369869e-09, 4.913612e-09, 
    3.328697e-09, 2.07921e-09, 9.876335e-10, 4.573499e-10, 4.025665e-10,
  1.686769e-08, 1.589162e-08, 1.48281e-08, 1.34106e-08, 1.052254e-08, 
    7.666511e-09, 5.002949e-09, 3.130409e-09, 2.290776e-09, 1.668607e-09, 
    1.45119e-09, 1.257322e-09, 1.030919e-09, 1.094953e-09, 1.038198e-09,
  1.831802e-08, 1.751765e-08, 1.609188e-08, 1.474333e-08, 1.206286e-08, 
    9.098471e-09, 6.121966e-09, 3.723115e-09, 2.515661e-09, 1.726414e-09, 
    1.586915e-09, 1.363859e-09, 1.065234e-09, 1.039585e-09, 1.137963e-09,
  1.881185e-08, 1.896658e-08, 1.792236e-08, 1.651436e-08, 1.374749e-08, 
    1.04477e-08, 7.432702e-09, 4.515344e-09, 2.892365e-09, 2.011641e-09, 
    1.707734e-09, 1.458037e-09, 1.198225e-09, 1.011113e-09, 1.049852e-09,
  1.897978e-08, 1.969221e-08, 1.921993e-08, 1.788785e-08, 1.570004e-08, 
    1.206706e-08, 8.717038e-09, 5.417871e-09, 3.452045e-09, 2.28278e-09, 
    1.902479e-09, 1.48981e-09, 1.257226e-09, 1.120755e-09, 1.014787e-09,
  1.963589e-08, 1.996875e-08, 2.084384e-08, 1.958107e-08, 1.757361e-08, 
    1.392245e-08, 1.011207e-08, 6.427967e-09, 4.219494e-09, 2.973758e-09, 
    2.092757e-09, 1.513944e-09, 1.220565e-09, 1.154147e-09, 9.371782e-10,
  2.029827e-08, 1.992998e-08, 2.106401e-08, 2.121615e-08, 1.98547e-08, 
    1.592652e-08, 1.133846e-08, 7.319736e-09, 5.015395e-09, 3.580845e-09, 
    2.361977e-09, 1.550134e-09, 1.306777e-09, 1.144775e-09, 1.009934e-09,
  2.168215e-08, 2.08795e-08, 2.132292e-08, 2.26956e-08, 2.157111e-08, 
    1.790194e-08, 1.280617e-08, 8.347477e-09, 5.755248e-09, 4.293836e-09, 
    2.998532e-09, 2.004392e-09, 1.42625e-09, 1.226821e-09, 1.069869e-09,
  2.525279e-08, 2.20297e-08, 2.168919e-08, 2.260448e-08, 2.351208e-08, 
    1.952543e-08, 1.438574e-08, 9.871282e-09, 6.883997e-09, 5.240052e-09, 
    3.770233e-09, 2.656189e-09, 1.757232e-09, 1.254267e-09, 1.16024e-09,
  2.885551e-08, 2.432893e-08, 2.166523e-08, 2.255199e-08, 2.390513e-08, 
    2.09075e-08, 1.547809e-08, 1.071205e-08, 7.577198e-09, 5.818581e-09, 
    4.358779e-09, 3.176577e-09, 2.125979e-09, 1.604066e-09, 1.276813e-09,
  3.07832e-08, 2.798258e-08, 2.347052e-08, 2.291683e-08, 2.436244e-08, 
    2.266428e-08, 1.610998e-08, 1.098109e-08, 7.580074e-09, 5.676976e-09, 
    4.404077e-09, 3.273712e-09, 2.322323e-09, 1.909427e-09, 1.50615e-09,
  4.626936e-09, 2.839023e-09, 2.136515e-09, 2.000919e-09, 1.773467e-09, 
    1.565735e-09, 1.160386e-09, 9.850045e-10, 1.140341e-09, 1.481251e-09, 
    1.574568e-09, 1.505405e-09, 1.435367e-09, 1.223562e-09, 1.339568e-09,
  5.392298e-09, 3.257927e-09, 2.264527e-09, 1.919017e-09, 1.732438e-09, 
    1.631253e-09, 1.350472e-09, 1.190878e-09, 1.107851e-09, 1.164793e-09, 
    1.398023e-09, 1.60315e-09, 1.758626e-09, 1.496241e-09, 1.415761e-09,
  6.946531e-09, 4.199844e-09, 2.845911e-09, 2.153964e-09, 1.750546e-09, 
    1.646321e-09, 1.541825e-09, 1.419891e-09, 1.218842e-09, 1.098031e-09, 
    1.087017e-09, 1.278839e-09, 1.458563e-09, 1.200448e-09, 1.086468e-09,
  9.026963e-09, 5.510287e-09, 3.636509e-09, 2.6518e-09, 1.995755e-09, 
    1.733511e-09, 1.643748e-09, 1.594923e-09, 1.470955e-09, 1.317949e-09, 
    1.071104e-09, 1.062021e-09, 1.017929e-09, 8.088469e-10, 4.559745e-10,
  1.050147e-08, 7.049023e-09, 4.423614e-09, 3.387282e-09, 2.505491e-09, 
    1.947559e-09, 1.751057e-09, 1.659542e-09, 1.513495e-09, 1.39203e-09, 
    1.259474e-09, 1.080911e-09, 8.041159e-10, 5.4658e-10, 2.452616e-10,
  1.106567e-08, 8.150865e-09, 5.380437e-09, 3.79847e-09, 3.148857e-09, 
    2.375876e-09, 2.036471e-09, 1.755516e-09, 1.579811e-09, 1.399919e-09, 
    1.279464e-09, 1.092047e-09, 7.823888e-10, 6.020444e-10, 4.296633e-10,
  1.13832e-08, 8.770485e-09, 6.491067e-09, 4.574784e-09, 3.512305e-09, 
    2.826144e-09, 2.349393e-09, 2.043538e-09, 1.829269e-09, 1.570223e-09, 
    1.38103e-09, 1.168301e-09, 9.01927e-10, 7.647136e-10, 7.27881e-10,
  1.117376e-08, 8.929077e-09, 7.473793e-09, 5.680963e-09, 4.272922e-09, 
    3.532433e-09, 2.838001e-09, 2.476044e-09, 2.281928e-09, 1.99586e-09, 
    1.739045e-09, 1.460721e-09, 1.023909e-09, 8.679282e-10, 9.200825e-10,
  9.97876e-09, 9.075474e-09, 8.840513e-09, 7.221749e-09, 5.481105e-09, 
    4.579004e-09, 4.008377e-09, 3.353821e-09, 2.911031e-09, 2.475707e-09, 
    1.992568e-09, 1.779996e-09, 1.309868e-09, 9.677655e-10, 8.080838e-10,
  9.611899e-09, 9.259642e-09, 9.062596e-09, 7.953354e-09, 6.8858e-09, 
    5.869192e-09, 5.08545e-09, 4.561179e-09, 3.900881e-09, 3.24333e-09, 
    2.616867e-09, 2.22515e-09, 1.7793e-09, 1.252448e-09, 8.755212e-10,
  3.84219e-09, 2.252841e-09, 1.457888e-09, 1.139822e-09, 7.874757e-10, 
    5.176871e-10, 5.814406e-10, 4.863591e-10, 4.259193e-10, 4.597216e-10, 
    2.541623e-10, 1.652818e-10, 7.577603e-11, 4.411111e-11, 1.051044e-10,
  4.708026e-09, 3.116286e-09, 1.894098e-09, 1.345767e-09, 1.003023e-09, 
    6.559271e-10, 6.197582e-10, 6.074525e-10, 4.750619e-10, 4.54837e-10, 
    3.388615e-10, 2.373209e-10, 1.348986e-10, 9.926738e-11, 1.090999e-10,
  5.925346e-09, 4.105098e-09, 2.511798e-09, 1.57921e-09, 1.16435e-09, 
    8.639458e-10, 6.88614e-10, 6.675328e-10, 6.064821e-10, 4.89174e-10, 
    3.957986e-10, 2.588144e-10, 1.980137e-10, 1.986389e-10, 2.16131e-10,
  7.678532e-09, 5.18878e-09, 3.193552e-09, 1.822884e-09, 1.227777e-09, 
    1.023306e-09, 7.827974e-10, 7.688861e-10, 7.402752e-10, 5.599555e-10, 
    4.399134e-10, 3.302604e-10, 2.541173e-10, 2.948176e-10, 3.421097e-10,
  1.068034e-08, 6.71754e-09, 3.820186e-09, 2.114119e-09, 1.387123e-09, 
    1.09983e-09, 9.348486e-10, 8.078589e-10, 7.958023e-10, 6.408734e-10, 
    5.062307e-10, 3.85224e-10, 3.010533e-10, 3.240433e-10, 4.044084e-10,
  1.317066e-08, 8.430412e-09, 4.879904e-09, 2.660442e-09, 1.700189e-09, 
    1.161119e-09, 1.051664e-09, 8.731336e-10, 8.519087e-10, 7.633111e-10, 
    6.581139e-10, 5.309219e-10, 3.782848e-10, 3.867603e-10, 3.935288e-10,
  1.559385e-08, 1.058338e-08, 6.244802e-09, 3.548472e-09, 2.16764e-09, 
    1.332379e-09, 1.066863e-09, 9.331723e-10, 8.840937e-10, 8.170016e-10, 
    7.652048e-10, 6.928591e-10, 5.012654e-10, 4.40239e-10, 3.98586e-10,
  1.758101e-08, 1.34702e-08, 8.043784e-09, 4.500241e-09, 2.742395e-09, 
    1.720015e-09, 1.221246e-09, 1.039987e-09, 1.008076e-09, 8.611875e-10, 
    7.973475e-10, 7.491089e-10, 6.438845e-10, 5.367877e-10, 4.921545e-10,
  1.896538e-08, 1.55716e-08, 9.954777e-09, 5.530768e-09, 3.40635e-09, 
    2.217591e-09, 1.442767e-09, 1.127596e-09, 1.109836e-09, 9.491892e-10, 
    8.231903e-10, 7.80818e-10, 7.166515e-10, 6.130478e-10, 5.482345e-10,
  1.946107e-08, 1.655835e-08, 1.158053e-08, 6.610029e-09, 4.058204e-09, 
    2.655725e-09, 1.720582e-09, 1.21724e-09, 1.110221e-09, 1.056291e-09, 
    9.447855e-10, 8.429167e-10, 8.15407e-10, 6.838536e-10, 6.056606e-10,
  3.01253e-09, 2.390625e-09, 1.815388e-09, 1.564072e-09, 1.086209e-09, 
    8.792898e-10, 7.607362e-10, 4.888087e-10, 3.482376e-10, 1.972258e-10, 
    2.501716e-10, 1.509507e-10, -1.214095e-10, -2.659748e-10, -1.028948e-10,
  3.374596e-09, 2.502364e-09, 1.957957e-09, 1.622338e-09, 1.182202e-09, 
    8.959061e-10, 8.278769e-10, 6.741723e-10, 4.419202e-10, 2.196096e-10, 
    7.830996e-11, 7.760298e-11, -7.868488e-12, -1.580627e-10, -1.780623e-10,
  3.772774e-09, 2.824339e-09, 2.151125e-09, 1.719124e-09, 1.214027e-09, 
    9.635212e-10, 7.695041e-10, 7.664465e-10, 5.84949e-10, 3.198405e-10, 
    9.984843e-11, 2.491785e-11, -5.358832e-11, -1.09649e-10, -1.271643e-10,
  4.380606e-09, 3.218632e-09, 2.375677e-09, 1.87802e-09, 1.308308e-09, 
    1.07693e-09, 8.965521e-10, 8.268567e-10, 7.892924e-10, 4.878073e-10, 
    2.2049e-10, 1.419076e-10, 8.902e-11, 4.411661e-11, 1.101662e-10,
  6.153924e-09, 3.544883e-09, 2.687489e-09, 2.03988e-09, 1.33257e-09, 
    1.051331e-09, 9.710301e-10, 9.516274e-10, 8.045309e-10, 6.488284e-10, 
    3.403054e-10, 2.875115e-10, 2.700173e-10, 2.807375e-10, 2.813915e-10,
  6.980812e-09, 4.540628e-09, 2.900167e-09, 2.304863e-09, 1.561811e-09, 
    9.868946e-10, 8.87715e-10, 7.829941e-10, 8.15794e-10, 8.023567e-10, 
    5.097112e-10, 3.609847e-10, 3.337765e-10, 2.894907e-10, 2.719355e-10,
  8.441831e-09, 5.928595e-09, 3.567797e-09, 2.657683e-09, 1.896211e-09, 
    1.181287e-09, 7.830186e-10, 6.90986e-10, 8.703384e-10, 8.446471e-10, 
    6.542033e-10, 3.920297e-10, 3.759132e-10, 3.19642e-10, 2.518268e-10,
  1.095945e-08, 7.779825e-09, 4.940442e-09, 3.186379e-09, 2.513675e-09, 
    1.438074e-09, 1.010473e-09, 8.559768e-10, 8.333518e-10, 9.896429e-10, 
    7.619881e-10, 5.039371e-10, 4.332038e-10, 4.122571e-10, 3.294089e-10,
  1.366773e-08, 1.005893e-08, 6.768696e-09, 3.943892e-09, 2.968727e-09, 
    1.963852e-09, 1.232309e-09, 1.090346e-09, 8.632316e-10, 9.752508e-10, 
    8.151321e-10, 6.484017e-10, 5.567381e-10, 5.138204e-10, 4.287313e-10,
  1.533278e-08, 1.293308e-08, 9.070077e-09, 5.222406e-09, 3.692236e-09, 
    2.745713e-09, 1.593259e-09, 1.207386e-09, 1.001155e-09, 9.509304e-10, 
    9.025982e-10, 7.488568e-10, 7.58652e-10, 6.574318e-10, 4.361975e-10,
  7.340334e-09, 3.992921e-09, 2.084594e-09, 1.12212e-09, 6.884671e-10, 
    7.416741e-10, 5.14046e-10, 2.226892e-10, 1.67366e-10, 2.769453e-10, 
    3.586548e-10, 4.005653e-10, 5.414109e-10, 6.253986e-10, 5.717147e-10,
  9.795988e-09, 5.08641e-09, 2.64104e-09, 1.313731e-09, 6.623505e-10, 
    6.957772e-10, 6.744228e-10, 4.679815e-10, 2.343297e-10, 2.264199e-10, 
    4.635548e-10, 4.755836e-10, 3.942008e-10, 4.338303e-10, 4.59115e-10,
  1.259327e-08, 6.66996e-09, 3.476012e-09, 1.596211e-09, 7.054828e-10, 
    6.273544e-10, 6.962754e-10, 6.195384e-10, 4.252289e-10, 3.59738e-10, 
    4.929524e-10, 6.303185e-10, 3.895426e-10, 2.67927e-10, 2.521006e-10,
  1.428076e-08, 8.862625e-09, 4.532428e-09, 2.051642e-09, 9.184076e-10, 
    6.378355e-10, 7.838875e-10, 7.288402e-10, 6.177519e-10, 6.001419e-10, 
    5.314495e-10, 7.504159e-10, 4.720647e-10, 3.343964e-10, 2.039513e-10,
  1.56668e-08, 1.091153e-08, 6.048849e-09, 2.790042e-09, 1.136033e-09, 
    6.832748e-10, 7.247083e-10, 7.560146e-10, 6.686722e-10, 8.172739e-10, 
    7.011627e-10, 6.076604e-10, 6.015509e-10, 3.998505e-10, 1.957908e-10,
  1.550366e-08, 1.232217e-08, 7.88893e-09, 3.724282e-09, 1.550168e-09, 
    8.79198e-10, 6.337299e-10, 7.415771e-10, 7.231238e-10, 8.026296e-10, 
    7.115502e-10, 5.816339e-10, 6.860051e-10, 5.751391e-10, 3.024113e-10,
  1.57044e-08, 1.340719e-08, 9.642169e-09, 5.017753e-09, 2.087908e-09, 
    1.08201e-09, 7.080538e-10, 7.150864e-10, 7.335217e-10, 6.556057e-10, 
    6.128604e-10, 5.894288e-10, 6.222908e-10, 5.972926e-10, 3.567084e-10,
  1.49843e-08, 1.365388e-08, 1.043258e-08, 6.375437e-09, 3.085681e-09, 
    1.4041e-09, 1.042182e-09, 7.436912e-10, 7.065392e-10, 6.502152e-10, 
    6.19268e-10, 5.941207e-10, 5.432905e-10, 5.226728e-10, 4.350238e-10,
  1.408637e-08, 1.373745e-08, 1.093701e-08, 7.281157e-09, 4.050267e-09, 
    1.949935e-09, 1.237467e-09, 1.050319e-09, 8.006009e-10, 5.583503e-10, 
    5.145045e-10, 5.416261e-10, 4.955618e-10, 5.036736e-10, 4.475265e-10,
  1.331874e-08, 1.344953e-08, 1.113288e-08, 7.71129e-09, 5.132107e-09, 
    2.658e-09, 1.609922e-09, 1.189056e-09, 1.143882e-09, 7.559314e-10, 
    4.414542e-10, 3.859391e-10, 3.992357e-10, 3.823116e-10, 3.970632e-10,
  2.149147e-08, 1.891283e-08, 1.534244e-08, 1.035861e-08, 6.988126e-09, 
    4.987502e-09, 3.404438e-09, 2.351296e-09, 1.274931e-09, 5.774516e-10, 
    2.660093e-10, 1.993697e-10, 1.779421e-10, 2.445422e-10, 3.018137e-10,
  2.33633e-08, 2.008583e-08, 1.657175e-08, 1.192412e-08, 7.988765e-09, 
    5.447967e-09, 3.676343e-09, 2.564659e-09, 1.418795e-09, 6.314746e-10, 
    2.990084e-10, 2.050354e-10, 1.820302e-10, 2.667697e-10, 4.34238e-10,
  2.465942e-08, 2.160304e-08, 1.803389e-08, 1.327125e-08, 9.122198e-09, 
    5.960639e-09, 3.985305e-09, 2.7623e-09, 1.579089e-09, 6.881831e-10, 
    3.284034e-10, 1.934761e-10, 1.584027e-10, 2.282031e-10, 4.001845e-10,
  2.572681e-08, 2.219939e-08, 1.934544e-08, 1.476899e-08, 1.02929e-08, 
    6.655861e-09, 4.264901e-09, 2.897514e-09, 1.762228e-09, 7.748509e-10, 
    3.49342e-10, 1.97652e-10, 1.486912e-10, 1.899852e-10, 3.522805e-10,
  2.658422e-08, 2.353328e-08, 2.053909e-08, 1.598368e-08, 1.139846e-08, 
    7.418437e-09, 4.711306e-09, 3.071765e-09, 1.959943e-09, 8.866726e-10, 
    3.758824e-10, 1.983442e-10, 1.393019e-10, 1.371332e-10, 3.501123e-10,
  2.420273e-08, 2.287302e-08, 2.106105e-08, 1.717346e-08, 1.23869e-08, 
    8.364758e-09, 5.008197e-09, 3.179316e-09, 2.090743e-09, 1.029518e-09, 
    4.199875e-10, 1.898052e-10, 9.304377e-11, 1.034715e-10, 2.368295e-10,
  2.582476e-08, 2.435766e-08, 2.166728e-08, 1.80114e-08, 1.319671e-08, 
    9.147694e-09, 5.669061e-09, 3.400689e-09, 2.19561e-09, 1.156738e-09, 
    4.681553e-10, 1.65508e-10, 1.062378e-10, 7.949023e-11, 1.494445e-10,
  2.621253e-08, 2.422669e-08, 2.209597e-08, 1.873327e-08, 1.407517e-08, 
    9.845145e-09, 6.097092e-09, 3.64887e-09, 2.350289e-09, 1.29742e-09, 
    5.247956e-10, 1.724271e-10, 1.369435e-10, 6.515695e-11, 9.706941e-11,
  2.539582e-08, 2.381141e-08, 2.206984e-08, 1.951289e-08, 1.469579e-08, 
    1.037079e-08, 6.602332e-09, 3.783749e-09, 2.347108e-09, 1.374005e-09, 
    5.822973e-10, 1.85462e-10, 1.194063e-10, 1.039062e-10, 1.068123e-10,
  2.40542e-08, 2.390445e-08, 2.186077e-08, 1.982508e-08, 1.4926e-08, 
    1.061049e-08, 7.082327e-09, 3.939515e-09, 2.351074e-09, 1.447647e-09, 
    6.581494e-10, 2.141856e-10, 1.038731e-10, 1.069202e-10, 1.39061e-10,
  2.548053e-08, 2.446496e-08, 2.1873e-08, 1.756228e-08, 1.486206e-08, 
    1.197313e-08, 9.244433e-09, 6.613416e-09, 4.898032e-09, 3.666278e-09, 
    2.490605e-09, 1.19332e-09, 2.748111e-10, 5.956866e-11, 2.12054e-10,
  2.620775e-08, 2.540994e-08, 2.285693e-08, 1.895148e-08, 1.52885e-08, 
    1.24384e-08, 9.50882e-09, 6.806873e-09, 4.903614e-09, 3.543834e-09, 
    2.36298e-09, 1.073101e-09, 1.927397e-10, 3.132675e-11, 2.952964e-10,
  2.665716e-08, 2.679079e-08, 2.363498e-08, 1.990539e-08, 1.583589e-08, 
    1.27861e-08, 9.814339e-09, 6.991225e-09, 4.849056e-09, 3.443636e-09, 
    2.265991e-09, 9.462066e-10, 1.576412e-10, 3.178308e-12, 3.718137e-10,
  2.658724e-08, 2.682879e-08, 2.462373e-08, 2.086361e-08, 1.635311e-08, 
    1.315398e-08, 1.001417e-08, 7.121652e-09, 4.768935e-09, 3.327969e-09, 
    2.174927e-09, 8.266629e-10, 1.515203e-10, 2.656233e-11, 4.428748e-10,
  2.605482e-08, 2.703614e-08, 2.530012e-08, 2.146564e-08, 1.683967e-08, 
    1.343518e-08, 1.029043e-08, 7.310322e-09, 4.663171e-09, 3.167383e-09, 
    2.083961e-09, 7.178648e-10, 1.649946e-10, 8.746408e-11, 4.546033e-10,
  2.517876e-08, 2.661275e-08, 2.626032e-08, 2.2068e-08, 1.739292e-08, 
    1.370013e-08, 1.034386e-08, 7.243045e-09, 4.484135e-09, 2.993351e-09, 
    1.949967e-09, 6.334994e-10, 1.563943e-10, 1.81821e-10, 4.741444e-10,
  2.462663e-08, 2.600969e-08, 2.714593e-08, 2.26696e-08, 1.773689e-08, 
    1.39797e-08, 1.054674e-08, 7.214142e-09, 4.300667e-09, 2.849465e-09, 
    1.806794e-09, 5.207031e-10, 9.587922e-11, 2.308281e-10, 4.230641e-10,
  2.496914e-08, 2.551089e-08, 2.721186e-08, 2.301959e-08, 1.838126e-08, 
    1.422068e-08, 1.053769e-08, 7.29628e-09, 4.325202e-09, 2.754186e-09, 
    1.621871e-09, 4.189764e-10, 5.284678e-11, 2.964636e-10, 4.014095e-10,
  2.496494e-08, 2.514846e-08, 2.684034e-08, 2.388913e-08, 1.878227e-08, 
    1.455039e-08, 1.051206e-08, 7.075138e-09, 4.121327e-09, 2.512223e-09, 
    1.447077e-09, 3.436487e-10, 6.912412e-11, 3.309793e-10, 3.408095e-10,
  2.538594e-08, 2.512168e-08, 2.630381e-08, 2.404671e-08, 1.92728e-08, 
    1.486813e-08, 1.035311e-08, 6.889278e-09, 3.894282e-09, 2.304988e-09, 
    1.2961e-09, 3.25954e-10, 1.025711e-10, 3.076968e-10, 3.113753e-10 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.2466774, 0.6143242, 0.0668168, 0.2301621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.4924844, 0.2132108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.600569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1560082, 0,
  1, 1, 0.7132517, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02739768, 0,
  0.6230268, 0.6280472, 0.3043983, 0.08344039, 0, 0.3148882, 0.01188002, 0, 
    0, 0, 0, 0.08803581, 0, 0, 0,
  0, 0, 0, 0, 0.01144353, 0.8597386, 0.8205094, 0.5086318, 0.1258651, 
    0.08909279, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.291879, 0.6933324, 1, 0.9996726, 0.6666086, 0.08008575, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.611689, 0.7180831, 0.4623523, 0.2838529, 0.02767258, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0.002817577, 0.8915156, 0.5654301, 0.7485356, 0.3018697, 0, 0, 0, 
    0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0.04916316, 0.5638732, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3486554,
  2.316188, 6.745579, 0.5592819, 0.3199724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  147.4583, 171.3604, 6.513342, 0.3383408, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03840884, 0.4204801, 0,
  316.1323, 305.6766, 15.46485, 0.007546596, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1807817, 1.695307, 0,
  309.9182, 276.4409, 123.1236, 0.0108671, 0, 1.460928, 0.05467265, 0, 0, 0, 
    0.009753421, 0.03281464, 0.7768181, 0.4781904, 0,
  365.1592, 241.1036, 8.988194, 1.559117, 0.4356286, 6.775464, 0.2077458, 
    1.032432, 0.002793631, 0.1432027, 0.862155, 4.338077, 0.2366837, 0, 0,
  0, 0, 0, 0, 0.1289662, 151.094, 22.45284, 14.93281, 5.254983, 2.574013, 
    0.002986824, 0.1528066, 0.0002596498, 0, 0,
  0, 0, 0, 0, 13.93511, 217.993, 380.8379, 455.4515, 234.498, 2.407733, 0, 0, 
    0, 0, 0,
  0, 0.0003258124, 0, 0, 414.0298, 282.8423, 143.9435, 10.21257, 0.1187258, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 1.536109, 363.0271, 340.0019, 397.2344, 11.61882, 0, 0, 0, 0, 0, 
    0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
