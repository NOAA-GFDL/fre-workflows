netcdf \00010101.atmos_daily.tile2.ps {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float ps(time, grid_yt, grid_xt) ;
		ps:_FillValue = 1.e+20f ;
		ps:missing_value = 1.e+20f ;
		ps:units = "Pa" ;
		ps:long_name = "Surface Air Pressure" ;
		ps:cell_methods = "time: mean" ;
		ps:cell_measures = "area: area" ;
		ps:time_avg_info = "average_T1,average_T2,average_DT" ;
		ps:standard_name = "surface_air_pressure" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:53:56 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile2.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile2.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 ps =
  101701.9, 101652.7, 101613.4, 101565.4, 101512.9, 101459.3, 101410.1, 
    101364.3, 101323, 101290.6, 101261.1, 101241, 101230.8, 101235.9, 101253.5,
  101720.6, 101687, 101660.5, 101627.4, 101585.4, 101541.7, 101500.7, 
    101461.7, 101427.3, 101398.9, 101375.5, 101355.4, 101345.4, 101346, 
    101360.9,
  101725.9, 101706.7, 101691.2, 101665.4, 101633.6, 101600.9, 101566.1, 
    101538.1, 101509.4, 101483.4, 101464.7, 101450.8, 101443.8, 101447, 
    101460.1,
  101716.5, 101708, 101703.7, 101691.3, 101672.3, 101647.8, 101622.8, 
    101596.1, 101572.9, 101554.2, 101540.7, 101525.5, 101523.9, 101525.6, 
    101532.2,
  101690, 101707.5, 101703, 101699.9, 101689.5, 101676.6, 101659.1, 101641.2, 
    101624, 101608.7, 101596, 101588.7, 101588, 101588.7, 101590.3,
  101637.8, 101677.1, 101692.4, 101703.1, 101698.3, 101698.1, 101685.6, 
    101673.2, 101656, 101645.4, 101633.9, 101630.1, 101625.5, 101616.4, 
    101615.1,
  101596.6, 101643.8, 101662.4, 101692.1, 101694.6, 101698.2, 101695.3, 
    101688.2, 101680.4, 101668.6, 101660.1, 101651.9, 101641.4, 101634.1, 
    101630.5,
  101570.9, 101620.5, 101640.6, 101664.2, 101681.7, 101699, 101702.1, 
    101692.2, 101682.4, 101674.6, 101666.9, 101655.8, 101647.8, 101634.9, 
    101624.4,
  101550.3, 101602.4, 101622.6, 101649.9, 101662, 101668.2, 101682.2, 
    101684.8, 101678.8, 101669.6, 101659.2, 101643, 101624, 101610.2, 101591.5,
  101550.3, 101574.7, 101597, 101634.6, 101653.1, 101659.4, 101654.4, 
    101648.4, 101644.7, 101630.8, 101612.4, 101594.2, 101573.9, 101543.1, 
    101521,
  101851.3, 101787.3, 101710.8, 101627.6, 101535.5, 101441.2, 101334.5, 
    101228.2, 101115.2, 100999.6, 100882.8, 100770.2, 100660, 100555.6, 
    100457.8,
  101875.2, 101820.4, 101756.3, 101685.6, 101605.2, 101520.5, 101424.1, 
    101325.9, 101221, 101117.2, 101008.2, 100902.5, 100797.8, 100697.3, 
    100602.6,
  101890.9, 101842.3, 101784.4, 101720.5, 101652, 101576.3, 101492.9, 101403, 
    101309.2, 101213.9, 101115.7, 101015.5, 100920.6, 100823.9, 100736.1,
  101889, 101847.6, 101804.9, 101748.6, 101686.8, 101619.5, 101545.3, 
    101467.4, 101382.4, 101294.5, 101206, 101117.1, 101028.1, 100941.6, 
    100857.7,
  101876.9, 101844.3, 101805.8, 101757, 101702.4, 101644.8, 101577.8, 
    101507.6, 101432.4, 101355.6, 101274.6, 101196.8, 101117.5, 101041.4, 
    100965,
  101852, 101824.3, 101795.8, 101759.2, 101710.3, 101661.7, 101603.1, 
    101542.6, 101474.4, 101405.9, 101334.4, 101264.4, 101193.7, 101123.3, 
    101055.3,
  101825.7, 101802.5, 101771.3, 101743.7, 101703.8, 101662.3, 101613.9, 
    101561.8, 101503.8, 101441.6, 101379.3, 101317.1, 101254.9, 101191.6, 
    101130.5,
  101782.5, 101760.8, 101748.6, 101725.9, 101693.4, 101658.5, 101616.1, 
    101571.2, 101519.3, 101466.5, 101411.4, 101356.2, 101300.2, 101243, 
    101186.7,
  101732, 101714.6, 101704, 101696.1, 101673.9, 101646.4, 101611.7, 101573.6, 
    101528.7, 101479.1, 101430.1, 101380.5, 101331, 101281.3, 101229.6,
  101678.7, 101657, 101653.4, 101664.4, 101646.9, 101627.5, 101599.3, 
    101566.2, 101528, 101488.8, 101443.1, 101397.5, 101350.9, 101303.2, 
    101258.9,
  101719.9, 101652.7, 101592, 101526.7, 101465.8, 101398.2, 101326, 101250.3, 
    101168.2, 101083.3, 100993.8, 100903.4, 100811.5, 100714.6, 100618.3,
  101754.8, 101703.8, 101660.6, 101603.9, 101542.6, 101478.2, 101410.1, 
    101341, 101267.6, 101188.5, 101105.3, 101019.9, 100932.9, 100849.1, 
    100764.8,
  101795.8, 101761.4, 101716.9, 101665.6, 101614, 101553.6, 101490.8, 101424, 
    101356.5, 101287.9, 101213.6, 101135.3, 101055.1, 100974.5, 100896,
  101808.1, 101790.4, 101759.6, 101718.1, 101676.4, 101625.9, 101568.9, 
    101508.4, 101445, 101380.5, 101315.9, 101249.1, 101178.4, 101106.9, 
    101034.5,
  101813.8, 101803.6, 101786.2, 101759.8, 101721.4, 101680.2, 101633.3, 
    101581.9, 101526, 101468.3, 101407.6, 101345.5, 101283, 101220.3, 101155.8,
  101800.3, 101805.3, 101797.3, 101782.2, 101756, 101721.9, 101683.2, 
    101640.7, 101592.9, 101544.5, 101492.4, 101438.8, 101383.5, 101327.4, 
    101271.1,
  101781.6, 101789.5, 101792, 101787.9, 101773.7, 101745.9, 101715, 101681.4, 
    101642, 101598.9, 101554.4, 101508.5, 101459.8, 101411.8, 101364.2,
  101749, 101766.3, 101774.5, 101776.6, 101767.2, 101756.3, 101731.1, 
    101705.5, 101674.2, 101641.4, 101602.7, 101564.1, 101524.1, 101481.2, 
    101440.1,
  101719.7, 101733.1, 101745.1, 101750.2, 101749.4, 101746.4, 101731.2, 
    101715.1, 101689.1, 101659, 101629.3, 101601.3, 101567.6, 101533.1, 
    101497.5,
  101677.9, 101696.1, 101705.3, 101717.9, 101721.9, 101722.2, 101713.1, 
    101702.2, 101685.1, 101666.9, 101642.7, 101617.9, 101591, 101564.8, 
    101536.1,
  101633.1, 101637, 101639.5, 101635.5, 101632.4, 101648.9, 101650.6, 
    101657.3, 101649.9, 101647.5, 101641.2, 101631.7, 101608.5, 101578.7, 
    101544.4,
  101633.4, 101654, 101661.1, 101666.3, 101665.8, 101667.4, 101676.6, 
    101686.1, 101687.5, 101686.5, 101674.3, 101661.1, 101645.9, 101623.2, 
    101597.2,
  101631.8, 101675.2, 101687.4, 101695.4, 101692.8, 101693.6, 101696.6, 
    101709.4, 101715.8, 101720.8, 101719.5, 101707.8, 101691.2, 101670.7, 
    101647.3,
  101615, 101665.1, 101693, 101706.1, 101708.4, 101713.6, 101717.8, 101721.7, 
    101730.6, 101737.7, 101741.2, 101739.4, 101728.6, 101715.4, 101694.1,
  101584.3, 101640.8, 101687.8, 101720.9, 101727.4, 101724.1, 101727.9, 
    101732.2, 101740, 101747.6, 101751.9, 101754.8, 101754.4, 101748.8, 
    101736.8,
  101552.7, 101612.2, 101662.8, 101696, 101727.7, 101729.5, 101731.9, 
    101736.5, 101742.3, 101746.3, 101751.9, 101755.6, 101756.1, 101760.3, 
    101760,
  101519, 101576.4, 101631.1, 101670.6, 101704.2, 101717.1, 101726, 101732.1, 
    101736.5, 101743.3, 101749, 101755.2, 101761.7, 101761.6, 101766.8,
  101484.1, 101543.4, 101594.4, 101635.8, 101669.2, 101693.8, 101711.7, 
    101722.6, 101730.4, 101733.7, 101740.7, 101746.7, 101755.3, 101760.7, 
    101764.9,
  101445.8, 101503.4, 101552.4, 101599.6, 101635.2, 101661.9, 101681.3, 
    101699.9, 101712.7, 101720.1, 101730, 101736.7, 101743.9, 101750.7, 
    101757.4,
  101415.9, 101464.3, 101501.7, 101549.6, 101586.9, 101618, 101641.1, 
    101662.6, 101679.8, 101694.5, 101707.4, 101717.9, 101726.1, 101735.3, 
    101745.7,
  101328.1, 101414.9, 101494.6, 101570.1, 101643.2, 101709.6, 101779.5, 
    101850.5, 101927.6, 102010.5, 102089.9, 102171.2, 102251.9, 102326.4, 
    102406.7,
  101320.1, 101407.7, 101486.2, 101560.7, 101631.1, 101699.8, 101768.9, 
    101841.7, 101924.4, 102011.8, 102089.1, 102161.1, 102239.8, 102310.2, 
    102388.9,
  101309.5, 101390.2, 101462.6, 101539.4, 101610.2, 101681.2, 101751.4, 
    101822.9, 101902.5, 101986.8, 102075.6, 102153.3, 102229.8, 102295.3, 
    102364.8,
  101284.6, 101365.5, 101439, 101511.7, 101578.8, 101647.1, 101715.9, 101790, 
    101867.6, 101948, 102035, 102117.6, 102191.3, 102266.4, 102336.6,
  101266.9, 101338.8, 101407.3, 101474.8, 101539.7, 101605.8, 101672.6, 
    101743, 101819.1, 101898.6, 101979.7, 102067.6, 102145.2, 102224.3, 
    102295.6,
  101238.7, 101310, 101376, 101438.7, 101498.8, 101557, 101618.4, 101686.2, 
    101758.6, 101835.6, 101910.6, 101989.3, 102073.7, 102154.6, 102237.4,
  101207.5, 101279, 101340, 101400.1, 101454.7, 101508.4, 101560.2, 101621.8, 
    101689.1, 101763.7, 101841.7, 101918.4, 101997.9, 102080.9, 102167.3,
  101178.2, 101246, 101303.5, 101360.8, 101410.4, 101458.9, 101502.9, 
    101553.4, 101615.2, 101681.8, 101754.9, 101831.3, 101911.4, 101994.8, 
    102080.8,
  101148.7, 101218.8, 101271.3, 101322.3, 101365.4, 101409.4, 101448.2, 
    101490, 101543.2, 101604.8, 101671.8, 101746.9, 101825.1, 101905.4, 
    101989.7,
  101118.5, 101186.2, 101237.3, 101286.9, 101321.2, 101359.8, 101395.9, 
    101429.4, 101470.4, 101522.4, 101584.5, 101652.3, 101732.1, 101816.1, 
    101901.8,
  101292.6, 101282.2, 101277.7, 101275, 101270.7, 101271, 101281.9, 101314.2, 
    101354.4, 101401.7, 101461.8, 101533.4, 101614.9, 101705.2, 101800,
  101250.1, 101258, 101259.3, 101274.4, 101289.9, 101310.4, 101327, 101354.1, 
    101392.6, 101447.5, 101512.5, 101586.1, 101665.7, 101753.8, 101851.1,
  101198.4, 101218.4, 101216.3, 101242.8, 101270.1, 101294.9, 101318.1, 
    101362.4, 101415.5, 101478, 101545.2, 101620.9, 101702.2, 101794, 101890.4,
  101127.7, 101136.6, 101146.9, 101194.9, 101238.3, 101286.4, 101319.4, 
    101368.8, 101420.4, 101482.6, 101554.6, 101635.8, 101722.4, 101811.6, 
    101910.8,
  101052.2, 101055, 101079.6, 101152.9, 101204.5, 101263.4, 101301.7, 
    101351.8, 101408.4, 101476.4, 101554.9, 101638.6, 101722.9, 101816.1, 
    101919.8,
  101017.1, 101014, 101054.8, 101124.4, 101183, 101234, 101280, 101336.1, 
    101398.8, 101471.7, 101551.3, 101637.5, 101726.7, 101820.5, 101914.1,
  101024.4, 101012.3, 101044.5, 101109, 101167.2, 101215.9, 101267.2, 
    101322.9, 101385.7, 101458.9, 101540.9, 101629.4, 101716.8, 101807.4, 
    101896.7,
  101053.9, 101040.6, 101060.8, 101106.4, 101151.6, 101206.5, 101258.9, 
    101308.1, 101371.2, 101447.5, 101525.6, 101614, 101700.9, 101785.8, 101874,
  101069.1, 101069.5, 101089.7, 101121.6, 101152.6, 101196.2, 101245.7, 
    101293.4, 101351.6, 101421.7, 101502.2, 101589.2, 101673.6, 101756.1, 
    101838.3,
  101081.1, 101088.9, 101106.2, 101121.2, 101152.7, 101197.8, 101234.3, 
    101282.7, 101332.8, 101401.9, 101478.3, 101560.2, 101644, 101724.1, 101800,
  101761.3, 101777.5, 101786.8, 101802.2, 101812.8, 101823, 101838.2, 101861, 
    101891.6, 101921.4, 101953.1, 101981.8, 102002, 101997.8, 101991.8,
  101682.3, 101675.6, 101673.1, 101681, 101691.6, 101707.7, 101725.8, 
    101750.1, 101775, 101818.9, 101866.1, 101893.1, 101929.1, 101955.7, 
    101957.9,
  101599.3, 101588.9, 101587.3, 101596.2, 101611.6, 101628, 101632.4, 
    101646.9, 101683.1, 101748.2, 101793.9, 101836.8, 101875.3, 101887.5, 
    101918.1,
  101525.9, 101507.5, 101506.1, 101501.5, 101498.9, 101515.5, 101516.1, 
    101532.2, 101566.9, 101635.8, 101721.4, 101767.1, 101801.5, 101831.4, 
    101847.6,
  101454.5, 101423.1, 101391.9, 101379.9, 101375.5, 101393.6, 101396, 
    101409.4, 101416.1, 101453.6, 101537.7, 101638, 101721.2, 101780.8, 
    101813.9,
  101389.5, 101336.5, 101282.5, 101282.4, 101292, 101306.3, 101321, 101331, 
    101356.1, 101423.2, 101508.8, 101569.4, 101635.5, 101700.6, 101759.1,
  101343.8, 101273.2, 101212.4, 101225.9, 101238.2, 101269.1, 101276.8, 
    101316.4, 101356.1, 101405.3, 101450.9, 101524.5, 101596.1, 101670.3, 
    101729.6,
  101311.1, 101229.8, 101175.7, 101214.1, 101213.2, 101244.7, 101256.2, 
    101289.5, 101332.9, 101391.2, 101457.8, 101520.3, 101577.6, 101635.9, 
    101700,
  101289.6, 101206.8, 101156.8, 101189.7, 101194.8, 101229.2, 101235.5, 
    101268.5, 101313, 101377.7, 101438.1, 101508.1, 101553.5, 101608.6, 
    101667.1,
  101285.2, 101197.7, 101156.1, 101177.3, 101178.4, 101206.5, 101222.1, 
    101240.7, 101276.2, 101351.9, 101413.1, 101480.6, 101525.3, 101579.7, 
    101630.5,
  101252.8, 101223.4, 101218.3, 101212.7, 101202.1, 101181.8, 101141.5, 
    101113.3, 101088.8, 101091.6, 101091.7, 101125.1, 101183.5, 101252.8, 
    101338.8,
  101230.5, 101202.1, 101198.5, 101191, 101180.9, 101164.2, 101120.3, 101080, 
    101061.7, 101091.3, 101132.5, 101171.6, 101224.7, 101282, 101360.7,
  101205.2, 101183.8, 101172.2, 101163.8, 101160.9, 101153, 101128.3, 101099, 
    101092.2, 101112.2, 101134.6, 101172, 101231.7, 101298.3, 101374.3,
  101185.1, 101164.4, 101149.4, 101142, 101141.7, 101135.6, 101117, 101099.3, 
    101105.8, 101123, 101151.2, 101197.7, 101255.6, 101317.6, 101383.1,
  101160.5, 101138.1, 101129.4, 101119.4, 101117.2, 101122.2, 101111, 
    101099.2, 101106.1, 101121.2, 101157.3, 101199.8, 101245, 101308.3, 
    101375.4,
  101138.3, 101124.6, 101104.6, 101102, 101093.5, 101090.5, 101096.7, 
    101097.2, 101103.7, 101132, 101166.3, 101212.3, 101250.8, 101304.4, 
    101359.1,
  101128.8, 101117.2, 101091.3, 101086.3, 101084.9, 101086.6, 101086.9, 
    101093.7, 101109.1, 101127.8, 101165.5, 101204.6, 101246.9, 101288, 
    101338.1,
  101120.9, 101094.8, 101081.5, 101079.4, 101075.4, 101085.4, 101091.7, 
    101096.4, 101114.2, 101136.4, 101165.7, 101204.3, 101244.8, 101278.9, 
    101326.7,
  101097.3, 101081.3, 101075.7, 101069.5, 101079, 101088.2, 101091.2, 
    101098.1, 101115.4, 101133.3, 101168.2, 101200.2, 101233.5, 101270.1, 
    101308.6,
  101073.4, 101064.3, 101061.6, 101051, 101064.4, 101072.7, 101080.3, 
    101091.8, 101112, 101132.9, 101166.4, 101197.3, 101233.9, 101262.5, 
    101308.7,
  101427, 101430.3, 101429.3, 101424.8, 101417.8, 101410, 101405.7, 101396.1, 
    101392.4, 101385, 101373.2, 101355.7, 101329.1, 101305.4, 101284.8,
  101451.1, 101448.2, 101449.3, 101448.8, 101444.2, 101437.7, 101438.7, 
    101431.3, 101426.7, 101417, 101401.1, 101382.2, 101351.6, 101321.5, 
    101298.2,
  101446.9, 101441.2, 101452.9, 101451.7, 101453.2, 101447.8, 101448.3, 
    101440.2, 101433.3, 101428, 101410.8, 101386.7, 101354.2, 101325, 101298.1,
  101430, 101424.8, 101440.2, 101437.4, 101436.2, 101438, 101442.1, 101438.8, 
    101430.7, 101423.6, 101402.8, 101370.5, 101343.4, 101314.3, 101287.5,
  101389.4, 101393, 101396.5, 101396.7, 101402.3, 101415.8, 101418.6, 
    101415.1, 101407.6, 101396.6, 101372.6, 101343.6, 101326.7, 101299.4, 
    101277.6,
  101345, 101355.7, 101349.9, 101355.7, 101365.1, 101376.8, 101383.2, 
    101382.4, 101377.7, 101358.7, 101334.5, 101313.9, 101290.6, 101271.2, 
    101259.2,
  101295.4, 101301.6, 101298.3, 101311, 101312.6, 101329.3, 101340.8, 101346, 
    101344.6, 101324.8, 101302.2, 101286.8, 101264.6, 101246.8, 101241.5,
  101247.9, 101255.7, 101250.1, 101254.5, 101260.4, 101273.7, 101283.8, 
    101295.7, 101297.4, 101283.5, 101265.6, 101252.3, 101234.2, 101229.1, 
    101237.4,
  101199.1, 101201.3, 101195.5, 101193.7, 101200.4, 101214.6, 101230.9, 
    101239.6, 101247.1, 101242.5, 101234, 101226, 101219.7, 101222.6, 101235.7,
  101158.7, 101155.5, 101151.6, 101154.5, 101162.1, 101173.9, 101184.8, 
    101194.9, 101199.6, 101200.8, 101199, 101210, 101210.1, 101219.9, 101240,
  101610.1, 101640.6, 101673.3, 101700.4, 101715.9, 101736.6, 101741.2, 
    101742.4, 101733.9, 101730.9, 101751.2, 101776.4, 101800.9, 101808, 
    101834.8,
  101572.9, 101619.5, 101656.4, 101687.2, 101706.9, 101713.3, 101723.7, 
    101727.8, 101742.7, 101773.5, 101790, 101809.5, 101813.3, 101829.9, 
    101852.2,
  101525.8, 101582.6, 101627.9, 101661.5, 101693.9, 101709.2, 101732, 
    101740.3, 101755.5, 101765.4, 101766.4, 101773.1, 101776.1, 101790.1, 
    101801.8,
  101475.3, 101535, 101584.7, 101621, 101658.2, 101679.1, 101700.9, 101713.8, 
    101725.1, 101732.1, 101732.6, 101730.4, 101728.9, 101733.3, 101735.4,
  101428.6, 101483.2, 101529.1, 101577.1, 101610.6, 101641.1, 101660.2, 
    101669.7, 101676.7, 101675.5, 101670.2, 101663.9, 101653.4, 101642.2, 
    101639.8,
  101384.1, 101434.2, 101472.4, 101519.1, 101552.2, 101582.6, 101598.9, 
    101615.4, 101620.3, 101612.4, 101610.4, 101590.4, 101563.4, 101546.2, 
    101553.7,
  101335.3, 101382.1, 101420, 101462.4, 101494.5, 101526.4, 101545.9, 101554, 
    101554.4, 101546.8, 101540.1, 101509.9, 101486.2, 101471.3, 101492.9,
  101280.5, 101326.1, 101359.8, 101400.2, 101429.3, 101455.6, 101471.7, 
    101483.7, 101487.5, 101482.1, 101473.4, 101451.2, 101429.5, 101436.5, 
    101460.8,
  101235.2, 101275, 101299.9, 101332.5, 101362.1, 101387.4, 101406.9, 
    101415.2, 101422.5, 101418.8, 101411, 101396, 101389.6, 101403.4, 101428.8,
  101186.8, 101219.5, 101244.1, 101272.3, 101293.7, 101312.2, 101328.5, 
    101339.2, 101346.8, 101351.9, 101346.9, 101344.8, 101349, 101372, 101408.3,
  101797.3, 101841, 101877.6, 101903.9, 101921.2, 101924.4, 101924.9, 
    101915.3, 101899.7, 101875.9, 101858.2, 101843.1, 101829.2, 101814.6, 
    101811.1,
  101765.1, 101807.2, 101843.8, 101864.8, 101881.1, 101886.7, 101886, 
    101875.8, 101855.4, 101839.9, 101828.7, 101813, 101805.7, 101784, 101777.9,
  101718.9, 101763.3, 101803.6, 101823.4, 101842.4, 101841.6, 101842.9, 
    101834.1, 101822.2, 101810.3, 101796.3, 101778.4, 101758, 101737, 101718.2,
  101674.7, 101718.4, 101756.7, 101781, 101798.9, 101803.6, 101802.7, 
    101794.5, 101785.7, 101772.6, 101754.3, 101739.5, 101708.6, 101678.5, 
    101631.1,
  101623.1, 101665.8, 101701.9, 101729.9, 101747.7, 101755.9, 101755.5, 
    101749, 101737.9, 101722.9, 101706.4, 101682, 101645.2, 101606.9, 101566.6,
  101575.6, 101611.6, 101639.9, 101666.2, 101684.5, 101698.8, 101699.3, 
    101690.4, 101679.9, 101662.8, 101643.1, 101609.8, 101581, 101549.6, 
    101528.8,
  101529.7, 101561.2, 101583.6, 101610.9, 101623.8, 101633, 101632.2, 
    101623.5, 101614, 101593, 101570.8, 101543.5, 101525.6, 101502.1, 101488.5,
  101477, 101506.2, 101529.6, 101546.4, 101556.4, 101559.9, 101558.9, 
    101549.4, 101536.1, 101517.7, 101496.4, 101479.1, 101458.1, 101444.6, 
    101457.6,
  101425.8, 101449.8, 101465.5, 101477.9, 101482.7, 101485.6, 101482.1, 
    101474.6, 101464, 101451.2, 101428.9, 101408.8, 101393.9, 101397.8, 
    101412.9,
  101372.5, 101392.3, 101402.6, 101413.7, 101417.8, 101417.3, 101412.1, 
    101403.4, 101391.7, 101373.4, 101354.5, 101343.6, 101349.6, 101359.4, 
    101397.9,
  100893.1, 100923, 101043.1, 101129.8, 101232.2, 101346.2, 101421.8, 
    101470.7, 101522.6, 101563.8, 101597.6, 101623.9, 101655.7, 101678.9, 
    101697,
  100874.9, 100909.3, 100994.2, 101073.7, 101171.6, 101260.7, 101320.2, 
    101377, 101427.5, 101468.3, 101500.7, 101528.8, 101558.3, 101577.2, 
    101591.9,
  100918.3, 100947.2, 101004.7, 101051.6, 101112.9, 101174.7, 101247, 
    101312.5, 101364.3, 101395.4, 101431.6, 101461.8, 101487.5, 101506.8, 
    101519.9,
  100957.5, 100973.2, 101008.2, 101043.7, 101086.8, 101135.4, 101193.7, 
    101240, 101285.9, 101329.6, 101361, 101390.7, 101411.5, 101429.7, 101441.4,
  100974.4, 100996.9, 101025.5, 101049.7, 101075.4, 101100.5, 101135.7, 
    101181.2, 101221.1, 101259.2, 101291.4, 101318.3, 101339.7, 101356.2, 
    101362.6,
  100979.4, 101004, 101030.4, 101045.8, 101063.2, 101079.7, 101103.4, 
    101132.3, 101162.5, 101193.7, 101220.9, 101242.1, 101259.6, 101278.3, 
    101293,
  100973.6, 100995.7, 101019.8, 101039.5, 101050.3, 101058.6, 101070.5, 
    101092.6, 101111.7, 101133.2, 101150.6, 101175.9, 101192.8, 101214.7, 
    101220,
  100962.2, 100985.8, 101005.8, 101017.6, 101020.6, 101028.8, 101035.6, 
    101046.3, 101058.4, 101074.2, 101093.7, 101118.9, 101136.8, 101159.4, 
    101178.8,
  100957.5, 100975.1, 100988.4, 100995.3, 100997, 100996.6, 100999, 101003.6, 
    101009.2, 101016.4, 101028.9, 101055.3, 101076.8, 101112, 101136.1,
  100950.1, 100965.7, 100971.5, 100971.8, 100966, 100961.5, 100955.6, 
    100955.7, 100959.9, 100966.7, 100984.4, 101015.5, 101043.1, 101090.1, 
    101128.2,
  100500.1, 100417.7, 100354.4, 100312.3, 100299.9, 100297, 100306.6, 
    100314.7, 100337.1, 100353.2, 100377, 100408.7, 100455.2, 100504.8, 
    100559.1,
  100559, 100484, 100422.8, 100383.1, 100362, 100350.4, 100354.7, 100350.4, 
    100357.3, 100372.5, 100393.5, 100416.8, 100447.7, 100487.2, 100530.3,
  100615, 100553.4, 100499, 100455.1, 100422.4, 100397.3, 100404.9, 100402.4, 
    100401.3, 100400.8, 100413.1, 100439, 100472.8, 100503.6, 100521.7,
  100671.8, 100611.5, 100565.9, 100520.6, 100487, 100466.4, 100457.7, 
    100442.7, 100436.9, 100440, 100450.4, 100472.7, 100498.7, 100523.4, 
    100538.7,
  100707.2, 100663, 100626.3, 100585.6, 100549, 100524.8, 100499.3, 100496.7, 
    100502.1, 100501.2, 100507.2, 100505.8, 100509.9, 100521.4, 100538.8,
  100725.3, 100702, 100671.4, 100640.3, 100605.1, 100577.8, 100560, 100543.4, 
    100528.4, 100525.6, 100528.8, 100547.7, 100562.4, 100581.6, 100603.6,
  100735.3, 100713.9, 100686.6, 100670.2, 100646.3, 100621, 100601.8, 
    100585.4, 100581.2, 100571.5, 100570.4, 100577, 100596.7, 100618, 100656.2,
  100761.1, 100733, 100719.2, 100692.3, 100667.9, 100647.9, 100631.4, 
    100620.9, 100612.8, 100609.2, 100616.7, 100630.5, 100656, 100685.6, 100728,
  100716.5, 100705.2, 100711.3, 100694.7, 100681.4, 100665, 100657.7, 
    100650.7, 100648, 100645.2, 100652, 100672.5, 100697.7, 100730.4, 100775.2,
  100734.2, 100718.8, 100713.3, 100693.1, 100682, 100664.3, 100661.3, 
    100649.3, 100652.5, 100661, 100679.3, 100704.4, 100738.6, 100776.4, 
    100820.7,
  101054.1, 101051.1, 101053.5, 101057.6, 101058.4, 101055.4, 101052, 
    101050.8, 101048.4, 101042.3, 101024.8, 101002.4, 100972.6, 100936.6, 
    100898.5,
  101069.7, 101065.7, 101065.4, 101065, 101069.4, 101070.2, 101070, 101068.1, 
    101064.9, 101058.5, 101052.5, 101035.5, 101013.1, 100978.8, 100950.8,
  101091, 101086.1, 101091.9, 101089.5, 101090.6, 101091, 101089.2, 101090.3, 
    101087.7, 101085.1, 101079.3, 101069.5, 101053.4, 101027.5, 101000.6,
  101120.6, 101121.2, 101125.4, 101118.9, 101115.5, 101115.2, 101111.5, 
    101110.2, 101110.6, 101107.4, 101099.1, 101092.2, 101080.4, 101060.7, 
    101044.1,
  101130.9, 101130.1, 101133.7, 101129.2, 101126.1, 101126.7, 101123.7, 
    101123.7, 101119.8, 101120, 101115.3, 101111.8, 101100.7, 101086.6, 
    101074.4,
  101129.3, 101130.4, 101128.8, 101125.3, 101126.1, 101125.2, 101126.2, 
    101122.9, 101121.7, 101116, 101108.6, 101106.7, 101101.2, 101096.2, 
    101087.9,
  101104.8, 101107.7, 101114.9, 101110.7, 101104.6, 101109.6, 101104.9, 
    101101.3, 101103, 101096.2, 101090.9, 101086.4, 101082.3, 101083, 101084.5,
  101085.8, 101088.6, 101088.1, 101084.2, 101078.3, 101077.4, 101073.3, 
    101072.8, 101068.5, 101061.7, 101058.4, 101058.6, 101063.7, 101066.2, 
    101074.2,
  101042.1, 101044.6, 101044.2, 101038.8, 101032.5, 101031.7, 101026.9, 
    101025.7, 101019, 101019.6, 101021.1, 101020.9, 101025.6, 101035.4, 
    101049.2,
  100996.7, 101003, 101002.7, 100996.2, 100994.4, 100987.3, 100978, 100975.7, 
    100978.8, 100974.2, 100979.8, 100982.2, 100997, 101019.3, 101043.7,
  101417.2, 101461.3, 101503.1, 101539.2, 101578.3, 101614.9, 101652.7, 
    101690, 101732.2, 101774.6, 101816.9, 101859, 101911.1, 101962.7, 102008.3,
  101420.3, 101463.2, 101507.1, 101546.2, 101581.9, 101621.1, 101657.9, 
    101699, 101737.4, 101779.7, 101823.1, 101870, 101923.9, 101968.2, 102015.1,
  101414.2, 101463.6, 101509.5, 101547.4, 101586.2, 101620.8, 101654.3, 
    101694.3, 101733.4, 101776.8, 101814, 101858.9, 101897.9, 101943.5, 
    101980.5,
  101393.6, 101441.2, 101492.6, 101535.2, 101572.7, 101606.6, 101637.6, 
    101675.1, 101710, 101751.7, 101785.1, 101827.5, 101858.9, 101902.4, 
    101937.4,
  101363.6, 101409.2, 101451.9, 101495.1, 101540.2, 101572.9, 101603.1, 
    101629.6, 101658, 101688.8, 101721.7, 101755.1, 101791.9, 101828.1, 101868,
  101336.2, 101377.5, 101415.3, 101448.6, 101482.9, 101515, 101541.5, 
    101565.2, 101591.5, 101617.3, 101644.4, 101673.3, 101701.4, 101728.9, 
    101764.5,
  101296.9, 101331.9, 101370.4, 101400.9, 101429.8, 101454.6, 101475.3, 
    101494.2, 101516.2, 101533.5, 101553.9, 101573.8, 101599.7, 101626.3, 
    101660.7,
  101265.4, 101293.3, 101321.2, 101346.8, 101372.6, 101391.6, 101411, 
    101423.2, 101440.7, 101455.2, 101471.6, 101488.9, 101510.7, 101534.5, 
    101568.8,
  101222.8, 101249.1, 101270.1, 101288.7, 101305.1, 101318.9, 101333.3, 
    101346.9, 101359.2, 101369.9, 101383.6, 101406.2, 101431.4, 101465.9, 
    101500.8,
  101179.9, 101199.5, 101215.1, 101228.8, 101237.8, 101247.9, 101258.1, 
    101267.4, 101278.7, 101294.6, 101316.5, 101340.4, 101367.3, 101399.9, 
    101437.6,
  101258.9, 101267.5, 101300.3, 101330.1, 101367.3, 101409.9, 101456.4, 
    101508.9, 101558, 101602.5, 101651.9, 101704.8, 101769.7, 101838.4, 
    101913.3,
  101261.5, 101289.6, 101328.9, 101363.6, 101401.1, 101436.5, 101471.9, 
    101504.9, 101538.3, 101587.8, 101638.5, 101691.7, 101755.1, 101820.7, 
    101888.7,
  101274.3, 101302.5, 101343.3, 101369.7, 101405.7, 101435, 101468.3, 
    101500.6, 101534.6, 101577.7, 101622.5, 101671.6, 101730.7, 101793.4, 
    101863.7,
  101281.4, 101304.3, 101345.4, 101370.5, 101405.8, 101429, 101456.1, 
    101482.1, 101509.6, 101552.6, 101598.8, 101647.9, 101703.5, 101764.2, 
    101828.6,
  101281.2, 101301.1, 101338.2, 101362.4, 101388.1, 101410.9, 101432, 
    101455.4, 101482.4, 101521.9, 101565.4, 101613.3, 101665.5, 101722.8, 
    101786.1,
  101270.1, 101289.4, 101322.4, 101343.8, 101364.5, 101383.8, 101397.9, 
    101416.2, 101448.9, 101487.6, 101531.2, 101581.1, 101632.7, 101684.6, 
    101742.9,
  101255.8, 101273.8, 101300.1, 101313.4, 101324.2, 101337, 101355.3, 
    101381.2, 101411, 101452.1, 101494.1, 101544.4, 101593.1, 101643.7, 
    101699.5,
  101236.1, 101250.7, 101268.7, 101280.1, 101288.4, 101295.6, 101312.4, 
    101337.1, 101370.2, 101409, 101455.8, 101502.6, 101553.3, 101607.2, 
    101656.4,
  101212.7, 101224.3, 101233.9, 101239, 101245.2, 101252, 101267.2, 101291.4, 
    101325.5, 101366.9, 101409.8, 101459.3, 101506.7, 101555.7, 101607.3,
  101186.5, 101191.2, 101195.2, 101195.1, 101193.6, 101199.5, 101214.2, 
    101238.3, 101272.5, 101316, 101358.3, 101402.5, 101450, 101497.6, 101543.3,
  101428.9, 101394.6, 101365.8, 101320.5, 101286.8, 101256.5, 101237.1, 
    101223.5, 101229.6, 101258.8, 101308.3, 101357.5, 101413.8, 101479.2, 
    101551.9,
  101408.2, 101376, 101343.2, 101310.6, 101287.7, 101263.8, 101259.9, 101274, 
    101297.3, 101331, 101369, 101416.2, 101473.5, 101538.2, 101599.6,
  101388, 101365.3, 101341, 101321.7, 101307, 101292.4, 101292.2, 101303.1, 
    101324.4, 101362.9, 101408.8, 101457.8, 101509.5, 101567.3, 101626.6,
  101372.9, 101352.4, 101344.1, 101317, 101312.8, 101310.2, 101316.5, 
    101331.7, 101363.1, 101400.8, 101439.9, 101482.3, 101532.1, 101587.2, 
    101642.8,
  101346.4, 101340.1, 101337.2, 101331.8, 101341.6, 101337.9, 101341.6, 
    101339.9, 101375.4, 101407.3, 101450.7, 101493.2, 101539.8, 101584.9, 
    101637,
  101334.5, 101336.4, 101342.9, 101349.5, 101345.8, 101333.2, 101347.8, 
    101353.9, 101388.7, 101417.4, 101457.2, 101492.5, 101536.2, 101578.8, 
    101621.8,
  101344.3, 101329.8, 101338.2, 101324.3, 101315.6, 101314.3, 101332.6, 
    101355.5, 101382.2, 101410.8, 101443.1, 101479.1, 101512.8, 101551.7, 
    101594.8,
  101327.7, 101308, 101315.8, 101302.4, 101299.2, 101310.9, 101324.2, 
    101341.7, 101366.1, 101393, 101419.2, 101450.8, 101485, 101517.8, 101552.1,
  101293.4, 101288.1, 101279.5, 101274, 101276.8, 101286.8, 101296.6, 
    101317.7, 101335.5, 101361.4, 101385.7, 101409.4, 101434.2, 101466.7, 
    101498.3,
  101264.3, 101255.2, 101249.3, 101247.4, 101245.3, 101253.5, 101262.4, 
    101278.4, 101292.6, 101312.9, 101334.6, 101357.4, 101380.8, 101404.6, 
    101432,
  101221.1, 101193.2, 101178.4, 101160.8, 101140.6, 101121.7, 101103.5, 
    101088.2, 101065.6, 101047, 101039.1, 101037.6, 101048.4, 101070.7, 
    101113.2,
  101237.9, 101217.2, 101205.9, 101189.3, 101169.7, 101152.2, 101136.7, 
    101117.9, 101097.3, 101091.3, 101095.1, 101102.3, 101118.1, 101150.2, 
    101190.4,
  101256.1, 101236.6, 101229.8, 101214, 101200.6, 101182.4, 101167.6, 
    101153.1, 101147, 101143.1, 101145.4, 101155, 101176, 101203.6, 101243,
  101265.6, 101256, 101254.3, 101239.5, 101224.7, 101210.4, 101197.5, 
    101186.4, 101178.6, 101177, 101184.1, 101198.4, 101218.9, 101249, 101294.5,
  101262.9, 101258.6, 101259.6, 101247.4, 101236.3, 101226.2, 101220.4, 
    101210.3, 101206, 101211.2, 101217.7, 101227, 101255.2, 101287.3, 101325.1,
  101250.9, 101254.1, 101252.7, 101252, 101245.2, 101234.6, 101226.1, 
    101219.4, 101218.3, 101221.7, 101224.1, 101251, 101276.6, 101306, 101340.3,
  101250.7, 101248.3, 101247.7, 101236.2, 101231.7, 101227.7, 101226.3, 
    101220.8, 101218.4, 101224, 101239, 101269.3, 101287.1, 101311, 101338.3,
  101223.4, 101226.9, 101230.3, 101221.6, 101224.2, 101223.8, 101208, 
    101212.3, 101214, 101229.9, 101243.4, 101255.4, 101274.5, 101296.1, 
    101317.3,
  101208.2, 101206.3, 101212.2, 101205.8, 101204.8, 101203, 101204, 101204.4, 
    101213, 101222.6, 101229.7, 101235.9, 101247.8, 101265.8, 101281.1,
  101178.2, 101180.8, 101190.3, 101183.8, 101183.7, 101180.7, 101186.6, 
    101191.8, 101198.3, 101194.7, 101198.1, 101199.9, 101205.7, 101215.3, 
    101230.5,
  101228.9, 101218.4, 101203.4, 101192.5, 101177.8, 101165.4, 101153.9, 
    101143.7, 101135.3, 101131.3, 101132.7, 101140.9, 101153.1, 101168.7, 
    101181.5,
  101248.9, 101238.3, 101234.3, 101232, 101224.2, 101215.5, 101207.6, 
    101203.5, 101199, 101199.7, 101205.9, 101215.5, 101224.2, 101232.5, 
    101249.3,
  101251.3, 101251.7, 101253.9, 101252.8, 101256.6, 101255.3, 101256.8, 
    101254.8, 101258.6, 101261.9, 101267.6, 101271.4, 101274.4, 101283.5, 
    101294.4,
  101244.5, 101249.3, 101262.9, 101270.3, 101274.9, 101280.7, 101285.4, 
    101288.9, 101294.5, 101295.3, 101299.7, 101297.8, 101299.4, 101307.6, 
    101329,
  101240.7, 101250.3, 101265.9, 101272.6, 101286.3, 101294.5, 101301.3, 
    101307, 101309.7, 101310.5, 101310.5, 101307.2, 101313.6, 101335.8, 
    101358.9,
  101231.7, 101244.7, 101262.6, 101270, 101285.7, 101295.2, 101302.1, 
    101305.5, 101303.3, 101310.6, 101315, 101304.1, 101330.5, 101343.9, 
    101361.4,
  101218.6, 101235.2, 101253.6, 101264.1, 101279.8, 101285.7, 101299.7, 
    101293.4, 101298.7, 101291.6, 101291.6, 101307.8, 101324.3, 101326, 
    101340.8,
  101205.2, 101224.5, 101244.7, 101259.2, 101270.4, 101281.3, 101287.7, 
    101282.4, 101274, 101279.7, 101278.6, 101280.3, 101288.4, 101295.1, 
    101291.6,
  101189.8, 101212.3, 101235.6, 101248.5, 101257.7, 101270.5, 101277.3, 
    101272.9, 101269.8, 101261.7, 101250.4, 101249.1, 101240, 101231.1, 
    101224.3,
  101173.5, 101201.2, 101225.2, 101242.2, 101253.8, 101257, 101256.5, 
    101252.2, 101247.3, 101232.4, 101216.9, 101197.9, 101174.2, 101154, 
    101133.5,
  102035.7, 102063.2, 102065.6, 102072.6, 102071.8, 102070.3, 102065.6, 
    102058.7, 102043.3, 102034.8, 102027.1, 102017.6, 102001.2, 101983.7, 
    101967.2,
  101975.4, 101999.3, 102004.7, 102015.5, 102013.6, 102014.5, 102003.9, 
    101995.5, 101989.8, 101980.3, 101963.2, 101948.6, 101940.4, 101930.5, 
    101927.1,
  101904.1, 101923.2, 101930.8, 101935.2, 101937.3, 101932.5, 101927.9, 
    101912.4, 101904.6, 101889.6, 101883.2, 101879.1, 101872, 101864.3, 
    101858.6,
  101831.9, 101846.1, 101854.8, 101859.5, 101859.2, 101852.1, 101842.7, 
    101833.1, 101826.7, 101818.5, 101806.9, 101794.5, 101784.5, 101786.1, 
    101786.3,
  101750.5, 101772.3, 101777.4, 101775.7, 101778.5, 101772.3, 101766.2, 
    101754.1, 101742, 101723.1, 101707.5, 101697.6, 101686.1, 101678.8, 
    101674.9,
  101685.6, 101694.8, 101697.4, 101701, 101701.3, 101696.2, 101686.9, 
    101674.9, 101657.7, 101639.8, 101620.5, 101598.1, 101580.9, 101570.4, 
    101563.9,
  101637.8, 101635.2, 101636.1, 101634.5, 101637.4, 101629.2, 101621.9, 
    101602.2, 101580.7, 101556.2, 101529.9, 101490.3, 101459.1, 101436, 
    101423.8,
  101599.8, 101597.6, 101592.7, 101589.2, 101585.8, 101576.6, 101566.2, 
    101538.1, 101510.5, 101471.6, 101420.7, 101367.9, 101317.8, 101279.6, 
    101258.7,
  101575, 101573.7, 101560, 101555, 101542.8, 101533, 101513.3, 101479.1, 
    101437, 101379.2, 101307.1, 101230, 101154.9, 101095, 101052.2,
  101552.8, 101550.3, 101537.2, 101527, 101509, 101493.1, 101463.4, 101424.6, 
    101365.6, 101290.1, 101195.2, 101086.6, 100979.5, 100886.1, 100826.8,
  101749.7, 101788.4, 101806.9, 101833.6, 101852, 101868.8, 101880.4, 
    101895.6, 101914.9, 101940, 101965.5, 101995, 102026.8, 102064, 102103.3,
  101700, 101729.1, 101743.2, 101758.1, 101767.2, 101776.8, 101785.2, 
    101795.3, 101803.9, 101818.1, 101834.1, 101859.3, 101889.1, 101926.1, 
    101964.4,
  101629.3, 101659.9, 101668.7, 101679.1, 101680.2, 101681.1, 101677.4, 
    101674.9, 101674.8, 101680.5, 101696.4, 101719.3, 101749, 101783.5, 101823,
  101565.3, 101592.4, 101599.2, 101597.1, 101587, 101575.3, 101561.9, 
    101549.2, 101540.9, 101542.1, 101551.2, 101571.5, 101604.4, 101640.2, 
    101677.4,
  101507.9, 101526.9, 101525.2, 101512.5, 101496, 101475.1, 101448.3, 
    101422.5, 101406.1, 101397.6, 101403.3, 101419.9, 101444.9, 101476.6, 
    101509.2,
  101448.8, 101464, 101457, 101436.4, 101407.9, 101374.1, 101336, 101295.7, 
    101262.8, 101241.3, 101238, 101248.3, 101271.6, 101307.5, 101350.9,
  101391.6, 101400.7, 101390.4, 101364.8, 101327.6, 101285.1, 101230.6, 
    101172.9, 101119.9, 101081.4, 101062.2, 101064.2, 101089.9, 101138.1, 
    101205.7,
  101349.5, 101349.9, 101337.5, 101303.6, 101257.9, 101201.5, 101131.5, 
    101051.2, 100969.9, 100904.3, 100869.4, 100864.2, 100898.3, 100966.5, 
    101059.5,
  101313.6, 101308.2, 101293.4, 101251.8, 101198.5, 101129.7, 101046.4, 
    100941.7, 100830.6, 100732.8, 100665.4, 100647.9, 100683.5, 100761.4, 
    100874.7,
  101282.6, 101271, 101256.3, 101211.6, 101151.6, 101073, 100975.9, 100850.7, 
    100709.5, 100568.1, 100452.4, 100396.5, 100413.1, 100511.7, 100654.6,
  101749.7, 101716.3, 101690.5, 101661.8, 101626.5, 101583.1, 101530.4, 
    101491, 101446.9, 101422, 101394, 101365.9, 101351.3, 101366.7, 101407.2,
  101673.9, 101639.4, 101600.8, 101560.5, 101518.8, 101472.9, 101425.6, 
    101379.1, 101341.2, 101317.6, 101299.2, 101309.2, 101320.5, 101333, 
    101339.4,
  101590.2, 101547.6, 101498.7, 101454.5, 101402.4, 101349.7, 101308.6, 
    101255.9, 101237.8, 101222, 101228.7, 101238.2, 101242.5, 101270.6, 
    101309.3,
  101508.1, 101468, 101407.1, 101351.3, 101290.5, 101234.8, 101174.4, 
    101135.8, 101112.8, 101098, 101112.9, 101125.4, 101144.3, 101181.6, 
    101236.2,
  101438.5, 101393.8, 101318.2, 101251, 101179.6, 101116.8, 101042.3, 
    101008.5, 100955.3, 100945.7, 100958.5, 100997.9, 101061.8, 101127.3, 
    101213.5,
  101374.1, 101324.2, 101238.5, 101162.1, 101081.1, 101003.3, 100919.8, 
    100855.6, 100779.7, 100773.7, 100787.1, 100861.3, 100952.4, 101039.7, 
    101150.3,
  101314.9, 101258.4, 101168.1, 101085.3, 100995.7, 100906.8, 100806.2, 
    100705.1, 100621.7, 100594, 100602.8, 100697.4, 100834.8, 100959.4, 
    101092.8,
  101252.4, 101197.5, 101111.2, 101022.8, 100930.2, 100830.3, 100713.9, 
    100580.9, 100479.1, 100420.3, 100414.9, 100524.2, 100697.7, 100860.7, 
    101008,
  101202.7, 101152.6, 101071.1, 100980.5, 100885.8, 100778.1, 100650, 100498, 
    100367.6, 100273, 100233.5, 100353.7, 100547.7, 100751.1, 100920.9,
  101154.5, 101114.2, 101041.8, 100955, 100859.9, 100752, 100619.6, 100458.9, 
    100308.6, 100178.5, 100092.5, 100189.9, 100408.8, 100646.9, 100829,
  102239.8, 102235.6, 102218.2, 102204.2, 102186.1, 102166, 102144.7, 102123, 
    102097.8, 102085.6, 102056.1, 102026.9, 102015.6, 102002.7, 101967.6,
  102164, 102152.5, 102129.3, 102111.5, 102087.7, 102059.6, 102032.9, 
    101996.2, 101970.2, 101935, 101917.9, 101912.3, 101904, 101874.6, 101862.5,
  102079.8, 102063.7, 102034, 102009.4, 101975.9, 101940.3, 101894.6, 
    101852.7, 101811.9, 101794.7, 101769.7, 101732.4, 101712.5, 101727.1, 
    101745.2,
  101990.7, 101971, 101937.7, 101905.2, 101861.2, 101815.8, 101759.4, 
    101718.5, 101674.5, 101616.7, 101552.6, 101577.4, 101622.9, 101632.4, 
    101625.6,
  101907.3, 101887.7, 101846.6, 101804.7, 101746.4, 101689.8, 101626.2, 
    101560.4, 101473.4, 101416.6, 101429.6, 101418.8, 101390.9, 101392.7, 
    101444.6,
  101832.9, 101807.2, 101756.7, 101702, 101637.3, 101568.9, 101488.8, 101395, 
    101311.3, 101305.6, 101264.1, 101232.6, 101192.9, 101234.3, 101277.7,
  101754.7, 101723.5, 101666.8, 101608.4, 101536.3, 101455.5, 101355.7, 
    101254.7, 101163.2, 101110.6, 101039.8, 101001, 100994.6, 101075, 101183,
  101678.9, 101645.7, 101582.4, 101519.7, 101441.7, 101350.3, 101241.8, 
    101130.2, 101023, 100909.5, 100841.1, 100893.5, 100972.4, 101076.4, 
    101158.7,
  101607.5, 101564.7, 101504, 101438, 101357.4, 101259.4, 101149.4, 101030, 
    100884.2, 100750.4, 100757.2, 100855.7, 100950.2, 101069.5, 101177.2,
  101535, 101490.1, 101434.3, 101366.4, 101284.9, 101190.2, 101079.5, 
    100949.4, 100788.1, 100675.4, 100716.9, 100828.9, 100945.9, 101073.4, 
    101185.8,
  101924.7, 101934.3, 101940.5, 101947.5, 101955.2, 101966.8, 101981.3, 
    101992.3, 101999.3, 101998, 101992.8, 101991.4, 101997.9, 102034.7, 
    102093.3,
  101856.5, 101865.9, 101865.4, 101869.3, 101873.6, 101882, 101890, 101898.2, 
    101905.3, 101908.2, 101901.2, 101882.9, 101853.6, 101839.7, 101885.4,
  101798.8, 101794.9, 101785.2, 101774.3, 101768.5, 101767.2, 101771.8, 
    101778.6, 101782.8, 101776.8, 101759.6, 101730.6, 101675.7, 101668.8, 
    101763.9,
  101739.8, 101724.5, 101704.7, 101684.9, 101666.9, 101654.4, 101651.9, 
    101663.6, 101678.2, 101689.5, 101682.4, 101660.2, 101592.4, 101521.2, 
    101590.8,
  101683.5, 101658.6, 101629.4, 101592.9, 101558.2, 101528.1, 101522.9, 
    101536.4, 101556.2, 101577, 101583.2, 101569.8, 101515.9, 101457.4, 
    101543.7,
  101633.7, 101600.9, 101557.5, 101508.7, 101457.1, 101415.3, 101404.3, 
    101420.1, 101455, 101492.6, 101517.9, 101523.7, 101477, 101487.9, 101560.5,
  101591.6, 101551.5, 101494.4, 101438, 101370.7, 101315.6, 101290.9, 
    101306.9, 101348.7, 101395, 101436.6, 101469, 101505.2, 101568, 101622.1,
  101550.3, 101507.4, 101440.4, 101377.6, 101301.6, 101236.1, 101198.9, 
    101212.4, 101254.6, 101313.6, 101379.5, 101454.4, 101508.9, 101567.6, 
    101631,
  101517, 101471.8, 101398.7, 101337, 101257.8, 101182.6, 101132.3, 101141.8, 
    101187.4, 101268.4, 101351.6, 101435.5, 101506.3, 101584.6, 101654.4,
  101486.9, 101440.8, 101367, 101303.3, 101230.9, 101151.1, 101092.8, 
    101098.5, 101146.9, 101235.6, 101324.9, 101413, 101492.4, 101571.5, 101646,
  101641.8, 101620.9, 101603.6, 101583.8, 101553.4, 101545.1, 101533.7, 
    101534, 101527.6, 101526.9, 101534.4, 101550, 101549.3, 101526.5, 101505.7,
  101619.5, 101599.9, 101571, 101550, 101525.6, 101484.6, 101444.9, 101414.2, 
    101397.5, 101407.8, 101433, 101458.6, 101469.5, 101461.1, 101479.8,
  101596.6, 101569.5, 101541.4, 101504.9, 101461, 101391.4, 101368.9, 
    101371.4, 101390.9, 101419.9, 101461.5, 101501.5, 101533.1, 101558.6, 
    101591.1,
  101577, 101544.5, 101518.3, 101477.5, 101404.1, 101346.3, 101339.9, 
    101345.4, 101381.3, 101423.1, 101468.7, 101513.9, 101553.9, 101590.7, 
    101631.8,
  101556, 101525.4, 101493.3, 101455, 101388.2, 101346.5, 101339.8, 101365.9, 
    101426.1, 101476.4, 101529.6, 101580.6, 101628.3, 101677.9, 101727.6,
  101545.9, 101507.7, 101477.9, 101443.3, 101377.4, 101346.8, 101349.4, 
    101397.4, 101458.3, 101512.6, 101571.4, 101626.5, 101676.1, 101727.4, 
    101776.5,
  101532.6, 101498.3, 101461.7, 101432.2, 101373.1, 101355.3, 101366.8, 
    101418.7, 101478.3, 101542.7, 101607, 101670.2, 101725.1, 101781, 101835.9,
  101520.4, 101486.2, 101448.2, 101418.7, 101373.1, 101352.4, 101373.4, 
    101427.3, 101486.3, 101552.4, 101619.2, 101687, 101746.2, 101807, 101861.2,
  101506.2, 101480.3, 101440.5, 101406.3, 101366.8, 101351.8, 101376.2, 
    101424.3, 101486, 101549.5, 101621.2, 101692.9, 101756.3, 101819.5, 
    101877.2,
  101485, 101467.9, 101426.4, 101395.8, 101357.1, 101347.6, 101364, 101412.4, 
    101472.4, 101535.5, 101607.4, 101681, 101746.1, 101812, 101871.7,
  101758.7, 101763.4, 101751.2, 101749.5, 101733.2, 101722.4, 101709.9, 
    101689.5, 101662.9, 101633.7, 101596.7, 101553.7, 101507.2, 101459.2, 
    101412.2,
  101768.9, 101770.7, 101759.4, 101759.3, 101748.3, 101734.2, 101723.3, 
    101696, 101662.6, 101635.4, 101598, 101564.6, 101524.7, 101482.5, 101441.8,
  101754.5, 101756, 101747.6, 101746.2, 101736.4, 101724.7, 101704.3, 101685, 
    101658.9, 101632.8, 101596.3, 101566.1, 101534.1, 101507.4, 101488.9,
  101733.3, 101732.3, 101731.6, 101724.1, 101711.6, 101702.3, 101680.2, 
    101655.2, 101629, 101600.8, 101577.6, 101563.5, 101547.6, 101535.8, 
    101523.4,
  101708.6, 101699.6, 101695.9, 101687.1, 101672.9, 101661.1, 101642.6, 
    101620.3, 101606.1, 101599.4, 101592.8, 101591.6, 101586.2, 101581.1, 
    101579.1,
  101674.4, 101662.1, 101659.5, 101645.4, 101631.8, 101622.1, 101607.9, 
    101596.3, 101580.7, 101572.5, 101578.9, 101590.7, 101600.4, 101612.7, 
    101622.2,
  101648.7, 101634.4, 101621.1, 101609, 101589.9, 101591.7, 101579.9, 
    101556.7, 101562.7, 101581.7, 101613.1, 101641.9, 101672, 101694.4, 
    101715.8,
  101615.4, 101601.9, 101583.7, 101566.3, 101554.4, 101549, 101527.1, 
    101546.7, 101576.1, 101604.2, 101640.5, 101673.9, 101708.2, 101740.3, 
    101770.4,
  101577.4, 101566.9, 101542.1, 101528.8, 101507.6, 101494.2, 101495.5, 
    101541, 101575.2, 101614.7, 101656.5, 101702.7, 101744.1, 101782.3, 
    101815.2,
  101544.3, 101534.9, 101508.3, 101485, 101464.5, 101451.8, 101484.9, 
    101533.2, 101568.2, 101615.2, 101661, 101705.9, 101748.9, 101790.2, 
    101832.9,
  101029.5, 101053.9, 101082.4, 101107.8, 101131.6, 101154.7, 101186.7, 
    101218.6, 101254.4, 101293.7, 101336.2, 101376.9, 101418.2, 101458.6, 
    101499.2,
  101049.6, 101077.2, 101100.7, 101123.6, 101144.6, 101171.6, 101207.6, 
    101242.9, 101280.6, 101323.4, 101363.9, 101404.5, 101445.9, 101486.7, 
    101520.2,
  101060.9, 101085, 101107.2, 101124.3, 101146.8, 101178.6, 101214, 101250, 
    101292.2, 101335.9, 101380.2, 101424.9, 101468.6, 101509.5, 101551.1,
  101062.2, 101087.6, 101111.2, 101116.7, 101138.8, 101175.4, 101215.6, 
    101255.2, 101298.9, 101341, 101383, 101425.2, 101466.2, 101505.4, 101540.5,
  101058.8, 101083.2, 101102, 101107.4, 101134.7, 101171.2, 101212.8, 
    101257.6, 101306.1, 101348.7, 101392.9, 101434.2, 101476.2, 101515.1, 
    101549.8,
  101057.4, 101075.2, 101088.3, 101092.5, 101130.4, 101170.9, 101217.9, 
    101264.4, 101311.2, 101356.6, 101405.4, 101449.6, 101493.5, 101529.8, 
    101567.2,
  101053.1, 101067.2, 101077.6, 101090.3, 101130.6, 101174.9, 101225, 
    101275.2, 101327.9, 101377.6, 101429.8, 101480.8, 101531.1, 101577.9, 
    101622.2,
  101048.5, 101058.8, 101069, 101086.8, 101130.5, 101177.1, 101229.7, 
    101286.1, 101339.1, 101391.7, 101448.1, 101503.5, 101553.7, 101600.8, 
    101643.4,
  101040.2, 101049.9, 101060.7, 101092.5, 101131.5, 101182.3, 101236.5, 
    101289.4, 101343.4, 101401.1, 101456, 101515.3, 101567.2, 101619.8, 
    101667.3,
  101036.4, 101042.5, 101057.9, 101084.2, 101127.7, 101173.2, 101227.8, 
    101283.4, 101339, 101394, 101453.2, 101509.8, 101563.1, 101613.9, 101661.9,
  101275.7, 101158.6, 101055.2, 100952.2, 100847.3, 100739.6, 100629.1, 
    100527.1, 100434.9, 100366.5, 100318.8, 100294.1, 100293.7, 100300.4, 
    100310.1,
  101267, 101162.8, 101082.9, 100993.3, 100896.2, 100793, 100695.1, 100599.1, 
    100524, 100472.9, 100438.7, 100425.4, 100424.7, 100431.6, 100458.7,
  101304.5, 101221.7, 101135.1, 101044.1, 100950.5, 100859.3, 100773, 
    100699.1, 100637.2, 100589.9, 100560.3, 100546.2, 100543.7, 100552, 
    100580.8,
  101316.4, 101232.6, 101158.9, 101079.7, 101002.3, 100921.3, 100845, 
    100777.2, 100724.5, 100687.5, 100665, 100654.4, 100656.1, 100666.1, 100695,
  101326.3, 101253, 101186.1, 101110.8, 101036.7, 100967.2, 100905.6, 
    100850.3, 100809.4, 100775.8, 100756.4, 100747.5, 100745.4, 100759, 
    100786.5,
  101314, 101250, 101184.8, 101121.4, 101060, 101001.7, 100949.6, 100906.4, 
    100871.2, 100845.3, 100829.7, 100823.4, 100826.5, 100839.3, 100866.9,
  101299.4, 101243.5, 101184.6, 101126, 101070.2, 101023.5, 100981.9, 
    100947.2, 100916.6, 100897.6, 100886.5, 100883.5, 100885.5, 100903, 
    100932.2,
  101271.4, 101218.6, 101166.8, 101116.8, 101071.1, 101034.2, 100998.7, 
    100971.9, 100950.2, 100936.5, 100926.4, 100925.6, 100939.6, 100958.4, 
    100983.4,
  101232.1, 101193, 101148.4, 101103.9, 101067, 101033.5, 101004.9, 100982.4, 
    100966.9, 100955.7, 100954.1, 100957.5, 100973.7, 100988.7, 101024.4,
  101193.9, 101158.2, 101122, 101086.1, 101053.4, 101025, 101000.4, 100983.4, 
    100969, 100962.5, 100964.8, 100977.1, 100996.3, 101014.5, 101057.4,
  102001.9, 102022.2, 102025, 102020.3, 102006.9, 101984.7, 101959.9, 
    101917.8, 101867, 101803.4, 101732.6, 101648.7, 101549.7, 101445.4, 
    101338.3,
  101981.7, 102000.4, 102005.9, 102002.9, 101988.9, 101970.2, 101942, 
    101904.1, 101853.4, 101793.4, 101725.7, 101647.8, 101554.9, 101454.8, 
    101350.4,
  101957.6, 101972.9, 101981.7, 101975.9, 101969.9, 101950.4, 101926.8, 
    101889.1, 101842.6, 101786.4, 101722.7, 101652.3, 101570.2, 101481.6, 
    101385.7,
  101930, 101944.8, 101955.5, 101953.6, 101942.1, 101922.2, 101893.5, 
    101859.7, 101815.4, 101762, 101702.3, 101636.5, 101562.8, 101485.7, 
    101392.8,
  101908.2, 101918.4, 101919.8, 101920.9, 101911.2, 101892.5, 101869.1, 
    101833, 101789, 101740.2, 101685, 101622.8, 101557.1, 101483.7, 101399.4,
  101884.5, 101894.5, 101893, 101888.3, 101877.9, 101863.1, 101840.1, 
    101806.8, 101768.2, 101719.6, 101666, 101607.7, 101543, 101471.4, 101391.3,
  101852.2, 101860.2, 101860.3, 101855.7, 101847, 101828.3, 101807.8, 
    101779.4, 101741.9, 101697, 101645.3, 101588.5, 101525.9, 101453.3, 
    101379.2,
  101813.7, 101823.4, 101817.1, 101814.2, 101802.2, 101789.4, 101769.4, 
    101743.8, 101707.6, 101663.7, 101613.6, 101557.7, 101492.4, 101426.5, 
    101351.1,
  101776.4, 101783.4, 101778.9, 101772.6, 101760, 101745.8, 101723.1, 
    101696.4, 101660.6, 101619.1, 101572.1, 101520.9, 101460.7, 101394.3, 
    101320.8,
  101741.4, 101739.5, 101731.2, 101724, 101711.6, 101695.1, 101670, 101640.1, 
    101605.7, 101565.7, 101520.4, 101469.4, 101414.3, 101348.9, 101274.2,
  101658.8, 101768.5, 101868.5, 101963, 102053.3, 102132, 102208, 102285.6, 
    102358.8, 102412.6, 102461.5, 102499.1, 102526.3, 102550.1, 102568.4,
  101634.4, 101742.5, 101846.2, 101940, 102027.4, 102105.4, 102175.7, 
    102241.4, 102311.9, 102379.3, 102427.6, 102468.5, 102499, 102518.2, 
    102531.1,
  101614.9, 101715.6, 101817.5, 101907.3, 101998.2, 102075.5, 102147, 
    102210.6, 102268.7, 102330.6, 102386.7, 102426.1, 102459.2, 102482.3, 
    102497.7,
  101584.4, 101682.9, 101781.8, 101869.3, 101956.4, 102036.5, 102106.2, 
    102173.1, 102229, 102279.5, 102333.9, 102380.5, 102412, 102433.3, 102445.9,
  101558.6, 101649.7, 101742.2, 101829.6, 101907.5, 101988.1, 102059.6, 
    102125.4, 102181.2, 102233, 102274.4, 102314.3, 102353, 102380.7, 102399.3,
  101528.9, 101613.9, 101696.3, 101778.9, 101855.6, 101930.4, 101997.4, 
    102064.9, 102121.8, 102173.5, 102221.2, 102256.1, 102288, 102310, 102326.5,
  101504.1, 101581, 101656.8, 101727.4, 101797.9, 101867.3, 101931.8, 
    101990.6, 102048.9, 102098.6, 102147.1, 102189.4, 102224.5, 102251.8, 
    102271.8,
  101476.7, 101548, 101615.4, 101674, 101738.2, 101796, 101859.9, 101917.5, 
    101970.5, 102021.6, 102068.1, 102107.6, 102143.7, 102174.4, 102197.9,
  101447.6, 101508.8, 101569.8, 101621.2, 101675.8, 101729.2, 101783.5, 
    101838.6, 101893.3, 101941.9, 101988.4, 102026.5, 102064.7, 102094.6, 
    102115.2,
  101422.6, 101474.6, 101524.3, 101572.4, 101619.6, 101665.1, 101711.7, 
    101761.6, 101814, 101861.1, 101910.2, 101949.1, 101982.5, 102011.5, 
    102033.9,
  101363.5, 101458.7, 101551.5, 101652.9, 101754.9, 101856, 101950.2, 
    102042.5, 102136.1, 102226.6, 102310.7, 102393.5, 102480.6, 102568.7, 
    102649.4,
  101350.5, 101450.3, 101545.4, 101642.1, 101739.2, 101838.9, 101931.3, 
    102022.1, 102114.2, 102202.8, 102290.4, 102374.7, 102458.1, 102540.5, 
    102625.3,
  101343.4, 101438.6, 101532.8, 101626.5, 101721.1, 101819.8, 101913.6, 
    102003.6, 102092.9, 102179.9, 102267.2, 102348.8, 102427.7, 102511.4, 
    102590.2,
  101317.2, 101412.4, 101506.5, 101600.6, 101691.9, 101786.6, 101878.4, 
    101968, 102057.5, 102141.4, 102225.3, 102307.1, 102387.9, 102461, 102540.5,
  101296.8, 101388.8, 101478.9, 101570.6, 101660.4, 101752.9, 101842.2, 
    101932.4, 102017.2, 102101, 102179.8, 102255.1, 102330.8, 102406.4, 
    102481.1,
  101270.7, 101356.7, 101444.3, 101534.1, 101619.9, 101708.1, 101794.8, 
    101883.8, 101968.2, 102049.4, 102124, 102197.3, 102269.3, 102336.4, 
    102405.1,
  101251, 101329.4, 101413.6, 101495.6, 101580.3, 101666.7, 101749.1, 
    101832.1, 101913.6, 101990.3, 102065.2, 102135, 102202.6, 102271.5, 
    102330.8,
  101230.5, 101300, 101378.1, 101457.4, 101536.2, 101614.4, 101695.1, 
    101772.8, 101848.7, 101923.4, 101993.1, 102062.5, 102126.8, 102195.1, 
    102255.8,
  101213.5, 101273.3, 101344, 101414.6, 101490.9, 101565.5, 101642.5, 
    101716.1, 101788.6, 101859.7, 101926, 101990.2, 102051.3, 102110, 102171.6,
  101194.1, 101243.7, 101302.2, 101364.3, 101438.8, 101508.3, 101581, 
    101653.2, 101717.8, 101785.1, 101848.6, 101908.9, 101971, 102028.1, 
    102082.2,
  101501.1, 101456.5, 101429.8, 101410.1, 101398.3, 101389.1, 101385.7, 
    101394.9, 101408.5, 101434, 101463.6, 101497.3, 101543.9, 101609.2, 
    101695.8,
  101481.8, 101456, 101445.2, 101433.2, 101428.2, 101430.7, 101440.3, 
    101450.1, 101463.6, 101484.3, 101514.1, 101555.6, 101611.6, 101683.1, 
    101764.5,
  101481.9, 101468.1, 101458.8, 101452.1, 101453.8, 101464.4, 101474.3, 
    101485.1, 101502.5, 101528.3, 101563.9, 101607, 101660.7, 101729.5, 
    101806.3,
  101465.6, 101461.7, 101462.9, 101464.2, 101471.5, 101482.3, 101497.7, 
    101516.3, 101533, 101561.1, 101603.1, 101648.3, 101701.2, 101767.2, 
    101844.7,
  101447.3, 101451.2, 101450.4, 101456.4, 101473.4, 101494.2, 101513.4, 
    101530.6, 101552.7, 101586, 101625.7, 101670.1, 101720.7, 101787.3, 
    101861.4,
  101416.1, 101420.9, 101433.5, 101452.4, 101475.7, 101497.7, 101514.2, 
    101540.1, 101563.6, 101592.2, 101629.3, 101676.3, 101729, 101794.7, 
    101866.2,
  101376.3, 101388.1, 101407.2, 101430.4, 101457.8, 101484.9, 101511.5, 
    101540.2, 101562, 101589.4, 101619, 101665.8, 101716.2, 101780.4, 101852,
  101337.9, 101342.2, 101367.6, 101403.6, 101437.3, 101471.3, 101494.4, 
    101527.3, 101543.1, 101569.1, 101594.1, 101641.4, 101691.9, 101757, 
    101826.3,
  101303.3, 101306.7, 101335, 101376.5, 101414.8, 101443.5, 101474.1, 
    101501.5, 101517.3, 101541.8, 101560.4, 101603.8, 101653.6, 101718, 
    101792.6,
  101266.6, 101274.8, 101300.3, 101342.2, 101379.3, 101409.7, 101438.4, 
    101467.2, 101481.2, 101501.3, 101517.6, 101559.5, 101609.5, 101672.6, 
    101743,
  102303.2, 102276.8, 102231.8, 102188.4, 102135.9, 102081.5, 102018.8, 
    101950.9, 101866.5, 101781.1, 101689.4, 101595.5, 101494.2, 101387.7, 
    101262.5,
  102271.7, 102234.4, 102193.8, 102153.4, 102106.4, 102054.9, 101989, 
    101918.4, 101839.9, 101758.9, 101667.5, 101575.5, 101458.3, 101341.5, 
    101234.4,
  102224.3, 102192.5, 102157.9, 102114.6, 102070, 102022, 101968, 101908.3, 
    101833, 101756.3, 101667.9, 101568.4, 101464.3, 101359, 101259.6,
  102169.6, 102141.7, 102106.1, 102066.4, 102023.3, 101977.6, 101922.7, 
    101863.8, 101798.9, 101723.8, 101644.9, 101552.1, 101455.2, 101349.8, 
    101257,
  102103, 102082.7, 102052.4, 102017.6, 101978.2, 101933.7, 101883.7, 
    101830.6, 101765.4, 101696, 101620.6, 101533.8, 101449.2, 101350.4, 
    101275.8,
  102031.3, 102011.6, 101976.3, 101945.5, 101910.9, 101875.6, 101828.8, 
    101775.1, 101717, 101648.4, 101582.6, 101504.7, 101423.1, 101342, 101278.7,
  101948.2, 101926.6, 101889.3, 101865.3, 101836.5, 101802.7, 101760.2, 
    101712.8, 101661.9, 101599.9, 101536.9, 101468.8, 101396.2, 101333.7, 
    101285.1,
  101863.7, 101844.6, 101804.8, 101779.9, 101748.1, 101713.4, 101680.8, 
    101642.2, 101596.3, 101539.1, 101481.8, 101420.2, 101367.9, 101324.5, 
    101287.5,
  101777.8, 101748.8, 101708.5, 101683.7, 101650.1, 101624.8, 101592.9, 
    101560.1, 101518, 101473.9, 101429.1, 101373.1, 101333.9, 101305.8, 101275,
  101672.3, 101645.3, 101608.7, 101583.3, 101555.4, 101533.5, 101503.4, 
    101477.5, 101444.2, 101408.8, 101362.9, 101327, 101303.9, 101276.1, 
    101275.4,
  102188.9, 102178.7, 102148.2, 102111.5, 102064.6, 102012.5, 101950.2, 
    101883.9, 101815.8, 101755.8, 101717.8, 101673.7, 101633.2, 101568.8, 
    101527.6,
  102164.5, 102154.8, 102132, 102103.1, 102064, 102016.4, 101960.3, 101892.8, 
    101823.2, 101751.4, 101699, 101649.9, 101606.2, 101548.7, 101490.8,
  102128, 102119.2, 102106.6, 102082.8, 102052.3, 102011.7, 101964.4, 
    101904.2, 101842.6, 101775.5, 101721.3, 101669.7, 101613.7, 101546.6, 
    101482.5,
  102085.4, 102077.5, 102071, 102050.6, 102030.5, 101999, 101957.5, 101900.8, 
    101835.4, 101768.9, 101711.9, 101660.7, 101608.9, 101551.4, 101488,
  102034, 102033, 102024.8, 102012.5, 101996.9, 101974.7, 101944.6, 101899.8, 
    101847.2, 101784.7, 101729.4, 101675.2, 101622.2, 101559, 101488.3,
  101984, 101983.8, 101976.7, 101968.2, 101955.2, 101938.4, 101914.7, 
    101879.3, 101836.8, 101785.1, 101728.2, 101677.2, 101624.2, 101561.1, 
    101494.1,
  101936.2, 101932.6, 101922.8, 101915.2, 101901.5, 101890.4, 101870.4, 
    101844.4, 101810, 101774.2, 101725.5, 101678.1, 101621.9, 101560.8, 101492,
  101877.3, 101873.5, 101862.4, 101852.3, 101840.8, 101829.7, 101811.1, 
    101792, 101760.4, 101731.3, 101692, 101650.3, 101602.3, 101543.2, 101477.2,
  101817.5, 101814.8, 101798.4, 101787.8, 101775.7, 101763.4, 101747, 101732, 
    101704.4, 101677.8, 101641.7, 101605.9, 101561.3, 101510.8, 101451,
  101762.3, 101752.8, 101731.9, 101722.9, 101704.9, 101690.8, 101672.2, 
    101654, 101629.9, 101606.4, 101579.6, 101548, 101509.9, 101460.4, 101412.2,
  101897, 101887.3, 101860, 101826.9, 101786, 101745.2, 101698.2, 101656.1, 
    101610.9, 101581.4, 101546.3, 101495.1, 101416.2, 101318.9, 101204.8,
  101882.1, 101869.1, 101850.6, 101821.6, 101786.3, 101748, 101705.2, 
    101665.6, 101620.6, 101578.6, 101540.4, 101500.9, 101446.5, 101363.9, 
    101276.8,
  101866.4, 101870.1, 101856.6, 101826.7, 101795.5, 101758, 101715.9, 
    101672.2, 101629, 101589.4, 101559.9, 101523.2, 101480.1, 101426.8, 
    101358.1,
  101837.8, 101851.7, 101847.5, 101824.7, 101797.4, 101763.9, 101727.1, 
    101685.4, 101644, 101600.3, 101560.6, 101531.3, 101500.7, 101462.2, 
    101417.3,
  101804.7, 101824.8, 101832.2, 101823.9, 101802.8, 101774.5, 101741.9, 
    101703.2, 101662.6, 101625.2, 101579.8, 101547.7, 101524.2, 101495.7, 
    101465,
  101765.1, 101793.6, 101805, 101805.8, 101794.1, 101776.1, 101751.5, 
    101716.5, 101682.6, 101644.9, 101602.8, 101568.4, 101540.3, 101519.1, 
    101494.8,
  101726.7, 101754.8, 101767.9, 101778.8, 101777.9, 101769.2, 101755.6, 
    101728.6, 101698.6, 101664.1, 101630.1, 101594.8, 101565.3, 101539.2, 
    101524.6,
  101680.6, 101711.6, 101727.1, 101741.7, 101747.1, 101750.7, 101746.4, 
    101732.1, 101711, 101680.4, 101651.2, 101619.1, 101591, 101562.6, 101546,
  101642.8, 101667.3, 101681.2, 101697.5, 101707.8, 101715.1, 101718.4, 
    101713.3, 101700.5, 101679.8, 101655.5, 101630.4, 101609.4, 101590, 
    101578.8,
  101602.8, 101620.6, 101631.2, 101644.7, 101653.9, 101664.1, 101670.4, 
    101673.1, 101670, 101658.9, 101645.9, 101634.2, 101615.6, 101602, 101586.2,
  101647.6, 101691.2, 101722.5, 101739.5, 101752.5, 101758.8, 101780.3, 
    101797, 101806.5, 101794.9, 101784.3, 101757.9, 101715.5, 101670.5, 
    101613.1,
  101603.5, 101645.9, 101688.8, 101707.2, 101730.4, 101740.1, 101757.3, 
    101771.3, 101781.9, 101777.4, 101762.4, 101735.3, 101703.8, 101663.3, 
    101615.4,
  101570, 101627.9, 101662.4, 101687.1, 101701.1, 101713.7, 101724.4, 
    101742.6, 101752.7, 101758.6, 101747, 101723.5, 101695.1, 101656.2, 101621,
  101534.1, 101593, 101635.1, 101658.5, 101683.5, 101696.2, 101703.5, 
    101714.9, 101724, 101730.9, 101729.1, 101712.3, 101686, 101658.2, 101620.6,
  101499.6, 101559.6, 101609, 101640.7, 101658.8, 101672.3, 101685.3, 
    101691.3, 101695.3, 101706.8, 101708.5, 101698.5, 101680, 101656.9, 
    101623.5,
  101461.8, 101529.1, 101578.5, 101614.8, 101638.2, 101655.4, 101667.7, 
    101676.5, 101687.5, 101690.5, 101691.5, 101682.3, 101667.6, 101650.5, 
    101617.8,
  101431.3, 101497.5, 101548.8, 101590, 101617.1, 101637, 101650.4, 101660.4, 
    101670.1, 101673.1, 101666.6, 101660.3, 101644.1, 101628.9, 101612.3,
  101402.6, 101465.3, 101513.9, 101558.5, 101590.1, 101614.1, 101628.6, 
    101638.4, 101649, 101649.1, 101644, 101635.8, 101627.1, 101612.1, 101594.8,
  101380, 101432.9, 101480.1, 101523.6, 101556.2, 101583.2, 101601.5, 
    101612.3, 101622.2, 101620.7, 101617.9, 101607.5, 101593.1, 101578.7, 
    101565,
  101356.2, 101398.8, 101440.5, 101479.1, 101512.2, 101540.5, 101559.1, 
    101572.4, 101580.2, 101583.2, 101580.3, 101575, 101572.8, 101556.5, 
    101540.4,
  100839.8, 100980.3, 101092.6, 101174.7, 101277.5, 101366, 101447.8, 
    101521.4, 101575.5, 101614.5, 101653.7, 101687.9, 101722.6, 101725.2, 
    101737,
  100793.7, 100959.9, 101062.8, 101168.2, 101258.5, 101344, 101428.7, 
    101506.7, 101568.7, 101607.8, 101636.1, 101660, 101699.3, 101718.4, 101725,
  100761, 100939.5, 101045.1, 101145.6, 101234.4, 101324.8, 101408.3, 
    101488.6, 101556.5, 101595.8, 101622.1, 101639.1, 101671.8, 101695.2, 
    101704.5,
  100766.3, 100922.5, 101033.5, 101141.7, 101233.1, 101310.6, 101387.2, 
    101462.2, 101533.8, 101582.2, 101607.1, 101620.6, 101646.7, 101672.2, 
    101684.5,
  100790.6, 100915, 101030.9, 101135.3, 101223.7, 101307.5, 101378.1, 
    101446.1, 101510.5, 101567.6, 101599.7, 101608, 101621.8, 101641.1, 
    101651.4,
  100825.3, 100919.5, 101028.3, 101127.1, 101218.5, 101294.2, 101363.5, 
    101425.2, 101484.1, 101534.5, 101571.7, 101584.3, 101597.6, 101612.8, 
    101623.3,
  100839.8, 100932.3, 101025.7, 101112.5, 101205.1, 101288, 101353.4, 
    101416.4, 101467.6, 101510.1, 101544.2, 101564.6, 101569.4, 101570.8, 
    101581.2,
  100862.5, 100935.1, 101020, 101105.6, 101180.1, 101252.1, 101322.7, 
    101384.4, 101438.2, 101481.2, 101517.5, 101538.6, 101550.2, 101551.5, 
    101547.4,
  100881.5, 100952.3, 101024.6, 101094.6, 101165.9, 101235.7, 101299, 
    101356.3, 101409.5, 101453, 101490.8, 101516.8, 101530.5, 101532.8, 
    101528.8,
  100891.4, 100950.5, 101016.5, 101081.9, 101140.7, 101201.7, 101261.9, 
    101317.1, 101368.5, 101417, 101454.2, 101489.3, 101507.8, 101517.6, 101516,
  100478.6, 100408.5, 100376.6, 100365, 100370, 100390.9, 100425.1, 100473.6, 
    100530.9, 100602.1, 100688.5, 100781.6, 100896.9, 101017.7, 101130.2,
  100560.5, 100501.1, 100467.5, 100447.9, 100449.7, 100468.8, 100509.4, 
    100559, 100623.1, 100693.9, 100776.9, 100866.3, 100979.2, 101094.6, 
    101199.4,
  100673, 100620.3, 100584.1, 100561.2, 100558.1, 100573.6, 100608.5, 
    100657.5, 100718.6, 100784.7, 100855.9, 100937.3, 101036.1, 101140.5, 
    101243.2,
  100778.9, 100733.1, 100700, 100675.1, 100670.4, 100684.2, 100716.5, 
    100758.6, 100813, 100874.2, 100940.7, 101016.3, 101100.4, 101199.4, 
    101293.4,
  100870.5, 100831.8, 100808.2, 100791, 100792, 100803.9, 100834.9, 100872.9, 
    100918.3, 100972.8, 101032.4, 101095.4, 101163, 101245.2, 101328.4,
  100942.3, 100911.1, 100897.9, 100889, 100894.7, 100910.4, 100938.6, 
    100974.1, 101013.8, 101061.3, 101114, 101171.3, 101228.4, 101296.2, 
    101372.2,
  100990.9, 100972, 100969.1, 100965.9, 100978.7, 100997.5, 101027.5, 
    101058.1, 101090.1, 101136.7, 101187.1, 101239.8, 101287.6, 101338.9, 
    101401,
  101016.2, 101010.9, 101008.6, 101016.2, 101031.1, 101056.2, 101084.4, 
    101123.6, 101152.4, 101191, 101236.5, 101290.4, 101335.3, 101388.8, 101435,
  101026.1, 101020.2, 101036.2, 101039.6, 101052.7, 101081.5, 101118.3, 
    101160.4, 101196.2, 101233.7, 101272.3, 101319.1, 101367.5, 101411.9, 
    101460.6,
  101036.9, 101017.9, 101025.6, 101037.4, 101066.5, 101098.1, 101133.1, 
    101169.1, 101200.1, 101241.5, 101284.8, 101335.6, 101386.6, 101438.5, 
    101483.4,
  101095.2, 101026.3, 100975.3, 100925.9, 100874.7, 100821.6, 100767, 
    100709.6, 100652, 100594.1, 100534.4, 100478.3, 100427.1, 100383.7, 
    100352.5,
  101157.9, 101098.9, 101056.5, 101009.7, 100964.9, 100919.8, 100873.8, 
    100826.2, 100778.3, 100728.1, 100681, 100634.2, 100590, 100551.5, 100526.1,
  101214.2, 101167, 101132.3, 101090.7, 101051, 101013, 100974.2, 100935.1, 
    100893.1, 100852.1, 100811.7, 100772.8, 100736.3, 100706.3, 100683.8,
  101257.9, 101223.6, 101192.9, 101158.3, 101126.9, 101092.9, 101060.1, 
    101027.2, 100992.5, 100958.8, 100925.3, 100892.8, 100863.3, 100839.9, 
    100822,
  101289.2, 101267.9, 101246.2, 101217.9, 101191.4, 101162.9, 101136.5, 
    101108.9, 101081.4, 101053.6, 101026.7, 101001.1, 100979.2, 100959.9, 
    100948,
  101305.3, 101292.6, 101280, 101259.6, 101238.6, 101217.4, 101195.8, 
    101174.7, 101154, 101132.7, 101111.2, 101089.6, 101070, 101055.9, 101047.9,
  101307.9, 101297.4, 101294.8, 101282.4, 101270.9, 101255.2, 101240.2, 
    101224.2, 101208.5, 101190, 101171.1, 101154.6, 101140.8, 101130.9, 
    101126.5,
  101294.3, 101293, 101296.4, 101288.4, 101281.2, 101269.8, 101261.8, 
    101249.6, 101236.4, 101223.1, 101206.8, 101194.8, 101185.3, 101182.3, 
    101187.5,
  101258, 101266.9, 101278, 101273.9, 101269.3, 101265.7, 101258.1, 101251.4, 
    101241.9, 101235, 101225.3, 101220.4, 101221.5, 101226.7, 101234.7,
  101229.9, 101243.8, 101251.8, 101249.2, 101245, 101239.7, 101240.2, 
    101240.8, 101241, 101236.4, 101228.5, 101226.2, 101233.4, 101248.1, 
    101271.4,
  102208.2, 102178.8, 102135.4, 102087.6, 102026.9, 101960.4, 101875.6, 
    101787.3, 101693.8, 101593.7, 101481.6, 101361.5, 101238.9, 101111.6, 
    100980.4,
  102187.7, 102165.4, 102127.9, 102088.6, 102035.4, 101976.5, 101909.1, 
    101831.2, 101744.7, 101652.8, 101553.4, 101448.3, 101335, 101220.4, 
    101103.4,
  102138.4, 102127.2, 102103.2, 102072.2, 102034, 101985.5, 101923.8, 
    101854.5, 101777.6, 101696.8, 101608, 101514.3, 101415.1, 101313.6, 
    101208.9,
  102088.3, 102077.5, 102063.7, 102040.5, 102013.6, 101975.2, 101924.2, 
    101864.4, 101798, 101725.7, 101648.4, 101565.5, 101477.4, 101393, 101302.1,
  102026.3, 102022.5, 102005.3, 101992.2, 101975.3, 101946.8, 101912.4, 
    101865.3, 101809, 101744.7, 101677.1, 101608.9, 101536.9, 101459, 101378.6,
  101962.7, 101962.5, 101942.8, 101938.6, 101925.5, 101905.5, 101879.9, 
    101846, 101802.8, 101753.2, 101698.2, 101638.6, 101574.6, 101511.4, 
    101442.4,
  101901.3, 101897.1, 101886.2, 101874.4, 101864.1, 101854.6, 101837.7, 
    101814.6, 101783.8, 101743, 101697.8, 101649.7, 101597.6, 101540.7, 
    101482.6,
  101832.6, 101830.9, 101827.6, 101819.3, 101808.5, 101798, 101784.6, 101769, 
    101742.7, 101711.5, 101675.3, 101634.3, 101590.8, 101543.9, 101494.9,
  101733.9, 101742.6, 101742.5, 101742.6, 101740.7, 101739.1, 101732.5, 
    101720.7, 101700.2, 101673.4, 101643.3, 101609.7, 101571.3, 101530.8, 
    101486.6,
  101641.8, 101659.6, 101666.3, 101670.5, 101665.2, 101667.6, 101665, 
    101658.6, 101646, 101628.9, 101604.6, 101573.8, 101539.4, 101503.5, 
    101467.6,
  102263.8, 102276.8, 102278.7, 102272.4, 102256.1, 102231.5, 102200.9, 
    102163.2, 102121.7, 102072.1, 102021.2, 101961.7, 101899.2, 101831.1, 
    101759.2,
  102267.2, 102273.8, 102276.1, 102280.2, 102273.2, 102261.5, 102243.5, 
    102217.2, 102182.9, 102140.1, 102094.9, 102040.5, 101988.3, 101930.3, 
    101868.7,
  102236.3, 102265.2, 102275.9, 102278.5, 102280.5, 102274.7, 102263, 102249, 
    102227.9, 102196.9, 102157.1, 102112.5, 102063.9, 102010.9, 101956.5,
  102199.5, 102234.8, 102251.5, 102262.9, 102272.1, 102272.2, 102269.1, 
    102257.7, 102244.1, 102225.6, 102199.3, 102164.1, 102122.9, 102077.9, 
    102030.1,
  102147.7, 102189.7, 102213.5, 102234.2, 102242.8, 102253, 102253.9, 
    102252.8, 102247, 102234, 102216.1, 102193.5, 102160.1, 102127.1, 102087.9,
  102089.6, 102127.5, 102155.1, 102185.7, 102200.1, 102214.6, 102223.4, 
    102228.3, 102227, 102220.6, 102209.7, 102195.7, 102177.4, 102152, 102123.9,
  102023, 102058.4, 102088.2, 102119.6, 102143.8, 102162.8, 102173.1, 
    102183.9, 102187.1, 102189.5, 102186.1, 102178.1, 102167.9, 102153.7, 
    102136.5,
  101969.2, 102000.2, 102025.7, 102056.7, 102082, 102106.1, 102119.9, 
    102131.3, 102136.4, 102140.4, 102140.2, 102141.7, 102135.3, 102130.5, 
    102119.5,
  101888.9, 101914.8, 101940.6, 101971.6, 101998.7, 102025, 102044.1, 
    102057.8, 102067.7, 102077.9, 102081.5, 102083.1, 102084.7, 102083.4, 
    102079.3,
  101809.3, 101836.6, 101854.1, 101883.3, 101907.4, 101933.6, 101954.7, 
    101975.6, 101990.1, 102002.7, 102011.1, 102018.4, 102022.1, 102024.1, 
    102021.8,
  101665.5, 101698.1, 101725.4, 101746.3, 101770.6, 101784.1, 101791.9, 
    101793.4, 101790.4, 101783.8, 101775.3, 101762.2, 101746.7, 101730.5, 
    101714.2,
  101649.4, 101689.8, 101728.1, 101752.6, 101781, 101806.9, 101826.3, 
    101837.9, 101845.7, 101849.7, 101846.8, 101842.5, 101838.1, 101831.7, 
    101823.6,
  101629.6, 101685.2, 101722.9, 101751.8, 101783.7, 101816, 101841.9, 
    101860.4, 101877.8, 101889, 101896.5, 101904.3, 101904.6, 101905.2, 
    101902.4,
  101606.2, 101657.4, 101700.4, 101735.6, 101770.8, 101799.4, 101833.1, 
    101863.3, 101888.5, 101910.2, 101926.3, 101940.1, 101950.8, 101961.1, 
    101965.6,
  101573, 101626.6, 101670.8, 101708.3, 101745.8, 101778.8, 101814, 101844.4, 
    101875.8, 101905.5, 101931.5, 101951.6, 101973.2, 101991.9, 102005.7,
  101539, 101582.2, 101634.1, 101668.7, 101705.7, 101741.5, 101776.3, 
    101811.3, 101848.1, 101878.3, 101906.2, 101932.5, 101968, 101995.8, 
    102013.6,
  101502.3, 101541.8, 101587.2, 101627, 101663, 101696.5, 101732, 101768.1, 
    101799.1, 101831.4, 101866.5, 101897.9, 101929, 101963.1, 101993.3,
  101460.2, 101499.1, 101539.7, 101575.6, 101610.1, 101644.8, 101677.7, 
    101713.7, 101746.7, 101779.2, 101813, 101848.4, 101884.5, 101920.1, 
    101953.4,
  101425.5, 101451.7, 101485.2, 101520.4, 101552.3, 101584.9, 101617.9, 
    101651, 101683.7, 101717.6, 101753.4, 101787.7, 101823.9, 101859.3, 
    101900.2,
  101380.4, 101400.5, 101429.2, 101459.6, 101491, 101522.5, 101553.4, 
    101587.3, 101617.9, 101651.3, 101682.6, 101718.3, 101752.8, 101791.1, 
    101829.6,
  101749.7, 101752.2, 101769.6, 101783.4, 101790, 101795.9, 101798.3, 
    101801.9, 101805.6, 101803.5, 101793.2, 101777.3, 101750, 101721.2, 
    101693.8,
  101754.1, 101768.3, 101781.5, 101791.9, 101801, 101809.1, 101813.1, 
    101812.7, 101810.9, 101804.8, 101799.8, 101791.4, 101780.9, 101764, 
    101742.6,
  101744.3, 101761.6, 101781.5, 101795.8, 101805.7, 101816.1, 101819.4, 
    101818.9, 101819.7, 101817.2, 101815.7, 101807.9, 101797.9, 101787.1, 
    101775.6,
  101727, 101740.9, 101760.6, 101774.2, 101789.3, 101801.9, 101811.6, 
    101818.4, 101823.3, 101824.8, 101825.3, 101824.1, 101819.5, 101813.6, 
    101806.8,
  101687.2, 101707.4, 101721.1, 101737.2, 101754.5, 101771.7, 101788, 
    101800.8, 101812.5, 101819.8, 101828.8, 101832.3, 101833.4, 101832.4, 
    101828.7,
  101645.9, 101665.6, 101675.6, 101693.4, 101710.3, 101732.3, 101750.7, 
    101769.8, 101784.6, 101801.5, 101812.9, 101820.5, 101830.5, 101831.5, 
    101832.1,
  101594.8, 101617.4, 101628.8, 101644.9, 101661.3, 101682.4, 101702, 
    101724.7, 101746.4, 101765.9, 101781.1, 101792, 101805.5, 101815.7, 
    101823.6,
  101545.7, 101557.4, 101571.8, 101588.5, 101606.8, 101628.8, 101647.2, 
    101669.1, 101685.4, 101705.8, 101725.6, 101741.6, 101757.9, 101773.8, 
    101792.2,
  101490.6, 101508.4, 101519, 101534.5, 101550.1, 101567, 101586.3, 101603.5, 
    101626.5, 101645, 101665.7, 101682.1, 101703.1, 101726.8, 101746,
  101427.1, 101444.2, 101456.9, 101472.2, 101487.6, 101507.9, 101528, 
    101543.1, 101559.3, 101574.9, 101593.3, 101611.1, 101635.3, 101658, 
    101682.9,
  101891.5, 101942.1, 101992.1, 102042.4, 102090.2, 102130.2, 102175, 
    102227.6, 102290.4, 102352.1, 102396.3, 102435, 102462.7, 102490, 102538.7,
  101867.9, 101924.1, 101969.6, 102015.6, 102061.7, 102105.1, 102150, 
    102192.9, 102234.7, 102283.6, 102335.7, 102384, 102431.9, 102468.7, 
    102504.7,
  101829.9, 101889.3, 101937.8, 101989.6, 102036.9, 102082.5, 102124.5, 
    102167.2, 102203.1, 102245.2, 102290.6, 102338.9, 102392.6, 102435.8, 
    102476.2,
  101783.5, 101840.3, 101894.4, 101948.5, 101993.1, 102041.8, 102085.4, 
    102131.2, 102170.7, 102207.2, 102245.7, 102290.9, 102339.3, 102387.5, 
    102429,
  101735.7, 101789.1, 101840.5, 101893.3, 101944.3, 101993.6, 102038.9, 
    102083.8, 102125.8, 102167, 102202.3, 102235.1, 102274.8, 102315.8, 102359,
  101682.6, 101731.2, 101778.9, 101830.9, 101880.2, 101931.7, 101978.8, 
    102027.2, 102073.1, 102114.2, 102154.5, 102189.8, 102223.3, 102254.4, 
    102285.3,
  101629.9, 101674.5, 101716.3, 101764, 101811.1, 101860.4, 101908.7, 101955, 
    102000.4, 102047.2, 102089.4, 102130.4, 102165.4, 102199, 102225.9,
  101574.7, 101611.9, 101648, 101693, 101737.1, 101782.7, 101826.8, 101873.7, 
    101922.4, 101972, 102020.6, 102066, 102107.4, 102145.5, 102176.5,
  101518, 101546.2, 101577.4, 101616.8, 101658.1, 101701.1, 101740.8, 101782, 
    101826.4, 101876.5, 101930.2, 101984.7, 102035.1, 102077.2, 102114.3,
  101457.1, 101476.9, 101502.9, 101535.4, 101572, 101609.2, 101647.1, 
    101684.5, 101726.6, 101774.1, 101828.1, 101881.9, 101937.2, 101988.2, 
    102031.4,
  101613.8, 101651.7, 101696.4, 101737.4, 101777.9, 101814.2, 101846.1, 
    101873.9, 101904.2, 101934.7, 101962.9, 101992.4, 102022.4, 102054.3, 
    102085.3,
  101571.7, 101612.6, 101665.5, 101709.8, 101755.4, 101796.4, 101834.6, 
    101868, 101900.9, 101938.3, 101976.6, 102016.4, 102050, 102084.2, 102112.6,
  101525.9, 101574.1, 101621.8, 101671.4, 101723, 101771, 101814.2, 101855.5, 
    101898.2, 101937, 101977.1, 102016.7, 102056.5, 102097.9, 102132.6,
  101469.6, 101519.6, 101571.4, 101619.4, 101670.9, 101721.8, 101774.9, 
    101827.4, 101872.5, 101917.1, 101962.8, 102008.1, 102046.6, 102090.3, 
    102129.7,
  101417.7, 101467.1, 101512.2, 101560.4, 101613.7, 101669, 101723.6, 
    101780.2, 101837.7, 101890, 101939.9, 101987.4, 102032.3, 102073, 102113.7,
  101364.1, 101408.9, 101454.9, 101498.1, 101546.5, 101599.6, 101660.8, 
    101723.8, 101781.9, 101840.6, 101897, 101953.7, 102003.6, 102049.4, 102089,
  101315.1, 101357.5, 101396.7, 101437.9, 101482.1, 101530.9, 101588, 
    101650.9, 101714, 101780.9, 101843.6, 101907.4, 101965.1, 102017.2, 102062,
  101262.2, 101303.6, 101340.4, 101379.2, 101414.6, 101459.3, 101512.4, 
    101575.6, 101639.7, 101708.5, 101778.3, 101847.1, 101910.5, 101968.1, 
    102020,
  101213.5, 101255.8, 101288.8, 101324, 101356.6, 101392.9, 101436.7, 
    101497.1, 101563.8, 101632.5, 101703.8, 101777.6, 101848.9, 101911.9, 
    101969.1,
  101161.6, 101209.5, 101239.4, 101276.3, 101303.5, 101334.4, 101368.7, 
    101418.4, 101484.2, 101558.5, 101631, 101703.1, 101777.5, 101841.4, 
    101904.9,
  101670.1, 101710.7, 101750.8, 101792.6, 101828.6, 101859.5, 101883.2, 
    101905.8, 101932.7, 101949.1, 101967.1, 101995.5, 102027.5, 102064, 
    102088.4,
  101604.5, 101646.1, 101677.3, 101721.5, 101763.2, 101802, 101838.4, 
    101864.3, 101882.2, 101903.2, 101925.5, 101952.5, 101978.8, 102006.6, 
    102038.7,
  101545.1, 101583.5, 101608.9, 101656, 101698.5, 101738.5, 101771.8, 
    101802.2, 101828.2, 101851.7, 101878.4, 101910.8, 101946.3, 101978.9, 
    102004.9,
  101491.8, 101524.2, 101555, 101595.3, 101636.7, 101687.6, 101726.4, 
    101766.4, 101800.6, 101829.2, 101863.6, 101900.7, 101939.8, 101973.5, 
    102003.3,
  101460.4, 101482.2, 101501.6, 101541.3, 101582.5, 101629.4, 101673.5, 
    101716.6, 101757.3, 101797.8, 101833.5, 101873, 101909.7, 101950.6, 101989,
  101422.3, 101445.6, 101467.3, 101493.2, 101528.2, 101573, 101618, 101664.1, 
    101702.7, 101745.1, 101784.9, 101830, 101875.1, 101923.6, 101968.9,
  101384.8, 101418.6, 101438.1, 101459.9, 101485.3, 101519, 101561.2, 
    101606.1, 101651.6, 101700.4, 101747.9, 101793, 101840.8, 101882.5, 
    101939.2,
  101332.4, 101382.4, 101406.8, 101434, 101446.8, 101472.5, 101504.8, 
    101546.2, 101593.4, 101640.4, 101690.8, 101744.1, 101798.8, 101846.1, 
    101895.8,
  101299, 101343.7, 101373, 101407.7, 101429.7, 101434.4, 101453.1, 101487.2, 
    101532.6, 101581.4, 101639.6, 101696.8, 101751.4, 101810.1, 101856.1,
  101274.3, 101319.7, 101352.2, 101377.5, 101404.1, 101418.9, 101422.4, 
    101431.4, 101471.2, 101522.1, 101585.2, 101643.9, 101707, 101762.8, 
    101822.6,
  101555.5, 101619.4, 101688.6, 101754.7, 101818.4, 101872.2, 101909.7, 
    101940.4, 101965.4, 101981.7, 102005.3, 102034.6, 102073.5, 102126, 
    102175.1,
  101495.8, 101561.6, 101623.7, 101682.4, 101737.8, 101790.9, 101836.9, 
    101870.9, 101895, 101907.4, 101913.5, 101928.2, 101957.6, 102006.6, 
    102066.1,
  101448.1, 101510.6, 101564.6, 101617.1, 101667.5, 101708.9, 101753.3, 
    101784.7, 101806.6, 101815.1, 101819, 101829.1, 101855.4, 101924.2, 
    102000.3,
  101406.4, 101453.9, 101505.1, 101557, 101606, 101647.3, 101692.8, 101732.1, 
    101761.4, 101778.5, 101782.5, 101775, 101781.2, 101821.9, 101916.7,
  101379.6, 101417.5, 101457.4, 101495.1, 101537.5, 101577, 101624.8, 
    101662.3, 101702.1, 101731.6, 101751, 101762.1, 101764.8, 101762.8, 
    101800.7,
  101340.4, 101387.4, 101422.7, 101450.5, 101485.6, 101519.7, 101557.6, 
    101601.1, 101649.9, 101686.8, 101717.9, 101733.1, 101742.1, 101754.8, 
    101772.6,
  101313.9, 101363.7, 101392.6, 101419, 101439, 101461.8, 101496, 101537, 
    101584.8, 101633.9, 101676.2, 101707.6, 101733.2, 101740.3, 101769.5,
  101285.2, 101334.9, 101374.8, 101397.7, 101407.9, 101418.9, 101441.8, 
    101475.8, 101525, 101583.4, 101633.5, 101679.9, 101704.3, 101738.9, 
    101756.4,
  101275.1, 101318.5, 101354.6, 101381.6, 101391.2, 101391.4, 101394.4, 
    101413.3, 101464.5, 101530.7, 101587.5, 101637.2, 101687.9, 101729.2, 
    101751.7,
  101262.1, 101308.4, 101341.9, 101364.5, 101385.1, 101381.9, 101374.2, 
    101374.6, 101398.7, 101472.7, 101536, 101606.8, 101652.1, 101702.7, 
    101747.8,
  100725.1, 100829.1, 100930.8, 101021, 101107.9, 101198.3, 101282.4, 
    101362.8, 101433.6, 101509.3, 101585.7, 101668.1, 101755.3, 101848.9, 
    101963.9,
  100724.9, 100825.1, 100921.6, 101006.2, 101086, 101171.6, 101259.5, 
    101344.8, 101415.9, 101483.3, 101551.5, 101622.7, 101698.6, 101788.7, 
    101888.3,
  100728.8, 100826.9, 100914.8, 100992.8, 101070.2, 101151.3, 101240, 
    101328.4, 101394.7, 101455.1, 101515, 101571.2, 101635.2, 101719.1, 
    101819.5,
  100743.1, 100831.6, 100913.5, 100985.2, 101053.7, 101126.8, 101207, 
    101300.7, 101374.5, 101435.9, 101491.7, 101539.4, 101582.6, 101641.6, 
    101732,
  100750.7, 100842.3, 100920.8, 100983.3, 101044.5, 101107.1, 101186, 101273, 
    101353, 101415.2, 101476, 101517, 101559.6, 101591.9, 101657.8,
  100757.6, 100850.4, 100930.3, 100988.8, 101040.2, 101093.6, 101160.5, 
    101245.1, 101325.2, 101393.1, 101458.5, 101504.1, 101549.2, 101571, 
    101607.4,
  100767.9, 100860.5, 100936.9, 100995.9, 101042, 101088.8, 101143.5, 
    101220.2, 101301.2, 101373, 101440.1, 101490.3, 101544, 101580.8, 101613.2,
  100786, 100874.9, 100947.7, 101006.3, 101047.8, 101087.3, 101131.5, 
    101198.9, 101280.1, 101355, 101421.4, 101488.7, 101527.9, 101579.1, 
    101608.6,
  100811, 100893.6, 100960.8, 101016.3, 101056.4, 101087.4, 101120.9, 
    101179.6, 101255, 101331.5, 101400.7, 101462.3, 101520, 101565.8, 101609.6,
  100839.1, 100917.1, 100979, 101025.4, 101065.3, 101091.2, 101105.6, 
    101159.7, 101227.4, 101305.2, 101375.5, 101443.2, 101500.1, 101549.1, 
    101596.5,
  101154.9, 101079.8, 101013.1, 100963.7, 100926.8, 100896.1, 100869.9, 
    100855.6, 100847.7, 100844.1, 100850.2, 100871.7, 100899.7, 100940, 100992,
  101152.4, 101086.9, 101036.7, 100994.2, 100960, 100927.5, 100897.9, 
    100884.9, 100882.3, 100893.9, 100915.5, 100950.1, 100984.3, 101027, 
    101078.4,
  101161.8, 101122.5, 101065.1, 101023.6, 100983.2, 100954.8, 100934.8, 
    100928.1, 100929.5, 100946.9, 100970.7, 101003, 101036.2, 101081, 101136.4,
  101164, 101124.8, 101064, 101024.3, 100987.2, 100960.5, 100942.4, 100937.6, 
    100946.6, 100969.8, 101001.9, 101042.8, 101090, 101141.1, 101197.1,
  101146, 101103.9, 101052.5, 101018.5, 100983.3, 100960.2, 100947.9, 
    100952.6, 100968.3, 100999.4, 101036.7, 101081.7, 101129.9, 101180.6, 
    101243.4,
  101126.4, 101084.8, 101041.5, 101008, 100976.4, 100957.5, 100953, 100956.4, 
    100976.3, 101011.5, 101056.6, 101110.4, 101167.4, 101229, 101294.5,
  101108.9, 101073.1, 101036.4, 101007.5, 100980.1, 100960.3, 100952, 100956, 
    100980.9, 101022.1, 101080, 101144.1, 101204.9, 101268.8, 101333.2,
  101092.6, 101069.5, 101040.6, 101012.4, 100987.2, 100966.7, 100955.2, 
    100962.6, 100993.8, 101044.8, 101104.8, 101169.4, 101233.7, 101298.1, 
    101363.3,
  101082.9, 101065.2, 101038.8, 101014.4, 100994.1, 100976.1, 100959.8, 
    100972.6, 101007, 101062, 101122.6, 101185.4, 101250.8, 101313.5, 101379.4,
  101077.3, 101066.2, 101042.5, 101021.7, 101003.1, 100985.7, 100970.9, 
    100986.1, 101020.2, 101072.3, 101129.5, 101193.9, 101257.4, 101318.3, 
    101383.6,
  102194.1, 102170.9, 102153.7, 102136.3, 102116.1, 102094.8, 102076.8, 
    102050.7, 102019, 101996, 101967.6, 101935.5, 101903.1, 101861.7, 101818.3,
  102149.1, 102123.4, 102105.7, 102081.4, 102060, 102036.3, 102010.7, 
    101980.5, 101957.7, 101930.2, 101899.2, 101868.4, 101836.7, 101798.6, 
    101756.3,
  102094.6, 102072.9, 102048.5, 102019.3, 101993, 101960.5, 101933.5, 
    101904.9, 101876.7, 101849.9, 101829, 101804.2, 101774.4, 101738.3, 
    101703.4,
  102045.9, 102017, 101983.5, 101948.3, 101914.9, 101884.6, 101850.5, 
    101813.2, 101791.3, 101768.9, 101749.2, 101725, 101694.5, 101668.4, 
    101641.1,
  101987, 101950.1, 101913.4, 101872.9, 101833, 101794.4, 101754.5, 101720.4, 
    101692.3, 101668, 101647.6, 101626.5, 101611, 101593.2, 101567.7,
  101928.9, 101888.4, 101842.8, 101794.6, 101746, 101697.3, 101645.1, 
    101610.8, 101571.7, 101556.9, 101547.7, 101542.2, 101529.1, 101511.6, 
    101493.9,
  101872.3, 101825.4, 101767.7, 101714.3, 101648.5, 101579.9, 101528, 101483, 
    101448.7, 101437.6, 101435.3, 101434.9, 101429.8, 101421.9, 101411,
  101819.3, 101762.8, 101697.5, 101633.6, 101551.3, 101480, 101416.4, 
    101357.8, 101310.1, 101304.4, 101328.8, 101345.1, 101347.2, 101358.4, 
    101359.4,
  101763.7, 101705.1, 101630.3, 101554.7, 101461.6, 101380.5, 101299, 
    101195.4, 101153.4, 101171.6, 101220.1, 101269.1, 101303.2, 101333.6, 
    101353.7,
  101713.4, 101646.6, 101569.3, 101488.7, 101386.9, 101298.4, 101203.3, 
    101110.2, 101089.3, 101130.9, 101199.8, 101240.6, 101288.1, 101322.4, 
    101361.8,
  102240.7, 102250.1, 102247.1, 102245.9, 102238.8, 102239.3, 102229.8, 
    102219.7, 102201.3, 102188, 102169.7, 102153, 102131, 102106.6, 102081.6,
  102212.5, 102212.2, 102216.7, 102223.3, 102225.9, 102223.9, 102216.8, 
    102216.7, 102215.2, 102204.3, 102191.7, 102172.6, 102150.1, 102128, 
    102110.6,
  102148.5, 102156.5, 102159.5, 102163.6, 102167.3, 102170.9, 102177.6, 
    102180.7, 102183.1, 102179.7, 102173.1, 102165.6, 102150.4, 102134.1, 
    102116.3,
  102086.2, 102091.5, 102092.5, 102100.5, 102105.7, 102115.5, 102124.6, 
    102134.8, 102139.4, 102139.4, 102136.5, 102128.3, 102121, 102108.8, 
    102092.8,
  102003.6, 102003.7, 101996.3, 102001.6, 102014.2, 102027.8, 102045.5, 
    102057.6, 102062.1, 102065.9, 102072.1, 102070.6, 102070.5, 102062.3, 
    102047.5,
  101926.7, 101916.8, 101907.7, 101916.9, 101921.3, 101931.5, 101940.9, 
    101952.3, 101966.1, 101980.3, 101983.6, 101984.9, 101987.2, 101986.8, 
    101983.9,
  101841.3, 101818.7, 101805.2, 101802.3, 101799.8, 101809.5, 101817.6, 
    101833.3, 101844.7, 101857.5, 101872.6, 101880.8, 101894.3, 101897.4, 
    101897.9,
  101755, 101727.8, 101703.6, 101688.6, 101681.3, 101685.6, 101696.6, 
    101719.5, 101742.9, 101761.6, 101776.2, 101787.4, 101798.2, 101806, 
    101810.2,
  101667.3, 101631.4, 101588.6, 101564.6, 101547.4, 101551.2, 101562.5, 
    101584, 101604.1, 101629.8, 101654.2, 101677.4, 101695.2, 101711.3, 
    101721.9,
  101582.7, 101537.7, 101480.8, 101451.5, 101432.6, 101444.4, 101463, 
    101492.5, 101519.9, 101552.4, 101577.8, 101602, 101625.1, 101649.8, 
    101669.9,
  102311.2, 102353, 102380.8, 102406.3, 102424.9, 102448.4, 102462.3, 
    102470.8, 102475.1, 102469.2, 102474, 102482.1, 102479.4, 102467.7, 
    102463.7,
  102281.7, 102319, 102348.9, 102378.9, 102402.3, 102423.5, 102440, 102457.8, 
    102474, 102482.8, 102481.1, 102482.4, 102479.9, 102490.9, 102493.4,
  102227.6, 102260.7, 102293.9, 102326.4, 102350.4, 102377.4, 102399.9, 
    102420.3, 102436, 102452.6, 102466.5, 102477.5, 102483, 102490.3, 102497.3,
  102168.4, 102202.4, 102232.3, 102261.8, 102288.9, 102317.2, 102340.2, 
    102362.6, 102384.2, 102403.7, 102419.7, 102435.2, 102448.3, 102456.5, 
    102464.4,
  102100, 102130.2, 102153.2, 102182.1, 102205.9, 102229.8, 102258.1, 
    102286.1, 102309.7, 102330.4, 102350.9, 102367, 102380.7, 102394.4, 
    102406.9,
  102028, 102061.7, 102091.5, 102117.7, 102137.3, 102163.2, 102182, 102203.9, 
    102223.8, 102244.2, 102263.5, 102282.2, 102301.6, 102319.1, 102339.8,
  101948.7, 101975.2, 101995.7, 102024.8, 102047.4, 102066.5, 102084.3, 
    102105, 102121.5, 102138.6, 102156.4, 102176.1, 102191.4, 102208.4, 102228,
  101869, 101897.7, 101910.9, 101934.2, 101949.5, 101973, 101990.2, 102005.2, 
    102020.7, 102036.5, 102053.1, 102068.3, 102087.2, 102107, 102128,
  101773.2, 101799.5, 101809.7, 101828.8, 101839.1, 101853.2, 101863.2, 
    101872.5, 101886, 101902.6, 101920.5, 101940.9, 101961.6, 101985.2, 
    102008.5,
  101687.5, 101707, 101710.6, 101725.3, 101732.5, 101744.2, 101749.1, 
    101758.3, 101767.7, 101782.5, 101801.6, 101823.8, 101851.6, 101882.7, 
    101920.1,
  102203.3, 102236.2, 102259.9, 102284.8, 102298.3, 102314, 102319.1, 
    102317.2, 102320.6, 102311.7, 102297.6, 102277.9, 102258.2, 102235, 
    102210.9,
  102151.4, 102180.7, 102207.7, 102234.4, 102254.8, 102272.6, 102286.9, 
    102297.3, 102306.6, 102314, 102315.1, 102310.4, 102301.9, 102281.5, 
    102269.3,
  102086.8, 102111.8, 102135.9, 102157.6, 102180.3, 102200.8, 102217.5, 
    102235, 102250, 102267.5, 102277.6, 102279.8, 102284.3, 102282, 102293.2,
  102029.6, 102044.3, 102061.6, 102080.7, 102102.5, 102123.4, 102144.2, 
    102164.9, 102184.2, 102201.3, 102215.9, 102231.6, 102248.6, 102253.4, 
    102258.6,
  101963.5, 101973.8, 101983.4, 101998.5, 102014.2, 102030.9, 102049.8, 
    102068.7, 102092, 102109.9, 102131.4, 102148, 102167.7, 102187.8, 102210.9,
  101885.7, 101895.9, 101900.4, 101909.3, 101918.8, 101931.7, 101947.2, 
    101965.1, 101984, 102005, 102027.9, 102051.7, 102074, 102097.2, 102121.9,
  101807, 101809.3, 101804.5, 101800.5, 101802.4, 101811, 101824.3, 101841.2, 
    101862, 101884.4, 101910.9, 101938.9, 101969.3, 102000.8, 102027.8,
  101725.8, 101712.8, 101701.1, 101691.8, 101691.3, 101692.6, 101700, 
    101710.3, 101730.9, 101757.4, 101788.5, 101822.1, 101855.8, 101893.5, 
    101926.4,
  101640, 101613.5, 101593.3, 101570.8, 101557.1, 101551.6, 101552.8, 
    101564.1, 101588.9, 101621.7, 101660.7, 101703.7, 101749.3, 101795.6, 
    101836.7,
  101549.4, 101509.2, 101477.6, 101443.2, 101420.6, 101407, 101406, 101420.5, 
    101452, 101492.3, 101544.1, 101597.7, 101656, 101708.7, 101764.2,
  102032.1, 102064.9, 102088.4, 102115.8, 102132.3, 102148.2, 102154.5, 
    102155.8, 102151.3, 102141.7, 102131.1, 102117.6, 102108.7, 102085.9, 
    102066.8,
  101976.8, 102009.8, 102031.8, 102062.8, 102085.3, 102106.3, 102123.1, 
    102135.3, 102141.7, 102143.8, 102138.3, 102122.2, 102110.1, 102083.8, 
    102063.2,
  101897.4, 101928.9, 101951.8, 101979.3, 102002.9, 102027, 102051.2, 
    102075.4, 102091.2, 102104.8, 102112.9, 102113.6, 102109.5, 102104.1, 
    102090.2,
  101827.9, 101847.6, 101865.5, 101889.2, 101913.5, 101937.1, 101964.8, 
    101989.9, 102013.8, 102031.1, 102045.6, 102056.8, 102075, 102080.5, 
    102072.7,
  101747.2, 101750.7, 101763.6, 101776.7, 101796.8, 101813.9, 101837.2, 
    101862.1, 101891, 101918.6, 101945.3, 101972, 101994, 102011, 102021.1,
  101655.7, 101647.1, 101652.8, 101659.7, 101673.9, 101690.2, 101712.5, 
    101739.4, 101767.5, 101796.3, 101824.2, 101852.4, 101879.3, 101903.5, 
    101925.2,
  101556.6, 101538.2, 101533.5, 101532.5, 101541.2, 101556.6, 101578, 
    101604.6, 101635.6, 101670.5, 101707.3, 101742.7, 101776.2, 101804.4, 
    101825.5,
  101457.9, 101432.3, 101413.5, 101406.9, 101410.7, 101424.5, 101446.1, 
    101472.7, 101504.5, 101541.1, 101578.7, 101618.5, 101652.6, 101688.7, 
    101715.2,
  101355.5, 101318.9, 101290.4, 101277.4, 101279.3, 101296.1, 101322, 
    101357.7, 101406.7, 101454.9, 101502.2, 101548.2, 101593.8, 101634.8, 
    101668.8,
  101249.4, 101209, 101172.7, 101156.8, 101158.5, 101173.6, 101203.6, 
    101249.9, 101297.6, 101344.5, 101391.2, 101440.1, 101490.4, 101551.3, 
    101610.7,
  101452.3, 101497.6, 101533.6, 101573, 101604.6, 101630.9, 101658.9, 
    101685.2, 101711.7, 101730.5, 101756.6, 101795.6, 101828, 101850.4, 
    101886.3,
  101436.9, 101474.5, 101511.6, 101547.4, 101585.4, 101620.4, 101651.8, 
    101680.7, 101708.6, 101736.6, 101758.5, 101784.2, 101811.8, 101831.1, 
    101875.1,
  101410.7, 101444.4, 101480.8, 101516.7, 101549.5, 101582.1, 101618.2, 
    101652.2, 101685.4, 101717.7, 101751, 101780.5, 101810.1, 101839.9, 
    101851.1,
  101374.3, 101405.2, 101434.9, 101466.6, 101501.3, 101532.2, 101566.7, 
    101603, 101639.5, 101676, 101713.6, 101751, 101787.9, 101821.3, 101848.8,
  101332.8, 101356.8, 101382.7, 101407.4, 101433.5, 101459.5, 101491.8, 
    101526, 101563.4, 101602.3, 101642.9, 101686.2, 101730.6, 101772.6, 
    101810.7,
  101282.5, 101296.6, 101315, 101335.1, 101358.8, 101384.5, 101412.7, 
    101446.1, 101481.8, 101521.5, 101562.7, 101606.2, 101651.5, 101695.8, 
    101743.3,
  101228.1, 101230.8, 101239.4, 101248.7, 101265.1, 101285.7, 101311.8, 
    101343.5, 101380.8, 101421.9, 101467.5, 101515, 101565.2, 101615.1, 101664,
  101166.3, 101158.4, 101156.4, 101157.1, 101166.7, 101182.1, 101205.8, 
    101236.2, 101275.8, 101320.6, 101370.8, 101421.9, 101475.2, 101528.3, 
    101580.6,
  101103.6, 101085.6, 101072, 101060.8, 101060.2, 101067.7, 101086.2, 
    101115.8, 101157.2, 101206.7, 101264.5, 101325.2, 101388.1, 101449.6, 
    101508.5,
  101037.5, 101006.7, 100979, 100954.6, 100940, 100939.2, 100951.2, 100979.2, 
    101022.8, 101078.6, 101148, 101220.3, 101297.9, 101373.5, 101443.7,
  101191.5, 101179.3, 101175.2, 101171.8, 101169.4, 101164.7, 101166.8, 
    101166.1, 101165.3, 101162, 101157.8, 101151.5, 101145.9, 101142.9, 
    101143.2,
  101205.3, 101189.3, 101197.1, 101195.5, 101198, 101199.2, 101202.9, 
    101209.3, 101212.2, 101215.6, 101217.5, 101220.4, 101224.2, 101232.4, 
    101243.6,
  101204.2, 101195.6, 101207.4, 101203.9, 101205, 101204.7, 101205.5, 
    101211.6, 101222.1, 101232, 101241.4, 101251.3, 101263, 101280.2, 101298.2,
  101191.1, 101171.8, 101181.6, 101174.3, 101178.3, 101178.1, 101186, 
    101191.3, 101201.6, 101215.2, 101234.6, 101256.4, 101279.7, 101307.5, 
    101334.8,
  101163.6, 101141.2, 101138.2, 101125.1, 101127.6, 101125.9, 101127.9, 
    101135.3, 101155.4, 101183, 101217.2, 101250, 101283.4, 101316.7, 101350.5,
  101128.3, 101094.5, 101084.5, 101060.7, 101051.3, 101035.4, 101042.4, 
    101062.6, 101095.3, 101133.6, 101175.4, 101220.9, 101265.9, 101309.8, 
    101352.4,
  101088.4, 101034.2, 101013.9, 100974.3, 100949.5, 100936.3, 100944.4, 
    100964.4, 101003.2, 101052.7, 101113.8, 101175.5, 101234.9, 101294.8, 
    101347.2,
  101038.7, 100978.7, 100940.2, 100878.8, 100843.5, 100815.9, 100811.7, 
    100835.6, 100883.8, 100944.2, 101017.7, 101097, 101178, 101250, 101322.5,
  100993.7, 100923.4, 100857.1, 100778.5, 100722.4, 100669.5, 100653.9, 
    100671.5, 100726.5, 100803.4, 100891.9, 100987.6, 101088.3, 101183.4, 
    101271.2,
  100953.1, 100872.3, 100784.7, 100690.8, 100605.1, 100525, 100478.5, 
    100480.4, 100539.6, 100638.4, 100754.4, 100857.8, 100974.8, 101085.3, 
    101198.5,
  101464.8, 101483.8, 101491.6, 101496.4, 101501.8, 101513, 101515.2, 
    101516.6, 101516.7, 101520.5, 101516.5, 101513.3, 101496.7, 101481.9, 
    101460,
  101433.3, 101440.2, 101446.7, 101446.3, 101443.7, 101441.1, 101449.1, 
    101458, 101466.1, 101468.5, 101465.6, 101459, 101452.4, 101442.8, 101432.3,
  101388.4, 101390.7, 101396.2, 101393.4, 101396.1, 101401, 101403.2, 101407, 
    101408.7, 101414.4, 101422.1, 101421.2, 101419, 101414.6, 101405.9,
  101344.3, 101340.1, 101340.6, 101337.6, 101333.7, 101326, 101323.2, 
    101326.8, 101327.8, 101330.2, 101330.9, 101337.1, 101344.9, 101348.4, 
    101351.9,
  101321.9, 101309.4, 101302.5, 101283.6, 101270, 101252.5, 101236.8, 
    101228.3, 101232.1, 101242.6, 101260.4, 101268.6, 101284.1, 101300, 
    101315.3,
  101297.2, 101274.8, 101253.2, 101221, 101194.4, 101160.1, 101133, 101120.1, 
    101119.8, 101129, 101143.8, 101164, 101190, 101211, 101234.2,
  101278.3, 101244, 101210.1, 101167.7, 101117.1, 101059.4, 101014.6, 
    100985.6, 100978.3, 100997.1, 101035, 101075.9, 101110.8, 101150.9, 
    101181.1,
  101254.8, 101209.8, 101163.2, 101101.8, 101032, 100958.8, 100884, 100824.9, 
    100807.8, 100842, 100908.9, 100983, 101038.9, 101089.9, 101133,
  101233.2, 101183.7, 101124.6, 101051.9, 100965.5, 100865.2, 100750.9, 
    100656.5, 100613.3, 100640.9, 100739.5, 100866, 100968.6, 101042.4, 
    101084.5,
  101217.6, 101156.9, 101083.7, 101003.1, 100903.1, 100785.4, 100633.4, 
    100488.8, 100361.6, 100375, 100539.9, 100709.5, 100866.3, 100982.3, 
    101046.7,
  101243.1, 101197.5, 101168.2, 101135, 101107.8, 101084.7, 101069.7, 
    101065.4, 101068.4, 101080.2, 101104.4, 101142.5, 101204.5, 101298.5, 
    101404.5,
  101261.7, 101222.1, 101195.3, 101156.2, 101124.7, 101096.7, 101078.4, 
    101065.1, 101054.9, 101055, 101060.9, 101079.2, 101121.8, 101192.7, 
    101275.4,
  101273.6, 101234, 101201.6, 101162.2, 101130.3, 101099.8, 101073.5, 
    101052.6, 101035.4, 101033.5, 101037, 101057.7, 101098.4, 101164.4, 
    101244.6,
  101271.1, 101233.9, 101196.5, 101152.9, 101115.8, 101081.1, 101047.1, 
    101020.8, 101006, 101007.2, 101018.4, 101043.5, 101081.6, 101137.4, 101204,
  101263.1, 101225.2, 101184.6, 101138.6, 101093.1, 101047.6, 101007.7, 
    100977.6, 100969, 100977.5, 100995.6, 101027.8, 101074.4, 101130.2, 
    101196.5,
  101247, 101209.9, 101162.9, 101107.6, 101052.5, 100997.2, 100947, 100918.8, 
    100914.2, 100923.9, 100954.9, 101000.5, 101053.1, 101107, 101171.3,
  101231.7, 101190, 101139.2, 101076.4, 101006.8, 100933, 100872.2, 100842, 
    100842.2, 100867.6, 100919.2, 100973.8, 101029.2, 101084.1, 101145.3,
  101215.3, 101171, 101114.6, 101043.7, 100956.4, 100861.2, 100782, 100742.7, 
    100757.4, 100808, 100873.2, 100942.7, 101008.6, 101068.8, 101127.8,
  101194.1, 101160.6, 101104.3, 101025.2, 100919.5, 100797.1, 100691.3, 
    100635.2, 100667.5, 100738.8, 100823.2, 100909.2, 100989.7, 101051.8, 
    101117.5,
  101188.5, 101152.6, 101098.5, 101016.8, 100901.2, 100754.4, 100611.5, 
    100528.4, 100559.3, 100654.3, 100760.6, 100863.3, 100961.6, 101036.1, 
    101107.8,
  101821.5, 101748.9, 101688.4, 101616.7, 101539.8, 101453.3, 101361.5, 
    101264.4, 101166.1, 101065.4, 100963.8, 100860.3, 100754.5, 100639, 
    100524.3,
  101834, 101761.3, 101705.9, 101639.2, 101570, 101489.7, 101407.7, 101319.6, 
    101229.1, 101136.1, 101038.5, 100940.1, 100836.1, 100728.3, 100623.6,
  101845.3, 101785.6, 101730.1, 101663, 101600.8, 101528.6, 101453, 101372.7, 
    101288.2, 101199.5, 101110.5, 101017.5, 100921.2, 100828.7, 100740.4,
  101849.3, 101796.2, 101737.7, 101675.9, 101616.4, 101549.9, 101477.4, 
    101398.4, 101317.4, 101233.9, 101146.5, 101061.1, 100978.8, 100900, 
    100826.5,
  101852.9, 101801.7, 101745.3, 101685.1, 101622.7, 101557.9, 101487.2, 
    101412.3, 101331.7, 101248.9, 101169.7, 101090.3, 101019.2, 100954.6, 
    100898.4,
  101850.8, 101798.8, 101744.8, 101684.6, 101618.5, 101554, 101479.8, 101401, 
    101323.2, 101246.4, 101168.5, 101095.5, 101037.7, 100986.3, 100937.7,
  101843.3, 101790.1, 101737.8, 101674.4, 101606.6, 101536.3, 101461, 101382, 
    101305.6, 101223.8, 101153.5, 101092.9, 101039.2, 100991, 100955.3,
  101825.5, 101773.1, 101720.8, 101654.2, 101582.5, 101509.1, 101429.8, 
    101349.7, 101268.6, 101188.9, 101124.4, 101065.8, 101019.6, 100983.7, 
    100944.5,
  101800.8, 101748.7, 101691.7, 101623.7, 101552.3, 101476.6, 101394.4, 
    101311.1, 101221.3, 101143.6, 101077.4, 101031.6, 100990.6, 100953.7, 
    100924.5,
  101765.5, 101715.7, 101657, 101589.3, 101516.8, 101442.4, 101358.1, 
    101269.4, 101171.4, 101085.3, 101016.7, 100986.2, 100945.1, 100924.9, 
    100909.2,
  102224.9, 102195.6, 102176, 102148.6, 102120.4, 102083.5, 102045.3, 
    102007.4, 101958.7, 101907.7, 101846.9, 101784, 101714.6, 101629.3, 
    101536.6,
  102218.7, 102202.5, 102190.6, 102162.4, 102142.2, 102107.4, 102068, 
    102027.1, 101983.7, 101932.4, 101873.9, 101806.2, 101738.5, 101666.9, 
    101581.3,
  102219.9, 102210.6, 102199.7, 102175.1, 102151.3, 102124.6, 102089.8, 
    102048.1, 102006.2, 101955.6, 101897.9, 101835.5, 101770.3, 101701.1, 
    101624.5,
  102206.6, 102201.6, 102189.8, 102173.7, 102156.9, 102130, 102095.4, 
    102059.9, 102016.9, 101969.1, 101915.8, 101852.1, 101786.6, 101723.4, 
    101651.7,
  102189.4, 102189.3, 102181.3, 102164.8, 102153.2, 102124.5, 102097.9, 
    102064.4, 102023.5, 101978.3, 101925.3, 101868.3, 101804.2, 101737.6, 
    101669.3,
  102167.5, 102169.3, 102158, 102149.1, 102137.4, 102119.1, 102088.9, 
    102056.8, 102019.9, 101975.4, 101926.2, 101869.6, 101808, 101739.8, 
    101670.4,
  102139.2, 102144.4, 102136.8, 102127.1, 102116.1, 102098.6, 102071, 
    102038.1, 101999.3, 101960, 101914.3, 101861.1, 101800.5, 101735.4, 
    101666.1,
  102112.7, 102117.4, 102104.8, 102093.9, 102079.9, 102061.9, 102039.5, 
    102007.8, 101972.4, 101935.2, 101889, 101838.4, 101781.8, 101716.5, 
    101657.1,
  102080.4, 102081.8, 102066, 102055.4, 102037.7, 102019.5, 101993.7, 
    101965.4, 101931.8, 101893.4, 101851, 101804.7, 101750.1, 101693.1, 
    101640.3,
  102041.5, 102037.2, 102021.9, 102009.2, 101988.9, 101967.3, 101944.5, 
    101917.9, 101884, 101850.7, 101811.2, 101765.1, 101713.4, 101664.9, 
    101612.8,
  102337.9, 102356.3, 102375.5, 102380.8, 102388.6, 102390.5, 102383.9, 
    102380.1, 102365.8, 102360.7, 102348.9, 102332.9, 102319.1, 102301.7, 
    102280.2,
  102316, 102350.6, 102378.4, 102390, 102398.3, 102406.2, 102403.9, 102396.6, 
    102390, 102378, 102367, 102354.1, 102331.4, 102318.8, 102302.8,
  102305.9, 102344.4, 102370.8, 102394, 102407.4, 102418.9, 102420.7, 
    102415.7, 102409.1, 102410.5, 102384.4, 102367.8, 102355.8, 102344.6, 
    102325.5,
  102279.3, 102320.6, 102356.8, 102382.9, 102399.6, 102412.9, 102416.4, 
    102420.9, 102417.1, 102413.9, 102398.2, 102381.9, 102368.5, 102349.3, 
    102335.7,
  102258.2, 102296.1, 102331.7, 102361.1, 102386.2, 102399.2, 102402.7, 
    102414.2, 102418.5, 102408.9, 102404.9, 102390.1, 102372.6, 102347.8, 
    102331,
  102232.9, 102268.5, 102298.9, 102329.5, 102352.1, 102370.8, 102379.6, 
    102388.8, 102394.4, 102388.8, 102383.6, 102370.5, 102357.2, 102341.9, 
    102321.6,
  102206.3, 102240.4, 102269.7, 102296.4, 102312.2, 102330.9, 102339.6, 
    102344.1, 102347.5, 102346.4, 102346.4, 102337.8, 102329.4, 102311.4, 
    102293.3,
  102176.6, 102201.4, 102225.2, 102251.8, 102269.4, 102286.4, 102292.7, 
    102294, 102299.7, 102302, 102300.8, 102297.1, 102289.9, 102276.4, 102262.5,
  102141.3, 102160.2, 102181.1, 102197.5, 102212.5, 102224.9, 102234.6, 
    102241.2, 102247.5, 102250.6, 102254.1, 102249.2, 102240.6, 102231.1, 
    102215.9,
  102100.4, 102115.9, 102132.9, 102144, 102155.1, 102166.6, 102173.5, 
    102179.5, 102184.5, 102190.6, 102191.8, 102188.7, 102181.2, 102172, 
    102159.1,
  102033.4, 102094.9, 102156.1, 102197.9, 102233.5, 102256.9, 102266.2, 
    102276.4, 102276.1, 102275, 102268.8, 102262.8, 102255.4, 102244.4, 
    102232.3,
  102009.5, 102073.9, 102138.7, 102191.8, 102234.4, 102276.5, 102302.1, 
    102323.1, 102326.6, 102330.9, 102322.2, 102311.5, 102302, 102291.6, 
    102278.8,
  102001.1, 102072.3, 102132.9, 102191.7, 102238.9, 102280.9, 102312.9, 
    102336.4, 102353.4, 102356.7, 102351.8, 102347.9, 102343.5, 102334.4, 
    102321.8,
  101978.9, 102046.9, 102108.9, 102166.2, 102215.2, 102264.7, 102308.6, 
    102340.8, 102362.9, 102376.4, 102370.7, 102371.1, 102371.1, 102367.6, 
    102359.9,
  101966.2, 102031.4, 102088.1, 102147.6, 102192.6, 102237.6, 102279.8, 
    102322.9, 102347, 102369.7, 102383.8, 102387, 102381.1, 102376.7, 102369.4,
  101947, 102006.5, 102059.4, 102110.1, 102158.4, 102201.1, 102236.8, 
    102274.4, 102300.8, 102328.8, 102344.2, 102358.9, 102367.3, 102372.5, 
    102364.4,
  101930, 101981.6, 102032.6, 102078.7, 102122.1, 102160.7, 102190.9, 
    102220.8, 102244.9, 102265.9, 102288.4, 102312.1, 102327.5, 102334.2, 
    102334.5,
  101905.6, 101947.7, 101996, 102039.4, 102078, 102113.8, 102146.2, 102177.3, 
    102202.5, 102223.5, 102240.8, 102259.1, 102271.6, 102280, 102285.3,
  101881.6, 101919.2, 101957.8, 101994.2, 102029.6, 102060.2, 102089.3, 
    102113.1, 102138.3, 102162.9, 102184.3, 102198.8, 102210.9, 102221.4, 
    102226.1,
  101857.2, 101886.8, 101922.6, 101952.4, 101982.3, 102008.1, 102033.8, 
    102058.4, 102080.8, 102102, 102117.5, 102131.4, 102142.4, 102155.3, 
    102161.8,
  101161.2, 101147.6, 101162.7, 101184.4, 101217, 101250.7, 101287.3, 
    101326.1, 101362.3, 101397.6, 101439, 101480.3, 101524.4, 101573.6, 
    101618.9,
  101195.3, 101207.3, 101228, 101249.1, 101280.5, 101320.7, 101365.9, 
    101413.9, 101457.2, 101504.1, 101547.6, 101589.6, 101632.9, 101668.9, 
    101701.9,
  101234.5, 101254.5, 101280.7, 101306.8, 101343, 101381.3, 101432.2, 
    101484.3, 101533.5, 101580.4, 101620.9, 101661.5, 101705.1, 101745.7, 
    101786.9,
  101270.9, 101300.1, 101331.8, 101362.1, 101397.8, 101435.4, 101484.4, 
    101536.6, 101589.9, 101643.2, 101688.3, 101727.5, 101769.5, 101810.8, 
    101846.2,
  101298.3, 101334.1, 101376.8, 101412.4, 101450.3, 101486.6, 101528.8, 
    101576, 101622.9, 101675.5, 101722.5, 101766.6, 101805.1, 101844.1, 
    101882.4,
  101319.2, 101360.8, 101408.8, 101448.2, 101488.8, 101527.6, 101565.6, 
    101605.3, 101642.8, 101690.4, 101737.4, 101781.9, 101821.2, 101858.9, 
    101888.9,
  101336.6, 101380, 101428.9, 101470.8, 101512.7, 101551.5, 101589.8, 
    101626.1, 101662.6, 101697.7, 101740.4, 101780.4, 101815.3, 101852.5, 
    101886.9,
  101351.2, 101395.2, 101443.4, 101485.8, 101526.6, 101565.8, 101601.1, 
    101635, 101670.6, 101705, 101743.8, 101780.3, 101810.2, 101840.6, 101865.9,
  101366.8, 101407.9, 101452.5, 101491, 101529, 101567.6, 101601.9, 101635.3, 
    101669.7, 101702.7, 101734.7, 101769.9, 101799.2, 101822.4, 101847.8,
  101385.7, 101420.2, 101461.3, 101492.6, 101528.1, 101565.9, 101598.6, 
    101631.2, 101664.8, 101693.7, 101721.4, 101752.6, 101781.5, 101803.4, 
    101823,
  101689.1, 101707.1, 101717, 101720.2, 101716.8, 101710.1, 101694.2, 
    101675.7, 101646.3, 101619.7, 101582.5, 101539.5, 101501.1, 101464.5, 
    101439.1,
  101666.4, 101679.1, 101690.4, 101700.2, 101700.4, 101694.6, 101680.7, 
    101659.5, 101633.5, 101603.9, 101571.1, 101536.9, 101509.5, 101482.3, 
    101460.7,
  101631.1, 101655, 101667.8, 101674.8, 101677.1, 101673.1, 101661.7, 
    101644.6, 101623.2, 101597.8, 101565.3, 101537.5, 101516.8, 101497.4, 
    101480,
  101587.3, 101611.9, 101627.7, 101636.3, 101644.8, 101643.1, 101635, 
    101624.9, 101608.3, 101589.5, 101567.4, 101549.7, 101535.4, 101526.1, 
    101517.8,
  101551.4, 101582, 101593.7, 101610.9, 101616.5, 101625.4, 101624.1, 
    101620.5, 101612.8, 101603.1, 101587.6, 101575.6, 101564.2, 101556.6, 
    101554,
  101503.6, 101548.1, 101559, 101576.7, 101586.2, 101598.9, 101605.2, 
    101612.5, 101614.3, 101608.7, 101605.5, 101600.8, 101598, 101594.5, 
    101594.5,
  101500.8, 101535.6, 101551.7, 101569.5, 101589.3, 101600.4, 101609.6, 
    101619, 101622.1, 101625.9, 101627.3, 101627.5, 101630.5, 101638.3, 
    101650.1,
  101520.6, 101535, 101570.6, 101582.8, 101597.8, 101612.4, 101622.6, 
    101632.5, 101641.2, 101649.6, 101657.5, 101666, 101678.8, 101691.9, 
    101710.7,
  101524.2, 101536.1, 101579, 101591.2, 101610.2, 101624.4, 101639.1, 
    101652.5, 101667, 101679.2, 101689.4, 101703.6, 101716.9, 101733.1, 
    101750.8,
  101520, 101536.3, 101577, 101589.6, 101609, 101626.3, 101644.7, 101660.4, 
    101674.2, 101689.9, 101706.3, 101722.5, 101739.9, 101755.3, 101773.1,
  101750.5, 101758.3, 101771, 101787.4, 101799, 101811.8, 101820.2, 101829.4, 
    101839, 101851.9, 101868.7, 101885.3, 101910, 101923.8, 101945.1,
  101754.2, 101774.6, 101793.8, 101809.7, 101823.5, 101838.9, 101853, 
    101865.6, 101876, 101889.7, 101907.8, 101927.1, 101941.2, 101952.4, 101967,
  101758.5, 101788.4, 101812.9, 101834, 101853.3, 101869.4, 101886.7, 
    101900.6, 101909.1, 101920.8, 101936.1, 101952.4, 101961.3, 101976.9, 
    101988,
  101765.8, 101793.3, 101822.1, 101846.3, 101867, 101884.8, 101900.5, 
    101917.2, 101924.5, 101936.2, 101949.8, 101967.5, 101981.5, 101987.5, 
    101990,
  101772.7, 101797.4, 101827.2, 101852.3, 101877.5, 101899.5, 101918.1, 
    101935.6, 101949.8, 101958.2, 101965.8, 101973, 101987.3, 101990.5, 
    102005.8,
  101776.8, 101800.7, 101834.6, 101855.2, 101880.8, 101899.1, 101918.9, 
    101936.2, 101945.8, 101956.9, 101970.4, 101978.6, 101984.6, 101987.2, 
    101992.3,
  101776.8, 101801.5, 101835.3, 101858.5, 101884.9, 101903.7, 101923.8, 
    101937.7, 101951, 101963.4, 101974, 101981, 101989.4, 101999.4, 102007.7,
  101775, 101797.4, 101827.9, 101849.8, 101873.3, 101895.5, 101915.8, 
    101936.9, 101955, 101969.1, 101983.5, 102000.1, 102015.3, 102025.7, 
    102043.5,
  101768.5, 101788.6, 101811.6, 101831.9, 101855.7, 101877.5, 101899.4, 
    101918.3, 101939.7, 101958.1, 101978.4, 101994.2, 102010.4, 102025.1, 
    102044.3,
  101755.8, 101768.8, 101790.9, 101807.4, 101827.1, 101845, 101864.5, 101885, 
    101905.9, 101924, 101941.9, 101959.5, 101979.1, 102000.1, 102024.5,
  102514.9, 102524.5, 102520.8, 102518.7, 102508.3, 102497.2, 102473.5, 
    102449, 102418, 102386.3, 102351.1, 102310.5, 102271.3, 102227, 102181.8,
  102458.6, 102463.5, 102470.3, 102472.5, 102470.7, 102462.8, 102448.6, 
    102430, 102407.1, 102383.4, 102352.8, 102318.4, 102283.2, 102245.5, 
    102208.5,
  102397.4, 102401.2, 102406.2, 102417.1, 102420.8, 102419.5, 102410.8, 
    102400.1, 102383.5, 102363.5, 102338.7, 102311.6, 102283.3, 102254.4, 
    102223.4,
  102322.4, 102334.5, 102338.5, 102348, 102353.1, 102360.4, 102362, 102355.8, 
    102345.9, 102331.4, 102310.4, 102286.1, 102263.5, 102239.4, 102212.8,
  102224.9, 102248.2, 102254.9, 102271.6, 102284.3, 102293.4, 102298.5, 
    102301.9, 102297.3, 102292.3, 102281.4, 102267.5, 102251.2, 102231.2, 
    102208.9,
  102177.3, 102182.3, 102192.1, 102200.9, 102217.1, 102228.9, 102241.3, 
    102245.6, 102253.1, 102253, 102247.1, 102241.4, 102229.5, 102215.4, 
    102196.7,
  102151.3, 102143.8, 102155.3, 102159.1, 102169.9, 102173.6, 102183, 
    102189.8, 102197.8, 102200.9, 102204.3, 102201.8, 102200.1, 102194.3, 
    102185.7,
  102118.8, 102111, 102124.6, 102124.2, 102134.2, 102135.7, 102147.1, 
    102152.2, 102160, 102164.4, 102168.5, 102173.5, 102177.9, 102184.2, 
    102186.8,
  102079.2, 102073.1, 102082.2, 102081.5, 102088.7, 102094.4, 102106.2, 
    102115.5, 102128, 102135.1, 102148.3, 102157.3, 102165.5, 102173.3, 102179,
  102021.2, 102014.1, 102016.1, 102017.6, 102023.9, 102034.2, 102044.8, 
    102057.4, 102072.4, 102081.8, 102093.4, 102103.3, 102116.6, 102130.1, 
    102143,
  102310.9, 102313.9, 102300.1, 102285.7, 102260.3, 102232.2, 102199.3, 
    102160.1, 102117.6, 102072.8, 102025, 101975.8, 101926.4, 101878.6, 
    101833.2,
  102288.7, 102306.5, 102302.2, 102295.7, 102282, 102262.9, 102238.1, 
    102209.8, 102178.8, 102147.8, 102112.7, 102074.3, 102035.1, 101998.8, 
    101960.9,
  102232, 102251.4, 102260.8, 102272.3, 102263.2, 102263.5, 102248.5, 
    102230.5, 102210.3, 102190, 102163.5, 102132.7, 102101.2, 102070.4, 
    102042.5,
  102159.5, 102185.4, 102198, 102215.5, 102227, 102235.5, 102228.3, 102224.4, 
    102211.7, 102194.4, 102179.4, 102163.2, 102143.2, 102122.4, 102098.9,
  102085, 102111.5, 102127.9, 102148.5, 102163.2, 102176.9, 102182.7, 
    102183.2, 102179.5, 102174.4, 102165.1, 102151.4, 102135.1, 102122.5, 
    102106,
  102035, 102046.3, 102061.1, 102080.3, 102099.5, 102115.2, 102120.1, 
    102126.8, 102130.9, 102135.3, 102130.5, 102127.3, 102122.3, 102116.6, 
    102104.4,
  102002.4, 101997.8, 102008.9, 102016.9, 102029, 102037.3, 102046.5, 
    102052.5, 102051.1, 102050.7, 102053.2, 102056, 102058.2, 102057.2, 
    102052.3,
  101959, 101957.3, 101967, 101972.1, 101982, 101988.7, 101995.3, 101999.2, 
    102007, 102011.7, 102014.9, 102021.4, 102025.9, 102031, 102031.6,
  101903.7, 101914.5, 101913.7, 101921.1, 101928.4, 101939.5, 101949.2, 
    101958, 101966.6, 101972.7, 101982.8, 101990.7, 101999.2, 102010, 102018,
  101839, 101844.9, 101841.5, 101849.5, 101854.6, 101863.1, 101876.3, 
    101886.4, 101903.2, 101914.8, 101926.7, 101943, 101955, 101964.4, 101969.9,
  102347.1, 102324.5, 102294.3, 102263, 102225.1, 102177.7, 102122.4, 
    102062.8, 101993, 101921.4, 101849.1, 101772.8, 101690.9, 101603.9, 
    101512.5,
  102336.9, 102332.5, 102312.4, 102283.1, 102252.9, 102218.2, 102170.5, 
    102119.8, 102060.8, 101997.5, 101928.7, 101855.9, 101781.5, 101703.8, 
    101623,
  102319.8, 102323.2, 102305.9, 102292.4, 102270.9, 102238.7, 102203.4, 
    102162.2, 102114.6, 102061.3, 102001.2, 101933.6, 101865.3, 101793.3, 
    101718.4,
  102287.1, 102296.1, 102287.9, 102288.2, 102269.9, 102250.9, 102224.2, 
    102192, 102151, 102106.3, 102056, 102000, 101935.3, 101871.1, 101802.8,
  102227, 102245.7, 102252.1, 102255.4, 102251.2, 102242.3, 102225.3, 102204, 
    102172.6, 102135.2, 102094.1, 102046.8, 101989.9, 101934.5, 101874.3,
  102146.4, 102182.2, 102194.4, 102209.4, 102216.2, 102215.4, 102205, 
    102190.6, 102170.2, 102144.2, 102110, 102073, 102030.2, 101980.6, 101929.1,
  102073.6, 102104.6, 102121.3, 102141, 102152.1, 102160.5, 102159.2, 102157, 
    102141.5, 102122.2, 102103.3, 102077.4, 102039.9, 102002.5, 101958.7,
  101988.7, 102018.3, 102034.8, 102057, 102069.3, 102080.4, 102086.9, 
    102085.5, 102085.9, 102077.9, 102063.9, 102043.6, 102025.8, 101998.6, 
    101966.3,
  101907.1, 101932.9, 101945.5, 101960.7, 101973.5, 101989.7, 102006.3, 
    102019.1, 102027, 102019, 102016.1, 102006.9, 101992.8, 101975.9, 101955.9,
  101817.4, 101836.2, 101844.3, 101860.9, 101873.3, 101890.3, 101909, 
    101930.4, 101943.5, 101952.5, 101953.5, 101951.7, 101946.3, 101934.2, 
    101923.1,
  102224.9, 102264.7, 102288.4, 102303, 102313.5, 102312.7, 102304.9, 
    102290.1, 102271.9, 102245.2, 102204, 102154.8, 102097.8, 102032.2, 
    101960.1,
  102203.1, 102241.1, 102269.2, 102289.5, 102305, 102313.7, 102317.1, 
    102310.3, 102300.9, 102280.4, 102251.9, 102212, 102163.4, 102109.9, 
    102048.2,
  102160.2, 102194.4, 102234.3, 102268.8, 102291.4, 102306, 102315.4, 
    102316.8, 102314.9, 102305.5, 102285.8, 102255.7, 102220, 102173.9, 
    102119.7,
  102119.9, 102156.3, 102188.8, 102227.3, 102255.3, 102278.3, 102297.3, 
    102308.7, 102314.2, 102313.9, 102302.2, 102283.4, 102256.9, 102223.1, 
    102182.1,
  102064.5, 102110.6, 102143.9, 102176.8, 102213.2, 102245.9, 102267, 
    102285.1, 102296.5, 102301.7, 102302.7, 102294.8, 102276.8, 102253.5, 
    102221.4,
  102003.4, 102048.4, 102086.2, 102121.9, 102155, 102191, 102217.9, 102246.2, 
    102264.6, 102278.2, 102281.5, 102282.3, 102277.9, 102262.8, 102238.9,
  101933.4, 101975.1, 102015, 102055.5, 102092.7, 102127.1, 102160.1, 
    102188.5, 102213.2, 102234, 102248.5, 102257.4, 102256.1, 102252.3, 
    102241.9,
  101853.7, 101889.9, 101924.6, 101968.9, 102014.4, 102058.6, 102096.9, 
    102131.9, 102162.5, 102187, 102205.7, 102216.8, 102221.5, 102223.3, 
    102220.1,
  101765.6, 101800.1, 101827.8, 101864.7, 101903.9, 101956.4, 102005.4, 
    102053.7, 102092.4, 102128.3, 102151, 102168, 102180.5, 102185.1, 102186.8,
  101667.9, 101699.9, 101715.3, 101752.7, 101794.2, 101841.2, 101886.3, 
    101943.4, 101995.8, 102047.8, 102086.7, 102115, 102131.1, 102141.3, 
    102146.6,
  101923.4, 101983.7, 102042.1, 102099.3, 102155.4, 102210.2, 102259.4, 
    102304.5, 102339.6, 102374.8, 102396, 102411.8, 102421.4, 102428.7, 
    102432.9,
  101892.5, 101945.5, 102003.9, 102057.1, 102116.1, 102172.8, 102226.2, 
    102277.7, 102327.1, 102371.4, 102398.9, 102419.1, 102433.2, 102447.5, 
    102458.4,
  101852.6, 101902.8, 101959.8, 102011.1, 102070.8, 102129, 102189.1, 
    102241.7, 102289.3, 102337.7, 102375.3, 102403.8, 102430.7, 102453.3, 
    102475.4,
  101805.2, 101847.7, 101899.2, 101940.7, 101994.1, 102045.8, 102109.8, 
    102165.6, 102228, 102279.2, 102328.5, 102369.9, 102407.6, 102440.1, 
    102466.5,
  101745.6, 101776.6, 101825.2, 101862.3, 101913.9, 101961, 102027.6, 
    102096.2, 102166.7, 102227.7, 102278.2, 102324.7, 102366.6, 102403.9, 
    102436.2,
  101674.1, 101693.3, 101736.5, 101766.5, 101805.4, 101863.7, 101929.1, 
    101996, 102062.4, 102131.7, 102198.5, 102247.2, 102291.6, 102332.1, 
    102376.1,
  101586.4, 101592.1, 101630.2, 101640.4, 101689.9, 101758.3, 101822, 
    101899.4, 101964.3, 102018.1, 102081.2, 102142.9, 102205.7, 102255.2, 
    102302.6,
  101491.3, 101480.3, 101496.4, 101492.7, 101565, 101636, 101709.9, 101772.4, 
    101848.4, 101901.6, 101970, 102032, 102096.1, 102154.2, 102209,
  101379.5, 101356.3, 101346.7, 101349.9, 101467, 101524.7, 101585.8, 
    101634.1, 101726.6, 101778.2, 101847.5, 101914.4, 101985.5, 102049.1, 
    102108,
  101269.5, 101243.2, 101211.3, 101273.9, 101355.6, 101403.5, 101424, 
    101493.3, 101592.8, 101647.8, 101732.7, 101808.8, 101887.1, 101953.2, 
    102016.9,
  101540.8, 101592.1, 101652.3, 101721.8, 101796.5, 101867.9, 101945.5, 
    102018.4, 102088.6, 102156.7, 102211, 102267, 102320.1, 102368.1, 102412,
  101451.3, 101476.3, 101525.8, 101593.5, 101674.3, 101758.9, 101847.7, 
    101928.5, 102007, 102082.7, 102151.6, 102214.3, 102277.2, 102335.8, 102394,
  101311.6, 101316.2, 101360.4, 101449.1, 101548, 101633.7, 101736.7, 
    101834.6, 101926.1, 102013.2, 102090.7, 102160.2, 102226, 102290.6, 
    102353.5,
  101175, 101146, 101166, 101255.8, 101378.5, 101489.2, 101611.5, 101725.8, 
    101828.8, 101923, 102007.3, 102080, 102153.3, 102227.8, 102296.5,
  101035, 100954.3, 100921.4, 100997.9, 101171.7, 101309.7, 101463.8, 
    101602.2, 101727.5, 101829.9, 101920.8, 101997.9, 102071.6, 102147.8, 
    102221.9,
  100936.4, 100782.1, 100691.6, 100725.9, 100916.5, 101110.1, 101292.5, 
    101458.3, 101604.5, 101722.4, 101824.8, 101912.4, 101990.4, 102065.9, 
    102140,
  100861.4, 100678.4, 100494.6, 100491.7, 100678.5, 100925.1, 101130.1, 
    101321.2, 101488.3, 101627.8, 101744.5, 101840, 101922, 101994.5, 102067.8,
  100815.2, 100642.8, 100372.9, 100327.3, 100485, 100738.3, 100978.9, 
    101190.3, 101373.9, 101533, 101669, 101776.3, 101868.7, 101940.7, 102013,
  100808.6, 100651.8, 100352.6, 100246.5, 100345, 100614.8, 100855.8, 
    101077.9, 101279.9, 101451.8, 101598.4, 101713.9, 101815.2, 101895.5, 
    101972.7,
  100845.8, 100689, 100408.6, 100242.1, 100307.9, 100548.5, 100770, 101000.1, 
    101206.2, 101383.1, 101537.9, 101661.2, 101772.9, 101861.3, 101937.8,
  100931.3, 100761.3, 100624.4, 100603.9, 100670.5, 100792.5, 100946.8, 
    101117.1, 101287.8, 101453.6, 101599.9, 101727.5, 101836.9, 101932.8, 
    102014.3,
  100872.2, 100731, 100589.5, 100621.8, 100712.8, 100867.6, 101028.4, 
    101194.5, 101352.3, 101497.3, 101630.4, 101746, 101853.1, 101944.9, 
    102024.9,
  100900.4, 100847, 100663.7, 100682.5, 100750.9, 100897.6, 101049.4, 
    101205.2, 101361.5, 101505.5, 101645.3, 101765.3, 101874.6, 101965.3, 
    102045.7,
  100967.6, 100899.1, 100737, 100736.7, 100826.2, 100966.1, 101122.8, 
    101269.2, 101416.4, 101547.6, 101675.5, 101788, 101893.6, 101986.2, 
    102069.7,
  101072.4, 100989, 100880.7, 100857.9, 100915.3, 101041.2, 101181.3, 
    101319.2, 101455.3, 101579.2, 101701.6, 101808.5, 101910.3, 102005.6, 
    102092.4,
  101162.2, 101100.2, 101029.5, 101005.3, 101045.5, 101152.5, 101271.3, 
    101395.7, 101516.6, 101631, 101739.6, 101832.4, 101928.6, 102021.8, 
    102111.4,
  101237.7, 101212.3, 101179.9, 101162.9, 101191.4, 101269.6, 101362, 101467, 
    101570.4, 101674.2, 101776.5, 101861.1, 101948.7, 102039.5, 102128.1,
  101301.4, 101303.8, 101304.3, 101300.5, 101332.3, 101390.5, 101454.7, 
    101538.8, 101629.3, 101721.4, 101810, 101887.5, 101973.6, 102057.2, 
    102142.9,
  101350.3, 101367.9, 101397.3, 101414.3, 101438.7, 101478.2, 101531.7, 
    101601.4, 101679, 101756.3, 101835, 101908.5, 101996.8, 102073.8, 102156.9,
  101398.2, 101424.8, 101460.5, 101485, 101511.7, 101551.2, 101596.2, 
    101657.9, 101720.1, 101786.4, 101855.2, 101924.2, 102014.1, 102092.1, 
    102172.8,
  101977.2, 101958.3, 101934.7, 101914.4, 101888.1, 101855.6, 101815.6, 
    101761.8, 101703.7, 101649.6, 101606.9, 101575.4, 101554.6, 101540.6, 
    101529.4,
  101967.4, 101965.1, 101962.1, 101954.9, 101941.6, 101925, 101898.2, 
    101862.6, 101826.6, 101792.8, 101763.8, 101737.4, 101717.7, 101703.3, 
    101691,
  101935.2, 101949, 101950.5, 101957.7, 101959.7, 101962, 101954.1, 101941.5, 
    101923.9, 101902.2, 101881.1, 101863.2, 101850.5, 101840.4, 101831.8,
  101901.7, 101937.6, 101954.3, 101973.9, 101990.4, 102005.6, 102014.5, 
    102014.6, 102008.2, 101997.5, 101986.5, 101979.6, 101972.2, 101967.1, 
    101963.3,
  101880.4, 101932.8, 101964.7, 101994.4, 102025.6, 102050.7, 102065, 
    102079.1, 102080.5, 102077.9, 102073.6, 102071.3, 102068, 102066.1, 
    102064.5,
  101875.4, 101920.6, 101969.2, 102006.3, 102044.8, 102075.3, 102101.9, 
    102124.3, 102138.8, 102138.1, 102140.9, 102146, 102148.9, 102148.4, 
    102152.7,
  101869.7, 101912, 101973.4, 102015.9, 102059.2, 102094.4, 102122.5, 
    102144.5, 102162.1, 102171.4, 102179.4, 102186.9, 102190.1, 102195.4, 
    102208.4,
  101868.6, 101910.3, 101978.8, 102021.6, 102068, 102103.5, 102135.1, 
    102163.1, 102180.9, 102196.3, 102204.2, 102216.2, 102228, 102242.8, 
    102260.9,
  101867.7, 101911.3, 101975.2, 102014.5, 102061.5, 102092, 102128, 102157.9, 
    102176.5, 102199.1, 102204.2, 102221.1, 102245.1, 102270.3, 102302.6,
  101863.2, 101912.9, 101969.6, 102007, 102049.3, 102083.3, 102118, 102140.5, 
    102160, 102180.2, 102200.5, 102238.3, 102275.4, 102305.1, 102338.5,
  102578.6, 102611.4, 102646.5, 102659.8, 102671.3, 102685.9, 102692.1, 
    102693.9, 102687.7, 102679, 102661.6, 102637.2, 102604.2, 102569.8, 
    102533.3,
  102505, 102554.5, 102591.6, 102618.9, 102640.3, 102647.2, 102652.6, 
    102662.1, 102664.7, 102660.1, 102654.8, 102635.2, 102612.6, 102583.5, 
    102551.2,
  102443.1, 102491.5, 102523.1, 102558, 102581.4, 102603.2, 102616.3, 
    102621.8, 102629.2, 102633.1, 102631, 102625.8, 102611.3, 102590.7, 
    102563.8,
  102360.2, 102415.2, 102462.8, 102502.9, 102528.6, 102552.2, 102567.1, 
    102583.1, 102590, 102599.5, 102603.1, 102596.8, 102588.2, 102578.4, 
    102557.4,
  102307.6, 102354.3, 102386.4, 102419.9, 102459.1, 102488.5, 102510.1, 
    102522.8, 102534.9, 102548.7, 102563, 102573, 102572, 102566.1, 102551,
  102283.1, 102308.1, 102352.8, 102385.4, 102418.9, 102442, 102460.5, 
    102479.6, 102511.4, 102528.3, 102529.2, 102536.5, 102542.6, 102541.9, 
    102539.7,
  102268, 102293.3, 102345.1, 102370.7, 102403.5, 102428.2, 102454.5, 
    102469.6, 102486, 102501, 102515.1, 102521, 102530.4, 102528.2, 102521.1,
  102232.6, 102263.7, 102301, 102332.2, 102363.7, 102392.5, 102421.1, 
    102448.3, 102471, 102480.2, 102493.1, 102510.8, 102515.5, 102516.4, 
    102514.5,
  102208.6, 102243.3, 102268.6, 102292.1, 102316.3, 102339.5, 102363.4, 
    102386.1, 102410, 102433, 102447.5, 102468.3, 102484.4, 102487.3, 102491.5,
  102173.1, 102205.6, 102227.8, 102244.5, 102268.6, 102291.9, 102317.8, 
    102339.5, 102365.9, 102392.3, 102417, 102442.1, 102459.1, 102474.9, 102485,
  102364.6, 102433.9, 102505.1, 102586.7, 102652, 102691.4, 102739.4, 
    102795.5, 102866.2, 102915.6, 102958.2, 102985.7, 103011.4, 103030.2, 
    103039.2,
  102332.3, 102395.8, 102472.5, 102537.3, 102599.1, 102667.8, 102729.7, 
    102773.7, 102811.6, 102849.2, 102913.4, 102955.6, 102994.5, 103019.7, 
    103050.5,
  102312.3, 102369.3, 102432.5, 102494, 102547.4, 102594.7, 102649.1, 
    102712.8, 102770.1, 102816, 102861.2, 102913.7, 102958.8, 103003.2, 
    103031.1,
  102296, 102348.9, 102400.4, 102448.2, 102503.2, 102555.8, 102597.3, 
    102636.3, 102680.4, 102743.7, 102801.6, 102846.5, 102894.5, 102939.2, 
    102982.5,
  102276.8, 102326.4, 102378.7, 102423.5, 102464.4, 102496.8, 102533.8, 
    102578, 102620.3, 102659, 102712.3, 102780.5, 102843.8, 102887.5, 102918.4,
  102255.1, 102303.7, 102350.4, 102394.4, 102439.9, 102474.4, 102505.9, 
    102529.2, 102559.9, 102591.3, 102636.7, 102685.4, 102735.2, 102802.6, 
    102868.1,
  102227.4, 102274.5, 102316, 102357.5, 102398.6, 102438.5, 102472, 102508.5, 
    102536.1, 102557.6, 102583, 102626.4, 102682.6, 102725.3, 102770.6,
  102205.1, 102244.9, 102284.4, 102323.5, 102361.5, 102395.8, 102430.1, 
    102464.1, 102497.2, 102532.7, 102556.8, 102577.6, 102609.4, 102652.6, 
    102707.3,
  102180, 102215.8, 102250.5, 102288.4, 102325.7, 102362.1, 102394.2, 
    102427.1, 102456.8, 102486, 102515.1, 102547.1, 102573.8, 102602.1, 
    102638.4,
  102145.9, 102181.2, 102213.4, 102248.1, 102285.5, 102318.6, 102358.1, 
    102390.6, 102428, 102456.7, 102485.1, 102506.6, 102532.4, 102555, 102582.6,
  101954.6, 102026.1, 102104.1, 102172.7, 102240.8, 102303.1, 102355.9, 
    102421, 102493.8, 102565.6, 102647.1, 102737, 102817.4, 102890.4, 102953.3,
  101988.1, 102058.5, 102133, 102196.4, 102258.2, 102314.9, 102372.5, 
    102434.2, 102491.6, 102557.4, 102632.7, 102718.3, 102807.4, 102889.1, 
    102962.7,
  102011.1, 102080.4, 102154.4, 102219.7, 102280.4, 102336, 102391.9, 
    102437.3, 102492, 102549.5, 102616, 102706.4, 102797.9, 102882, 102946.6,
  102031.6, 102098.7, 102170.5, 102232.8, 102289.9, 102345.9, 102395.9, 
    102443.5, 102496.9, 102547.3, 102603.7, 102679.9, 102767.5, 102857.5, 
    102930.9,
  102044.4, 102109, 102179.4, 102242.5, 102299.5, 102350.1, 102400.1, 
    102446.3, 102489.6, 102539.7, 102597.7, 102662.3, 102740.1, 102819.8, 
    102901.4,
  102053.2, 102117.7, 102178.5, 102241.1, 102296.8, 102344, 102392.4, 
    102438.3, 102482.9, 102526, 102578.3, 102637, 102710.3, 102789.7, 102864.8,
  102057.6, 102116.7, 102173.9, 102230.4, 102286.1, 102334.4, 102377.4, 
    102419.3, 102461.8, 102508.9, 102555.7, 102615.1, 102673.4, 102740.7, 
    102814.1,
  102057.4, 102109.6, 102163, 102209.8, 102258.9, 102304.4, 102354.4, 
    102398.7, 102439.2, 102479, 102524.6, 102577.3, 102635.8, 102695, 102757.3,
  102051.2, 102095.8, 102145.3, 102189.7, 102236.2, 102277.9, 102319.9, 
    102362, 102407.7, 102446.7, 102487.6, 102528.2, 102581.8, 102637.6, 
    102696.9,
  102037.2, 102076.7, 102119.3, 102160.2, 102203.3, 102243.6, 102285.9, 
    102325.6, 102367.1, 102406.7, 102447.8, 102483.7, 102528.2, 102574.7, 
    102629.2,
  101747.7, 101747.5, 101764.1, 101790.8, 101820.5, 101853.1, 101890.4, 
    101928.1, 101970.8, 102023.3, 102082.5, 102140.7, 102204.1, 102267.8, 
    102334.9,
  101786.4, 101809.6, 101842.6, 101874.1, 101909.6, 101953.2, 101998.1, 
    102037.9, 102082.8, 102131.7, 102181.9, 102237.8, 102299.2, 102367.1, 
    102437.8,
  101823.8, 101855.6, 101887.8, 101929.5, 101972.4, 102013.9, 102054, 
    102092.7, 102142.4, 102197, 102251.5, 102310.5, 102374, 102441.9, 102511.1,
  101855.1, 101892.9, 101931.7, 101979.7, 102026, 102066.5, 102107.1, 
    102149.2, 102196.6, 102250.6, 102301.7, 102360.8, 102425.5, 102496.3, 
    102562.3,
  101874.6, 101916.9, 101964, 102009.6, 102053.4, 102091.2, 102134.4, 
    102178.2, 102224.6, 102276.9, 102332.9, 102394.1, 102460.8, 102526.6, 
    102593.7,
  101894.2, 101936, 101985.7, 102027, 102073.1, 102112.7, 102155.9, 102196.7, 
    102244, 102292.5, 102348.2, 102409.1, 102470.7, 102536.5, 102609.2,
  101908.8, 101940.2, 101993.2, 102031.4, 102076.3, 102117.4, 102157.6, 
    102200.7, 102244.7, 102293.3, 102346.5, 102405.5, 102466.4, 102531.4, 
    102597.4,
  101912.1, 101940.7, 101992.6, 102028.3, 102072, 102111.1, 102152, 102195.1, 
    102237.4, 102280.1, 102331.4, 102384.7, 102443.3, 102505.6, 102569.9,
  101901, 101933.1, 101978.8, 102013.8, 102054.7, 102095.1, 102133.1, 
    102174.1, 102215.2, 102258.2, 102302.8, 102351.3, 102407.1, 102464.1, 
    102525.8,
  101884.7, 101921.8, 101956.9, 101992.4, 102027, 102065.9, 102104.6, 
    102142.4, 102184.1, 102223.8, 102267.7, 102310.6, 102361.2, 102413.1, 
    102469,
  102867, 102840.7, 102805.4, 102766.2, 102731.1, 102696.3, 102656.5, 
    102619.6, 102581.1, 102542.2, 102502, 102463, 102427.8, 102395.1, 102369,
  102811.9, 102781, 102748.2, 102716.7, 102683.6, 102646.9, 102611.3, 
    102577.1, 102540, 102507.2, 102476.8, 102448.6, 102425.6, 102407.5, 
    102395.4,
  102750.5, 102725.3, 102687.8, 102648.6, 102615.3, 102585.9, 102556.3, 
    102524, 102496.2, 102472.4, 102450.4, 102430.4, 102415.3, 102406.9, 
    102404.1,
  102681.4, 102647.1, 102610, 102576.5, 102549.4, 102523.9, 102495.9, 
    102474.7, 102447.8, 102428.2, 102412.4, 102405.8, 102406, 102413.4, 
    102427.7,
  102613.2, 102567.7, 102537.2, 102502.7, 102477.2, 102451.1, 102427.9, 
    102408.8, 102393.9, 102391, 102388.6, 102392.7, 102410.1, 102429.2, 
    102452.9,
  102536.6, 102492.5, 102458.6, 102435.8, 102413.3, 102388.3, 102375.7, 
    102370.2, 102365.8, 102370.1, 102384.8, 102411.2, 102424.8, 102447.2, 
    102483.7,
  102444.6, 102426.3, 102391.3, 102368.4, 102347, 102333.2, 102334.2, 
    102341.9, 102350.8, 102369.9, 102386.4, 102408, 102436.4, 102465.7, 
    102497.7,
  102376.3, 102359, 102321.6, 102308.5, 102300.6, 102311.3, 102310, 102325.1, 
    102340.7, 102358.9, 102381.3, 102407.5, 102435.3, 102463.8, 102499.5,
  102311.5, 102283.2, 102260.8, 102258.2, 102260.1, 102269, 102278.3, 
    102292.3, 102309.9, 102331.4, 102355.8, 102381.1, 102415.5, 102448.8, 
    102486.8,
  102242, 102218.5, 102209.1, 102206.9, 102210.6, 102215.6, 102224.3, 
    102237.1, 102257, 102280.8, 102311.9, 102342.2, 102380.7, 102416, 102459.1,
  102944.7, 102952, 102946.5, 102942.1, 102935, 102924.8, 102913.2, 102899.7, 
    102879.3, 102852.6, 102825.9, 102801.7, 102769, 102735, 102699,
  102904.9, 102908.1, 102907.4, 102912.6, 102910.7, 102904.4, 102895.1, 
    102881.8, 102864.2, 102843.5, 102822.9, 102799.9, 102773.1, 102744, 
    102718.4,
  102823.6, 102845.6, 102838.6, 102844.4, 102839.4, 102834.4, 102829, 
    102822.6, 102814.7, 102799.5, 102784.9, 102767.5, 102749.3, 102729.4, 
    102705.6,
  102749.8, 102770.4, 102764.1, 102768.1, 102765.1, 102767.5, 102761, 
    102756.2, 102749, 102739.6, 102726.4, 102713.2, 102699.6, 102687.8, 
    102673.5,
  102667.8, 102663.3, 102665.8, 102666, 102661.4, 102656.8, 102653.7, 
    102654.6, 102654, 102642.9, 102633.1, 102624.5, 102617.8, 102607.8, 
    102593.9,
  102585.5, 102559, 102568.9, 102565.9, 102563.3, 102558.5, 102556.4, 
    102547.9, 102541.8, 102539.6, 102541.6, 102538.8, 102535.9, 102535.3, 
    102544.2,
  102488.9, 102465, 102465.3, 102451.2, 102440.6, 102437.1, 102437.4, 
    102438.2, 102439.9, 102449.6, 102455.2, 102465.1, 102478.2, 102484.1, 
    102488.6,
  102392.1, 102374.7, 102354.2, 102350.7, 102350.4, 102357.7, 102364.4, 
    102370.7, 102381.3, 102392, 102410.5, 102423.4, 102436.4, 102466.8, 
    102489.4,
  102297.2, 102296.6, 102273, 102276.2, 102276.6, 102284, 102289.3, 102302.4, 
    102320.6, 102338.9, 102357, 102382.9, 102404, 102419.7, 102439.1,
  102223.2, 102224.4, 102198.8, 102200, 102195.7, 102203.6, 102217.4, 
    102233.8, 102253.2, 102277.6, 102302.4, 102328.9, 102354.1, 102384.6, 
    102406.1,
  102674.8, 102725.2, 102742.5, 102766.4, 102780, 102784.2, 102787.4, 102781, 
    102770.1, 102746.2, 102719.9, 102693.2, 102667.5, 102634.1, 102602.4,
  102640.9, 102674, 102696.2, 102715.7, 102731.4, 102744.8, 102756, 102757.4, 
    102749.5, 102728.8, 102715.2, 102691.3, 102664.8, 102634.6, 102605.6,
  102573.3, 102609.6, 102640.3, 102665, 102684.4, 102702.1, 102713.5, 
    102718.9, 102715.7, 102704.4, 102695.3, 102674.7, 102658, 102633.3, 
    102605.5,
  102486.8, 102531.4, 102565.5, 102602.1, 102627.3, 102638.9, 102650.7, 
    102654.3, 102661.7, 102659.2, 102655, 102643.3, 102634, 102612.7, 102593.3,
  102390.3, 102439.3, 102466, 102493.3, 102524.7, 102547.8, 102569, 102582.2, 
    102592.6, 102596.6, 102598.1, 102597.1, 102595.7, 102585.4, 102566.8,
  102301.8, 102349.4, 102380.7, 102416.8, 102439.1, 102462, 102479.2, 
    102497.2, 102508.6, 102521.3, 102526.9, 102529.7, 102529.9, 102528.1, 
    102523.6,
  102220.6, 102252.9, 102276.4, 102305.4, 102324.8, 102349, 102371.5, 
    102385.5, 102400.8, 102414, 102428.1, 102436.8, 102451.3, 102456.1, 
    102456.5,
  102149.7, 102174.9, 102190.3, 102212.4, 102232.2, 102251.8, 102268.5, 
    102284.7, 102301.6, 102314, 102330.8, 102346.6, 102348, 102362.1, 102366.7,
  102081.3, 102095.9, 102108.4, 102127.8, 102145.1, 102163.8, 102182.2, 
    102202.8, 102218.9, 102235, 102249.3, 102261.7, 102274.7, 102285.3, 
    102290.8,
  102019.4, 102026.9, 102039.2, 102056.1, 102074.4, 102097.2, 102114.8, 
    102136.8, 102156.9, 102175.2, 102191.9, 102204.8, 102216.9, 102225.1, 
    102230.7,
  102278.3, 102359.7, 102431.4, 102500.1, 102552.9, 102586.8, 102612.4, 
    102630.2, 102643.9, 102655.2, 102653.8, 102647.5, 102633.4, 102613, 
    102584.6,
  102203.6, 102294.7, 102363.2, 102425.9, 102481.9, 102530.2, 102562, 
    102586.3, 102606.9, 102612, 102618.7, 102611.5, 102597, 102578.6, 102556.4,
  102121, 102193.5, 102270.3, 102351.2, 102406.9, 102465.8, 102509.5, 
    102540.8, 102567.5, 102581.5, 102584.1, 102579.2, 102576.7, 102567.9, 
    102552.2,
  102079.6, 102150.4, 102191.3, 102264.6, 102325.4, 102378.7, 102422.7, 
    102463.7, 102502.6, 102528.8, 102544.6, 102551.8, 102549.8, 102547.2, 
    102536.9,
  101979, 102050.1, 102110.6, 102174.9, 102232, 102292.4, 102345.5, 102393.8, 
    102431.9, 102464.8, 102487.4, 102507.2, 102520, 102523.3, 102514.1,
  101895.6, 101968, 102035.5, 102087, 102139.1, 102190.6, 102239.7, 102292.6, 
    102340, 102380.9, 102415, 102437.7, 102462.3, 102472.1, 102475.8,
  101828.3, 101885.2, 101933.1, 101991, 102042.3, 102095.7, 102143.7, 
    102193.3, 102238.3, 102282.6, 102326, 102361.2, 102387.9, 102407.8, 
    102419.6,
  101785.9, 101825.3, 101871.7, 101917.6, 101957.7, 102001.8, 102049.7, 
    102093, 102142.6, 102191.3, 102235.6, 102269.8, 102302.6, 102325.6, 
    102348.1,
  101732.9, 101777, 101808.8, 101847.2, 101887.7, 101924.7, 101961.5, 
    102003.4, 102042.6, 102086.6, 102130.1, 102173.4, 102210.2, 102241.2, 
    102264.8,
  101688.8, 101714.4, 101743.2, 101778.2, 101814.5, 101856, 101892.9, 101930, 
    101969.3, 102006.4, 102040.6, 102075.8, 102108.6, 102141.5, 102167.9,
  102143.7, 102247.6, 102298.2, 102355, 102400.5, 102443, 102476.6, 102505.7, 
    102538, 102561.2, 102567.2, 102551.8, 102533.4, 102510.8, 102470.1,
  102023.3, 102131.8, 102211.5, 102286.6, 102337.2, 102383.3, 102418.3, 
    102449.5, 102476.1, 102501.2, 102524.7, 102526.2, 102519.1, 102486.9, 
    102454.2,
  101929.3, 102014, 102104.9, 102192.2, 102258.1, 102309.7, 102356.8, 
    102393.6, 102423, 102448.8, 102465.6, 102477.9, 102478.6, 102463.1, 
    102440.2,
  101812.3, 101893.5, 101980.7, 102061.6, 102147.6, 102217.8, 102270.8, 
    102319.7, 102360.6, 102392.8, 102414.8, 102424.9, 102433.2, 102429, 
    102422.6,
  101738.7, 101825, 101887.9, 101967.9, 102029.9, 102107.9, 102170.9, 
    102237.4, 102280.4, 102322.7, 102355.1, 102376.1, 102385.9, 102396.1, 
    102390.2,
  101606.7, 101704, 101782.7, 101867.6, 101922, 101997.6, 102049.3, 102121.6, 
    102177.1, 102227.9, 102265, 102297.2, 102323.5, 102340.4, 102349.5,
  101530.3, 101604, 101686.9, 101759.1, 101825.8, 101895.9, 101959.5, 102019, 
    102077.9, 102135.1, 102181.3, 102220, 102246.4, 102267.2, 102277.2,
  101455.9, 101517.5, 101568.8, 101644.5, 101715.4, 101785.6, 101857.1, 
    101918.8, 101981.4, 102036.4, 102088.8, 102130.1, 102164.4, 102191.7, 
    102211,
  101409.4, 101446, 101501.9, 101550.9, 101616.5, 101681.2, 101752.4, 
    101810.7, 101879.1, 101938.6, 101993.1, 102043.2, 102082, 102110.8, 
    102136.1,
  101372.8, 101394, 101428.7, 101468.6, 101527.2, 101583.1, 101648.1, 
    101713.5, 101775.9, 101838.1, 101897.5, 101945.8, 101993.5, 102028.2, 
    102057.7,
  102217.8, 102280.2, 102326.7, 102378.9, 102419.8, 102458.2, 102483.6, 
    102509.2, 102524.5, 102539.3, 102536.6, 102531.5, 102516.4, 102502.3, 
    102483,
  102094.4, 102166.4, 102214.5, 102279.3, 102330.1, 102385, 102426.5, 
    102459.8, 102480.9, 102494.9, 102501.8, 102509.3, 102507.3, 102505.1, 
    102491.1,
  101979.5, 102055.9, 102114.1, 102180.1, 102235.2, 102290.3, 102338.6, 
    102379.9, 102410.7, 102430.4, 102445, 102455.5, 102461.5, 102468.3, 
    102461.4,
  101844.9, 101895.9, 101963.9, 102048, 102115.8, 102180.6, 102238, 102287.6, 
    102325.7, 102352, 102374.6, 102391.4, 102405.7, 102412.2, 102407.1,
  101712.7, 101790.4, 101829.2, 101897.8, 101973.8, 102053.1, 102121, 
    102179.5, 102230.5, 102267.2, 102292.9, 102314.1, 102329.2, 102341.7, 
    102346.3,
  101604.3, 101738.1, 101765.6, 101811.3, 101848.4, 101913.1, 101982.3, 
    102058.2, 102112.8, 102162.3, 102197.9, 102228.8, 102251.7, 102274.6, 
    102288.8,
  101416.5, 101528.2, 101614.5, 101683.4, 101707.3, 101773.9, 101835.6, 
    101917, 101984.1, 102049.6, 102091.7, 102126.9, 102155.4, 102181.8, 
    102208.2,
  101248.8, 101328.5, 101422.4, 101519.7, 101569.5, 101633.4, 101693.6, 
    101783.4, 101853.9, 101923.7, 101977.8, 102023, 102057, 102088.9, 102117.4,
  101122.1, 101166, 101235.7, 101328.8, 101412.2, 101483.8, 101547.2, 
    101637.1, 101725.9, 101799.3, 101866, 101915.2, 101958.7, 101993.1, 
    102029.1,
  101109.4, 101098.8, 101130.5, 101180.8, 101261.3, 101341.7, 101418, 
    101489.9, 101587.4, 101664.7, 101740.6, 101802.3, 101851.3, 101889.3, 
    101928.6,
  101992.5, 102031.1, 102059.5, 102088.6, 102111.9, 102135.8, 102151.1, 
    102167.4, 102171.9, 102177.6, 102175.5, 102170.5, 102174.2, 102175.8, 
    102173.4,
  101915.9, 101943.8, 101974.8, 102014.1, 102046.5, 102082.4, 102112, 
    102138.8, 102152.4, 102165.9, 102170.6, 102172.4, 102174.6, 102176.2, 
    102172.2,
  101820.2, 101855.6, 101882, 101917.2, 101950.5, 101987.2, 102015.4, 
    102048.1, 102076.6, 102102.2, 102121.2, 102142.7, 102154.2, 102173.5, 
    102179,
  101721.5, 101749.9, 101775.9, 101810.5, 101843.9, 101882.2, 101924.8, 
    101962.2, 101992.7, 102020.9, 102045.6, 102071.6, 102095.8, 102121.5, 
    102134.8,
  101614.9, 101630, 101653.2, 101685.6, 101719.9, 101755.2, 101782.2, 
    101819.3, 101859.4, 101899.5, 101937.8, 101972.9, 102004, 102035.4, 
    102057.7,
  101510.7, 101515.4, 101519.3, 101552.1, 101582.6, 101629.9, 101684, 
    101725.8, 101761.7, 101794, 101824.7, 101858.9, 101891.8, 101925.9, 
    101956.7,
  101409.3, 101426, 101431.5, 101446.9, 101450.2, 101450, 101471.8, 101508.7, 
    101562.9, 101619.1, 101672.9, 101721.2, 101766.7, 101808.8, 101845.7,
  101302.5, 101316.6, 101335.5, 101376.9, 101387.1, 101402.2, 101426.7, 
    101455.2, 101491.3, 101530.4, 101561, 101601, 101640.9, 101686.6, 101724,
  101147.5, 101161, 101186.1, 101206.4, 101211.4, 101225.3, 101240.4, 
    101277.1, 101310.6, 101354.6, 101399.9, 101447.8, 101492.2, 101535, 
    101573.7,
  101019.9, 101015.4, 101025.9, 101026.1, 101048.7, 101086, 101097.9, 
    101123.6, 101160.2, 101203.7, 101240.9, 101285.7, 101328.1, 101375.6, 
    101419.3,
  101428.4, 101410.5, 101381.4, 101358.3, 101327.4, 101294.8, 101265.3, 
    101235, 101205.6, 101187.4, 101166.5, 101147, 101136.9, 101136.5, 101144.4,
  101446, 101427.3, 101403, 101387.8, 101367, 101350.1, 101322.3, 101296.7, 
    101265.6, 101249.6, 101220.3, 101197.7, 101184.6, 101175.3, 101169.5,
  101445.4, 101424, 101398.8, 101379, 101355.4, 101333, 101306.7, 101286.3, 
    101258.4, 101233.8, 101211.4, 101195.4, 101178.9, 101165.4, 101154.5,
  101432.5, 101414.9, 101395.4, 101374.9, 101346.2, 101322.1, 101292.5, 
    101265.5, 101236.9, 101206.8, 101175.7, 101150.3, 101128.1, 101106.2, 
    101097.1,
  101412.9, 101394.9, 101370.7, 101343, 101314, 101280.7, 101242.6, 101204.2, 
    101168.4, 101135.5, 101110, 101083.4, 101054.8, 101035.7, 101015.5,
  101389.9, 101367.1, 101344.2, 101311.1, 101276.7, 101240.5, 101201.1, 
    101163.2, 101124.2, 101079.6, 101030.7, 100980, 100937, 100906.2, 100880.2,
  101361.4, 101332.5, 101307.3, 101269.9, 101230.6, 101183.7, 101135.3, 
    101078.9, 101015.3, 100953.9, 100907.3, 100872.8, 100848.6, 100829.5, 
    100810.5,
  101337.9, 101305.1, 101273.6, 101228.2, 101181, 101129.5, 101079, 101022.7, 
    100981, 100934.7, 100893.7, 100840.2, 100772.5, 100714.1, 100670.7,
  101303.1, 101269.9, 101225.8, 101177.5, 101127.9, 101077.4, 101027.4, 
    100968.6, 100905.9, 100835.2, 100765.6, 100696.4, 100644, 100585.8, 
    100532.7,
  101272.9, 101236.4, 101193.1, 101142.6, 101090.5, 101035.7, 100977, 
    100904.6, 100830.8, 100750.4, 100671, 100599.3, 100523.2, 100470.9, 100423,
  101558.3, 101496.6, 101430.9, 101361.1, 101285, 101202.9, 101114, 101017.9, 
    100919.6, 100814.4, 100712.5, 100611.7, 100504.8, 100400, 100299.3,
  101575.2, 101516.1, 101456.3, 101390.9, 101318.8, 101241.3, 101158.9, 
    101073.9, 100983, 100889.9, 100792.9, 100695.1, 100597.8, 100501, 100409.1,
  101597.5, 101544.8, 101489.9, 101428.6, 101359.8, 101288.5, 101211.9, 
    101133.5, 101051.3, 100961.5, 100872.7, 100780.3, 100688.5, 100594.9, 
    100503.7,
  101619.2, 101567.7, 101515.9, 101460.3, 101401, 101333.5, 101263.5, 
    101192.5, 101117.1, 101036.5, 100953.7, 100868.1, 100781.1, 100694.8, 
    100608.9,
  101640.1, 101593.3, 101545.6, 101494.5, 101438.9, 101378.9, 101316, 
    101247.3, 101177.3, 101101.8, 101023.8, 100945.5, 100865.8, 100785.3, 
    100705.6,
  101657.2, 101617.1, 101574.2, 101525, 101474.3, 101418.7, 101363.5, 101301, 
    101234.4, 101164.8, 101093.1, 101019.1, 100945, 100868.4, 100793.9,
  101670.2, 101633.2, 101597, 101552.1, 101503.8, 101453.3, 101401.7, 
    101344.7, 101281.7, 101215.9, 101147.9, 101079.8, 101009, 100937.2, 
    100865.7,
  101679.1, 101646.6, 101616.1, 101573.7, 101531.5, 101481.5, 101432.5, 
    101379.3, 101321.9, 101260.9, 101197.2, 101131.6, 101063.3, 100994.4, 
    100926.3,
  101677.9, 101652.8, 101626.9, 101589, 101550.1, 101504.4, 101458.5, 
    101407.7, 101354.7, 101298.3, 101236.8, 101172.3, 101108.9, 101044.9, 
    100979.7,
  101667.6, 101650.1, 101630.7, 101596.7, 101561.1, 101518.1, 101475.2, 
    101427, 101377.6, 101324, 101269.1, 101209, 101148.4, 101089.2, 101029.3,
  102300.4, 102348, 102383.5, 102410.3, 102421.3, 102424.8, 102428.8, 
    102430.5, 102423.3, 102402, 102367.9, 102323.3, 102283.4, 102226.5, 
    102161.3,
  102272.8, 102320.8, 102360.9, 102399.8, 102420.4, 102428.8, 102427.3, 
    102432.8, 102429.6, 102413.8, 102386.9, 102351.8, 102308.5, 102260.9, 
    102202.8,
  102241, 102291.4, 102326.2, 102367.2, 102395.3, 102418.7, 102427.4, 
    102427.6, 102428.1, 102422.3, 102401.8, 102372.3, 102336.7, 102295.5, 
    102241.7,
  102207.6, 102258, 102293.9, 102331.4, 102366.7, 102390.3, 102402.4, 
    102410.9, 102416.2, 102413, 102399.6, 102375.6, 102344.7, 102313.8, 
    102270.4,
  102173.6, 102224.4, 102257.9, 102296.6, 102325.5, 102350.5, 102365, 
    102388.4, 102392.6, 102392.2, 102383.2, 102372, 102351.8, 102328.3, 
    102287.4,
  102137.9, 102181, 102220.5, 102257, 102285.9, 102310.7, 102329.8, 102351.8, 
    102361, 102365.3, 102361.3, 102348.2, 102332.9, 102313.2, 102287.4,
  102109.8, 102141.4, 102171.8, 102200.4, 102228.6, 102256.8, 102276.8, 
    102296.5, 102312.2, 102322.1, 102322.9, 102319.8, 102311.4, 102297.3, 
    102273.8,
  102075.1, 102103.1, 102128.4, 102151.7, 102178.4, 102197.2, 102221.9, 
    102237.3, 102252.9, 102267.7, 102273.8, 102277.2, 102274.3, 102256, 
    102242.1,
  102049, 102067.2, 102088.6, 102103.4, 102121.9, 102140, 102161.1, 102178.6, 
    102191.2, 102206.2, 102213.9, 102223.4, 102227.3, 102219.7, 102204.4,
  102026.2, 102037.7, 102047.1, 102057.9, 102067.5, 102078.7, 102094.3, 
    102112.8, 102128, 102137.8, 102144.9, 102159.7, 102166.1, 102161.1, 
    102154.9,
  101582.2, 101675.1, 101769.2, 101859.7, 101946.9, 102030.9, 102110.5, 
    102192.1, 102272.9, 102348.3, 102415.9, 102479.2, 102539, 102600.4, 102648,
  101597.1, 101687.2, 101783, 101875, 101963.3, 102046.2, 102129.1, 102212.1, 
    102295.6, 102371.8, 102446.1, 102513.1, 102580.1, 102644.4, 102699.6,
  101612.6, 101699.8, 101796.5, 101886.7, 101974.2, 102057, 102140.4, 
    102221.1, 102304.5, 102384.9, 102462.5, 102537.2, 102608, 102672.9, 
    102734.9,
  101619, 101705.7, 101798.8, 101885.9, 101971.8, 102052, 102134.4, 102216.3, 
    102299.5, 102378.8, 102458.1, 102537.2, 102610.1, 102683, 102747.6,
  101628.5, 101709.5, 101800.5, 101881.3, 101967, 102044.2, 102121, 102199.7, 
    102279.5, 102360.5, 102439.5, 102515, 102593, 102670.6, 102742.6,
  101631.1, 101708.1, 101794.6, 101867.4, 101948.5, 102023.9, 102101, 
    102178.2, 102252.9, 102330.3, 102409.7, 102486.6, 102559.8, 102636.3, 
    102711.9,
  101640, 101709, 101784.7, 101854.3, 101925.7, 102000.4, 102076.4, 102146.6, 
    102220.4, 102295.7, 102371.1, 102449.8, 102524.9, 102601.2, 102674.6,
  101642.9, 101706.2, 101770.6, 101828.9, 101896.5, 101964.2, 102035.4, 
    102109.8, 102181, 102253, 102327.8, 102403.8, 102474.6, 102551.3, 102627.3,
  101649.5, 101699.9, 101755.1, 101805.3, 101859.6, 101922, 101986.2, 
    102055.1, 102128.7, 102202.4, 102273.9, 102350.5, 102424.7, 102496.7, 
    102566.9,
  101650.3, 101688.8, 101733.1, 101774.8, 101817.7, 101869.5, 101926, 
    101991.3, 102061.5, 102135.9, 102212.8, 102284.8, 102358.4, 102434, 
    102504.7,
  100935.2, 100951.2, 100976.1, 101006.3, 101042.3, 101090.3, 101149.1, 
    101214.3, 101289.9, 101371, 101458.4, 101548.5, 101646.4, 101747.9, 
    101852.2,
  100956.8, 100995.6, 101040, 101084.9, 101140.5, 101200.9, 101263.3, 
    101328.5, 101398.7, 101473.3, 101554.7, 101641.6, 101735.8, 101833, 
    101934.5,
  100993.9, 101041, 101090.9, 101141.8, 101195.4, 101256, 101320.1, 101391.1, 
    101465.3, 101542.8, 101626.9, 101715.7, 101807.5, 101903.4, 102004.2,
  101025.6, 101079.9, 101139.2, 101193.5, 101249, 101309.5, 101370.3, 
    101443.1, 101516.2, 101593.4, 101679.4, 101764, 101855.5, 101951.9, 
    102048.4,
  101064.2, 101116.8, 101179.5, 101228, 101278.7, 101333.7, 101396.3, 
    101467.8, 101542.4, 101621.9, 101708.3, 101796.4, 101888.6, 101983.3, 
    102081,
  101097.9, 101146.4, 101205.3, 101249.7, 101299, 101353.4, 101411.8, 
    101480.2, 101553.8, 101631.9, 101718.2, 101806.9, 101900.7, 101997, 
    102093.2,
  101128.1, 101169.7, 101225.4, 101265.1, 101310.3, 101357, 101411.1, 
    101477.3, 101551, 101628.9, 101714.4, 101807.7, 101901.5, 101996.7, 
    102093.8,
  101150.1, 101190.1, 101235.4, 101268.1, 101308.8, 101354.8, 101403.5, 
    101466.4, 101537.1, 101615.5, 101700.4, 101792.2, 101885.4, 101981.9, 
    102074.6,
  101171.5, 101207.1, 101243.3, 101271.5, 101306.2, 101343.2, 101387.7, 
    101443.6, 101514.2, 101591.5, 101675.6, 101766.8, 101856.4, 101952.6, 
    102048.3,
  101185.8, 101219, 101243.9, 101265, 101292.5, 101328.2, 101372.1, 101420.1, 
    101483.7, 101561.1, 101638.9, 101724.6, 101817.9, 101912.6, 102015.8,
  102260.2, 102182.1, 102123, 102060.7, 102000.7, 101937.8, 101866.9, 
    101791.9, 101709.1, 101626.2, 101534.7, 101439.2, 101355.3, 101273, 
    101199.5,
  102195.4, 102130.2, 102079, 102014.1, 101951.4, 101887.9, 101818.2, 
    101748.9, 101678.6, 101606.5, 101530.8, 101444.7, 101359.3, 101278.6, 
    101209,
  102156.9, 102102.7, 102047.1, 101981, 101922.7, 101862.4, 101799.5, 
    101731.1, 101660.8, 101591.1, 101514.8, 101444.1, 101370, 101301.1, 
    101241.3,
  102103.5, 102052.4, 101990.8, 101931.6, 101878.6, 101820.2, 101759.7, 
    101700.2, 101639.9, 101577.3, 101512.7, 101441.9, 101375.2, 101313.4, 
    101260.9,
  102038, 101991.5, 101931.3, 101882.3, 101829.9, 101776.2, 101720.7, 
    101665.7, 101607.3, 101548.6, 101491.4, 101435.6, 101380.5, 101330.8, 
    101288.6,
  101971.6, 101942.3, 101891.3, 101842.6, 101793.5, 101743.2, 101691.1, 
    101641, 101589.5, 101538.3, 101488.3, 101438, 101391, 101346.8, 101311.7,
  101911.7, 101880, 101833.5, 101789.3, 101744.5, 101697.1, 101649.2, 
    101603.1, 101555.1, 101508.9, 101467.2, 101431.8, 101397.1, 101364.9, 
    101339.2,
  101851.4, 101810.5, 101777, 101741, 101700.5, 101657.1, 101610, 101569.4, 
    101527.3, 101492.6, 101459.9, 101428.9, 101399.9, 101374.3, 101358.1,
  101776.2, 101737.1, 101707.1, 101671.6, 101632.7, 101598.1, 101561.8, 
    101527.6, 101494.2, 101463.9, 101439.2, 101419.7, 101403.1, 101387.8, 
    101381.9,
  101680.5, 101653, 101625.6, 101597.9, 101569.9, 101541.2, 101511, 101482.2, 
    101451.7, 101432.6, 101416.4, 101404, 101397.7, 101393.6, 101398.3,
  102729.5, 102721.2, 102713.7, 102700.7, 102686.8, 102664.6, 102634.2, 
    102590.8, 102544.3, 102492.3, 102427.3, 102359.9, 102282.8, 102203.7, 
    102127.6,
  102673.2, 102683.6, 102676.2, 102674.6, 102669.5, 102651.7, 102629.7, 
    102596.8, 102552.7, 102507.2, 102446, 102381, 102311.9, 102238.2, 102162.2,
  102634.7, 102646.6, 102642.6, 102642.8, 102637, 102628.8, 102609, 102576.6, 
    102544.9, 102500.3, 102446.1, 102389.8, 102325.6, 102258.6, 102188.2,
  102585.2, 102600, 102597.2, 102600.6, 102598.4, 102597.7, 102578.8, 102556, 
    102519.4, 102474.9, 102434.4, 102380.3, 102324.6, 102260.7, 102197.4,
  102535.8, 102546.4, 102549.8, 102558, 102554.4, 102551.3, 102535, 102513.1, 
    102477.4, 102443.6, 102403.1, 102353.6, 102301.8, 102244.5, 102187.6,
  102480.8, 102489.5, 102491.5, 102493.6, 102490.4, 102489.5, 102477.6, 
    102458.2, 102427.9, 102396.4, 102351, 102305.2, 102255.8, 102205.9, 
    102158.7,
  102394, 102413.7, 102417.1, 102420.5, 102413.8, 102407.4, 102393.4, 102376, 
    102349.3, 102320.5, 102283.8, 102245.1, 102199.2, 102157.5, 102113.5,
  102319.1, 102329.8, 102323.1, 102326.3, 102322.5, 102316.6, 102307.2, 
    102288.2, 102266.9, 102238.7, 102205.8, 102167.4, 102125, 102086.7, 
    102049.6,
  102230.8, 102242.2, 102241, 102240.6, 102235.1, 102225.9, 102212, 102196.6, 
    102178.9, 102152.1, 102122.6, 102091.5, 102060.2, 102026.9, 101989.6,
  102169.8, 102152.9, 102151.6, 102148.7, 102144.9, 102138.1, 102129.9, 
    102116, 102095.3, 102071.8, 102048, 102012.7, 101976, 101940.5, 101908.6,
  102346.2, 102419.4, 102473.5, 102502.6, 102510.9, 102517, 102518.2, 102508, 
    102494.1, 102479.7, 102452.5, 102416.3, 102379.7, 102335.1, 102282,
  102291.3, 102362.9, 102436.3, 102496.7, 102529, 102530.4, 102529.8, 
    102520.6, 102507.1, 102489.1, 102469.2, 102439.6, 102402.1, 102359.4, 
    102310.4,
  102251.4, 102321.6, 102391.2, 102453.3, 102501, 102537.2, 102553.9, 
    102547.8, 102532.5, 102510.8, 102486.9, 102459.1, 102424.7, 102385.6, 
    102342.6,
  102192.5, 102264, 102337.3, 102405.7, 102457.9, 102499.9, 102530.5, 
    102550.2, 102555.4, 102530.5, 102504.6, 102475.8, 102446.8, 102411.9, 
    102371.1,
  102137.6, 102216.7, 102284.6, 102349.9, 102407.3, 102458.2, 102496.2, 
    102527.7, 102543.1, 102538.8, 102524.3, 102496.1, 102467.3, 102434.2, 
    102397.1,
  102064.4, 102144, 102213.5, 102280.4, 102334.5, 102386.5, 102434.5, 
    102473.5, 102507.8, 102522.5, 102522.2, 102506.7, 102483.7, 102452.8, 
    102418.9,
  102016.9, 102084, 102158, 102222.1, 102272, 102313.3, 102363.1, 102403.8, 
    102440.3, 102472, 102488.1, 102490.1, 102475, 102457.4, 102429.3,
  101953.2, 102035.5, 102094.3, 102153.6, 102198.6, 102237.8, 102280.2, 
    102327.3, 102364.8, 102398.2, 102426.4, 102442.4, 102445.3, 102433.9, 
    102422.2,
  101870.2, 101985.8, 102050.7, 102123.7, 102156.9, 102187.1, 102216.9, 
    102262, 102297.8, 102329.7, 102355.5, 102374.9, 102388.6, 102394.7, 
    102392.1,
  101767.8, 101872.7, 101943.1, 102024.4, 102078, 102119.8, 102151.9, 
    102193.9, 102231.2, 102262.5, 102287.9, 102308.7, 102325.5, 102337.6, 
    102341.7,
  101458.6, 101541.8, 101625.1, 101711, 101800.9, 101889.8, 101975.9, 
    102052.8, 102126.5, 102187.5, 102245.3, 102295.6, 102339.6, 102389.4, 
    102416.7,
  101471.3, 101549.6, 101624.2, 101706.1, 101792.1, 101884.5, 101970.6, 
    102052, 102122.6, 102190.1, 102246.7, 102296.7, 102337.7, 102384.7, 
    102419.6,
  101471.1, 101554.6, 101633.9, 101713.8, 101796.4, 101881.9, 101969.6, 
    102049.7, 102127.8, 102191.4, 102247.1, 102296.2, 102339.9, 102377.9, 
    102412.9,
  101453.1, 101533.6, 101611, 101687.2, 101767.3, 101856.6, 101944.4, 
    102029.1, 102109.6, 102180.7, 102242, 102290.5, 102334.2, 102376.3, 
    102409.1,
  101429.2, 101505.4, 101583.4, 101661.8, 101738, 101823.2, 101914.6, 101999, 
    102082.6, 102163.1, 102231.9, 102281.1, 102322.1, 102361.5, 102396.8,
  101407.7, 101478.6, 101560, 101639, 101710.4, 101784.8, 101870.7, 101959.7, 
    102044.9, 102127.4, 102204.6, 102266.5, 102307.8, 102341, 102373.6,
  101366, 101449.1, 101528.8, 101613.2, 101686.2, 101752.1, 101825.5, 
    101914.8, 101999.6, 102084.2, 102164.2, 102232.9, 102285.5, 102327.6, 
    102348.9,
  101300.7, 101410, 101484.6, 101577.3, 101658.4, 101730.3, 101790.6, 
    101870.1, 101958.3, 102039, 102118.9, 102192, 102249.3, 102297.7, 102326.5,
  101250.9, 101366.1, 101433.5, 101523.2, 101600, 101681.1, 101745.8, 
    101824.7, 101906.1, 101988.6, 102064.4, 102137.5, 102204, 102255.9, 
    102292.8,
  101223.9, 101319.8, 101414.8, 101488.1, 101565.1, 101643.5, 101709.8, 
    101772.8, 101851.4, 101933.8, 102006.5, 102080.5, 102146, 102205.4, 
    102251.5,
  101223.4, 101156.6, 101095.2, 101047.6, 101007, 100976.1, 100957.9, 
    100961.2, 100985.9, 101041.2, 101121.6, 101211.9, 101309.4, 101411.9, 
    101515,
  101245.4, 101185.8, 101134.7, 101089.2, 101049.1, 101019.4, 100999.4, 
    101003.9, 101033.4, 101088.6, 101161.7, 101245.7, 101342.2, 101449.8, 
    101555.7,
  101271.9, 101212.5, 101162.7, 101118.3, 101081.1, 101057.5, 101044.5, 
    101051.3, 101074.6, 101129.8, 101203, 101299.9, 101402.5, 101502.4, 
    101601.3,
  101290.2, 101240.4, 101194, 101145.9, 101110.9, 101082.6, 101070.5, 
    101080.2, 101114.5, 101176.3, 101256.8, 101347.3, 101442.8, 101537.2, 
    101632.2,
  101294.8, 101255.3, 101212.9, 101167.4, 101134.8, 101104.5, 101093.7, 
    101106.1, 101141.7, 101199.5, 101278.9, 101376.8, 101477.8, 101568.7, 
    101655.5,
  101279.8, 101248.2, 101221.6, 101186.3, 101157.7, 101133.4, 101125.1, 
    101137.5, 101172.6, 101228.8, 101308.9, 101405.9, 101501.7, 101589.4, 
    101675.6,
  101260.9, 101231, 101211, 101184.6, 101170.7, 101157.1, 101156.7, 101172.2, 
    101203.3, 101247.1, 101319.4, 101414.9, 101511.7, 101608.4, 101691.3,
  101223, 101192.6, 101179.3, 101159.3, 101160.6, 101160.6, 101160.4, 
    101174.3, 101207.3, 101265.2, 101338.4, 101426.7, 101516.1, 101612.2, 
    101700.9,
  101191.9, 101166.1, 101142.3, 101116.2, 101113.6, 101118.1, 101138.5, 
    101170.8, 101218.3, 101277, 101341.8, 101425.3, 101513.8, 101607.8, 101698,
  101154.3, 101128.9, 101105, 101075, 101071.4, 101074.9, 101099.1, 101141.3, 
    101186.1, 101245.5, 101336.1, 101429.8, 101517.1, 101600.9, 101680.7,
  100899.3, 100867, 100859.2, 100846, 100841.2, 100838.5, 100834, 100832.2, 
    100833.4, 100836.8, 100837.9, 100831.2, 100817.9, 100806.2, 100799.1,
  100974.1, 100954.6, 100951.5, 100945.5, 100935.9, 100924.6, 100919.5, 
    100914.8, 100907.6, 100894, 100878.7, 100865.9, 100850.1, 100836.3, 
    100831.3,
  101033.8, 101021.5, 101016.2, 101010, 100995, 100981.4, 100969.8, 100968.2, 
    100958.2, 100945.4, 100928.8, 100914, 100887.9, 100878.1, 100865.4,
  101068.3, 101067.7, 101072.6, 101061.8, 101042.4, 101032.6, 101016.9, 
    101001.8, 100986, 100963.2, 100945.7, 100919.5, 100907.3, 100884.1, 100879,
  101093, 101094.9, 101089.7, 101076, 101060.4, 101042.9, 101029.5, 101017.1, 
    101000.7, 100986.5, 100952, 100934.4, 100899.9, 100889.2, 100942,
  101086.4, 101089.4, 101084.8, 101078.4, 101068.1, 101049.9, 101032.2, 
    101012.5, 100989.5, 100949.4, 100928, 100908.2, 100882.6, 100937, 101005.3,
  101074.9, 101078.9, 101073.2, 101067.3, 101049.7, 101037.3, 101020.7, 
    100995.9, 100969.7, 100950.5, 100936.4, 100878.3, 100890.9, 100951.1, 
    101043.7,
  101039.2, 101051.1, 101047.2, 101043.8, 101031.2, 101010.7, 100983.4, 
    100957.1, 100929.6, 100902.2, 100854.1, 100848, 100877.2, 100928, 101004,
  101013.4, 101022.5, 101014.9, 101009, 100994.4, 100987.6, 100957.2, 
    100928.8, 100890.2, 100844.3, 100819.9, 100817.6, 100814.5, 100848.1, 
    100945.6,
  100976.2, 100971.3, 100974.9, 100976.1, 100957.2, 100942.3, 100909.8, 
    100873.8, 100830.6, 100778.1, 100752.7, 100737.6, 100762.3, 100806.5, 
    100909.8,
  101210.8, 101159.3, 101081.8, 101015.3, 100943.9, 100868.9, 100797.9, 
    100735.5, 100683.6, 100638.8, 100600.3, 100566.4, 100540.8, 100516.2, 
    100478.5,
  101223.4, 101174.8, 101108.4, 101049, 100977.7, 100909, 100842.3, 100782.2, 
    100729.1, 100689.2, 100653.4, 100617, 100578.9, 100540.8, 100526.5,
  101251.5, 101189, 101135.2, 101090.2, 101030.3, 100971.1, 100908.4, 
    100846.3, 100791.1, 100739, 100695.4, 100658.2, 100622.7, 100593.2, 
    100543.5,
  101270, 101201.1, 101151, 101103.6, 101060.8, 101010.4, 100956.8, 100902.7, 
    100848.1, 100793.9, 100747.8, 100701.3, 100661, 100619.7, 100552.9,
  101288.6, 101223.4, 101178.1, 101128.6, 101084.7, 101039.2, 100996.3, 
    100948.5, 100898, 100844.6, 100795.5, 100747.9, 100707.2, 100651.1, 
    100599.5,
  101303, 101241, 101194.6, 101143.1, 101100.4, 101054.1, 101016.4, 100978.2, 
    100931.3, 100883.8, 100835, 100788.7, 100736.4, 100678.4, 100618.3,
  101305.4, 101248.2, 101203.1, 101153.9, 101107.8, 101060.9, 101023.3, 
    100982, 100946.6, 100905.9, 100864.6, 100828.5, 100775.4, 100703.7, 
    100642.1,
  101295.7, 101240.5, 101197.4, 101149.2, 101102.1, 101056.7, 101019.2, 
    100986.7, 100954.8, 100919.6, 100883.3, 100835.5, 100779, 100729.8, 
    100686.9,
  101276.3, 101221.9, 101176.2, 101123, 101074.2, 101027.3, 100986.6, 
    100949.3, 100923, 100896.3, 100868.2, 100852.2, 100833.7, 100782.6, 
    100722.7,
  101237.9, 101181.4, 101137.3, 101082.1, 101033.3, 100997.2, 100972.6, 
    100961.8, 100950.3, 100937.4, 100926.3, 100895.3, 100859.9, 100830, 100794,
  102590.3, 102544.4, 102494.8, 102443.3, 102374.5, 102302.4, 102227, 
    102147.8, 102063.7, 101973.4, 101882.3, 101783, 101687.2, 101587.6, 
    101501.4,
  102600.2, 102557.9, 102508.5, 102458.9, 102393, 102325.6, 102251, 102171.8, 
    102089.4, 101997.3, 101903.3, 101807.6, 101710.3, 101614, 101516.6,
  102604.8, 102561.3, 102516.3, 102471.7, 102408.8, 102345.3, 102272.4, 
    102192.2, 102109.4, 102018.4, 101924.1, 101825.5, 101726.8, 101626.7, 
    101530.6,
  102599.3, 102560, 102519, 102476.3, 102416.4, 102354.8, 102283.7, 102204.3, 
    102122.5, 102035.2, 101943, 101846.6, 101747.1, 101645.6, 101543.3,
  102592.7, 102555.9, 102516.8, 102473, 102419.6, 102360, 102290.9, 102212, 
    102131.5, 102047.9, 101957.7, 101860.1, 101760.2, 101656.3, 101551.9,
  102580, 102544.8, 102505.5, 102462.8, 102412.2, 102354.9, 102286.6, 
    102210.9, 102135, 102053.4, 101962.3, 101865, 101764.2, 101663.3, 101559.8,
  102562.4, 102528.8, 102490.3, 102446.9, 102398.8, 102342.3, 102275.8, 
    102205.7, 102128.7, 102048.6, 101958.7, 101863.6, 101761.2, 101657.6, 
    101553.4,
  102539.5, 102507, 102467.1, 102423.6, 102375.1, 102316.9, 102254.2, 
    102185.1, 102112, 102033.5, 101944.7, 101850.4, 101748.5, 101645, 101538.1,
  102513.1, 102482.4, 102441, 102397.2, 102346.8, 102290.4, 102226.8, 
    102161.2, 102091.9, 102012.4, 101921.9, 101831.3, 101729.7, 101628.4, 
    101521.5,
  102482.8, 102448.1, 102405.5, 102360.5, 102310.3, 102254.3, 102194, 
    102131.5, 102065.6, 101986, 101900.7, 101809.7, 101711, 101603.8, 101507.9,
  102960.8, 103012, 103050.6, 103082.6, 103091, 103092.1, 103072, 103049.4, 
    103025.3, 102990.1, 102946.7, 102896, 102844.3, 102790.4, 102738.7,
  102970.2, 103013.7, 103054, 103088.7, 103105.4, 103106, 103101.6, 103086.5, 
    103063.1, 103034.2, 102997, 102951, 102901.5, 102853.5, 102802.9,
  102958.9, 103001.8, 103044.1, 103072.8, 103095.7, 103110.2, 103113.5, 
    103111.4, 103095.3, 103072, 103037.7, 102998.4, 102951.2, 102905.5, 
    102856.5,
  102944.1, 102988.8, 103032.2, 103062.2, 103082.7, 103101.3, 103109.2, 
    103111.6, 103104.9, 103086.2, 103062.8, 103025.2, 102986.4, 102944.9, 
    102901.5,
  102922.8, 102962.7, 103000.8, 103033.4, 103059.4, 103080.6, 103091.7, 
    103096.3, 103092.7, 103083.3, 103066.8, 103042.5, 103010.7, 102973.8, 
    102935.1,
  102901.2, 102936.6, 102969, 102997.5, 103024, 103043.1, 103055.9, 103062.2, 
    103064.7, 103059.9, 103049.4, 103030.5, 103007.6, 102981.6, 102946.3,
  102872.5, 102903.1, 102933, 102958.5, 102979.7, 102996.9, 103008.6, 
    103016.4, 103021.9, 103020, 103013.9, 102999.2, 102979.7, 102956.5, 
    102926.5,
  102832.6, 102858.6, 102883.2, 102909.7, 102930.9, 102945.3, 102956.2, 
    102964.9, 102969.5, 102969.6, 102962.5, 102950.3, 102932.2, 102914.6, 
    102884.1,
  102791.9, 102809.9, 102829.2, 102848.3, 102866.5, 102883.3, 102895, 
    102907.9, 102912.3, 102911, 102903.2, 102889.4, 102876.6, 102856.4, 102828,
  102745, 102761.6, 102775.1, 102787.2, 102801.7, 102813.2, 102827, 102838.1, 
    102841.1, 102835, 102826, 102818.2, 102804.3, 102785.2, 102754.4,
  102529, 102601.1, 102673.7, 102733.4, 102795.8, 102850.6, 102903.7, 
    102952.1, 102994.1, 103025.6, 103051.1, 103067.9, 103085, 103096.5, 103104,
  102552.8, 102624.2, 102693.4, 102753.9, 102818.9, 102874.8, 102931.5, 
    102984.5, 103027.6, 103060.5, 103085.5, 103101.2, 103114.6, 103131.3, 
    103135.7,
  102551.8, 102623, 102694.2, 102758.5, 102823.2, 102882, 102939.9, 102993.7, 
    103040.4, 103080, 103100.4, 103121.1, 103128.5, 103142, 103152.8,
  102547.5, 102618.4, 102689.1, 102754.5, 102817.3, 102877.2, 102935, 
    102992.7, 103043.6, 103082.7, 103112.2, 103132.4, 103146.5, 103157.7, 
    103151.5,
  102535.2, 102602.8, 102667.5, 102729.8, 102793.1, 102856, 102916.5, 
    102973.9, 103028.7, 103071.4, 103107.7, 103132.7, 103145.5, 103155.6, 
    103148.2,
  102517.5, 102580.7, 102643.8, 102704.2, 102761.6, 102819.3, 102877.2, 
    102935, 102989.8, 103041.1, 103084.1, 103117.7, 103142.6, 103153.3, 
    103164.1,
  102494, 102549.8, 102605.4, 102665.3, 102720.2, 102778.8, 102833.3, 102889, 
    102941.9, 102990.4, 103036.5, 103074.1, 103106, 103133.4, 103150.8,
  102466.4, 102515.6, 102563.6, 102617.9, 102671.2, 102724.9, 102779.7, 
    102833, 102886, 102934.7, 102980.9, 103018.7, 103053.4, 103085.4, 103110.9,
  102432.3, 102473.1, 102513.9, 102559.8, 102609.3, 102662.1, 102715.5, 
    102767.5, 102819.8, 102865.7, 102908.8, 102948.8, 102988.9, 103020.8, 
    103048.4,
  102390.5, 102425.5, 102460.7, 102499.3, 102539.7, 102585.6, 102634.2, 
    102685.8, 102742.5, 102790.8, 102833.3, 102872.2, 102908.5, 102942, 
    102970.8,
  102126.8, 102169.7, 102225.1, 102275.8, 102325.8, 102377.1, 102433.5, 
    102480.4, 102530.9, 102579.5, 102621.5, 102661.1, 102695.7, 102727.6, 
    102756.9,
  102152.2, 102210, 102275.1, 102331.4, 102385.3, 102442, 102492.6, 102538.7, 
    102595.3, 102641, 102685.7, 102725.5, 102764.5, 102798.5, 102825.3,
  102156.3, 102215.6, 102283, 102342.4, 102403.8, 102469.9, 102527.7, 
    102579.4, 102632.3, 102677, 102719.9, 102764.9, 102806.1, 102845.9, 102872,
  102157.8, 102216.9, 102288.1, 102353.6, 102419.7, 102482.7, 102540, 
    102592.6, 102641.1, 102688.2, 102734, 102781.6, 102829, 102871.7, 102899.3,
  102143.6, 102204.7, 102279.3, 102342.2, 102408.9, 102473, 102533.7, 
    102583.3, 102632.3, 102679.6, 102729.5, 102775.1, 102824, 102871.1, 
    102911.7,
  102126.5, 102188.1, 102259.5, 102322.2, 102389.5, 102451.8, 102508.6, 
    102558.2, 102608.6, 102659.7, 102709.9, 102755.9, 102802.5, 102847.2, 
    102893,
  102104.5, 102162.8, 102228.8, 102291.5, 102354.9, 102415.6, 102476.6, 
    102525.7, 102574.6, 102623.8, 102676, 102722.3, 102769.2, 102812, 102857.5,
  102078.7, 102133.9, 102195.1, 102251.6, 102311.8, 102370.2, 102428.5, 
    102483.7, 102532, 102578.2, 102626.9, 102676, 102721.1, 102765, 102810.4,
  102047.9, 102098.4, 102154.9, 102208.6, 102263.2, 102316.7, 102373.4, 
    102427.7, 102478.8, 102524.4, 102569.1, 102615.5, 102658.5, 102700.7, 
    102741.2,
  102012.6, 102060.5, 102111, 102159.6, 102208.9, 102254.9, 102304.3, 
    102357.9, 102413, 102460.8, 102508.2, 102553.1, 102597.3, 102637.5, 
    102677.3,
  101774.3, 101761, 101885.1, 101959, 102032.8, 102083.9, 102135.6, 102181.4, 
    102225.2, 102260.3, 102291.6, 102318.1, 102339.8, 102358.9, 102381.2,
  101785.1, 101837, 101929.7, 101987.5, 102057.9, 102118.5, 102180.5, 
    102231.9, 102270.7, 102304.7, 102336.2, 102363.5, 102389.2, 102415.3, 
    102437.1,
  101790.6, 101868, 101936.2, 102001, 102071.4, 102128.9, 102185.1, 102236.1, 
    102279.9, 102317.9, 102356.8, 102387, 102415.7, 102447.1, 102474.8,
  101851, 101912.7, 101969, 102030.7, 102088.9, 102140, 102193.5, 102238, 
    102283.7, 102323.1, 102363.6, 102397.7, 102429.3, 102461.3, 102493.9,
  101880.3, 101928.7, 101978.8, 102031, 102085, 102133.7, 102186.4, 102228, 
    102270.4, 102318, 102354.1, 102393.9, 102425.8, 102461, 102494.1,
  101904.6, 101943, 101983.3, 102027.1, 102078.2, 102124.8, 102168.8, 
    102213.4, 102252.5, 102292.9, 102332.2, 102368.8, 102407.1, 102443.5, 
    102473.5,
  101905.9, 101938.5, 101976, 102014.4, 102058, 102096.9, 102140.8, 102184.2, 
    102224.1, 102264, 102302.8, 102340.4, 102375.8, 102409.1, 102437.9,
  101898.8, 101929.2, 101960.4, 101992.8, 102031.6, 102068.9, 102109.9, 
    102154.9, 102191.1, 102230.7, 102264.8, 102301.5, 102333.4, 102365.6, 
    102395.7,
  101878.6, 101912, 101938.4, 101966.9, 102001, 102036.8, 102073.9, 102116.2, 
    102154.1, 102190.3, 102226, 102260.9, 102290.1, 102318, 102340.4,
  101857.5, 101887.6, 101912.7, 101939.6, 101968.1, 102000.7, 102030.9, 
    102072.7, 102111.8, 102148.3, 102178.3, 102211.2, 102241, 102265.4, 
    102283.9,
  101665.1, 101469.9, 101299.2, 101138.8, 101014, 100940.1, 100952.8, 101093, 
    101249.1, 101420.5, 101548.2, 101645.9, 101728.5, 101796.3, 101850.6,
  101694.6, 101528.3, 101394.2, 101262.9, 101153.6, 101081.1, 101096.4, 
    101183, 101287, 101423, 101550.2, 101664.2, 101750.8, 101821.7, 101876.7,
  101774.5, 101631.2, 101511.2, 101382.8, 101278.1, 101200, 101189.7, 
    101235.1, 101328.3, 101437.8, 101550.6, 101654.9, 101736.2, 101807.3, 
    101865.2,
  101821.6, 101699.4, 101598.4, 101498.9, 101413.1, 101337.3, 101315.9, 
    101338.5, 101395.2, 101475.3, 101569.9, 101668.2, 101747.9, 101810.2, 
    101866.9,
  101859.2, 101764.4, 101673.6, 101591, 101515.7, 101449.2, 101420.5, 
    101418.7, 101457, 101519.8, 101595.5, 101676.8, 101740.8, 101797, 101848.7,
  101893.8, 101814, 101735.8, 101664.9, 101597.9, 101545.5, 101513, 101509.4, 
    101519.7, 101565.2, 101618.5, 101686.1, 101744.2, 101794.3, 101830.8,
  101914.6, 101853.4, 101781.1, 101720.6, 101661.3, 101613.5, 101581.9, 
    101565.3, 101571.5, 101600.3, 101642.7, 101698.2, 101745.7, 101786.1, 
    101816,
  101929, 101875.9, 101820.6, 101767, 101714.1, 101671.1, 101641, 101620.9, 
    101622.5, 101637.8, 101673.3, 101711.4, 101749.6, 101785.5, 101805.8,
  101927, 101880.5, 101841.2, 101793, 101747.4, 101710.8, 101680.4, 101661.7, 
    101662.9, 101674.9, 101697.9, 101729.8, 101755.9, 101780, 101800,
  101914.5, 101877.9, 101847.7, 101804.9, 101771.9, 101738.6, 101713.4, 
    101699.7, 101693.1, 101707.5, 101721.2, 101746.1, 101767, 101786.9, 
    101795.4,
  101741, 101588.8, 101413.3, 101206.5, 101001.8, 100820.1, 100704.2, 
    100735.9, 100836.6, 100965.3, 101155.4, 101346.5, 101465.8, 101577.4, 
    101664.7,
  101724.3, 101598, 101443.5, 101248.5, 101054, 100855.4, 100734.5, 100713.1, 
    100736.8, 100819.4, 100961.2, 101148.6, 101311.3, 101449.8, 101570.2,
  101768.8, 101664.3, 101530.7, 101355.2, 101165, 100948.4, 100764.1, 
    100663.3, 100670.3, 100706.1, 100804.8, 100966, 101162.8, 101329.7, 
    101476.6,
  101785.2, 101706.2, 101591.2, 101449.6, 101290.2, 101104.1, 100915.7, 
    100769.5, 100711.6, 100706.6, 100774.8, 100865.2, 101024.4, 101187.8, 
    101361.9,
  101788.2, 101742.8, 101656.5, 101551.9, 101409.6, 101257.3, 101086, 
    100924.5, 100811.2, 100771.5, 100793.7, 100865.7, 100980.6, 101114.8, 
    101267.3,
  101804.5, 101758.8, 101692.8, 101616.6, 101506.1, 101388.5, 101253.2, 
    101117.4, 100996.8, 100923.3, 100895, 100927.5, 100998, 101103.1, 101222.5,
  101821.3, 101785.6, 101731.5, 101668.8, 101581, 101489.4, 101383.5, 
    101273.1, 101166, 101083.7, 101038.5, 101039.2, 101072.4, 101136.4, 
    101225.5,
  101832.2, 101801.6, 101758.5, 101706.8, 101639.4, 101563.7, 101481.2, 
    101395.3, 101305.8, 101229.7, 101174.7, 101150.5, 101160.4, 101196, 
    101255.3,
  101833.4, 101812, 101779.9, 101732.3, 101676.7, 101616.9, 101551.6, 101481, 
    101408, 101341.7, 101292.1, 101262.6, 101253.3, 101267.2, 101309.7,
  101811.5, 101800.1, 101790.3, 101753.6, 101704.8, 101658.3, 101604.5, 
    101543.7, 101481.9, 101431.4, 101377.4, 101347.5, 101332.7, 101338.3, 
    101365.7,
  101471.8, 101432.3, 101419.2, 101410.1, 101400.3, 101384.4, 101373.7, 
    101376.3, 101394, 101442, 101518.1, 101630.1, 101763.8, 101890.8, 102015.6,
  101475.8, 101432.1, 101398.7, 101362.7, 101342.7, 101318.8, 101296, 
    101276.4, 101270.7, 101291, 101339, 101431.4, 101560.8, 101709.4, 101844.3,
  101513.6, 101446.1, 101394.2, 101346.1, 101312.3, 101276, 101239.1, 
    101201.3, 101175.5, 101164.3, 101184.2, 101232.6, 101350.5, 101488.6, 
    101659.5,
  101569.7, 101510.3, 101441.3, 101378.9, 101328.2, 101282.2, 101238.8, 
    101196.3, 101175, 101146.1, 101143.6, 101153.3, 101238.1, 101352.5, 
    101483.8,
  101620.5, 101573.6, 101516.9, 101443.7, 101375.5, 101315, 101261.4, 
    101210.7, 101176, 101145.2, 101122.8, 101134.1, 101172.2, 101287.2, 
    101423.5,
  101629.7, 101605.8, 101582, 101535.1, 101470.2, 101400.2, 101331.8, 
    101271.9, 101223, 101183.2, 101163.4, 101157.1, 101199.1, 101272.6, 
    101385.9,
  101635.2, 101619.8, 101611.3, 101588.5, 101548.4, 101495.4, 101437.8, 
    101371.5, 101313.7, 101267.9, 101241.7, 101236.6, 101261.9, 101324.8, 
    101404.2,
  101621.2, 101643.5, 101619.9, 101614.3, 101593.9, 101558.2, 101515.2, 
    101467.4, 101422.4, 101384.3, 101356.8, 101347.5, 101362.6, 101396.4, 
    101441.2,
  101544.2, 101644.8, 101658.7, 101635.3, 101614.9, 101596, 101566.2, 
    101528.7, 101498.4, 101471.7, 101450.8, 101439.3, 101442.7, 101455.9, 
    101481.7,
  101487.5, 101567.5, 101633.1, 101661.3, 101635.7, 101616.9, 101601.7, 
    101581.8, 101556, 101536.4, 101520.6, 101509.5, 101507.2, 101514.2, 
    101528.3,
  101717, 101708.5, 101709.2, 101720.2, 101728.8, 101745, 101770.9, 101811.8, 
    101864.7, 101922.7, 101983.4, 102063, 102142.9, 102234.7, 102314,
  101688.9, 101686.8, 101670.5, 101668.1, 101663.6, 101668.6, 101675.1, 
    101694, 101715.2, 101759.3, 101816.3, 101888.9, 101962.7, 102037.1, 
    102117.2,
  101674.6, 101671.4, 101639.4, 101626.6, 101603.6, 101583.9, 101567.9, 
    101564.2, 101571.8, 101599.7, 101637.9, 101700.6, 101794.2, 101890.4, 
    101983.5,
  101655.8, 101657.1, 101634.8, 101629.5, 101592, 101574.8, 101545.8, 101522, 
    101508.5, 101493.4, 101511, 101555.1, 101621.1, 101703.7, 101798.6,
  101672.2, 101657, 101633.8, 101627.7, 101588.5, 101565.1, 101527.9, 101498, 
    101489.1, 101476.7, 101473.5, 101475.4, 101520.2, 101598.4, 101682.1,
  101668, 101658.2, 101656.8, 101635.5, 101602.2, 101570.6, 101536.6, 
    101497.6, 101480.4, 101461.9, 101448.6, 101436.9, 101466.2, 101525.5, 
    101591.7,
  101635.6, 101650.4, 101662.9, 101647, 101626.4, 101588.9, 101554.8, 
    101513.3, 101482.3, 101459.5, 101440.4, 101430.1, 101445, 101504.1, 
    101563.6,
  101589, 101635.1, 101634.6, 101646.6, 101643.9, 101621, 101595.1, 101550.4, 
    101512.4, 101482.1, 101457.1, 101446.8, 101460.5, 101496.8, 101539.2,
  101517.3, 101591.7, 101628.2, 101636.1, 101642.6, 101640, 101617.8, 
    101594.2, 101558.1, 101526.6, 101499.8, 101486.6, 101489, 101508.4, 101536,
  101497.8, 101502.8, 101563.5, 101619.7, 101630.8, 101644.1, 101636, 
    101619.5, 101598.8, 101574.3, 101548.1, 101529.2, 101523.3, 101526.3, 
    101536.8,
  101726.9, 101752.4, 101788.6, 101824.1, 101857, 101901.1, 101950.5, 
    102002.6, 102061.3, 102115.3, 102156.6, 102192, 102210.5, 102218.2, 
    102221.8,
  101696.3, 101727.3, 101757.6, 101776.3, 101802.2, 101832.4, 101871.8, 
    101916.2, 101959.5, 102001.6, 102041.5, 102072.7, 102094.6, 102108.3, 
    102104.2,
  101679.7, 101710.1, 101731.4, 101738.7, 101749.5, 101766.8, 101788.7, 
    101825, 101867.9, 101910.7, 101949.3, 101984.1, 102005.2, 102003.7, 
    101988.4,
  101655, 101702.1, 101729.1, 101733.4, 101733.3, 101733.2, 101739.8, 
    101752.6, 101773.4, 101802.8, 101834.7, 101869, 101891.4, 101915.1, 101903,
  101641.3, 101683.4, 101715.9, 101727.9, 101723.1, 101715.2, 101709.5, 
    101711.7, 101717.3, 101725.3, 101750.2, 101773.4, 101805.8, 101814.7, 
    101825.5,
  101608.9, 101657.7, 101695.1, 101717.5, 101715.8, 101713.2, 101700.1, 
    101691.8, 101690.3, 101681.1, 101676.4, 101684, 101713, 101730.7, 101749.2,
  101574.5, 101632.5, 101674.4, 101696, 101690.1, 101698.6, 101687.6, 
    101673.6, 101663.7, 101651.3, 101634.3, 101635.5, 101648.2, 101667.9, 
    101675.4,
  101537.3, 101603, 101642.1, 101679.8, 101702.7, 101700.7, 101678, 101665.2, 
    101651.2, 101633.5, 101607.4, 101595.5, 101592.5, 101611.8, 101619.7,
  101516.7, 101569.7, 101612.5, 101638.7, 101672.3, 101683.4, 101681.6, 
    101662.8, 101640.5, 101625.3, 101600.3, 101579.2, 101564.1, 101573, 
    101576.7,
  101502.7, 101535.5, 101580.1, 101614.4, 101634.1, 101661.6, 101667.1, 
    101664.5, 101647.2, 101631.7, 101600.7, 101578.2, 101553.9, 101546.6, 
    101559.6,
  101415.2, 101395.7, 101419.8, 101459.9, 101527, 101579.8, 101630.2, 
    101689.8, 101735.3, 101755.3, 101751.9, 101737.4, 101725.4, 101696.3, 
    101674.4,
  101419.7, 101417.2, 101445, 101477.4, 101541.4, 101590.8, 101633.7, 
    101676.5, 101726.8, 101755.4, 101756.9, 101722.8, 101695.1, 101645.2, 
    101619,
  101431.2, 101439.5, 101455.3, 101481.3, 101542, 101599.3, 101635, 101675.2, 
    101726.9, 101754.8, 101756.6, 101721.2, 101681.2, 101625.8, 101584.8,
  101441.7, 101452.2, 101462.5, 101484.9, 101535.2, 101604.1, 101639.1, 
    101673.4, 101707.2, 101750.4, 101754.3, 101729.2, 101670.1, 101609.1, 
    101551.1,
  101452.2, 101463.7, 101474.1, 101493.8, 101534.7, 101600.5, 101643.9, 
    101674.1, 101698.4, 101731.2, 101752.2, 101735.2, 101685.7, 101619.1, 
    101552.1,
  101445.3, 101470.3, 101480, 101502.5, 101539, 101592.3, 101636.6, 101665.9, 
    101687.7, 101703.5, 101728.8, 101732, 101699.5, 101635.4, 101566.4,
  101427.6, 101463.7, 101489.5, 101510, 101543, 101585.8, 101636.4, 101657, 
    101679.8, 101686.8, 101706, 101711.3, 101702.8, 101659.3, 101594.3,
  101408.9, 101456.5, 101492, 101522.5, 101553.5, 101591.8, 101623.4, 
    101658.7, 101666.9, 101675.9, 101687.5, 101689.7, 101688.8, 101666.9, 
    101620.2,
  101404.2, 101450.9, 101492.7, 101518.8, 101558.9, 101591.6, 101636.1, 
    101666.1, 101666.9, 101677, 101672.3, 101670.4, 101671.5, 101665, 101634.3,
  101415.2, 101460.7, 101501.5, 101525.9, 101557, 101583, 101612.6, 101646.3, 
    101665, 101690.8, 101668.1, 101664.7, 101653.7, 101649.9, 101630.2,
  102074, 102012.3, 101947.5, 101886.8, 101816.8, 101754.2, 101688.1, 
    101626.2, 101569.2, 101514.8, 101460.5, 101403.9, 101350.9, 101313.7, 
    101283,
  102098.3, 102036.3, 101977, 101916, 101839.6, 101766.5, 101709.4, 101654.5, 
    101595.9, 101536.2, 101483, 101429.9, 101392.4, 101348.3, 101321.8,
  102130.1, 102060.3, 102000.8, 101931.1, 101847.5, 101780.9, 101718.2, 
    101663.6, 101603.2, 101543, 101492.1, 101440.1, 101407.8, 101366.7, 
    101346.5,
  102147.3, 102079.2, 102020.2, 101945.5, 101856, 101785.8, 101725.7, 
    101668.4, 101602.8, 101549.2, 101502.3, 101461.8, 101431, 101392.4, 
    101375.9,
  102162.3, 102089.6, 102024, 101949.1, 101847.4, 101764.3, 101711.8, 
    101664.3, 101616, 101564.5, 101517.3, 101476.6, 101447.5, 101410.3, 
    101396.7,
  102160.8, 102095.8, 102028.1, 101946.3, 101840.8, 101754.6, 101707.4, 
    101661.8, 101617, 101570.6, 101534.5, 101503.3, 101472.7, 101439.3, 
    101419.7,
  102145.7, 102085.5, 102009.3, 101923.9, 101826.8, 101726.4, 101661.7, 
    101647.8, 101612.4, 101570.7, 101550.8, 101523, 101493.8, 101468.3, 
    101442.4,
  102133.2, 102076.2, 101999.2, 101916.6, 101824, 101733.1, 101639.2, 
    101587.1, 101579.4, 101561.4, 101553.4, 101533.8, 101514.9, 101494, 
    101464.4,
  102113.2, 102056, 101983.8, 101905.3, 101816.5, 101730.7, 101627.2, 
    101542.3, 101505.6, 101519.1, 101546.4, 101545.8, 101532.5, 101517.2, 
    101490.5,
  102084, 102027.2, 101953, 101883.8, 101809, 101729.4, 101631.8, 101541.2, 
    101473.8, 101444.5, 101492.7, 101545.9, 101549.5, 101542, 101528.5,
  102056.5, 102039.6, 102015, 101983.4, 101954.6, 101925.9, 101898.3, 
    101868.2, 101828.1, 101791.6, 101744.2, 101695, 101637.7, 101574.4, 
    101509.6,
  102073.6, 102056.3, 102029.2, 102004.1, 101973.4, 101941.1, 101910.1, 
    101879.4, 101841.2, 101800.7, 101748.5, 101693.4, 101630.5, 101561.1, 
    101486.4,
  102085.4, 102063.4, 102040.6, 102012.6, 101978.6, 101945, 101911, 101878.3, 
    101842.4, 101799.9, 101749.2, 101688.3, 101618.4, 101546.2, 101460.7,
  102085.1, 102065, 102043.3, 102016.5, 101984.4, 101949.4, 101915.5, 
    101878.7, 101840.9, 101796.3, 101742.5, 101678.2, 101600.7, 101520.7, 
    101426.1,
  102083.3, 102061.1, 102042.8, 102013.7, 101982.7, 101948.4, 101913.1, 
    101874.1, 101832.6, 101786.7, 101734.8, 101667, 101583.1, 101496.3, 
    101394.9,
  102078.6, 102061.4, 102039.6, 102010.5, 101981.3, 101947.2, 101910.8, 
    101871.6, 101823.8, 101776.4, 101719.5, 101647.8, 101562.1, 101462.9, 
    101358.1,
  102077.9, 102059, 102034.8, 102006.9, 101977, 101943.4, 101905.3, 101861.5, 
    101813, 101763, 101706.9, 101632.3, 101544.3, 101442.5, 101327.9,
  102079.7, 102058.3, 102031.4, 102000, 101970.8, 101935.1, 101893.4, 
    101852.1, 101801.4, 101749.6, 101690.1, 101615.5, 101525.4, 101429.8, 
    101310.6,
  102078.7, 102052.8, 102023.7, 101992.2, 101958.4, 101921.2, 101880.8, 
    101836.2, 101789.6, 101735.6, 101675, 101599.1, 101509.6, 101421.1, 
    101315.1,
  102077.9, 102047.5, 102016.2, 101980.6, 101948.8, 101905.9, 101863.5, 
    101820.9, 101774.7, 101719.1, 101658.8, 101581.7, 101499.2, 101416.4, 
    101327,
  101657.8, 101677.9, 101702.9, 101720.3, 101734.7, 101747.7, 101758.5, 
    101772, 101779.9, 101779.6, 101776.1, 101769.8, 101762.2, 101753.8, 
    101747.4,
  101705.9, 101719.7, 101739, 101758.5, 101778.9, 101795.7, 101809.2, 101829, 
    101837.3, 101834, 101827.1, 101817, 101807, 101800.4, 101787.7,
  101735.7, 101748.8, 101775.3, 101796.3, 101819.1, 101835.4, 101850, 
    101868.5, 101870.3, 101866.1, 101858.2, 101848.3, 101837.9, 101831.6, 
    101829.5,
  101752.6, 101767.9, 101792.8, 101814.8, 101836.8, 101860.6, 101882, 
    101885.2, 101893.8, 101882.2, 101875, 101866.4, 101857.8, 101858.7, 
    101843.7,
  101763.1, 101786.6, 101810.1, 101829.8, 101851.1, 101879.3, 101896.2, 
    101901.5, 101899.5, 101891.8, 101877.9, 101874.3, 101863.5, 101856.9, 
    101834.6,
  101773, 101793, 101815.7, 101834.5, 101852.1, 101868.9, 101882.2, 101892.5, 
    101898.5, 101889.8, 101878.7, 101869.5, 101859.4, 101842.8, 101807.9,
  101766, 101794.5, 101818.7, 101839.3, 101852.4, 101865.7, 101877, 101883.3, 
    101882.1, 101880, 101870.8, 101858.2, 101836.8, 101810.2, 101770.1,
  101766.7, 101792.4, 101812.2, 101828, 101840.9, 101852.5, 101860, 101866, 
    101869.4, 101866.1, 101856.8, 101840.1, 101810.1, 101771.9, 101725.6,
  101762.9, 101792.3, 101806.9, 101825.4, 101832.2, 101836.6, 101848, 
    101853.4, 101857.5, 101851.8, 101840.5, 101818, 101784.5, 101740.1, 
    101698.8,
  101764.2, 101783.6, 101804.5, 101814.8, 101823.5, 101828.3, 101830, 
    101837.6, 101839.9, 101836.1, 101825, 101799.9, 101768.1, 101720.1, 
    101687.2,
  101366.8, 101316.4, 101282.6, 101251.7, 101222.4, 101195.1, 101174.4, 
    101164.1, 101157.5, 101167.9, 101182.3, 101202.4, 101222.7, 101248.9, 
    101274.4,
  101449.7, 101413, 101388.6, 101362.7, 101334.9, 101313.7, 101296.3, 
    101288.2, 101291.6, 101299.9, 101314.6, 101332.7, 101354.5, 101387.3, 
    101418.7,
  101535.3, 101506.2, 101488.1, 101470.6, 101450.1, 101432.9, 101420.9, 
    101413.4, 101413.7, 101420.1, 101430.6, 101446.2, 101464.8, 101495.3, 
    101522.1,
  101578, 101565.5, 101557.7, 101552.4, 101542.6, 101533.6, 101528, 101525, 
    101526.8, 101534.4, 101545.1, 101557.5, 101576.5, 101607.5, 101632,
  101630.7, 101631, 101634.5, 101632.7, 101631.3, 101626.9, 101626.5, 
    101623.6, 101628.6, 101631.5, 101642.7, 101655.3, 101673.8, 101696.6, 
    101713.4,
  101670.1, 101679.6, 101690.9, 101696.4, 101698.6, 101700.9, 101704.9, 
    101704.8, 101713.6, 101718.2, 101733, 101740, 101760.2, 101770.1, 101772,
  101709.6, 101725, 101743.9, 101751.4, 101756.4, 101762, 101766.2, 101771.1, 
    101778.9, 101787.9, 101805.2, 101815.6, 101823.4, 101812.9, 101816,
  101741.9, 101763.8, 101782.5, 101791.3, 101802.5, 101810, 101816.6, 
    101823.8, 101835.8, 101846.6, 101861.7, 101869.4, 101861.4, 101854.1, 
    101839.9,
  101770.1, 101794.7, 101816, 101831.3, 101845.2, 101854.3, 101859.8, 
    101867.7, 101880.3, 101889.3, 101898.3, 101898.2, 101890.4, 101877.7, 
    101866.2,
  101801.3, 101822.1, 101845.9, 101861.4, 101876.7, 101884.9, 101890.2, 
    101896.8, 101906.9, 101925.2, 101937.7, 101934.9, 101923, 101905.7, 
    101897.1,
  101530.8, 101481.3, 101454.2, 101429.5, 101397.7, 101367.3, 101327.6, 
    101284.6, 101233.2, 101184.9, 101136.9, 101084.5, 101023.8, 100960.3, 
    100892.1,
  101587.3, 101552.6, 101516, 101485, 101444.4, 101405.2, 101368.1, 101332.8, 
    101294.9, 101245.4, 101193.8, 101142.5, 101087.6, 101033, 100971.9,
  101660.3, 101614.8, 101579.2, 101550.6, 101514.8, 101476.2, 101437.8, 
    101394.4, 101354.5, 101311.6, 101264.9, 101214.4, 101162.4, 101113.2, 
    101062.1,
  101717.2, 101681.5, 101648.3, 101618.1, 101585.1, 101546.3, 101506.7, 
    101464.6, 101425.6, 101385.2, 101340.8, 101294, 101246.8, 101196.6, 
    101153.3,
  101759.8, 101737.1, 101711.1, 101683.3, 101651.7, 101615.5, 101581.1, 
    101543.2, 101502.8, 101462.2, 101417.2, 101372.8, 101330.7, 101291.9, 
    101250.1,
  101789.5, 101784.4, 101765.9, 101749.8, 101719.2, 101692.5, 101659.6, 
    101627.2, 101588.7, 101553, 101514, 101473.9, 101430.2, 101392.3, 101357.3,
  101807.1, 101819.5, 101818, 101807.8, 101786.9, 101763.4, 101735.6, 
    101706.6, 101673.8, 101642.7, 101608.4, 101575.6, 101538.9, 101501.1, 
    101472.9,
  101818.8, 101833.3, 101853.2, 101856.5, 101849, 101830.1, 101809.1, 
    101783.3, 101763.5, 101738.1, 101711.2, 101683.7, 101653.6, 101624.2, 
    101597,
  101827.7, 101863.6, 101887.8, 101896.2, 101894, 101886.7, 101874.8, 
    101858.7, 101842.9, 101826.3, 101809.1, 101785, 101763.1, 101739, 101717,
  101860.5, 101882.8, 101920.6, 101936, 101943.8, 101943, 101935.2, 101924.6, 
    101915.1, 101903.4, 101890.3, 101875.4, 101861.2, 101845.3, 101830.3,
  101531.7, 101444.4, 101373.9, 101300.3, 101223.7, 101154.1, 101083.4, 
    101020, 100957.9, 100894.8, 100838, 100789.3, 100740.6, 100699.8, 100657.9,
  101582.4, 101526.4, 101465.9, 101403.2, 101340.2, 101273.1, 101211.3, 
    101150, 101095.2, 101039.9, 100989.7, 100944, 100905.2, 100864.7, 100820.3,
  101639.7, 101589.3, 101536.6, 101488.5, 101432.9, 101376.8, 101323, 
    101271.4, 101222.5, 101173.7, 101129, 101085, 101047.5, 101013, 100978.9,
  101682.8, 101640.6, 101605.6, 101568.2, 101519.7, 101471.9, 101422.2, 
    101375.1, 101330.3, 101288.1, 101244.6, 101206.5, 101172, 101141, 101112,
  101718.2, 101683.8, 101653.9, 101625.4, 101582.9, 101541.1, 101503, 
    101461.9, 101423.7, 101387.6, 101353.2, 101317.3, 101286.1, 101259.5, 
    101231.6,
  101750.3, 101724.5, 101701.6, 101678, 101645.7, 101613.2, 101579.2, 
    101546.1, 101511.4, 101480.7, 101450.1, 101424.6, 101392.2, 101365.6, 
    101340.3,
  101777.7, 101763.5, 101749.7, 101733.3, 101706.2, 101680.5, 101649.7, 
    101622.2, 101592.2, 101566, 101540.4, 101515.6, 101491, 101470.9, 101449.5,
  101798.6, 101796.6, 101790.2, 101779.7, 101766.8, 101748, 101728.1, 
    101700.3, 101678.6, 101655.2, 101633.9, 101615.1, 101594, 101570, 101550.4,
  101821.2, 101830.8, 101831.9, 101829.7, 101821.2, 101807, 101789.8, 
    101772.8, 101759, 101740.4, 101722, 101705.1, 101690, 101671.3, 101660.5,
  101854.5, 101864.7, 101875, 101877.6, 101879.1, 101873.5, 101863.7, 101851, 
    101837.9, 101826.7, 101815.2, 101801.2, 101789.3, 101773.9, 101761.3,
  102132.5, 102077.1, 102030.9, 101971, 101906.1, 101833.7, 101760.6, 
    101679.5, 101593.3, 101505.5, 101415.7, 101321.8, 101230.6, 101143, 
    101056.7,
  102166.8, 102132.7, 102096.1, 102048.7, 101990.2, 101927, 101856.8, 
    101783.3, 101708.4, 101632.9, 101551.2, 101467.9, 101384.1, 101299.2, 
    101215.4,
  102199.8, 102179.4, 102146.8, 102110.9, 102063.4, 102006.8, 101945.8, 
    101884.5, 101814.6, 101744.9, 101670.3, 101596.5, 101518.7, 101442.7, 
    101370.2,
  102228.6, 102205.4, 102185.4, 102163.4, 102123.4, 102080.8, 102028.1, 
    101972.4, 101913.1, 101851.4, 101788.5, 101719, 101648.9, 101575.6, 
    101504.2,
  102243.2, 102223, 102212.2, 102191.4, 102153.9, 102115.9, 102075.4, 
    102024.9, 101971.7, 101917.4, 101860.3, 101800.8, 101739.8, 101677.4, 
    101615.3,
  102242.7, 102223.7, 102221.2, 102206.6, 102186.2, 102151.6, 102113.3, 
    102074.9, 102030.5, 101982.6, 101930.6, 101877.7, 101821, 101764.8, 
    101707.9,
  102237.8, 102229, 102226.9, 102211.4, 102191.6, 102166.4, 102132.9, 
    102095.5, 102057.2, 102013.7, 101971.5, 101921.6, 101872, 101820.8, 
    101773.1,
  102223.9, 102220.6, 102214, 102209.1, 102195, 102169.2, 102138.6, 102103.6, 
    102069.6, 102029.9, 101993.9, 101950.9, 101905.4, 101858.6, 101812.4,
  102197.7, 102202, 102196.9, 102198.7, 102184.7, 102159.1, 102134.7, 
    102101.6, 102073.9, 102034.5, 102000.2, 101962, 101922.4, 101881.9, 
    101840.4,
  102169.7, 102183.9, 102182.3, 102174.7, 102166.3, 102143.9, 102118.7, 
    102090.5, 102069.3, 102036.6, 102003.5, 101969, 101933.6, 101895.4, 
    101859.2,
  102055.2, 102061, 102069.3, 102055, 102037.6, 102010.3, 101974.4, 101928.1, 
    101874, 101817.8, 101754.4, 101683.6, 101613.8, 101542.4, 101475.2,
  102103.5, 102119.1, 102132.9, 102127.6, 102113.9, 102089.1, 102056.9, 
    102018.6, 101974.4, 101924.4, 101866.6, 101802.9, 101735.5, 101669, 
    101596.1,
  102139.3, 102168.9, 102190, 102194, 102185.7, 102168.2, 102141.6, 102106.4, 
    102065.8, 102018.3, 101966.9, 101909.4, 101846.3, 101779.7, 101715,
  102166.4, 102197.4, 102227.8, 102240.9, 102242.1, 102237.3, 102219, 
    102190.5, 102154.5, 102112.6, 102065.1, 102013, 101953.8, 101893.9, 
    101829.9,
  102184.3, 102222.4, 102256.5, 102273.9, 102279.5, 102278, 102268.9, 
    102251.1, 102221.9, 102187.8, 102142.6, 102096.5, 102043.2, 101986.8, 
    101926.2,
  102197.9, 102236.8, 102273.6, 102296.5, 102311.2, 102317.8, 102310.3, 
    102299.6, 102277, 102253.2, 102218.5, 102176.8, 102129.5, 102074.7, 
    102020.1,
  102212.3, 102242, 102283.5, 102308, 102330.5, 102340.3, 102342.2, 102332.9, 
    102314.5, 102293.8, 102267.3, 102232.9, 102193.4, 102149.6, 102099.3,
  102216.7, 102248.8, 102283.1, 102314.4, 102337.3, 102350.5, 102366.4, 
    102363, 102351.5, 102333.7, 102311.9, 102285.4, 102249.3, 102207.3, 102162,
  102216.9, 102248.4, 102274.4, 102306.9, 102329.4, 102349.8, 102362.8, 
    102363, 102358.6, 102355, 102342.5, 102319.6, 102292, 102259.8, 102217.5,
  102210.4, 102247.4, 102264.8, 102293.8, 102314.9, 102327.4, 102350.1, 
    102358.6, 102364.1, 102364.9, 102357.1, 102343.4, 102319.2, 102292.3, 
    102261.3,
  101556.2, 101572.9, 101596.1, 101610.1, 101617.9, 101616.2, 101604.1, 
    101593, 101583.1, 101569.7, 101542.3, 101511.6, 101490.6, 101461.6, 
    101423.7,
  101640.5, 101665.2, 101693, 101717.3, 101727.2, 101734, 101730.3, 101719.3, 
    101705.2, 101687.7, 101668.1, 101639.2, 101595.8, 101553.4, 101508.3,
  101710.3, 101740.3, 101775.7, 101803.7, 101822.2, 101836.5, 101839.9, 
    101837, 101826.4, 101814.7, 101794.6, 101767.1, 101726.9, 101678.2, 
    101625.2,
  101775, 101808.9, 101849.1, 101878.5, 101904.9, 101923.5, 101937.4, 
    101941.5, 101939.2, 101928.3, 101911.2, 101885.4, 101852.9, 101807.7, 
    101758.7,
  101829.4, 101869.4, 101914.1, 101945.6, 101973.8, 101999.7, 102015.2, 
    102027.1, 102031, 102029, 102018.9, 101996.7, 101969.4, 101929, 101883.9,
  101877.7, 101923, 101968.3, 101999.3, 102031.8, 102058.7, 102081, 102099.7, 
    102109.4, 102114.8, 102111.6, 102097.6, 102077.1, 102043.4, 102001.9,
  101921, 101963.7, 102007.8, 102040, 102077.1, 102100.8, 102130.9, 102150, 
    102170.7, 102178.5, 102184, 102177.9, 102161, 102134.2, 102098.5,
  101955.3, 101997.3, 102039.6, 102074.4, 102113.2, 102138.4, 102169.3, 
    102195.5, 102223.6, 102238.6, 102248.9, 102247, 102235.5, 102215.1, 
    102186.3,
  101982.8, 102026.5, 102067.2, 102100.4, 102133.7, 102160.8, 102193.1, 
    102224, 102258, 102276, 102288.7, 102295.2, 102287.8, 102271.5, 102249,
  102002.4, 102042.4, 102083, 102115.7, 102146.2, 102177, 102204, 102244.4, 
    102282.5, 102294.9, 102318.2, 102327.2, 102325.4, 102316.9, 102299.8,
  101152.9, 101169.9, 101191.6, 101209, 101220.2, 101219.1, 101210, 101201.8, 
    101191.3, 101171.2, 101154.3, 101138.1, 101108, 101070.2, 101035.8,
  101238.7, 101265.4, 101301.7, 101327.8, 101345.7, 101358.1, 101364.7, 
    101366.4, 101361.3, 101357, 101346, 101322.8, 101299.4, 101271.9, 101241.5,
  101306.8, 101347.1, 101395.2, 101431.3, 101458.8, 101482.3, 101497.7, 
    101505.1, 101507.4, 101509.9, 101506.9, 101498.5, 101480.3, 101456.7, 
    101431.9,
  101370.6, 101418.1, 101472.4, 101513.4, 101555.5, 101588.1, 101610.7, 
    101626, 101636.2, 101646.9, 101650.8, 101650.3, 101642.7, 101629.4, 
    101605.8,
  101425.4, 101480.4, 101547.8, 101596.4, 101644.5, 101677.5, 101705.1, 
    101725.5, 101744.6, 101762.2, 101775.9, 101785.3, 101787.4, 101780.4, 
    101769.8,
  101475.5, 101533.8, 101609.2, 101657.8, 101710.6, 101746.6, 101777.7, 
    101804.8, 101829.8, 101858, 101878.3, 101897, 101906.2, 101910.9, 101911.2,
  101516.9, 101578.2, 101659.2, 101708.5, 101764.5, 101798.7, 101836.1, 
    101867.7, 101905.3, 101938.3, 101962.7, 101989.2, 102009, 102026.6, 
    102033.4,
  101557.3, 101620.8, 101698.1, 101750, 101800.3, 101836.6, 101879.4, 
    101915.9, 101958, 101994.2, 102028.4, 102065.2, 102093.5, 102119.3, 
    102130.1,
  101597.8, 101658.2, 101728.2, 101780.1, 101825.4, 101862.4, 101907.6, 
    101941.9, 101988.7, 102033.8, 102077.4, 102117.2, 102152.7, 102183.2, 
    102199,
  101636.8, 101693.4, 101753.5, 101804.1, 101841.3, 101878.2, 101919.1, 
    101958, 102007.1, 102055.8, 102104.1, 102148.7, 102190.8, 102220.6, 
    102248.3,
  101657.4, 101575.8, 101526.9, 101471.6, 101436.8, 101404.6, 101378.7, 
    101343.2, 101311.7, 101280.3, 101237.3, 101188.5, 101124.7, 101055.1, 
    100987.2,
  101697.6, 101621.9, 101579.6, 101529.4, 101494.9, 101459.3, 101432.5, 
    101409.9, 101383.8, 101349.4, 101313.5, 101272.3, 101225.7, 101174.2, 
    101111,
  101744.7, 101689.6, 101648.9, 101601.1, 101563.4, 101526.3, 101495.2, 
    101468.7, 101444.3, 101418.4, 101392.3, 101360.5, 101321.7, 101277.6, 
    101228.4,
  101775.7, 101735, 101699.2, 101660.4, 101630.8, 101600.2, 101578.2, 
    101552.8, 101529.2, 101502.7, 101479.1, 101453.9, 101426.3, 101396.4, 
    101362.2,
  101789, 101765.1, 101735.6, 101710.6, 101686.6, 101664.7, 101645.9, 
    101626.1, 101604.2, 101582.1, 101559.7, 101540.4, 101523.8, 101502.3, 
    101478.6,
  101778.9, 101776.8, 101761.9, 101747.6, 101733.2, 101722.1, 101708.9, 
    101692.9, 101676.6, 101660.2, 101644.4, 101631.9, 101616.9, 101603.8, 
    101591.7,
  101764.5, 101771.1, 101776.2, 101773, 101768.8, 101760.3, 101751.6, 101740, 
    101731.8, 101725.1, 101717, 101711.8, 101704.6, 101698.1, 101689.7,
  101733.8, 101763.4, 101776.6, 101787.7, 101787.4, 101786.2, 101781.2, 
    101776.7, 101777.3, 101778.6, 101781, 101783.2, 101787.7, 101788.6, 101789,
  101696.1, 101739.9, 101768.1, 101787.1, 101796.2, 101796.2, 101796.7, 
    101802.6, 101813.5, 101821, 101833.6, 101842.6, 101854.5, 101861.8, 
    101870.2,
  101675.5, 101727.8, 101762.6, 101786.4, 101799.9, 101806.8, 101812.1, 
    101821.9, 101835, 101850.8, 101868.9, 101886.2, 101908.8, 101923.4, 
    101940.7,
  102583.9, 102665.7, 102732.3, 102806.6, 102877.2, 102942.2, 103007.8, 
    103071, 103133.4, 103188.4, 103229.7, 103261.2, 103284, 103307.6, 103322.8,
  102522.2, 102574.7, 102641.7, 102707, 102774.4, 102833.4, 102903.8, 
    102973.2, 103040.8, 103097.2, 103142.3, 103176.9, 103203.3, 103220.6, 
    103231.9,
  102483.2, 102508.9, 102560.1, 102609.4, 102669.8, 102732.6, 102791.8, 
    102856.8, 102922.2, 102982.1, 103035.5, 103075.8, 103105.9, 103128.4, 
    103142.4,
  102454, 102467.1, 102498.9, 102537, 102582.5, 102630.6, 102687.3, 102744.7, 
    102806.9, 102864.1, 102916.9, 102964.7, 103002.5, 103026.5, 103037.9,
  102434.2, 102432.2, 102444.7, 102466.9, 102501.3, 102537.8, 102581.4, 
    102630.9, 102684.8, 102739.2, 102791.8, 102840, 102879, 102906.9, 102925.2,
  102406.2, 102404.2, 102412.3, 102415.9, 102429.5, 102454.8, 102487.9, 
    102529.5, 102574.4, 102619, 102670.8, 102714.3, 102753, 102792.4, 102812.9,
  102378.8, 102376.1, 102373.7, 102370.2, 102379.6, 102388.3, 102403.8, 
    102427.8, 102462.9, 102499, 102543.7, 102581.3, 102625.4, 102663.6, 
    102692.4,
  102341.4, 102333.4, 102333.1, 102328.2, 102326.4, 102325.7, 102335.4, 
    102352.2, 102375.7, 102401.7, 102432.3, 102467, 102501.4, 102534.8, 
    102563.6,
  102292.8, 102288.1, 102285.5, 102276.4, 102267.1, 102263.1, 102265.1, 
    102270.4, 102281.8, 102298.3, 102323.4, 102352.4, 102384.1, 102413.5, 
    102440.4,
  102229.5, 102234.7, 102224.5, 102219.4, 102210.8, 102197.6, 102190.4, 
    102195.2, 102203.5, 102215.6, 102239.6, 102266, 102286.6, 102308.6, 
    102330.3,
  102301.5, 102421.8, 102526.7, 102624, 102724, 102821, 102911.8, 103001.1, 
    103093.7, 103181.8, 103262.8, 103342.7, 103419.3, 103491.6, 103551.5,
  102203.1, 102334.5, 102446.5, 102557.2, 102658.1, 102753.6, 102846, 
    102937.4, 103023.4, 103113.8, 103200.7, 103280, 103351, 103425, 103493.3,
  102136.9, 102274.7, 102386.1, 102492, 102589, 102688.8, 102777.8, 102867.3, 
    102956.4, 103047.1, 103132.3, 103214.2, 103286.6, 103356.5, 103422,
  102062.1, 102189.9, 102302.5, 102414.6, 102512, 102610.3, 102698.7, 
    102787.6, 102869.6, 102958.5, 103042.1, 103127.5, 103201.7, 103273.9, 
    103341.4,
  102020.1, 102130.8, 102237.7, 102344.1, 102439.1, 102528.1, 102617.5, 
    102702.7, 102786.9, 102870.1, 102951.6, 103033.8, 103109.8, 103176.2, 
    103242.9,
  101983, 102066.6, 102166.8, 102263.5, 102353.9, 102444, 102524.9, 102609.4, 
    102689.3, 102767.3, 102850.4, 102927.3, 103005, 103074.9, 103139.1,
  101956.4, 102019.8, 102106.6, 102188.6, 102275.5, 102358.1, 102436.5, 
    102513.4, 102589.7, 102665.2, 102739.5, 102813.6, 102887.9, 102957.4, 
    103024.7,
  101930, 101972.2, 102040, 102110.8, 102188.9, 102266.2, 102339.6, 102418.9, 
    102492.4, 102559.9, 102634.5, 102701.5, 102766.8, 102831.9, 102891.2,
  101900.7, 101932.4, 101982.4, 102037.9, 102100.4, 102171.9, 102244.8, 
    102311.4, 102387, 102456.5, 102523.4, 102590.6, 102653.7, 102710.4, 
    102766.9,
  101867.1, 101894.6, 101925.2, 101964.2, 102012.6, 102072, 102141.2, 
    102212.4, 102270.5, 102344.8, 102405.8, 102472.3, 102531.9, 102587.8, 
    102641.7,
  100920.6, 101036.5, 101210, 101412.9, 101615.1, 101814.8, 101991.9, 
    102151.3, 102299.9, 102437, 102567.2, 102690.9, 102811.4, 102923.7, 
    103028.7,
  100920.1, 101006.3, 101180.1, 101363.2, 101554, 101745.7, 101921.6, 102090, 
    102242.4, 102385.6, 102518.6, 102647.6, 102768.5, 102882.2, 102988.5,
  100999.3, 101055.1, 101171, 101317.2, 101482.6, 101660.6, 101839, 102011.9, 
    102167.9, 102314.6, 102457.4, 102591.6, 102717.4, 102835.8, 102946.3,
  101123.2, 101152.6, 101225.4, 101337.3, 101483.3, 101634.6, 101794, 
    101952.8, 102105.9, 102252.1, 102392.1, 102527.5, 102657, 102775.1, 
    102882.3,
  101251.7, 101267, 101321.6, 101401.6, 101514.3, 101638.7, 101781.4, 
    101920.2, 102063.9, 102195.5, 102328.4, 102460.4, 102588.9, 102708, 102817,
  101351.2, 101362.1, 101407.4, 101471.7, 101568.1, 101675.3, 101792, 
    101903.7, 102023.9, 102146.3, 102269.8, 102392.4, 102513.4, 102633.9, 
    102739.1,
  101427.5, 101436.7, 101476.9, 101527.4, 101610.1, 101702.4, 101804.5, 
    101894.8, 101995.3, 102097.7, 102210.8, 102325, 102438, 102549.6, 102656.1,
  101479.9, 101485.9, 101520.2, 101565.7, 101637.3, 101710, 101793.9, 
    101873.5, 101959.5, 102050.3, 102153.6, 102259.2, 102361.7, 102468, 102568,
  101519.4, 101529.1, 101556.9, 101587.8, 101641.5, 101695.8, 101777.7, 
    101839.5, 101921.2, 101999.5, 102089.6, 102187.8, 102284, 102380.7, 
    102477.7,
  101549.6, 101556.4, 101579.8, 101604.4, 101643.3, 101685.8, 101740.4, 
    101801.7, 101865.3, 101942.8, 102022.6, 102112.5, 102201, 102295.5, 
    102386.1,
  101551.2, 101391.8, 101211.5, 101041.2, 100907.8, 100827.6, 100803.7, 
    100843, 100941.1, 101091.9, 101277.8, 101470.2, 101660.8, 101849.5, 
    102037.9,
  101578.8, 101439.2, 101287.2, 101140.5, 101026.5, 100954.5, 100927.3, 
    100949.8, 101030.8, 101167.5, 101333.6, 101509.1, 101696.9, 101876.2, 
    102055,
  101653.4, 101538.6, 101412.7, 101277, 101170, 101095.3, 101058.9, 101065.2, 
    101123.4, 101232.3, 101373.6, 101534.7, 101710.9, 101892.2, 102064.7,
  101704.4, 101619.7, 101513.1, 101399.6, 101311.8, 101244.1, 101205.2, 
    101201.5, 101242.5, 101332.4, 101447.2, 101587.5, 101748, 101914.9, 
    102075.7,
  101750.9, 101686.8, 101603.5, 101518.4, 101437.7, 101374.1, 101330.4, 
    101318, 101343, 101407.2, 101498.5, 101617.4, 101766.3, 101926.6, 102075.9,
  101793.8, 101735.9, 101672.9, 101599.5, 101530.1, 101476.1, 101436, 
    101422.9, 101438.9, 101487.7, 101553.4, 101645.9, 101768.2, 101915.9, 
    102061.5,
  101832.7, 101776.3, 101723.9, 101663.4, 101603.2, 101554.1, 101514.3, 
    101498.2, 101506.5, 101527.4, 101577.9, 101652.3, 101761.8, 101896.5, 
    102036.5,
  101853.5, 101806.9, 101759.1, 101703.7, 101654.1, 101607.1, 101575.6, 
    101557.5, 101553, 101567.9, 101604.9, 101663.1, 101754.1, 101877.1, 
    102001.5,
  101867.1, 101824.3, 101782.2, 101734.7, 101687.7, 101647.4, 101606.1, 
    101589.6, 101581.9, 101581.8, 101611.3, 101667.7, 101759.3, 101864.3, 
    101974.9,
  101867.1, 101831.7, 101793.1, 101751.4, 101709.3, 101672.1, 101636.9, 
    101611.5, 101594.4, 101593.8, 101617.1, 101670, 101752.5, 101852.2, 
    101953.7,
  102426.1, 102352.3, 102274.4, 102189.8, 102089.8, 101983.3, 101857.4, 
    101714.9, 101555.9, 101388.5, 101218.6, 101056, 100916.1, 100799.6, 
    100715.5,
  102379.2, 102321.9, 102259.4, 102177, 102081.2, 101978, 101858.8, 101727.7, 
    101579.1, 101418.6, 101253.6, 101101.1, 100965.2, 100855, 100764.6,
  102354.7, 102310.7, 102244.8, 102167.1, 102077.3, 101982.8, 101876, 
    101752.7, 101617.2, 101464.9, 101306.8, 101156.5, 101016.5, 100906.2, 
    100818,
  102322.2, 102287.7, 102226.9, 102158.2, 102080.5, 101992.1, 101892.7, 
    101779.8, 101656.5, 101519, 101371.8, 101229.5, 101090.5, 100979.2, 
    100893.6,
  102291.2, 102266.3, 102212.2, 102152.1, 102076, 101997, 101908.2, 101808.8, 
    101697, 101573.7, 101439.1, 101304.4, 101172, 101054.5, 100971.1,
  102270.5, 102238.3, 102198.9, 102143.3, 102072.6, 102003.2, 101920.3, 
    101830.2, 101731.7, 101623.1, 101505.5, 101382.8, 101258.7, 101143.5, 
    101062.5,
  102251.1, 102214, 102174.2, 102133.5, 102067.1, 102003.7, 101930.7, 
    101848.4, 101759.3, 101664, 101561.9, 101453.1, 101343.8, 101236, 101158.1,
  102238.3, 102193.6, 102150.8, 102116.6, 102063, 102000.9, 101934.5, 
    101859.8, 101782.8, 101696.7, 101607.7, 101513.4, 101421.1, 101323.9, 
    101251.8,
  102225.8, 102177.9, 102133.2, 102093.8, 102050.6, 101995.5, 101934, 
    101867.3, 101797.4, 101722.6, 101643, 101561.3, 101479.3, 101399, 101329.8,
  102212, 102163.4, 102119.2, 102076.8, 102040.2, 101987.7, 101930.4, 
    101872.8, 101812.7, 101742.4, 101671.1, 101597.1, 101522.8, 101448.8, 
    101391.6,
  102858.2, 102830.2, 102775.7, 102718.5, 102643.5, 102553.7, 102450.1, 
    102337.4, 102215.1, 102081.8, 101941.2, 101795.3, 101636, 101460, 101274.3,
  102824.1, 102789.8, 102728.4, 102659.7, 102576.8, 102485.4, 102380.4, 
    102265.6, 102138, 102002.1, 101856.2, 101707.6, 101544.8, 101360, 101153.4,
  102790.7, 102759.9, 102703.9, 102635.3, 102546, 102446.8, 102335, 102209.8, 
    102077.6, 101935.6, 101786.7, 101636.1, 101480.3, 101298.5, 101098.9,
  102745, 102715.3, 102659.5, 102592.3, 102505.8, 102406.7, 102295.7, 
    102171.1, 102038.7, 101892, 101747.4, 101590.8, 101440.9, 101267, 101073.9,
  102705.2, 102685.4, 102631.6, 102567.5, 102484, 102386.6, 102271.4, 
    102147.6, 102006.8, 101863.1, 101707.8, 101559, 101408.2, 101244.6, 
    101081.1,
  102666.8, 102647.9, 102601.1, 102540.8, 102459, 102368.4, 102257, 102134.4, 
    102000.8, 101857.9, 101704.1, 101553, 101404.1, 101250.5, 101098.6,
  102629.6, 102615.3, 102569.2, 102515.3, 102441.9, 102357.2, 102250.1, 
    102130, 101999.1, 101860, 101717.3, 101566.7, 101417.2, 101279.3, 101142,
  102586.2, 102578.1, 102533, 102486.2, 102416.2, 102341.9, 102241.8, 
    102130.1, 102007.1, 101874, 101734.1, 101594.3, 101447, 101311.6, 101189.3,
  102550.3, 102539.8, 102498.1, 102455.3, 102391.7, 102322.8, 102232.6, 
    102134.1, 102016.5, 101896.4, 101763.1, 101631.2, 101496.7, 101365.6, 
    101248.9,
  102513.2, 102497.6, 102460.6, 102415.7, 102363.3, 102298.1, 102218.7, 
    102130, 102029.7, 101916.2, 101798.9, 101677.7, 101555.3, 101432.8, 
    101321.8,
  102118.3, 102142, 102142.5, 102130.4, 102096.7, 102036.5, 101963.7, 
    101858.5, 101731.9, 101560.3, 101367.3, 101154.8, 100933.2, 100741.5, 
    100628.4,
  102132.5, 102160.1, 102162.7, 102142.7, 102107.1, 102043.4, 101964.9, 
    101860.1, 101732.9, 101572.6, 101384.3, 101161.2, 100908.5, 100687.9, 
    100534.5,
  102148.4, 102176.6, 102180.7, 102164.6, 102125.2, 102066.6, 101990.8, 
    101891.2, 101760.7, 101601.1, 101417.2, 101208, 100934.2, 100684.7, 100486,
  102162.2, 102193.5, 102195.4, 102188.1, 102145.3, 102086, 102007.7, 
    101916.2, 101796.5, 101651.3, 101475.3, 101281.3, 101039.1, 100773.9, 
    100550.7,
  102182.7, 102211.5, 102212.4, 102207.3, 102170, 102116.4, 102042.6, 
    101954.1, 101843.7, 101712.2, 101549.3, 101377, 101171.6, 100930.1, 100710,
  102192.4, 102221.8, 102229, 102220.9, 102189.9, 102142, 102072.1, 101988.7, 
    101889.8, 101772.7, 101630.2, 101472, 101295, 101097.1, 100900.9,
  102207.3, 102232.9, 102244, 102235.8, 102207.6, 102167.8, 102107.4, 
    102028.2, 101937, 101829.6, 101709.9, 101570.6, 101416, 101252.7, 101090.3,
  102213, 102244.5, 102256, 102251.8, 102224.3, 102188, 102134.4, 102061.9, 
    101980.2, 101883.5, 101776.5, 101660, 101527.5, 101390.6, 101253.8,
  102223.3, 102252.4, 102262, 102260.3, 102239.1, 102202.9, 102158.9, 
    102095.2, 102020.4, 101935.5, 101838, 101737.2, 101623.2, 101510.1, 
    101393.7,
  102233.9, 102259.3, 102268.8, 102267.2, 102246.1, 102216, 102175, 102123, 
    102058.3, 101981.1, 101895.2, 101804.9, 101706.9, 101607.4, 101505.8,
  101714.2, 101709.1, 101704, 101697.7, 101685.9, 101666.9, 101634.7, 
    101598.9, 101563.2, 101546.5, 101526.2, 101496.3, 101448.9, 101404.3, 
    101348.8,
  101746.5, 101762.2, 101771.6, 101776.7, 101774.9, 101769.3, 101751.4, 
    101720.5, 101684.3, 101652.4, 101617.6, 101582.7, 101535.8, 101484, 
    101427.3,
  101784.7, 101814.7, 101834.4, 101853.4, 101857.7, 101859.6, 101853.5, 
    101831.3, 101796.9, 101757.8, 101721.1, 101682.7, 101634.9, 101577.8, 
    101518.6,
  101821.4, 101858.1, 101889, 101921, 101937.1, 101951.3, 101949.5, 101936.4, 
    101909.5, 101871.2, 101830.5, 101786.5, 101736.7, 101677.8, 101612.9,
  101849.8, 101900.7, 101945.3, 101982.5, 102004.3, 102025.5, 102034.5, 
    102029.9, 102011.8, 101981.2, 101940.4, 101896.2, 101846.5, 101788.6, 
    101720.2,
  101874.7, 101936.6, 101991.3, 102032.6, 102066.9, 102094.9, 102110.9, 
    102111.7, 102101.5, 102078.9, 102047.2, 102005.1, 101954.7, 101896.5, 
    101833,
  101903.6, 101968.4, 102031.2, 102077.6, 102117.2, 102148, 102169.4, 
    102176.5, 102176, 102158.4, 102136.1, 102098.8, 102053.8, 101999.9, 
    101935.4,
  101930.4, 102001.4, 102069, 102115.8, 102162.9, 102195.1, 102216.9, 
    102227.7, 102232, 102224.7, 102207.8, 102181.7, 102140.4, 102093.9, 
    102037.4,
  101965.2, 102033.3, 102105.1, 102153.8, 102204.5, 102234.6, 102253.5, 
    102270.3, 102277.7, 102280.3, 102267, 102249, 102213.2, 102176, 102123.8,
  102000.8, 102068.2, 102139.7, 102189.5, 102241.5, 102267.8, 102287.3, 
    102304, 102319.7, 102327.3, 102320.5, 102303.3, 102274.6, 102240.9, 
    102196.1,
  101396.2, 101406.4, 101436.3, 101460.5, 101493.9, 101519.7, 101541, 
    101561.5, 101575, 101576.1, 101568, 101555.1, 101532, 101502.3, 101467.7,
  101445.4, 101471.5, 101499.8, 101530.3, 101561.1, 101595.6, 101624.5, 
    101644.1, 101652.8, 101654.8, 101651.7, 101641.3, 101623.9, 101593.4, 
    101556.4,
  101501.9, 101544.4, 101574.6, 101611.3, 101640.6, 101674.2, 101704.6, 
    101729.2, 101740.6, 101742.5, 101736.4, 101721, 101699.6, 101678.3, 
    101651.2,
  101548.8, 101602.7, 101641.6, 101683.9, 101720.9, 101752, 101777.3, 
    101793.6, 101806.3, 101811.4, 101810.8, 101799, 101778.4, 101754.9, 
    101726.3,
  101598, 101656.3, 101711.9, 101758.9, 101799.3, 101833.2, 101861.1, 101881, 
    101894.7, 101895.2, 101887.2, 101875.8, 101860.8, 101842, 101817.9,
  101639.5, 101704.8, 101768.8, 101820.1, 101867.6, 101905.9, 101934.7, 
    101960.4, 101975.4, 101984.9, 101982.7, 101972.7, 101952.2, 101931.8, 
    101906.1,
  101682, 101752, 101819.1, 101877.1, 101928.5, 101967.1, 101999.1, 102029.9, 
    102049.2, 102062.7, 102065, 102062.1, 102049.6, 102032.9, 102009.4,
  101722.4, 101793.8, 101867.7, 101927.5, 101980.3, 102019.3, 102059, 
    102092.3, 102112.9, 102130.7, 102140.7, 102142.4, 102137.7, 102123.3, 
    102106.9,
  101767.1, 101838, 101913.5, 101969.1, 102026.9, 102068.1, 102109.8, 
    102140.4, 102164.4, 102185.8, 102198.8, 102203.9, 102203.7, 102196.2, 
    102187.1,
  101812, 101880.1, 101953.7, 102005.4, 102064.6, 102105.9, 102144.5, 
    102171.9, 102200.6, 102225.8, 102240.7, 102256.7, 102264, 102264.1, 
    102261.9,
  101692.9, 101643.3, 101588.2, 101531.5, 101467, 101400.6, 101337.6, 
    101277.5, 101229.9, 101192.2, 101168.2, 101157.1, 101138.2, 101106.4, 
    101065.3,
  101748.6, 101697.5, 101640.5, 101580.8, 101517.2, 101456.1, 101397.7, 
    101356.2, 101319.8, 101289.2, 101264.8, 101236.7, 101208.5, 101184.9, 
    101172.2,
  101797.9, 101747, 101690.6, 101639.6, 101581.6, 101525.2, 101471.4, 
    101423.2, 101390.6, 101368.6, 101347.9, 101324.6, 101314.8, 101300.9, 
    101290.5,
  101830.2, 101780.4, 101724, 101672.1, 101617, 101572.3, 101543.7, 101521, 
    101494.5, 101459.2, 101431.5, 101413.8, 101406, 101398.5, 101384.8,
  101849.5, 101808.4, 101763.8, 101728.9, 101689.6, 101663.1, 101634.1, 
    101601.1, 101563.3, 101529.1, 101508.9, 101497.8, 101492.5, 101487.9, 
    101486.4,
  101863.2, 101835.8, 101798.2, 101765.1, 101733.8, 101706.7, 101680.9, 
    101658.8, 101634.6, 101612.5, 101594.1, 101582.4, 101572.2, 101574.1, 
    101573.7,
  101865.6, 101841.7, 101817.4, 101793.6, 101766.3, 101743.7, 101728.2, 
    101713.7, 101692.3, 101678.7, 101668.6, 101662.1, 101656.2, 101656.9, 
    101664.2,
  101851.1, 101841.7, 101824.4, 101809.2, 101789.3, 101771.6, 101760.8, 
    101747.2, 101744.5, 101738.6, 101737.7, 101738.2, 101738.3, 101743.8, 
    101751.9,
  101821.3, 101829.1, 101821.8, 101811, 101801.3, 101788.6, 101781, 101777.4, 
    101780.6, 101784.8, 101795.3, 101806.1, 101813.7, 101820.3, 101832.4,
  101788.6, 101807.8, 101810.9, 101811.2, 101808.6, 101799.9, 101795.5, 
    101795.9, 101810.9, 101823.3, 101838.7, 101856.4, 101868.2, 101884.5, 
    101902,
  101872.1, 101796, 101732.7, 101673.4, 101612, 101554.5, 101497.9, 101446.3, 
    101401.1, 101361.2, 101327.5, 101298.5, 101273.5, 101254.4, 101245.5,
  101957.6, 101902.1, 101849.6, 101798.6, 101745.3, 101691.3, 101640.7, 
    101591.9, 101550.6, 101508.9, 101474, 101441.1, 101412.5, 101396.6, 
    101384.4,
  102028.2, 101980, 101938.8, 101899, 101852.7, 101808.4, 101764.1, 101720.6, 
    101679.4, 101637.3, 101603.8, 101568.8, 101538, 101517.9, 101505.8,
  102078, 102044.5, 102014.5, 101985.5, 101948.4, 101907.8, 101871, 101830.7, 
    101791, 101755.4, 101715.1, 101683.4, 101650.4, 101625, 101608.2,
  102115.7, 102092.7, 102072.1, 102046.1, 102020.3, 101988.2, 101952.2, 
    101917.6, 101881.6, 101845.9, 101807.8, 101770.4, 101735.6, 101708.9, 
    101685.4,
  102141.8, 102123.8, 102114.2, 102092.6, 102069.7, 102044.9, 102014.7, 
    101984.6, 101950.3, 101915.3, 101877.8, 101835.8, 101798.8, 101770.6, 
    101749.6,
  102161.5, 102146.5, 102139, 102123.2, 102100.7, 102080.5, 102059, 102030, 
    102000.3, 101967.9, 101928, 101884, 101849.9, 101819.9, 101792.9,
  102171.5, 102157, 102154.4, 102137.6, 102117.8, 102095.3, 102070.6, 
    102042.6, 102016.9, 101992.1, 101958.4, 101930.4, 101896.7, 101873.9, 
    101838,
  102170.8, 102162, 102157.1, 102137, 102120.7, 102093, 102068.7, 102050.5, 
    102031.9, 102011.5, 101986.5, 101960.2, 101929.5, 101906.5, 101870.8,
  102157.5, 102150, 102143.1, 102125.3, 102110.5, 102080.6, 102058.4, 102039, 
    102022.7, 101997.8, 101988.9, 101967.2, 101943.3, 101920, 101894.2,
  102477.1, 102457.2, 102439, 102409.2, 102371.3, 102328.9, 102280.1, 
    102225.4, 102150.4, 102074.4, 101988.4, 101894.2, 101793.5, 101685.9, 
    101568.3,
  102486.5, 102479.1, 102468.4, 102443.3, 102410.7, 102370, 102319.6, 
    102270.4, 102207.9, 102138, 102060.8, 101976.7, 101879.1, 101775.3, 
    101666.4,
  102507.1, 102507.6, 102494.8, 102475, 102449.7, 102410.1, 102362.8, 
    102312.2, 102253.9, 102189.7, 102116.2, 102038.3, 101952.7, 101856.5, 
    101757.8,
  102518.5, 102520.9, 102514.6, 102496.8, 102471.7, 102443.2, 102402.4, 
    102359, 102306.6, 102247.4, 102180.8, 102108.4, 102026.9, 101938.9, 
    101846.6,
  102534, 102528, 102522.4, 102508.8, 102484, 102459.3, 102426.6, 102386.7, 
    102338.5, 102285.4, 102225.8, 102159.8, 102086.2, 102008.2, 101923.6,
  102545.6, 102534.9, 102525.3, 102515.6, 102496.1, 102474.5, 102443.8, 
    102407.9, 102367.2, 102315.9, 102265.3, 102205.7, 102138.7, 102068.8, 
    101994.2,
  102547.8, 102534.1, 102522.1, 102508.4, 102492.1, 102472.4, 102448.2, 
    102416.5, 102379.6, 102341.1, 102295.1, 102244.2, 102183.4, 102120.4, 
    102054.8,
  102536.8, 102524.7, 102510.4, 102496.8, 102481.5, 102461.7, 102439.3, 
    102413.2, 102385.4, 102352.1, 102312.4, 102269.7, 102218.5, 102162.3, 
    102102.3,
  102523.5, 102513.3, 102494.9, 102478.4, 102462.8, 102442.7, 102422.6, 
    102403.7, 102377.5, 102354.6, 102320.1, 102283.8, 102239.9, 102192.1, 
    102140.2,
  102502, 102491.1, 102473.8, 102460.4, 102442.9, 102424, 102408.8, 102389, 
    102371.4, 102344.3, 102315.7, 102285.6, 102248.9, 102208.3, 102163.6,
  101468.6, 101469.6, 101491.1, 101511.1, 101539.6, 101582.8, 101618.7, 
    101667.6, 101718.3, 101764, 101807.1, 101845.6, 101881.5, 101916.1, 101940,
  101539.1, 101550.8, 101573.8, 101599.9, 101634.8, 101676.8, 101715.5, 
    101765.2, 101814.6, 101861.2, 101902.4, 101937.9, 101973, 102004.4, 
    102029.9,
  101617.5, 101644.1, 101663.8, 101694.6, 101727.8, 101768.4, 101810.3, 
    101857.7, 101903.2, 101949.1, 101985.9, 102022.3, 102053.5, 102085.3, 
    102108.4,
  101684.2, 101706.3, 101727.4, 101761.5, 101796.9, 101844.5, 101883.9, 
    101937.1, 101985, 102026.9, 102065, 102101.8, 102136.4, 102158.2, 102178.5,
  101728.9, 101754.7, 101786.1, 101824.8, 101861.7, 101905.3, 101945.3, 
    101998.5, 102043.6, 102087.9, 102127.3, 102164.5, 102196.3, 102222.9, 
    102239.7,
  101775.1, 101799.1, 101833.6, 101871, 101913.5, 101954.4, 101999.9, 
    102047.7, 102095.8, 102138, 102176.3, 102212, 102241.2, 102271.6, 102292.1,
  101801.9, 101829.9, 101871.1, 101904.1, 101947.5, 101983.3, 102029.4, 
    102080.4, 102131.8, 102176.6, 102213.5, 102249.8, 102277.4, 102302.6, 
    102327.1,
  101827.4, 101861.7, 101904.8, 101935.5, 101974.6, 102010.6, 102053.9, 
    102107.7, 102158.1, 102202.2, 102239.6, 102275.6, 102298.1, 102325.1, 
    102349.9,
  101849.9, 101886.6, 101927.4, 101960.9, 101993.8, 102023.8, 102068.5, 
    102116.1, 102165, 102214.9, 102251.4, 102287.1, 102308.7, 102335.9, 
    102358.6,
  101869.4, 101907.4, 101948.6, 101981.5, 102014, 102040.9, 102076.1, 102112, 
    102160.2, 102203.3, 102247, 102283.2, 102307.6, 102331.7, 102354.1,
  101649.9, 101603.2, 101588, 101559.8, 101530, 101484.6, 101433, 101376.4, 
    101312.2, 101239.3, 101170.9, 101106.9, 101057.1, 101016, 100975.3,
  101654.6, 101628.3, 101609.6, 101585.6, 101550.8, 101516.8, 101471.5, 
    101418.6, 101368.5, 101314.9, 101264.8, 101210.9, 101163.7, 101121.4, 
    101080.7,
  101636.4, 101623.6, 101605.3, 101587.6, 101566.1, 101539, 101509.9, 
    101465.4, 101421.1, 101373.2, 101330.8, 101287.1, 101251.8, 101217.6, 
    101191.8,
  101644.3, 101630.3, 101609, 101599.4, 101582.5, 101558.4, 101537.9, 
    101509.3, 101480.6, 101443.6, 101416.3, 101385.8, 101363.1, 101331.9, 
    101304.4,
  101642, 101623.7, 101615.6, 101601.3, 101586.4, 101575.3, 101559.3, 
    101544.1, 101527.4, 101505.4, 101481.5, 101460.4, 101440.6, 101422.9, 
    101408.4,
  101638.9, 101630.4, 101618.2, 101616, 101602.6, 101593.2, 101581.4, 
    101570.3, 101563.2, 101552.6, 101547.2, 101540.9, 101529.7, 101517.9, 
    101506.7,
  101625.7, 101617.7, 101613.7, 101606.8, 101596.7, 101594.9, 101589, 
    101591.2, 101585, 101591.6, 101594.7, 101594.5, 101594.5, 101598.8, 
    101600.7,
  101621.1, 101642, 101628.6, 101632.8, 101628.1, 101622.4, 101620.5, 
    101623.3, 101625.3, 101631.8, 101642.6, 101652.4, 101669.5, 101683.2, 
    101701,
  101582.2, 101612.7, 101612.1, 101619.5, 101630.3, 101631, 101636.2, 
    101646.3, 101658.5, 101666.7, 101672.8, 101686.1, 101699.2, 101717.4, 
    101736.4,
  101555.6, 101590.8, 101611.5, 101629.5, 101634, 101638.9, 101645.7, 101659, 
    101666.1, 101682.5, 101702, 101722, 101747.9, 101775.5, 101800.3,
  102193.7, 102185, 102185.5, 102193.2, 102194.7, 102189.5, 102183.1, 
    102178.5, 102163.5, 102148.6, 102141.4, 102130.8, 102107.5, 102080.5, 
    102044.9,
  102162.1, 102157.5, 102149.8, 102170, 102168.6, 102164.8, 102163.7, 
    102161.3, 102157.9, 102150.4, 102140.7, 102131.3, 102113.2, 102097.8, 
    102076.3,
  102131, 102114.6, 102111.1, 102124.5, 102143, 102144, 102135.8, 102135.9, 
    102133.9, 102134.2, 102127.7, 102125.7, 102122.6, 102106.2, 102082.4,
  102093.5, 102077.3, 102074.5, 102089.4, 102099.3, 102115.1, 102113.5, 
    102116.4, 102121.9, 102118.8, 102119.1, 102117.2, 102115.8, 102104.3, 
    102089.2,
  102055.4, 102045.9, 102033, 102037.1, 102054, 102066.7, 102069.1, 102083.9, 
    102094.4, 102100.3, 102103.5, 102098.9, 102098.3, 102090.6, 102076,
  102019.7, 102010.2, 102000.8, 102008.6, 101997.4, 102000.1, 102012.2, 
    102030.5, 102046, 102061.5, 102074.9, 102079.9, 102083, 102083.5, 102075.9,
  101992.4, 101974, 101965.4, 101952.7, 101941.1, 101939.6, 101944.6, 
    101960.1, 101978.1, 101997.9, 102016.1, 102026, 102036.5, 102043.5, 
    102040.3,
  101947.8, 101936.6, 101919.8, 101896, 101856.8, 101844.4, 101848, 101869.1, 
    101885.8, 101912.5, 101935.8, 101957, 101976, 101990.8, 101999.8,
  101918.4, 101892.2, 101862.1, 101824.8, 101786.1, 101768.4, 101764.3, 
    101780, 101788.8, 101814.9, 101833.3, 101863.1, 101889.2, 101909.8, 
    101922.2,
  101879, 101843.2, 101814.7, 101768.9, 101715.5, 101681.3, 101673, 101684.7, 
    101694.3, 101734.5, 101754.6, 101780.8, 101786.1, 101812.8, 101843.7,
  102036.2, 102089, 102118, 102150.6, 102175.6, 102193.9, 102208.9, 102227.2, 
    102240.8, 102254.8, 102248.6, 102249, 102244.4, 102255.7, 102252.5,
  102007, 102051.8, 102084.6, 102114.6, 102140.9, 102166.2, 102186.4, 102207, 
    102219.9, 102241.4, 102267.2, 102288.3, 102288, 102301.9, 102310.8,
  101972, 102020.7, 102056.5, 102091.7, 102118.5, 102142.5, 102167.3, 
    102178.7, 102200.4, 102228.5, 102249.3, 102269.9, 102285.2, 102295.3, 
    102296.5,
  101935.4, 101982.4, 102019.7, 102052.2, 102074.4, 102103.4, 102129.5, 
    102154.7, 102179.5, 102201.1, 102225.5, 102247.9, 102272.8, 102280.1, 
    102292.9,
  101901.9, 101945.9, 101983.6, 102019.5, 102045.7, 102075, 102094.7, 
    102120.1, 102138.5, 102155.3, 102171, 102189.1, 102196.9, 102195.5, 
    102190.9,
  101870.6, 101906.7, 101947.2, 101979, 102006.5, 102029.5, 102049.9, 
    102066.3, 102081.6, 102095.6, 102102.3, 102101.1, 102100.8, 102102.4, 
    102104,
  101835.7, 101870.9, 101906.1, 101937.5, 101972.2, 101987.5, 102002.5, 
    102012.1, 102017.4, 102017.3, 102008.7, 102002.6, 101997.2, 101993.4, 
    101994.6,
  101822.1, 101838.2, 101864.3, 101885.1, 101909.1, 101927.5, 101933, 
    101942.1, 101934.1, 101932, 101913.1, 101902.3, 101879.9, 101866.9, 
    101869.7,
  101808.9, 101810.3, 101831.3, 101847.9, 101861.6, 101876.1, 101872, 
    101870.8, 101858.2, 101840, 101805.4, 101780, 101732.6, 101727.3, 101743.6,
  101768.9, 101787.3, 101797.5, 101800.6, 101806, 101806.6, 101802.3, 
    101790.9, 101758.3, 101704.5, 101664.8, 101631.5, 101616.4, 101615.3, 
    101598.7,
  101709.5, 101760.6, 101806.5, 101839.6, 101868.1, 101894.5, 101907.2, 
    101920.6, 101935.1, 101939.8, 101926.1, 101921.5, 101896.8, 101874.2, 
    101858.5,
  101728.4, 101775.3, 101831.8, 101867.3, 101888.4, 101906.2, 101926, 
    101941.8, 101949.3, 101962, 101961, 101952.3, 101930.6, 101909.7, 101889.2,
  101711.7, 101755.2, 101820.2, 101861.7, 101905.4, 101927.5, 101944.8, 
    101952, 101963.4, 101981, 101980.2, 101976.9, 101947, 101922.4, 101898.3,
  101696.4, 101738.7, 101805, 101849.1, 101892.9, 101921.4, 101942.8, 
    101963.6, 101978.4, 101987.8, 101984.8, 101973.5, 101949.6, 101917.6, 
    101890.6,
  101646.6, 101690.1, 101754.8, 101819.9, 101876.9, 101916, 101942.8, 
    101962.3, 101976.8, 101977.8, 101972.2, 101956, 101929.6, 101890.2, 
    101849.3,
  101618.8, 101662, 101687.4, 101757.4, 101809.8, 101876.1, 101912.5, 101942, 
    101957.3, 101956.9, 101944.6, 101919.9, 101883.1, 101840.2, 101792.9,
  101520.8, 101640.8, 101649.7, 101725.7, 101760.4, 101824.4, 101877.4, 
    101913.8, 101928.5, 101929, 101913.5, 101881.5, 101835.3, 101782, 101717.5,
  101295.6, 101493.8, 101540.1, 101635.8, 101684.1, 101760.3, 101814.3, 
    101864.1, 101894.7, 101891.9, 101867.1, 101828.2, 101779.8, 101718.5, 
    101630.8,
  101081.2, 101310.5, 101430.9, 101552, 101622, 101702.7, 101762, 101828.1, 
    101843.5, 101863.3, 101848.3, 101804.6, 101738.9, 101657.5, 101559.1,
  100973.7, 101110.9, 101290.4, 101450.2, 101543.8, 101643.5, 101704.7, 
    101773.8, 101810.6, 101815.9, 101785.4, 101753.8, 101699.8, 101609.1, 
    101514.5,
  101485.8, 101503.9, 101540, 101570.8, 101608.3, 101638.9, 101659.6, 
    101678.7, 101694.5, 101706.6, 101715.6, 101720.6, 101726.1, 101727.1, 
    101725,
  101550.5, 101567.2, 101612.8, 101639.1, 101669, 101695.2, 101723.5, 
    101751.8, 101773.6, 101790.8, 101805.5, 101817.8, 101823.7, 101826.4, 
    101823,
  101571.3, 101580.9, 101618.6, 101650.3, 101687.4, 101719.2, 101749.4, 
    101779.8, 101806.8, 101829.8, 101849.4, 101865.6, 101875, 101879.9, 
    101884.5,
  101577.4, 101592, 101624.2, 101660.4, 101691.4, 101725.8, 101762, 101797.8, 
    101832, 101860.2, 101886.2, 101902.7, 101920.7, 101924.5, 101922.5,
  101563.8, 101566.9, 101592.1, 101625.8, 101664.1, 101702.4, 101740.5, 
    101776.5, 101813.5, 101847.7, 101874.3, 101900.3, 101925.5, 101945, 
    101946.6,
  101526.3, 101545.2, 101548.4, 101575, 101609, 101654.7, 101699.7, 101748.4, 
    101788.9, 101827.3, 101860.8, 101887.2, 101911.9, 101930.5, 101937.1,
  101470.1, 101494.2, 101486.1, 101518.3, 101549, 101588.5, 101633.8, 
    101683.5, 101733.4, 101779.7, 101818.8, 101851.4, 101874.3, 101891.1, 
    101894.7,
  101346.9, 101382.8, 101377.1, 101424.5, 101451.7, 101500.2, 101553, 
    101616.8, 101670.2, 101727.4, 101774.4, 101819.2, 101847.9, 101866.4, 
    101869.4,
  101201.4, 101221.7, 101241, 101282.8, 101333.9, 101409.7, 101465.7, 
    101527.8, 101582.8, 101643.3, 101697.2, 101743.9, 101778.4, 101803.6, 
    101813.4,
  101138.8, 101073.6, 101086.8, 101142.4, 101181.9, 101266.5, 101354.9, 
    101438.7, 101512.3, 101585.4, 101643.9, 101703.2, 101752, 101769.7, 
    101784.8,
  101473.1, 101440.5, 101416.8, 101397, 101376.6, 101363.8, 101352.9, 
    101345.6, 101342.1, 101345.2, 101350.5, 101364, 101384.3, 101409.2, 
    101437.8,
  101531.4, 101499.5, 101484.2, 101469.9, 101461.7, 101450.4, 101441.4, 
    101435.4, 101435.7, 101441.9, 101452.1, 101471.6, 101501, 101535.7, 
    101566.1,
  101581.6, 101555.7, 101542.3, 101531.9, 101519.2, 101510.6, 101507.3, 
    101508.2, 101511, 101521.5, 101534, 101557, 101585.2, 101616.6, 101646,
  101621.3, 101605.1, 101593.2, 101583.1, 101574.7, 101570.2, 101566.3, 
    101567.8, 101571.6, 101581.2, 101596.6, 101619.5, 101648.2, 101679, 
    101704.8,
  101659.3, 101651, 101640.4, 101626.3, 101615.4, 101608.4, 101602.5, 101601, 
    101605.7, 101616.1, 101631.4, 101652.6, 101678.4, 101708.2, 101731.6,
  101681.4, 101670.4, 101660.6, 101649.1, 101638, 101627.6, 101619.8, 
    101615.9, 101621.2, 101630.6, 101649.6, 101667.6, 101687.3, 101713, 101731,
  101695.8, 101676.8, 101666.6, 101651.2, 101636.7, 101620.5, 101616.3, 
    101611, 101612.3, 101624.1, 101651.9, 101659.9, 101679.9, 101702, 101719.1,
  101694.5, 101669.8, 101655.7, 101635.3, 101615.1, 101602, 101592.9, 
    101592.7, 101597.3, 101604, 101621.2, 101633.4, 101658.3, 101669.9, 
    101686.5,
  101685.8, 101657.2, 101634.7, 101605.3, 101577.3, 101569.7, 101578.3, 
    101567.6, 101576.5, 101581.8, 101591.7, 101604.6, 101614.1, 101629.7, 
    101643,
  101672.1, 101635, 101606.1, 101567.4, 101541.8, 101538.4, 101533.8, 
    101535.8, 101540.1, 101551.5, 101550.6, 101561.6, 101564.4, 101577, 101598,
  102020.6, 102093.6, 102119.5, 102145.6, 102137.9, 102110.5, 102081, 102052, 
    102008.5, 101962.6, 101904, 101841.9, 101773, 101699.4, 101626.4,
  102027.6, 102053.7, 102072, 102075, 102085.9, 102087.1, 102076.3, 102050.4, 
    102012.9, 101973.5, 101923.6, 101870, 101808.2, 101743.4, 101677,
  102019, 102013.8, 102050.2, 102062.7, 102069.7, 102058.9, 102046.7, 
    102027.4, 102001.8, 101972, 101936.4, 101888.4, 101838.6, 101786.9, 
    101731.9,
  102001.5, 101998, 102016.8, 102023.1, 102031.9, 102032.3, 102026.6, 
    102019.2, 101993.9, 101968, 101941, 101907.2, 101860.6, 101815.4, 101772.3,
  101993.5, 102008.2, 102010.1, 102011.6, 102021.2, 102014.8, 102010.1, 
    102002.4, 101986, 101968.6, 101948.1, 101920.5, 101885.7, 101843.3, 
    101805.8,
  101985.6, 102004.2, 102015.3, 102019.9, 102023, 102017, 102010, 102000, 
    101980.9, 101967.6, 101951.7, 101928.8, 101904, 101871.5, 101837.9,
  101971.5, 101993.2, 102011.1, 102021, 102029.1, 102023.3, 102018.2, 102006, 
    101995.6, 101977.6, 101961.9, 101943.3, 101917.9, 101888.6, 101857.3,
  101945.1, 101963, 101999.6, 102000, 102022.6, 102028.9, 102035.6, 102020.5, 
    102012.5, 101992.1, 101978.3, 101960.4, 101949.3, 101928.1, 101896.2,
  101922.4, 101940.7, 101970.5, 101964, 101985.8, 102004.3, 102015.8, 
    102014.7, 102009.4, 102020.5, 102000.8, 101981.6, 101966, 101947.2, 
    101920.4,
  101881, 101900.6, 101920.6, 101918.8, 101937.6, 101966, 101991.1, 101999.6, 
    102015.9, 102025.5, 102018.3, 102004.9, 101986.1, 101977.5, 101950.5,
  102449.6, 102549.7, 102611, 102652.7, 102673.6, 102703.4, 102711.6, 
    102713.3, 102695.8, 102657.8, 102610.6, 102543.5, 102464, 102381.4, 
    102298.8,
  102415.8, 102497.3, 102536.6, 102576.1, 102633.2, 102647.2, 102661.5, 
    102654.9, 102635.6, 102610.3, 102568, 102512.8, 102443.8, 102364.7, 
    102280.8,
  102351.9, 102436.7, 102503.3, 102546, 102571.5, 102601.1, 102614.5, 
    102613.9, 102606.4, 102581.2, 102545.5, 102497.1, 102436.3, 102366.7, 
    102289.3,
  102311.8, 102366.2, 102430.4, 102487, 102516.6, 102542.3, 102548.8, 
    102563.9, 102551.8, 102541.7, 102514.4, 102472.6, 102424.2, 102365.2, 
    102298.7,
  102255, 102301.6, 102355.4, 102414.1, 102458.8, 102493.3, 102513.3, 
    102527.7, 102520.8, 102499.9, 102485.1, 102453.1, 102412.4, 102361.1, 
    102305.3,
  102185, 102242.3, 102289.6, 102335.2, 102380.1, 102412.9, 102444.5, 
    102460.6, 102463.6, 102456.8, 102450, 102423.1, 102394.9, 102354.9, 
    102308.6,
  102117.2, 102159.6, 102209.8, 102256.9, 102313.7, 102341.2, 102366.3, 
    102386.3, 102395.2, 102401.8, 102402.9, 102385.1, 102370.5, 102333.9, 
    102296.5,
  102056.2, 102083.8, 102141.4, 102186.8, 102231.7, 102276.5, 102313.1, 
    102325.4, 102336.5, 102339.3, 102340.9, 102332.2, 102318.7, 102302.6, 
    102277,
  102002, 102008.1, 102053, 102114.8, 102179.4, 102213.1, 102236.4, 102257.1, 
    102274.5, 102289.2, 102286.4, 102280.7, 102270.2, 102253.8, 102233,
  101968.9, 101970, 102011.6, 102081.3, 102154.7, 102176.4, 102194.8, 
    102228.5, 102252.2, 102266.8, 102266.1, 102251, 102231.3, 102217.1, 
    102201.7,
  102644.4, 102721.8, 102783.1, 102832.1, 102862.5, 102886.6, 102897.1, 
    102898.3, 102894.1, 102876.8, 102851.7, 102818.7, 102777.1, 102731.8, 
    102684.2,
  102606.5, 102672.4, 102717.8, 102768.6, 102814.3, 102837.1, 102846.6, 
    102846.1, 102834.3, 102812.3, 102781.7, 102737.7, 102690.7, 102632.5, 
    102560.8,
  102549.6, 102620.9, 102677.4, 102719.4, 102754.5, 102771.2, 102779.5, 
    102778.4, 102771.3, 102752.1, 102718.2, 102669.6, 102605.2, 102526, 
    102428.4,
  102482.4, 102553.9, 102605.4, 102651.4, 102683.7, 102713.9, 102722.3, 
    102720.2, 102709.7, 102688, 102651.1, 102601.7, 102537.5, 102457.4, 
    102364.8,
  102405.1, 102482.8, 102530.8, 102579.6, 102610.4, 102633.9, 102649.1, 
    102654.9, 102644.9, 102625.3, 102594, 102544.3, 102482.3, 102409.4, 
    102325.6,
  102322.5, 102395.3, 102448, 102496.6, 102530.6, 102560.3, 102577.4, 
    102584.6, 102583.2, 102566.9, 102538.9, 102495.1, 102439.1, 102373.4, 
    102300.2,
  102234.9, 102297.5, 102349.4, 102394.9, 102430, 102460.8, 102489.2, 
    102504.4, 102507.9, 102500.2, 102479.6, 102441.3, 102396.5, 102339.7, 
    102274.2,
  102166.9, 102216.2, 102262.6, 102305.8, 102345.1, 102378.1, 102403.2, 
    102422.9, 102432.2, 102432.8, 102419, 102392.9, 102353.7, 102306.6, 
    102251.9,
  102088.5, 102129.4, 102165.5, 102191.1, 102223.2, 102260.8, 102297.5, 
    102323, 102345.4, 102350.8, 102348.7, 102329.8, 102307.1, 102269, 102219.4,
  102028.4, 102049.6, 102081.6, 102112.8, 102136, 102155.6, 102191.4, 
    102217.8, 102247.2, 102259.2, 102265.6, 102260.4, 102243.8, 102214.8, 
    102181,
  102763.4, 102829.9, 102872.9, 102914.7, 102947.7, 102975.8, 102994.7, 
    103008.9, 103025.2, 103037.8, 103048.7, 103055.9, 103048.5, 103040.3, 
    103029.2,
  102712.4, 102775.2, 102820.7, 102860.6, 102891.2, 102918.9, 102938.1, 
    102953.9, 102969.1, 102974.7, 102979.9, 102973.9, 102958.8, 102935.3, 
    102908.8,
  102649.1, 102709.6, 102755.8, 102797.3, 102824.1, 102849.9, 102868.7, 
    102885.3, 102893.8, 102895.2, 102888.6, 102871.7, 102843.1, 102811.2, 
    102776.9,
  102584, 102643.1, 102690.9, 102730.3, 102758.3, 102782.8, 102800, 102814.3, 
    102817.7, 102812.6, 102794.2, 102769.3, 102733.6, 102696, 102654.4,
  102512.2, 102568.5, 102615.2, 102654, 102681.5, 102706.7, 102723.5, 
    102735.5, 102735.8, 102725.2, 102701.4, 102668.5, 102628.9, 102584.4, 
    102537.8,
  102442, 102496.2, 102539.6, 102577.9, 102605.4, 102627.3, 102641.9, 
    102652.6, 102653, 102640.4, 102613.2, 102574.1, 102529.5, 102484.1, 
    102430.6,
  102367.6, 102422.1, 102463.9, 102500.1, 102526.4, 102546.2, 102559.8, 
    102568.6, 102567, 102555.4, 102526.9, 102486.7, 102440.2, 102388.5, 
    102327.3,
  102290, 102344.8, 102381.1, 102418.4, 102444.3, 102464.3, 102478.6, 102485, 
    102483.3, 102471.9, 102444.5, 102403.3, 102355, 102297.9, 102232.8,
  102220.2, 102268.1, 102301, 102338.6, 102362.4, 102385.4, 102398, 102403.6, 
    102402.1, 102389.3, 102364.5, 102327, 102276.2, 102213.8, 102142.4,
  102138, 102183.2, 102217.8, 102255.4, 102277.2, 102304, 102315.3, 102323.2, 
    102319.6, 102310.4, 102288, 102249.8, 102199.7, 102135.4, 102064.1,
  102501.3, 102587.3, 102657.5, 102721.7, 102786.4, 102830.2, 102867.1, 
    102893.8, 102907.6, 102911.1, 102899.9, 102889.5, 102879.7, 102864.3, 
    102843,
  102486.4, 102562.6, 102632.7, 102694.4, 102753.5, 102798.2, 102836.6, 
    102860.6, 102867.4, 102866.8, 102850.5, 102835.9, 102815.3, 102786.8, 
    102756.3,
  102464.4, 102539, 102609.4, 102668.2, 102718.9, 102757, 102781.8, 102802.9, 
    102809, 102804.1, 102786.9, 102767, 102739.8, 102702.6, 102659.3,
  102436, 102507.2, 102574.5, 102632.8, 102682.7, 102717.7, 102738.6, 
    102753.8, 102753.9, 102747.9, 102727.2, 102701.6, 102662.9, 102614.5, 
    102556.5,
  102408.1, 102475.6, 102535.6, 102591.8, 102638.5, 102672.8, 102689, 
    102697.2, 102692.7, 102683.2, 102659.7, 102626.1, 102579.2, 102521.8, 
    102452.6,
  102375.8, 102442.2, 102493.6, 102549.8, 102589.5, 102621.3, 102636.4, 
    102643.2, 102634.7, 102622, 102592.1, 102549, 102497.9, 102433.6, 102350.1,
  102344, 102405.4, 102449.4, 102497.2, 102533.1, 102562.5, 102575.6, 
    102582.5, 102570.7, 102552.2, 102518.4, 102478.3, 102420.8, 102346.9, 
    102251.2,
  102310.8, 102366.9, 102404.4, 102449.4, 102478.2, 102504.7, 102517.9, 
    102521.2, 102510.6, 102486.8, 102453.2, 102409.2, 102344, 102266.8, 102166,
  102279.4, 102324.1, 102357.8, 102396.2, 102422.2, 102447.2, 102457.8, 
    102460.2, 102446.4, 102421.3, 102388.4, 102341.1, 102277.2, 102194.5, 
    102090,
  102242.5, 102279.6, 102310.9, 102340.1, 102364.7, 102386.2, 102395.5, 
    102391.5, 102380.8, 102359.5, 102324.6, 102275, 102210.6, 102128.9, 
    102025.7,
  102227, 102297.4, 102377.8, 102443.1, 102505.6, 102541.9, 102573.1, 
    102586.8, 102592.9, 102590, 102578.3, 102573.7, 102563.1, 102561.7, 
    102549.2,
  102273.8, 102337.4, 102404.6, 102453.8, 102507.4, 102552.7, 102587.3, 
    102595.3, 102585.6, 102579.2, 102564.4, 102543.2, 102525.7, 102508, 102479,
  102288.7, 102346.9, 102424.1, 102480.1, 102531.2, 102552.1, 102577.6, 
    102587.6, 102572.9, 102561.6, 102536.5, 102515.9, 102487.9, 102456.4, 
    102413.4,
  102304.4, 102362.7, 102430.4, 102476.3, 102527.6, 102554.3, 102570.4, 
    102578.4, 102556.5, 102531.5, 102502.8, 102474.6, 102438.9, 102395.9, 
    102344.8,
  102306.1, 102363.7, 102427.5, 102483.3, 102519.3, 102541.6, 102545.9, 
    102552.6, 102533.8, 102504.7, 102467.2, 102432.5, 102387.4, 102338.7, 
    102281.7,
  102305.5, 102358.8, 102418.9, 102469.8, 102508.7, 102532, 102527.6, 
    102530.8, 102506.8, 102478.3, 102432.1, 102382.6, 102330.3, 102274.3, 
    102211,
  102297.1, 102348.1, 102404.2, 102448.9, 102486.7, 102503.7, 102502.8, 
    102500.5, 102473.2, 102439.2, 102388.7, 102338.3, 102279.5, 102220, 
    102146.5,
  102290.6, 102333.4, 102387.1, 102429.3, 102458.3, 102471.1, 102476.7, 
    102470.6, 102435.4, 102400.1, 102346.6, 102292.4, 102230, 102159.2, 
    102081.6,
  102283.6, 102316.9, 102364.1, 102404.1, 102436.9, 102449.3, 102444.3, 
    102434.8, 102406.6, 102364.6, 102309.4, 102253, 102184.1, 102108.9, 
    102022.8,
  102271.6, 102304.2, 102337.5, 102363.9, 102390.7, 102409.1, 102412.7, 
    102406, 102378, 102336, 102279.3, 102217, 102142.5, 102058, 101967.7,
  101830.2, 101795.2, 101774.4, 101752.9, 101745.2, 101737.8, 101754.8, 
    101768.6, 101771.4, 101782.6, 101795.3, 101814.3, 101838.3, 101866.7, 
    101899.6,
  101898.3, 101874.8, 101875.2, 101864.7, 101859.5, 101858.4, 101864.1, 
    101879.7, 101889.6, 101900.9, 101919.9, 101933.6, 101947.3, 101960.8, 
    101964.6,
  101956.9, 101954.9, 101959.6, 101956, 101949.8, 101958.6, 101974.8, 
    101984.2, 101992.7, 102000.4, 102003.5, 102012.4, 102016.4, 102015.8, 
    102011.2,
  102012.3, 102023.1, 102035, 102045, 102045, 102059.9, 102068.1, 102082.8, 
    102089.5, 102086.8, 102091.3, 102087.4, 102089.7, 102076, 102050.6,
  102063.3, 102085.6, 102102.7, 102114.9, 102129.6, 102146, 102148.4, 
    102153.5, 102167.5, 102162.7, 102157.2, 102147.2, 102141.8, 102118.8, 
    102078,
  102105.4, 102137.1, 102161.7, 102179.2, 102201.4, 102216.3, 102222.6, 
    102223.8, 102236.9, 102227, 102216.3, 102196.7, 102176.6, 102145.5, 
    102096.9,
  102144.2, 102180.8, 102206.4, 102231.4, 102257, 102266.8, 102277.9, 102293, 
    102289.2, 102270.2, 102252.8, 102233.9, 102201.7, 102165.3, 102112.8,
  102179.6, 102211.2, 102241.5, 102270.4, 102293.5, 102301.2, 102319.7, 
    102332.8, 102319.6, 102301.7, 102282.7, 102253.5, 102216.8, 102177.9, 
    102119.3,
  102211.8, 102238.7, 102267.2, 102293.9, 102317.2, 102333.2, 102345.1, 
    102367.7, 102349.1, 102316.6, 102288.8, 102258.2, 102228.1, 102180.3, 
    102123.3,
  102235.9, 102259, 102290, 102311.6, 102338.9, 102367.4, 102387.8, 102388.2, 
    102357.4, 102332.9, 102306.6, 102276.4, 102241.3, 102194.6, 102128.2,
  102056.5, 102011.2, 101924.9, 101837.7, 101738.5, 101653.7, 101562.3, 
    101485, 101411.4, 101358.1, 101311.5, 101275.6, 101255, 101231.8, 101226.2,
  102103.5, 102043.6, 101957.1, 101893, 101805.8, 101725.3, 101644.8, 
    101571.3, 101501, 101437.1, 101381.6, 101337.1, 101306, 101297.1, 101302,
  102107.6, 102052.2, 101992.6, 101928.3, 101850.1, 101773.6, 101695.7, 
    101626.4, 101562.8, 101506.7, 101460.3, 101418, 101396.2, 101369.5, 
    101378.8,
  102120.5, 102066.6, 102025.2, 101970.4, 101903.4, 101835.8, 101766.6, 
    101696, 101629.5, 101571.9, 101528.5, 101492.3, 101463.7, 101453.7, 
    101452.9,
  102121.3, 102085.1, 102041.5, 101997.6, 101945, 101882.2, 101821.5, 
    101758.5, 101696.7, 101639.6, 101589.4, 101558.8, 101537.7, 101532.6, 
    101533.9,
  102131.4, 102096.6, 102064.4, 102029.2, 101983.2, 101931.7, 101881.5, 
    101821.9, 101768.3, 101714.4, 101666.4, 101626.1, 101603.4, 101603.2, 
    101605.9,
  102141.2, 102122.1, 102092.2, 102058.9, 102017.1, 101975.5, 101929.4, 
    101881.7, 101834.4, 101789.3, 101747.4, 101717.9, 101688.9, 101684.3, 
    101692.9,
  102152.2, 102141.4, 102119.7, 102094.3, 102056.2, 102022.3, 101980.9, 
    101940, 101906.2, 101870.5, 101837.5, 101813.8, 101793, 101783.2, 101792.3,
  102169.1, 102167, 102147.9, 102128.7, 102099.8, 102068.7, 102037.2, 
    102008.9, 101978.6, 101954.6, 101930.7, 101914.3, 101896, 101892.3, 
    101891.8,
  102200.8, 102189.9, 102178.4, 102162.4, 102141.4, 102120.6, 102092.1, 
    102073.7, 102057.1, 102038.2, 102023.5, 102008.2, 102003.3, 101998.5, 
    102000.6,
  102177, 102109, 102006.4, 101908.1, 101801, 101713.1, 101621.9, 101520.7, 
    101433.4, 101345.4, 101303.7, 101301.3, 101333.7, 101400.1, 101488.7,
  102215.1, 102167.6, 102083.6, 102001.4, 101904.2, 101806.7, 101718, 
    101632.5, 101568.5, 101509.9, 101466.7, 101447.7, 101469.8, 101517.9, 
    101579.6,
  102259.7, 102225, 102170.5, 102102.4, 102017.2, 101929.6, 101846.1, 
    101766.3, 101694, 101635.5, 101595.8, 101579.9, 101590.5, 101621.1, 
    101669.3,
  102292.7, 102258, 102226.5, 102174.5, 102111.2, 102038.8, 101968.8, 
    101898.6, 101835.4, 101784.7, 101749.5, 101730.7, 101733.3, 101750.5, 
    101787.1,
  102282.3, 102287.4, 102275.7, 102237.1, 102195.4, 102140, 102079.5, 
    102019.7, 101967.1, 101916.2, 101883.1, 101862, 101856.1, 101864.2, 
    101883.3,
  102279.8, 102283.3, 102285.9, 102270.7, 102247.6, 102211.7, 102169.4, 
    102121.9, 102079.9, 102043.5, 102014.2, 101990.1, 101975.9, 101973, 
    101973.7,
  102252, 102282, 102288.3, 102288.6, 102273.8, 102252, 102223.8, 102195.9, 
    102162.8, 102131.4, 102104.5, 102082.9, 102069.1, 102054.6, 102046.7,
  102249.7, 102279.2, 102274.2, 102282.5, 102289.3, 102279.5, 102260.7, 
    102237.4, 102214.2, 102190.3, 102168.4, 102152.1, 102135.4, 102119, 
    102104.6,
  102223, 102246.4, 102278.5, 102282.1, 102275.6, 102286.5, 102280.2, 
    102261.9, 102238.5, 102221.1, 102200, 102181.9, 102163.6, 102149.6, 
    102138.2,
  102221, 102227.6, 102263.5, 102262.9, 102271.2, 102275.5, 102272.7, 
    102272.7, 102262.6, 102243.4, 102230.9, 102216.7, 102203.3, 102189.3, 
    102175.6,
  101842.9, 101879.2, 101897.4, 101908, 101918.4, 101911.6, 101875.1, 
    101805.5, 101720.4, 101614.2, 101487.7, 101355.7, 101236.5, 101138.5, 
    101064.8,
  101864.7, 101903.2, 101929.8, 101943.1, 101945.4, 101943.4, 101933.9, 
    101893.8, 101824.1, 101738, 101638, 101537.2, 101434.7, 101352, 101291.9,
  101885.4, 101929, 101966.6, 101987.7, 101989.4, 101985.4, 101974.9, 
    101959.4, 101923, 101860.3, 101783.5, 101702.3, 101623.5, 101547.4, 
    101481.4,
  101897.4, 101946.8, 101995.7, 102024.1, 102038.4, 102034.8, 102019.4, 
    102002.2, 101980.1, 101948.5, 101902.1, 101841.6, 101776, 101713.5, 
    101655.9,
  101903.1, 101960.2, 102007, 102046.9, 102075.4, 102084.3, 102081, 102061, 
    102040.2, 102011.9, 101981.8, 101943.4, 101898.4, 101850.7, 101802.7,
  101905.7, 101964.6, 102015.2, 102059.6, 102095.6, 102117.5, 102121.2, 
    102114, 102096.6, 102076.9, 102050.5, 102024.8, 101989.7, 101958.2, 
    101928.4,
  101910.9, 101958.6, 102011.1, 102054.4, 102105.3, 102140.2, 102155.4, 
    102160.2, 102154.8, 102139.1, 102121, 102100.8, 102075.7, 102052.6, 102029,
  101919.5, 101963.5, 102011, 102048.5, 102091.9, 102127.8, 102161.2, 
    102182.3, 102194.6, 102190, 102180, 102170.2, 102155.7, 102139, 102122.5,
  101928.7, 101969.6, 102007.1, 102042.4, 102082.3, 102119.1, 102153.2, 
    102192.3, 102206.1, 102216.1, 102219, 102215.9, 102209.8, 102200.9, 102191,
  101939.6, 101980.8, 102012.3, 102040.3, 102069.4, 102114.5, 102141.6, 
    102192.6, 102223.1, 102232.6, 102238.4, 102248.1, 102252.7, 102256.6, 
    102249,
  101580.4, 101559.1, 101531.1, 101517.1, 101505.9, 101501.9, 101498.7, 
    101503.9, 101505.8, 101511.8, 101515.5, 101512.3, 101510.3, 101503.4, 
    101481.8,
  101631.9, 101621.9, 101609.4, 101602.9, 101598.1, 101598.9, 101603.2, 
    101613.1, 101620.3, 101632, 101636.6, 101640.7, 101639, 101630.7, 101614.4,
  101684.8, 101679, 101674.9, 101675.2, 101679.2, 101686, 101701.3, 101715.8, 
    101732.7, 101744, 101754.2, 101762.9, 101761.7, 101758.6, 101749.8,
  101721.7, 101722.6, 101728.6, 101733.5, 101742.6, 101757.5, 101778.7, 
    101800.6, 101819.2, 101836.8, 101851.4, 101862.2, 101867.3, 101869.1, 
    101861.1,
  101755.3, 101761.8, 101773.1, 101784.9, 101799.8, 101816.7, 101840.9, 
    101868.8, 101894.1, 101919.6, 101937.3, 101951.9, 101962.7, 101968.5, 
    101969.9,
  101780.3, 101790.8, 101808, 101823.5, 101843.6, 101865.3, 101890.3, 
    101914.9, 101944.3, 101972.8, 101995.9, 102014.1, 102030.1, 102041.8, 
    102051.9,
  101802, 101815.6, 101835.5, 101857.5, 101877.2, 101900.7, 101923.4, 
    101950.9, 101978.2, 102008.4, 102036.8, 102059.9, 102082.5, 102103.2, 
    102120.2,
  101811, 101831.7, 101856.1, 101878.5, 101897.8, 101917, 101941.9, 101967.4, 
    101996.9, 102026.1, 102058.3, 102082.9, 102113.1, 102138.5, 102165.8,
  101821.9, 101843.1, 101870, 101897.9, 101913.5, 101932.7, 101949.8, 
    101975.2, 101998.7, 102028, 102056.6, 102087.4, 102131.1, 102161.6, 
    102198.2,
  101832.3, 101857.2, 101884.2, 101911.9, 101926.1, 101939.6, 101958.1, 
    101967.6, 101991.6, 102019.4, 102050, 102082.5, 102122.1, 102160.6, 
    102200.4,
  102680.1, 102648, 102606.6, 102568.5, 102524.8, 102480.3, 102428.3, 
    102377.7, 102320.9, 102259.3, 102182.1, 102097, 102007.1, 101914, 101819.1,
  102673.8, 102640.6, 102598.9, 102561, 102518.7, 102477.3, 102433, 102381.8, 
    102330.7, 102273.8, 102206.4, 102133.3, 102054.9, 101981, 101899.8,
  102658, 102630.4, 102593.2, 102551.9, 102513.9, 102473.5, 102434.5, 
    102387.6, 102336.8, 102283.9, 102225.7, 102168.3, 102098.2, 102030.8, 
    101960.5,
  102643, 102617.1, 102581.5, 102541.4, 102502.3, 102465.3, 102422.4, 
    102384.9, 102341.1, 102293.5, 102241.8, 102191.5, 102134.8, 102082.5, 
    102023.7,
  102616.2, 102598.2, 102563.7, 102528.2, 102488.3, 102451.3, 102412.8, 
    102375.7, 102333.3, 102293.4, 102250.1, 102208.1, 102160.4, 102117.9, 
    102065.8,
  102593.8, 102573.5, 102543.5, 102507.8, 102472.5, 102437.3, 102397.3, 
    102362.9, 102329.4, 102292, 102252.7, 102218, 102174.2, 102136.3, 102094.5,
  102567, 102541.2, 102512.8, 102484.4, 102449.6, 102418, 102380.7, 102346.3, 
    102309.7, 102278.7, 102247.1, 102214.3, 102179.8, 102148.8, 102114.6,
  102535.3, 102508.1, 102482.5, 102451.9, 102425.6, 102396.4, 102364.4, 
    102331.4, 102300.8, 102268.7, 102238.6, 102210.5, 102178.4, 102146.3, 
    102118.1,
  102497.5, 102470.6, 102447.1, 102417.2, 102391.7, 102367, 102341.5, 
    102316.1, 102287.2, 102254.7, 102227.8, 102196.8, 102168.1, 102138.9, 
    102110.4,
  102457.8, 102436.2, 102411.2, 102383, 102358, 102335.3, 102315.1, 102295.1, 
    102268.8, 102242.8, 102215.4, 102189.6, 102162.1, 102135.2, 102104.5,
  102502.4, 102560.5, 102601.1, 102649.1, 102678, 102699.6, 102706.4, 
    102681.7, 102641.4, 102594.2, 102537.4, 102472, 102398.5, 102317.7, 
    102218.7,
  102510.6, 102554.3, 102585.2, 102636.2, 102676, 102714.5, 102718, 102710.8, 
    102683.2, 102645.8, 102596.6, 102542.6, 102478.5, 102399.9, 102312.8,
  102501.3, 102540.3, 102569, 102623.7, 102672.1, 102705.6, 102727.3, 
    102731.7, 102717.8, 102696.6, 102656.1, 102607.6, 102552.9, 102488.5, 
    102411,
  102494.2, 102523.6, 102549.8, 102590, 102645.9, 102690, 102719, 102732.5, 
    102734.3, 102715.1, 102689.3, 102652.8, 102609.6, 102554.7, 102491.9,
  102476.7, 102500.8, 102528.4, 102552.4, 102600.6, 102655.3, 102692.2, 
    102716.5, 102729.6, 102723.5, 102712.1, 102687.7, 102657, 102608.7, 
    102552.7,
  102463.4, 102479.6, 102503.9, 102516.3, 102550.5, 102592.4, 102631.7, 
    102675.5, 102699.3, 102708.3, 102709.3, 102700.8, 102675.4, 102646.3, 
    102598.5,
  102448.1, 102454.4, 102477.4, 102481.4, 102501.2, 102536.8, 102577.3, 
    102609.2, 102646.3, 102665.3, 102673.4, 102674.8, 102666.7, 102649.4, 
    102614.1,
  102422.3, 102431.3, 102446.2, 102448.6, 102454.4, 102475.6, 102511.2, 
    102553.3, 102586.5, 102617, 102632.3, 102640.8, 102635.7, 102625, 102602.7,
  102399.6, 102406.4, 102410.1, 102414.4, 102428.4, 102434.9, 102454.3, 
    102482.8, 102514.8, 102549.6, 102574, 102584.6, 102587.5, 102582.5, 
    102573.1,
  102379.7, 102375.4, 102380.1, 102374.6, 102377.6, 102384.8, 102400.5, 
    102423, 102450.2, 102477.4, 102496.6, 102515.4, 102530.6, 102534.8, 
    102527.9,
  101264.2, 101323.4, 101386.5, 101476, 101581.4, 101692.9, 101773.4, 
    101850.4, 101907.7, 101960.2, 101993.4, 102012.2, 102033.7, 102070.7, 
    102061.9,
  101283.8, 101358.2, 101428.2, 101515.2, 101613.4, 101707.3, 101780.5, 
    101869.2, 101941.2, 101997.8, 102027.9, 102057.6, 102068.8, 102074.4, 
    102082.1,
  101320.6, 101393, 101452.9, 101532.5, 101622.6, 101723.4, 101809.4, 
    101892.4, 101963.3, 102029.3, 102074.9, 102101.2, 102114.2, 102120.4, 
    102112.1,
  101338.4, 101412.9, 101476.7, 101544.1, 101621.6, 101717.5, 101797.5, 
    101885.5, 101965, 102034, 102092.8, 102135.6, 102152.8, 102155.6, 102150.2,
  101360.8, 101431.6, 101493.4, 101548.1, 101617.9, 101708, 101792.6, 101880, 
    101956.1, 102031.8, 102106.5, 102161.1, 102199.4, 102202.6, 102192.7,
  101378.9, 101441.5, 101502.2, 101552.9, 101607.7, 101689.2, 101769.3, 
    101860.8, 101940.3, 102002, 102083.8, 102150.1, 102204.2, 102235.7, 
    102237.1,
  101397.3, 101461, 101512.9, 101555.7, 101596.9, 101667.9, 101763.2, 
    101837.6, 101922.1, 101981, 102053.4, 102124.2, 102189.3, 102240.6, 
    102266.2,
  101427.2, 101482.2, 101523.2, 101559.4, 101591.2, 101645.2, 101727.5, 
    101809, 101892.8, 101955, 102021.7, 102090.8, 102153.3, 102206.5, 102244.2,
  101453.8, 101498.9, 101539.4, 101568.4, 101595.9, 101632, 101710.8, 
    101777.4, 101859.7, 101922.3, 101986.6, 102058.5, 102114.6, 102172.6, 
    102218.1,
  101487.8, 101524.6, 101556.5, 101580.5, 101605.4, 101641, 101696.3, 
    101749.8, 101818.5, 101895.4, 101948.1, 102015.6, 102071.2, 102123.4, 
    102166.6,
  101046.9, 100989.5, 100955.9, 100932.1, 100918.1, 100914.6, 100923, 
    100946.3, 100985.6, 101040.5, 101111.4, 101187.8, 101276.8, 101364.8, 
    101448.3,
  101121.1, 101062.7, 101034, 100999.5, 100987.4, 100986.4, 101006.4, 
    101027.9, 101072.8, 101130.5, 101206.5, 101292.1, 101390.4, 101485.3, 
    101571,
  101185.1, 101135.3, 101100.5, 101075.3, 101063.7, 101066.5, 101069.3, 
    101108.9, 101155, 101228.7, 101292.6, 101388.5, 101468.1, 101560.5, 
    101643.9,
  101228.2, 101180.1, 101146.4, 101111.8, 101105.8, 101104.8, 101129.2, 
    101167.3, 101225.8, 101295.8, 101360.2, 101441.6, 101535.7, 101633.8, 
    101721.5,
  101259.3, 101205.2, 101180.1, 101174.8, 101175.1, 101187, 101196, 101223.2, 
    101261, 101330.7, 101405.4, 101489.2, 101581, 101677, 101770.1,
  101265.4, 101218.9, 101179.2, 101171.9, 101155.6, 101181.6, 101187.6, 
    101228.1, 101276.7, 101353.9, 101430.7, 101517.8, 101615.8, 101711.5, 
    101809.6,
  101254.2, 101197, 101133.4, 101111.1, 101098.6, 101125.4, 101141.4, 
    101213.4, 101273.2, 101356, 101442.2, 101536.3, 101630.3, 101728.4, 
    101828.9,
  101255.3, 101185.4, 101110.1, 101079.1, 101063.1, 101073.6, 101105.1, 
    101178, 101260.2, 101344.5, 101436.1, 101540, 101637, 101735.5, 101836.3,
  101305.2, 101235, 101159.5, 101119.7, 101087.9, 101092.1, 101116.3, 
    101184.7, 101258.9, 101351.9, 101431.4, 101544.7, 101635.5, 101733, 
    101828.7,
  101378.7, 101303.2, 101231, 101192.8, 101149.4, 101144.5, 101158.2, 101209, 
    101267.1, 101343, 101432.2, 101522.7, 101621.8, 101723.8, 101818,
  101892.6, 101795.5, 101692.7, 101603.4, 101516.2, 101446, 101381.8, 
    101329.1, 101274.9, 101226.2, 101176.9, 101124.5, 101078.5, 101034.6, 
    101000.4,
  101940, 101841.4, 101741.6, 101653.1, 101566.3, 101493.4, 101424.9, 
    101371.3, 101321.5, 101275.8, 101230.7, 101189.1, 101147.5, 101112.4, 
    101087.1,
  101980.8, 101883.3, 101785.3, 101690, 101602.2, 101522.5, 101454.2, 
    101397.9, 101346.4, 101303.7, 101262.4, 101228.5, 101203, 101182.7, 
    101168.4,
  102016, 101918.6, 101820.5, 101723.8, 101632.8, 101551.1, 101478.9, 
    101415.8, 101365.2, 101322.7, 101286.8, 101253.1, 101226.2, 101209.4, 
    101200.7,
  102049.2, 101953.2, 101852.2, 101754.5, 101662.5, 101578.4, 101499.6, 
    101434.9, 101381.5, 101327, 101294.8, 101264.6, 101238.2, 101231.7, 
    101235.5,
  102076.3, 101982.4, 101881, 101783.9, 101690, 101599.9, 101515.7, 101442.1, 
    101372.8, 101326.9, 101272.6, 101224.3, 101215.3, 101230.9, 101257.8,
  102103.9, 102011.5, 101909.7, 101813.5, 101718.6, 101621.8, 101525.2, 
    101426.3, 101339.4, 101278.4, 101222, 101203.3, 101199.2, 101228.7, 
    101280.2,
  102128.4, 102037.8, 101939.4, 101843.5, 101746.8, 101646.9, 101539.6, 
    101424, 101313.3, 101250.5, 101191.3, 101181.1, 101169.3, 101208.7, 
    101274.6,
  102153.3, 102064.7, 101969.7, 101874.8, 101777.2, 101674.3, 101564.4, 
    101451, 101341.3, 101270.5, 101221.6, 101195, 101180.7, 101202.1, 101280.3,
  102173.7, 102092.7, 101998.8, 101907, 101808.2, 101709.4, 101606, 101498.1, 
    101399, 101321, 101271.3, 101242.7, 101217.1, 101226.4, 101287.5,
  102429.9, 102356.8, 102280.5, 102203.1, 102125.7, 102043.4, 101959.5, 
    101870.9, 101778.8, 101683.8, 101590.2, 101494.7, 101400.9, 101305.6, 
    101212,
  102493.9, 102428.1, 102359.5, 102288.4, 102211.3, 102134.5, 102052, 
    101969.3, 101883, 101795.8, 101707, 101618.3, 101533.5, 101446.2, 101358.3,
  102552.3, 102492.9, 102430, 102362.3, 102290, 102215.9, 102140.1, 102061.1, 
    101980.3, 101897.2, 101814.3, 101729.7, 101646.8, 101566, 101482.6,
  102597.2, 102542.3, 102486.9, 102423.9, 102358.2, 102288.5, 102216.6, 
    102141.9, 102065.2, 101987.2, 101907.6, 101829, 101748.6, 101670.7, 
    101592.7,
  102632.8, 102582.1, 102530.6, 102472.6, 102412.2, 102346, 102278.5, 
    102207.6, 102135.2, 102060.5, 101984.8, 101908.2, 101831.7, 101754.7, 
    101676.2,
  102654.9, 102606.8, 102560.3, 102506.7, 102450.3, 102388.9, 102325.3, 
    102257.2, 102188.9, 102117.4, 102045, 101969, 101890.1, 101812.5, 101738.3,
  102666.2, 102620.9, 102576.5, 102525.4, 102473.6, 102415.4, 102353.8, 
    102288.4, 102222.4, 102154.9, 102083.2, 102008.9, 101929, 101850.1, 
    101773.6,
  102666.9, 102622.5, 102579.4, 102530.8, 102482.2, 102425.8, 102366, 
    102303.7, 102238.9, 102172.5, 102102.5, 102029.2, 101947, 101865.2, 
    101784.8,
  102659.8, 102614.9, 102570.9, 102522.4, 102475.9, 102420.4, 102362.5, 
    102303.4, 102240.7, 102175.5, 102106.5, 102036.5, 101956.4, 101867.8, 
    101777,
  102642.1, 102597.1, 102552.8, 102503.6, 102455.3, 102401.2, 102347.7, 
    102290.3, 102225.2, 102163.1, 102101.1, 102035.6, 101960.4, 101865.6, 
    101764,
  102403.1, 102367.8, 102321.1, 102264.4, 102196.2, 102118.2, 102031.1, 
    101934.1, 101820.9, 101695.2, 101558.1, 101417.8, 101263.6, 101109.3, 
    100954.8,
  102439.9, 102395.4, 102354.9, 102303.9, 102248, 102176.6, 102095.4, 
    102003.2, 101904.2, 101798.7, 101679.6, 101550.8, 101413.3, 101268.6, 
    101120.2,
  102486.8, 102437.7, 102399.7, 102349.2, 102291.3, 102229.1, 102157.3, 
    102078.9, 101988.6, 101886.6, 101774.9, 101657.7, 101534.6, 101405.7, 
    101268.6,
  102520.6, 102483.3, 102442.5, 102395.2, 102344.4, 102286.6, 102218.8, 
    102148.7, 102068.2, 101981.5, 101886.4, 101782.6, 101669.6, 101551.7, 
    101427.6,
  102553.4, 102522.4, 102484.9, 102440.5, 102388.4, 102335.3, 102272.4, 
    102203.4, 102132.1, 102052.4, 101964.9, 101873.6, 101773.8, 101669.7, 
    101557.4,
  102577.5, 102552.9, 102521.2, 102480.4, 102436.6, 102383.6, 102327.1, 
    102263.3, 102194.8, 102124.1, 102046.7, 101963.2, 101873.4, 101780.3, 
    101681.8,
  102590.1, 102567.7, 102544.5, 102513, 102474.4, 102428.1, 102373.5, 
    102313.1, 102251.2, 102183.6, 102112.3, 102039.7, 101956.9, 101872.1, 
    101782.9,
  102588.1, 102577, 102558.9, 102531.9, 102500.6, 102461.2, 102414.8, 102361, 
    102303.1, 102241.4, 102175.6, 102106.3, 102032.9, 101954.7, 101873.9,
  102584.1, 102576.7, 102560, 102540.5, 102511.7, 102478.4, 102439.9, 
    102395.9, 102344.9, 102288.7, 102227.6, 102165.8, 102097.9, 102026.4, 
    101951.4,
  102578.8, 102565.1, 102550.8, 102538.2, 102511, 102486.2, 102455, 102419.2, 
    102376.1, 102327.7, 102273.5, 102215.3, 102154.9, 102089.1, 102020.9,
  102543.8, 102605.3, 102630.4, 102666.9, 102676.6, 102680.9, 102677.4, 
    102660.9, 102627.8, 102593.1, 102543.3, 102479.6, 102404.5, 102317.1, 
    102216.2,
  102562.9, 102604.4, 102636.6, 102669.8, 102698.8, 102708.1, 102703.5, 
    102696.3, 102668.6, 102640.1, 102596.9, 102544, 102476.4, 102396.2, 
    102302.6,
  102591.4, 102604.7, 102646.6, 102684.2, 102708.1, 102727.3, 102730.9, 
    102729.5, 102710.5, 102679.3, 102644.1, 102595.1, 102537.9, 102470.2, 
    102382,
  102611.9, 102622.7, 102644.8, 102678.5, 102709.2, 102734.7, 102748.7, 
    102747.9, 102733.9, 102718.5, 102681.6, 102644.9, 102591.7, 102529, 
    102457.7,
  102623.1, 102640, 102658.8, 102671, 102707.8, 102731.5, 102745, 102754.6, 
    102750.8, 102728.9, 102713.6, 102670.8, 102632.2, 102574.5, 102509.8,
  102631.9, 102646.8, 102665.2, 102671.5, 102695.7, 102719.6, 102739.8, 
    102751.8, 102755.7, 102746.4, 102725.9, 102701.7, 102657.2, 102611.5, 
    102554.4,
  102635.7, 102649.7, 102666, 102677.7, 102680.5, 102695.6, 102722.9, 
    102742.1, 102745.1, 102749.9, 102734.9, 102710.9, 102680.2, 102635.3, 
    102589.2,
  102627.5, 102644.7, 102663.4, 102671.4, 102677.3, 102680.2, 102698.7, 
    102723.9, 102737.7, 102737.8, 102735.6, 102719, 102695.6, 102656, 102608.6,
  102622.3, 102637.7, 102655.2, 102664.2, 102667.2, 102669.9, 102683, 
    102696.8, 102710.6, 102720.3, 102723.4, 102712.2, 102693.2, 102663, 
    102626.5,
  102609.2, 102629.7, 102643.9, 102651, 102656, 102662.2, 102670.3, 102678.9, 
    102687.6, 102701.9, 102699.9, 102697.2, 102681.8, 102660.5, 102627,
  102324.8, 102358.5, 102386.1, 102405.8, 102427.2, 102447.9, 102459.3, 
    102467.9, 102457.1, 102452.6, 102441.3, 102409.8, 102361.9, 102302.8, 
    102243.3,
  102368.8, 102404.9, 102428.6, 102453.5, 102474.4, 102493.6, 102507.2, 
    102516.7, 102516.8, 102510.4, 102493.4, 102472, 102440.2, 102381.8, 
    102313.3,
  102403.4, 102441.4, 102468.5, 102498.1, 102523.3, 102552.1, 102570, 
    102587.2, 102593.1, 102587.3, 102568.7, 102537.5, 102504.6, 102463.1, 
    102401.9,
  102437, 102471.8, 102506.6, 102538.9, 102561.6, 102587.4, 102604.7, 
    102624.8, 102639.2, 102646.8, 102641.5, 102624.5, 102590.9, 102541.7, 
    102487.3,
  102453.9, 102500.6, 102530.5, 102566.1, 102592.9, 102614.1, 102641.2, 
    102665.6, 102689.1, 102706.5, 102707.5, 102698.4, 102673.1, 102634.6, 
    102582.7,
  102478, 102519.7, 102551.4, 102593.9, 102618.1, 102634.7, 102661.2, 
    102688.5, 102717.5, 102748.2, 102759.3, 102756.8, 102744.8, 102716, 
    102673.1,
  102496.8, 102532.9, 102574.8, 102607.6, 102627.2, 102651, 102678.6, 
    102710.6, 102746.2, 102769.8, 102799.8, 102797, 102793.4, 102777.9, 
    102746.3,
  102512.5, 102541.8, 102581.2, 102611.7, 102638.3, 102654.6, 102678.9, 
    102714.1, 102757.7, 102795, 102808.7, 102836.9, 102829.7, 102825.7, 102802,
  102529.3, 102551.4, 102596.2, 102619.3, 102638.5, 102659.6, 102684.8, 
    102719, 102766.6, 102799.6, 102825.7, 102839.9, 102844.4, 102851.4, 
    102841.9,
  102538, 102559.3, 102596.5, 102618.1, 102643.6, 102660.2, 102684.7, 102712, 
    102755.7, 102799.5, 102821.1, 102840.5, 102848.9, 102859.9, 102858.2,
  101728.1, 101740.4, 101772.3, 101796.2, 101822.9, 101848.8, 101875.9, 
    101907.4, 101934.1, 101961.8, 101985.3, 102009.1, 102041.7, 102076.6, 
    102105.4,
  101800.2, 101821.8, 101855.1, 101884, 101913.2, 101943.8, 101975.3, 
    102004.5, 102031.2, 102061.3, 102086.5, 102110.8, 102142.2, 102175.5, 
    102198.1,
  101879.7, 101906.2, 101945.9, 101973.1, 102001.9, 102036.3, 102066.5, 
    102100.1, 102134.9, 102159.3, 102184.9, 102213.3, 102236.1, 102264.5, 
    102296,
  101949, 101982.3, 102017.1, 102053.8, 102085.8, 102120.9, 102151.4, 
    102184.2, 102213.2, 102242.3, 102274.3, 102305.5, 102334.1, 102360.4, 
    102381.5,
  102011.2, 102051.2, 102086.2, 102125.5, 102157.4, 102186.2, 102216.8, 
    102249.5, 102283.3, 102314.6, 102357.5, 102396.6, 102430.1, 102455.2, 
    102475.4,
  102067.6, 102103.1, 102146.3, 102182.4, 102220.8, 102250.6, 102279.8, 
    102315.3, 102342.9, 102383.1, 102434.7, 102472.9, 102504.7, 102539, 
    102560.3,
  102113.6, 102150.4, 102196.5, 102233.1, 102269.1, 102300, 102332.1, 
    102367.8, 102399.1, 102447.4, 102495.9, 102536.5, 102575.4, 102611, 
    102631.9,
  102159.7, 102195.6, 102238.9, 102273.8, 102305.9, 102337.6, 102370, 
    102410.4, 102444.5, 102501.8, 102552.5, 102593.9, 102628.9, 102668.1, 
    102694.7,
  102201.8, 102228.7, 102274.9, 102310.3, 102340.7, 102372.8, 102407.9, 
    102446.3, 102488.2, 102544.8, 102591.2, 102628.5, 102668.7, 102710.1, 
    102740.4,
  102235.4, 102265.9, 102306.1, 102339.2, 102368.9, 102398.4, 102432.4, 
    102467.2, 102516.7, 102562.1, 102614.6, 102657.3, 102699, 102738.7, 
    102776.4,
  101832.4, 101756.3, 101667.7, 101590.1, 101510.5, 101432.8, 101365, 
    101298.8, 101229.2, 101186.8, 101138.3, 101088.2, 101067.6, 101032.1, 
    101026.5,
  101862, 101785, 101705.8, 101634.6, 101557.8, 101486.5, 101409.3, 101344.6, 
    101294.2, 101231.5, 101185.4, 101155.3, 101133.4, 101126.9, 101143.8,
  101890.7, 101818.4, 101744.8, 101675.4, 101609.6, 101541.1, 101479.7, 
    101417.4, 101366.7, 101321.4, 101288.7, 101261.1, 101247.6, 101252.2, 
    101282.1,
  101920.7, 101855.7, 101785.8, 101730.9, 101664.3, 101608.6, 101548.1, 
    101487.6, 101435.4, 101395, 101361.8, 101352.9, 101352.8, 101373.9, 101409,
  101948.5, 101888.3, 101825.8, 101774.3, 101720.3, 101667.9, 101612.7, 
    101570.8, 101528.5, 101495.5, 101475.1, 101467.1, 101475.5, 101501.7, 
    101542.6,
  101973.7, 101919, 101867, 101820.4, 101773.7, 101729.3, 101685.5, 101641.1, 
    101608, 101586.1, 101572.5, 101578.7, 101590.7, 101622, 101658.3,
  101993.7, 101950.6, 101902.1, 101863.8, 101822.3, 101782.8, 101750, 
    101721.6, 101689.5, 101679.1, 101670.6, 101680.4, 101698, 101740, 101777.6,
  102000, 101978.5, 101930.8, 101901.3, 101862.4, 101828.4, 101794.6, 
    101774.1, 101755.6, 101752.6, 101755.6, 101774.7, 101804.3, 101827.2, 
    101873.8,
  102013.6, 101992.5, 101954.5, 101931.1, 101894.6, 101869.4, 101842.1, 
    101826.8, 101814.9, 101818, 101831, 101851.9, 101878.3, 101910.1, 101955.3,
  102029.1, 102004.4, 101977.3, 101956.3, 101928.5, 101901, 101885, 101866.5, 
    101852.2, 101862.1, 101887.7, 101911.4, 101938.8, 101972.1, 102025,
  102573.7, 102612.7, 102628, 102632.6, 102625.1, 102606.5, 102577.8, 102537, 
    102477.2, 102415.6, 102333.4, 102247.2, 102147.4, 102047.9, 101942.1,
  102584.8, 102619, 102634.9, 102642.1, 102631.3, 102615, 102585.2, 102554.8, 
    102502.2, 102444.3, 102366.9, 102283.1, 102189.1, 102089.5, 101981.6,
  102581.9, 102615, 102634, 102643.2, 102637.6, 102623.5, 102596.9, 102564.7, 
    102516.5, 102466.3, 102395.5, 102313.9, 102224, 102125.7, 102012.6,
  102575.6, 102608.2, 102627.4, 102640.5, 102634.1, 102621.5, 102601.6, 
    102568.6, 102523.6, 102474.4, 102411.4, 102335, 102245.4, 102146.7, 
    102034.2,
  102568.1, 102599.4, 102609, 102627.9, 102622.1, 102612.7, 102591.2, 
    102566.4, 102526.6, 102476.1, 102417.4, 102343.7, 102256.3, 102157.6, 
    102047.7,
  102561, 102584.9, 102590.9, 102599.5, 102603.4, 102594.1, 102574.5, 
    102549.3, 102515.2, 102466.9, 102413.1, 102341.3, 102256.2, 102163, 
    102055.5,
  102538.9, 102562.8, 102570.3, 102573.9, 102567.8, 102565.8, 102546.7, 
    102526.1, 102491.4, 102451.6, 102398.9, 102331.5, 102249.8, 102160.5, 
    102058.9,
  102511.8, 102534.3, 102543.4, 102545.5, 102533.5, 102527.7, 102517.8, 
    102498.4, 102467.7, 102428.5, 102378.3, 102314.3, 102238.3, 102154.7, 
    102063.5,
  102482, 102502.4, 102503.2, 102508.2, 102500.8, 102487.9, 102481.3, 
    102461.9, 102436.4, 102398.6, 102351.5, 102292.2, 102224.8, 102151.5, 
    102059.4,
  102453.3, 102466.4, 102465.4, 102470.6, 102461.5, 102452.5, 102438.1, 
    102425, 102398.1, 102365, 102321.4, 102270.4, 102209.8, 102147.4, 102071.1,
  101875.2, 101953.4, 102033, 102110.9, 102187, 102263.7, 102336.1, 102393.3, 
    102437.3, 102474.4, 102495.9, 102501, 102497.8, 102480.3, 102452.8,
  101934.3, 102013.2, 102095.8, 102173.3, 102250.3, 102324.2, 102394.9, 
    102451.6, 102495.9, 102534.1, 102554.7, 102569.9, 102564.3, 102553.4, 
    102520.1,
  101972.6, 102048.3, 102129.8, 102212.6, 102291.8, 102364.4, 102437.3, 
    102498.5, 102539.3, 102586.6, 102609.6, 102629.2, 102630.2, 102617.7, 
    102597.1,
  101996.9, 102075, 102158.4, 102240.1, 102317, 102389.4, 102463.7, 102527.3, 
    102578, 102616.9, 102649, 102669.3, 102680.8, 102677.2, 102652.8,
  102012.8, 102083.4, 102165.5, 102237.7, 102322.4, 102396.7, 102468.6, 
    102538.5, 102593, 102634, 102672.5, 102692.7, 102708.8, 102712.4, 102704.9,
  102015.8, 102085.7, 102165.7, 102234.9, 102313.9, 102386.6, 102459.9, 
    102527.3, 102590.7, 102635.3, 102674.6, 102702.9, 102721.1, 102732.2, 
    102728.6,
  102014.8, 102079, 102153, 102216.7, 102288.6, 102363.5, 102437.4, 102505.6, 
    102569.1, 102620.7, 102665.3, 102696.4, 102721.3, 102743.2, 102744.6,
  102020.2, 102070.8, 102137, 102191.4, 102257.6, 102323.3, 102404.8, 
    102473.8, 102538.2, 102592.8, 102639.7, 102678.4, 102709.7, 102732.1, 
    102739.1,
  102029, 102065.4, 102125, 102167.5, 102225.5, 102283, 102350.6, 102422.5, 
    102488.9, 102551.1, 102604.7, 102647.2, 102680.5, 102704.3, 102718.2,
  102042.3, 102069.1, 102114.4, 102149.9, 102195.7, 102246.9, 102302.4, 
    102364.6, 102430.3, 102492.9, 102549.1, 102599.2, 102638.5, 102671.5, 
    102694.2,
  101586.1, 101489.4, 101398.1, 101326.1, 101270.2, 101239, 101229.5, 
    101204.9, 101244.9, 101262.6, 101352.6, 101418.3, 101533.8, 101670.4, 
    101805.1,
  101554.2, 101480.9, 101410.5, 101352.6, 101293.5, 101259.4, 101232.3, 
    101230, 101286.1, 101267.5, 101413.1, 101492.6, 101627.7, 101748.4, 101872,
  101568.2, 101488.8, 101411.9, 101346.6, 101283.3, 101261.8, 101240.5, 
    101255.9, 101277.5, 101343.7, 101423.9, 101505, 101648.6, 101794.6, 
    101932.4,
  101571.9, 101489.4, 101421.6, 101372.5, 101310.9, 101278.8, 101248.5, 
    101273.5, 101274, 101369.9, 101430.7, 101567.6, 101697.6, 101840.3, 101974,
  101599.8, 101507.7, 101429.9, 101381.5, 101327.4, 101294.4, 101270, 
    101296.7, 101288.3, 101355.7, 101439.6, 101572.7, 101695.6, 101850.8, 
    101990.3,
  101623.2, 101529.2, 101447.9, 101398.1, 101340.9, 101302, 101278.7, 
    101291.3, 101309.7, 101357.2, 101441.8, 101556.9, 101693.9, 101847.3, 
    101992.7,
  101660.5, 101567, 101486.8, 101417.2, 101358.1, 101312, 101288.3, 101293.7, 
    101321.1, 101364.4, 101429, 101543.5, 101687.4, 101834.3, 101973.7,
  101698.4, 101610.9, 101520.2, 101448.9, 101380.4, 101333.1, 101302.9, 
    101305, 101336.4, 101375.6, 101429.3, 101543.3, 101680.4, 101815, 101950.3,
  101732.3, 101642.8, 101557.3, 101482.6, 101408.7, 101363.6, 101327.5, 
    101325, 101350.4, 101380, 101435, 101543.5, 101666.4, 101784.6, 101919.7,
  101766.2, 101677.2, 101593.1, 101512.5, 101443.6, 101402.2, 101361.8, 
    101361.4, 101366.4, 101392.1, 101448.7, 101526.8, 101630.4, 101752.4, 
    101892.1,
  102089.2, 102009.9, 101911.6, 101792.4, 101666, 101520.3, 101378, 101217.1, 
    101126.5, 101042.8, 101027.2, 101026.6, 101103.4, 101222.5, 101376.2,
  102037.6, 101953.9, 101862.7, 101739.5, 101611, 101440.1, 101273, 101088, 
    100982.2, 100879.2, 100860.6, 100886.5, 100974.3, 101112.7, 101284.9,
  102019.2, 101933.5, 101824.8, 101693.2, 101554.8, 101384, 101200.5, 
    101005.2, 100884.8, 100772.1, 100765.7, 100780.4, 100857.3, 100990.3, 
    101156.1,
  101999, 101906.5, 101800.5, 101675, 101530.7, 101361.8, 101173.7, 100963, 
    100815.2, 100702.5, 100702.3, 100736, 100810.6, 100927.5, 101075.1,
  101989.7, 101891.1, 101782.8, 101655.9, 101510.1, 101342.1, 101176.5, 
    100977, 100826.7, 100702.5, 100699.6, 100721.8, 100798, 100890.1, 101014.5,
  101980.4, 101878.8, 101771.1, 101647.4, 101506.8, 101340.2, 101174.2, 
    100997, 100846.8, 100731, 100725.3, 100737.6, 100810.8, 100880.6, 100984.3,
  101979.7, 101870.4, 101760.4, 101636.5, 101496.3, 101336.8, 101175.1, 
    101015.6, 100869.9, 100763.6, 100744.1, 100745.3, 100826.5, 100878.4, 
    100962.1,
  101973.9, 101863.5, 101755, 101633.2, 101497.3, 101341.9, 101173.1, 
    101016.2, 100874.4, 100774, 100751.2, 100750.5, 100826, 100880.7, 100946.5,
  101976.9, 101863.9, 101747, 101633.1, 101496.8, 101346.9, 101188.8, 
    101023.1, 100888.1, 100758, 100727.4, 100751.8, 100816.3, 100877.7, 
    100931.3,
  101973.4, 101865.7, 101750.3, 101641.4, 101504.7, 101370.1, 101203.1, 
    101043.7, 100879.4, 100744.7, 100718.3, 100750.3, 100814.5, 100870, 
    100927.5,
  100844.4, 100822.8, 100792.8, 100755.7, 100698.7, 100632, 100539.1, 
    100471.9, 100436, 100410.2, 100407.5, 100418, 100423.1, 100481.2, 100507.8,
  100922.2, 100900.4, 100865.9, 100820.2, 100764.8, 100696.3, 100592.4, 
    100526, 100488.6, 100460.8, 100446.4, 100451.3, 100479.7, 100505.9, 
    100515.1,
  100987.6, 100972.6, 100944.9, 100902.6, 100843.9, 100773.6, 100664.2, 
    100590.3, 100539.4, 100511.8, 100495.6, 100492.4, 100517.6, 100505.1, 
    100551,
  101062.8, 101050.8, 101021.9, 100985.6, 100923.6, 100861.9, 100746, 100661, 
    100598.1, 100568.6, 100541.1, 100523.8, 100542.2, 100543.9, 100592.7,
  101124.1, 101117.9, 101095.7, 101065.2, 101002.5, 100948.3, 100847, 
    100746.3, 100667.8, 100627.2, 100596.8, 100559.9, 100577.7, 100577.4, 
    100614.8,
  101182.6, 101177.2, 101160.5, 101138.4, 101085, 101032.3, 100944.1, 
    100843.9, 100753.5, 100700, 100657.1, 100605.5, 100607.5, 100611, 100641.2,
  101221.2, 101232.7, 101218.6, 101197.5, 101157.3, 101105.8, 101035, 
    100938.4, 100846.6, 100772.8, 100713.5, 100665.4, 100646.7, 100651.6, 
    100668.7,
  101265.8, 101278.5, 101273.3, 101256.4, 101224.1, 101178.1, 101116.6, 
    101036.3, 100936, 100860.4, 100778.8, 100727.5, 100697, 100701.9, 100718.9,
  101310.5, 101319.1, 101324.4, 101312.1, 101287.7, 101251.3, 101193, 101129, 
    101033.4, 100949.2, 100844.2, 100791.3, 100765.7, 100764.3, 100785.6,
  101369.8, 101370.5, 101376.5, 101371.5, 101347.9, 101319.4, 101268.6, 
    101213.4, 101121.4, 101046.8, 100925.9, 100872.8, 100841, 100848.9, 
    100867.7,
  100659, 100591.3, 100532.3, 100476.4, 100422.1, 100382.1, 100350.6, 100334, 
    100322.6, 100311.4, 100301.5, 100292.6, 100282.8, 100274.3, 100273.5,
  100797.5, 100743.3, 100687.7, 100636.1, 100583.8, 100543.2, 100514.8, 
    100495.5, 100482.4, 100473.8, 100462.3, 100451.3, 100440.8, 100433.5, 
    100433.4,
  100930.2, 100883.2, 100836.2, 100792.2, 100744.8, 100704.1, 100674, 
    100656.1, 100644.7, 100635.6, 100630.3, 100620.4, 100612.1, 100607.4, 
    100602.9,
  101042.6, 101000.8, 100964.4, 100928.9, 100889.8, 100854.4, 100827.7, 
    100808.9, 100798.3, 100792.1, 100789, 100785.4, 100780.8, 100775, 100777.1,
  101136.8, 101105, 101077, 101050, 101018.4, 100987.4, 100964.9, 100950.2, 
    100940.2, 100937.1, 100935.4, 100939.1, 100939.1, 100940.8, 100943.3,
  101210.1, 101189.6, 101165.5, 101146.8, 101122.9, 101099.9, 101081.5, 
    101071.3, 101065.2, 101065.2, 101068.6, 101077, 101084.5, 101094, 101101.9,
  101265.6, 101257.7, 101236.9, 101226.1, 101206.2, 101189.1, 101177.1, 
    101170, 101169.6, 101174.3, 101183.4, 101196.2, 101212, 101228.4, 101244.8,
  101316.2, 101311.5, 101295.5, 101291, 101272.6, 101264.3, 101257, 101260.6, 
    101266.8, 101280.1, 101293.9, 101314, 101333.7, 101358.3, 101378.8,
  101356.3, 101357.6, 101351.1, 101350, 101338.3, 101334.9, 101337.9, 
    101345.4, 101361.2, 101377.9, 101398.9, 101421.9, 101449.4, 101476.6, 
    101503,
  101409.4, 101412.5, 101409.4, 101412, 101408.9, 101414, 101421.3, 101438.3, 
    101454.2, 101479.2, 101507.5, 101535.6, 101566.5, 101595, 101622.8,
  101368.6, 101333, 101304.5, 101276.8, 101242.1, 101214.9, 101180.6, 
    101153.9, 101125.5, 101102.5, 101077.4, 101058.1, 101039.1, 101023.4, 
    101007.4,
  101485, 101463, 101439.3, 101420.4, 101393.2, 101371, 101347.5, 101323.4, 
    101300.4, 101272.9, 101248.8, 101228.3, 101209.2, 101193.5, 101180.3,
  101581.3, 101567.8, 101553.6, 101547.8, 101532.6, 101515.7, 101499.6, 
    101479.7, 101461.6, 101437.3, 101416.5, 101395.9, 101375.4, 101357.8, 
    101341.4,
  101661.6, 101661.4, 101658.5, 101660.7, 101652.2, 101641.8, 101630.8, 
    101619.2, 101604.5, 101586.8, 101568.2, 101548.4, 101527.8, 101508.9, 
    101492.5,
  101721.5, 101736.3, 101741.6, 101749.4, 101747.8, 101745.1, 101741, 
    101734.9, 101726.9, 101717.1, 101703.9, 101689.4, 101670.9, 101653.3, 
    101635.4,
  101767, 101787, 101799.9, 101815.3, 101822.5, 101827.3, 101829, 101830.7, 
    101828.3, 101824.7, 101816.2, 101805.9, 101790.6, 101774.9, 101759.6,
  101799.1, 101822.3, 101844.7, 101865.6, 101877.3, 101891.7, 101899.6, 
    101906.6, 101910.4, 101912.5, 101909.8, 101903.2, 101891.6, 101878.7, 
    101866.7,
  101827.1, 101846.1, 101874.8, 101901.2, 101920.4, 101943.5, 101958.5, 
    101970.9, 101980.7, 101985.7, 101988.1, 101985.1, 101979.7, 101970.8, 
    101963.3,
  101854.6, 101870, 101902.4, 101933.4, 101956, 101983.9, 102004.9, 102023.9, 
    102036.3, 102045.8, 102049.6, 102052, 102052.9, 102052.1, 102051.9,
  101878.2, 101899, 101933.4, 101964.5, 101993.3, 102021.5, 102044.6, 
    102062.5, 102076.4, 102091.6, 102102.7, 102108.7, 102113, 102119.3, 
    102128.9,
  101159.8, 101157.9, 101162.1, 101168, 101176.9, 101188.1, 101202.3, 
    101215.9, 101231.5, 101244.4, 101256.4, 101263.5, 101275.6, 101283.2, 
    101291.7,
  101249.1, 101251, 101265.9, 101278, 101291.6, 101305.7, 101325.2, 101343.8, 
    101364.4, 101383.8, 101403.1, 101419.1, 101436.6, 101449.7, 101460,
  101334.4, 101343.5, 101362.3, 101380.5, 101398.8, 101421.7, 101446, 
    101472.7, 101502.4, 101529.8, 101554, 101575.1, 101595.2, 101613, 101629.8,
  101406.2, 101424.2, 101448.1, 101471, 101493.4, 101523.7, 101553.9, 
    101588.2, 101621.6, 101656.3, 101687.3, 101717.4, 101742.5, 101764.9, 
    101785.3,
  101472.5, 101500.3, 101526.5, 101556.2, 101588.9, 101625.2, 101662.1, 
    101702.4, 101742.5, 101781.7, 101817.8, 101851, 101880.3, 101907.6, 
    101931.9,
  101532.3, 101568.6, 101599.3, 101634.2, 101673.9, 101712.1, 101757.5, 
    101799.8, 101842.9, 101884.4, 101925.4, 101963.4, 101998, 102029.9, 
    102059.1,
  101593, 101628, 101668, 101708.4, 101751.6, 101796.5, 101842.8, 101886.9, 
    101932.5, 101975.1, 102020, 102060.6, 102099.8, 102134.2, 102166,
  101656.5, 101682.6, 101734.2, 101778, 101825.6, 101873.1, 101918.5, 
    101962.4, 102009.4, 102053.4, 102099.3, 102141.3, 102181.7, 102217.5, 
    102247.6,
  101714, 101739, 101800.2, 101845.3, 101896.1, 101944.1, 101984.1, 102027.3, 
    102071.3, 102114.5, 102163.6, 102204.4, 102245.2, 102279, 102315.8,
  101761.9, 101796.8, 101860.8, 101905.1, 101957.5, 102000.7, 102038.3, 
    102073.7, 102116.5, 102158.8, 102211.8, 102252.8, 102291.7, 102327.6, 
    102365.2,
  100923, 100909.2, 100901.6, 100900.1, 100906.4, 100916.7, 100934, 100957.1, 
    100985, 101016.8, 101053.2, 101087.1, 101127.7, 101164.5, 101204.8,
  101025.2, 101014.1, 101016.7, 101021.1, 101028.5, 101041.5, 101063.9, 
    101093.2, 101124.8, 101157.3, 101197.7, 101237.3, 101276.7, 101320.2, 
    101364.6,
  101116.6, 101111.3, 101121.5, 101128.9, 101143.2, 101162.5, 101190.9, 
    101220.9, 101260.3, 101303.8, 101345.9, 101389.6, 101433.1, 101477.3, 
    101523,
  101180.1, 101184.2, 101202.6, 101216.1, 101238.1, 101265.5, 101301.1, 
    101340.3, 101384, 101429.5, 101474, 101518.7, 101562.6, 101607.6, 101651.1,
  101231.4, 101251, 101269.7, 101294.9, 101327.3, 101363.3, 101403.6, 
    101447.8, 101495.8, 101541.7, 101585.8, 101631.4, 101676.7, 101721.4, 
    101761.9,
  101266.7, 101301.2, 101324.8, 101363.8, 101403.8, 101448.2, 101493.1, 
    101537.4, 101581.1, 101623.7, 101666.9, 101711.6, 101754.4, 101795.9, 
    101843.4,
  101304.5, 101352.5, 101383.9, 101428.6, 101473.8, 101518.6, 101560.3, 
    101603.6, 101646.8, 101685.5, 101727.4, 101771.6, 101814, 101859.7, 
    101899.1,
  101353.1, 101396.2, 101434.9, 101483.7, 101529.4, 101576.2, 101616.7, 
    101657.6, 101695.4, 101729.7, 101770.5, 101812.5, 101856.8, 101898.1, 
    101941.8,
  101401.5, 101431.9, 101489, 101534.4, 101583.3, 101624.6, 101663.2, 101697, 
    101729.9, 101752.3, 101790.1, 101832.5, 101882.9, 101921.6, 101953.9,
  101444.6, 101476.2, 101536.1, 101578.3, 101629.2, 101667.7, 101700.2, 
    101722.5, 101740.1, 101756.8, 101792.9, 101840, 101892.2, 101918.7, 
    101962.2,
  100780.2, 100783.6, 100788.8, 100799.2, 100818.1, 100845.1, 100880.8, 
    100924.8, 100972.6, 101024.5, 101080.4, 101142.5, 101206.7, 101271.9, 
    101335,
  100866.1, 100874.4, 100888.1, 100901.5, 100920.7, 100944.1, 100976.6, 
    101020.5, 101072.8, 101129.5, 101193.6, 101259.8, 101329.3, 101399.7, 
    101462.1,
  100946.6, 100955.3, 100972.9, 100989, 101006.7, 101033.6, 101077.5, 101127, 
    101183.8, 101248.4, 101312.1, 101382.9, 101449.7, 101505.9, 101556.5,
  100997.8, 101018.2, 101040.1, 101058.4, 101080.9, 101114.7, 101158.7, 
    101214.8, 101277.3, 101344.5, 101413, 101480.7, 101540.3, 101594.6, 
    101644.1,
  101042.6, 101066.3, 101090.4, 101120.3, 101151.1, 101192.7, 101243.2, 
    101301.6, 101367.1, 101434.6, 101502.7, 101569.8, 101623.1, 101673.1, 
    101722.3,
  101075.2, 101109.9, 101140.7, 101177.1, 101217.8, 101262.6, 101315.1, 
    101376.6, 101444.6, 101511.3, 101580.4, 101638, 101687.2, 101740.5, 
    101786.9,
  101111.2, 101154.4, 101186.4, 101229.9, 101280.1, 101329.8, 101388.5, 
    101451.7, 101516.1, 101580.2, 101646.5, 101693.3, 101747.9, 101799.5, 
    101843.1,
  101154.4, 101192, 101239.2, 101293.2, 101345, 101399.6, 101459.3, 101519.8, 
    101581.1, 101645.3, 101698.5, 101751.2, 101801.5, 101849.6, 101892.5,
  101204.5, 101237.1, 101297.8, 101349.1, 101412, 101466.8, 101526.2, 
    101581.4, 101640.5, 101697.5, 101753.5, 101801.4, 101848.7, 101895.4, 
    101939.5,
  101257.3, 101294.4, 101355.7, 101412.4, 101475.6, 101528.4, 101582.7, 
    101631.9, 101690.6, 101742.6, 101796.2, 101844.2, 101892.5, 101936.4, 
    101974.3,
  101227.8, 101185.3, 101148.3, 101117.3, 101091.8, 101077.3, 101069.8, 
    101074.5, 101065.5, 101051.2, 101043, 101045.4, 101055.4, 101086.1, 
    101139.2,
  101299.1, 101259.3, 101219.3, 101184.1, 101155, 101134.5, 101128.1, 
    101106.9, 101086.8, 101075.1, 101072.5, 101092.2, 101144.1, 101200.9, 
    101259.1,
  101370.1, 101332.9, 101294, 101260.5, 101232.8, 101207, 101185.7, 101164.7, 
    101151.8, 101142.3, 101160.7, 101203.6, 101234.7, 101287, 101361.6,
  101400.5, 101366.3, 101332.3, 101299.6, 101273.5, 101245.4, 101219.1, 
    101200, 101195.8, 101211.8, 101231.9, 101241.4, 101293.2, 101379.5, 
    101468.7,
  101431.5, 101389.5, 101359.2, 101327.5, 101301.2, 101283.3, 101266.1, 
    101256.5, 101257.7, 101249.1, 101269.7, 101331.2, 101409.7, 101485.7, 
    101570.7,
  101428.8, 101391, 101364.1, 101334.1, 101304.5, 101291.3, 101273.6, 
    101264.7, 101264.9, 101300.2, 101363.3, 101434, 101504.9, 101584.7, 
    101664.2,
  101413.4, 101395.8, 101365.8, 101334.4, 101301.7, 101283.3, 101280.3, 
    101299, 101335.9, 101390.5, 101454.5, 101526.9, 101600.5, 101675.4, 
    101746.1,
  101396.8, 101381.7, 101350.7, 101326.9, 101313.2, 101316.7, 101331.7, 
    101366.3, 101412.7, 101470.3, 101541.3, 101612.6, 101682.7, 101751, 
    101822.3,
  101430.2, 101400.9, 101378.5, 101365.7, 101366.1, 101377.6, 101404, 
    101439.5, 101487.1, 101547.7, 101620.8, 101685.3, 101751.2, 101819.6, 
    101886.2,
  101493, 101450.4, 101432.6, 101421, 101429.1, 101443.8, 101473.2, 101511.4, 
    101563.4, 101624.1, 101689.2, 101750.9, 101815.8, 101875, 101940.3,
  101555.1, 101490.6, 101424.3, 101365.9, 101306.1, 101242.5, 101182.9, 
    101124.2, 101073.8, 101026, 100983.6, 100941.6, 100890.8, 100858.5, 
    100842.7,
  101655.3, 101602.1, 101535.2, 101481.3, 101419.2, 101360.5, 101300.3, 
    101245.4, 101190.5, 101139.5, 101089.8, 101039.9, 101009.4, 100977.6, 
    100923.2,
  101771.5, 101709.5, 101644.2, 101590.7, 101530.6, 101472.9, 101416.7, 
    101365.1, 101313.6, 101268.2, 101214.4, 101172.5, 101125.2, 101067.2, 
    101030.2,
  101880.6, 101818.1, 101754.6, 101704.3, 101645.9, 101589.5, 101534.8, 
    101483.1, 101430.6, 101377.8, 101331.7, 101285, 101230.8, 101191.4, 101156,
  101982.3, 101927.6, 101866.5, 101816.2, 101757, 101701.3, 101643.5, 
    101592.2, 101544.2, 101494, 101441.4, 101390.8, 101343.1, 101295.6, 
    101254.5,
  102064.8, 102020.7, 101966.9, 101919.2, 101861.4, 101804.1, 101747.9, 
    101695.4, 101644, 101589.6, 101538, 101485.9, 101439.3, 101399.9, 101377.4,
  102141.2, 102095.5, 102053.2, 102007.6, 101954.1, 101900.9, 101845.6, 
    101790.8, 101736.4, 101681.1, 101631, 101585.3, 101545.1, 101516.4, 
    101493.8,
  102205.9, 102162, 102122.7, 102080.3, 102028.6, 101977.6, 101927.6, 
    101873.4, 101820.3, 101766.9, 101718.4, 101677.5, 101646.3, 101622.5, 
    101606.9,
  102250.4, 102214.7, 102180.2, 102141.4, 102096.2, 102045.4, 101997.5, 
    101943.6, 101891.7, 101839.5, 101796.8, 101759.6, 101730.5, 101713.3, 
    101697.3,
  102290.7, 102257.1, 102224.3, 102187, 102145, 102099.5, 102047, 101997.3, 
    101945.4, 101899.8, 101857.8, 101825.4, 101799.7, 101780.6, 101768.2,
  101474.9, 101381.8, 101292.3, 101209.6, 101127.5, 101055.9, 100986.4, 
    100912.6, 100849.2, 100789.6, 100738.1, 100683.4, 100630.6, 100571.9, 
    100511.7,
  101621.3, 101550.7, 101475.8, 101398.3, 101313.1, 101233.6, 101157.8, 
    101090.7, 101020.2, 100953.3, 100888.2, 100828.7, 100766.5, 100705.7, 
    100654.3,
  101760.7, 101698.8, 101630.8, 101566.6, 101492.2, 101418.4, 101344.3, 
    101270.9, 101201.4, 101132.6, 101068.2, 101003.5, 100943.3, 100882.1, 
    100821.5,
  101879.9, 101827, 101776.2, 101725, 101659.6, 101591.6, 101523.2, 101454.8, 
    101389.1, 101322.8, 101260.8, 101197.4, 101133.2, 101071.8, 101011.2,
  101977.4, 101941.2, 101901.9, 101859.7, 101802.9, 101745.6, 101686.5, 
    101625.2, 101562, 101501.2, 101441.4, 101383.9, 101323.6, 101264.8, 101207,
  102050.8, 102029.9, 102006, 101976.9, 101932, 101886.4, 101835, 101781.7, 
    101726, 101669.7, 101613.7, 101558.9, 101503, 101448.4, 101393.9,
  102113.1, 102101.1, 102089.7, 102068.4, 102037, 102001.8, 101959.6, 
    101916.2, 101869.6, 101822.1, 101771, 101720.1, 101668.3, 101616.4, 
    101567.2,
  102163.6, 102158, 102157.1, 102143.4, 102119.1, 102093.5, 102060.3, 
    102026.7, 101989.5, 101951.1, 101907.9, 101862.7, 101815.7, 101768.7, 
    101721.9,
  102210.4, 102211.3, 102215.3, 102207, 102188.8, 102170.4, 102145.2, 
    102120.3, 102091.6, 102060.4, 102024.7, 101985.1, 101944.4, 101901.3, 
    101859.1,
  102253.7, 102259.5, 102265.1, 102261.1, 102250, 102235, 102215.2, 102192.8, 
    102168.9, 102143.7, 102118.2, 102086.7, 102051.7, 102015.7, 101978.2,
  101255, 101216.6, 101191.5, 101155.9, 101114.2, 101081.5, 101042.5, 
    101000.6, 100961.4, 100926.2, 100892.9, 100854.2, 100808.4, 100750.6, 
    100693.4,
  101371.6, 101351.9, 101334.3, 101307.6, 101272.5, 101237, 101203.5, 
    101167.2, 101127.3, 101081.8, 101033.6, 100986, 100940.8, 100894.5, 
    100835.5,
  101481.1, 101473.6, 101462.3, 101449.6, 101422.8, 101391.4, 101358.7, 
    101326.4, 101291.5, 101251.8, 101202, 101152.3, 101095, 101038.1, 100977.2,
  101568.1, 101572.8, 101569.9, 101567.2, 101546.6, 101527.3, 101502.9, 
    101474.2, 101443, 101409.2, 101370.4, 101325.4, 101268.7, 101213.4, 
    101151.2,
  101625.9, 101649.2, 101656.1, 101662.7, 101651.9, 101643.7, 101627.2, 
    101607.7, 101582.4, 101553.7, 101516.6, 101480.1, 101429.8, 101374.3, 
    101313.9,
  101669.1, 101707.1, 101720.3, 101736.4, 101738, 101741.6, 101733.9, 
    101722.1, 101704.7, 101683.7, 101654.3, 101621.5, 101580.2, 101532.3, 
    101478,
  101705, 101745.4, 101770.4, 101794.4, 101806.2, 101817.4, 101815.8, 101815, 
    101806.8, 101796.1, 101775.4, 101749.3, 101714.9, 101671.8, 101625.3,
  101734.6, 101782.2, 101817.4, 101848.2, 101873.3, 101889.8, 101897.7, 
    101903.6, 101901.6, 101897.9, 101886.2, 101866.9, 101840.7, 101807.8, 
    101765.3,
  101778.9, 101820.1, 101868.1, 101907.1, 101941, 101962.8, 101977.9, 
    101987.4, 101990, 101988.7, 101983.3, 101972.1, 101953.2, 101927.5, 
    101893.4,
  101825.8, 101865.2, 101923.7, 101964.4, 102003.6, 102032.6, 102050.2, 
    102058.4, 102061.9, 102065.6, 102065.5, 102060.3, 102048.9, 102031.7, 
    102006.1,
  101612.3, 101587, 101569.8, 101545.9, 101512.7, 101475.5, 101426.6, 
    101377.4, 101323.4, 101266.1, 101199.8, 101129.3, 101052.4, 100973.8, 
    100890.9,
  101605.1, 101587.2, 101579, 101557.6, 101540.5, 101513.5, 101479, 101444.7, 
    101401.7, 101353.1, 101299.4, 101237.8, 101171.7, 101103.7, 101030.1,
  101609.5, 101592, 101590.3, 101580.1, 101570.4, 101552.6, 101529.3, 
    101501.5, 101468.8, 101431.6, 101389.8, 101339.9, 101284.5, 101223.3, 
    101157.6,
  101631.7, 101613.4, 101611.6, 101598.8, 101591, 101580.8, 101568.7, 
    101550.8, 101531.5, 101504.5, 101474.2, 101439.5, 101396.5, 101350.4, 
    101300.9,
  101651, 101638.1, 101633.4, 101624.8, 101623.6, 101622.8, 101621, 101613.3, 
    101602.3, 101586.4, 101564.2, 101539.3, 101507.5, 101469.5, 101427.6,
  101672.3, 101668.7, 101660, 101656.2, 101658.5, 101665.4, 101672.3, 
    101677.8, 101683, 101679.1, 101670.3, 101655.4, 101633.1, 101605.4, 101571,
  101684.1, 101690.8, 101684.4, 101688.5, 101700, 101716.4, 101735.6, 101749, 
    101762.6, 101769, 101769.7, 101765.1, 101752.4, 101731.7, 101708.5,
  101696.4, 101709, 101712, 101729.1, 101747.1, 101768.7, 101793.5, 101821.9, 
    101840.8, 101857.8, 101865.6, 101869.9, 101867.3, 101858.7, 101841.9,
  101716.9, 101737, 101751.2, 101775.7, 101803.1, 101830.7, 101865.9, 
    101894.7, 101916.3, 101934.6, 101950, 101961.9, 101967.9, 101965.5, 
    101958.9,
  101751.7, 101776.1, 101798.7, 101828.5, 101862, 101896.4, 101933.7, 
    101960.4, 101985.5, 102010.5, 102035.5, 102056.9, 102069.5, 102073.5, 
    102071.5,
  103335.2, 103345.1, 103343.9, 103345.1, 103324.9, 103301.9, 103256.6, 
    103209.3, 103147, 103074.9, 102991.4, 102900.2, 102802, 102693.3, 102577,
  103260.4, 103294.3, 103311.9, 103319.3, 103305.1, 103291.4, 103257.2, 
    103219.2, 103169.3, 103113.7, 103044.3, 102966.7, 102879.4, 102778.8, 
    102672.8,
  103198.7, 103243.2, 103261.5, 103271.5, 103271.2, 103264.3, 103244.6, 
    103215.6, 103173.8, 103125.9, 103070.6, 103002.5, 102930, 102845.8, 
    102748.9,
  103120.5, 103167.3, 103193.9, 103214.5, 103217.9, 103221.3, 103205.2, 
    103186.3, 103158.5, 103126.8, 103083.2, 103029, 102968.2, 102897.2, 
    102814.6,
  103043, 103087.8, 103110.1, 103136.9, 103146.8, 103153.4, 103144.9, 
    103135.8, 103117.1, 103092.4, 103061, 103019.7, 102970, 102912.4, 102844.9,
  102960.5, 103003.6, 103031.5, 103051.8, 103060.8, 103069.3, 103070.5, 
    103068.4, 103057, 103044.7, 103022, 102990.8, 102955.7, 102910.1, 102855.3,
  102873.4, 102914.4, 102935, 102958, 102967.4, 102976.7, 102981.3, 102985.9, 
    102985.8, 102979.2, 102963.1, 102938.4, 102913.7, 102878.7, 102834.6,
  102791.3, 102829, 102845.7, 102864.9, 102875.5, 102886.9, 102896.9, 
    102903.2, 102907.5, 102905.6, 102900.5, 102889.1, 102867.5, 102837, 102803,
  102715.4, 102749.5, 102760.8, 102780.2, 102788.9, 102802.8, 102813.6, 
    102824, 102830.5, 102835.5, 102832.9, 102826.5, 102823, 102802.6, 102771.8,
  102645.3, 102677.6, 102686, 102705.4, 102711.3, 102721.6, 102732, 102744.5, 
    102752.1, 102763.1, 102774.4, 102781.1, 102782.2, 102771, 102753.2,
  103281.4, 103371.7, 103458.2, 103535.8, 103592.1, 103639.2, 103666.9, 
    103691.1, 103686.6, 103652.9, 103605.9, 103552.3, 103497.3, 103431.7, 
    103365,
  103233.1, 103331.5, 103425.3, 103503.3, 103574.1, 103625.8, 103660.4, 
    103687.7, 103702.6, 103691.7, 103657.5, 103608.9, 103558.2, 103497, 
    103428.4,
  103184.5, 103284.4, 103383.5, 103469.1, 103540.4, 103605.5, 103651, 103682, 
    103705.2, 103715.8, 103695.9, 103657.9, 103609.8, 103555, 103490.9,
  103121.4, 103228.8, 103325.2, 103418.4, 103497.5, 103568.2, 103622.2, 
    103664, 103691.5, 103709.4, 103713.7, 103690.3, 103654.2, 103605.7, 
    103548.3,
  103048.6, 103168.3, 103255.3, 103354.4, 103431.1, 103512.8, 103578, 
    103631.1, 103669.1, 103694.5, 103709.5, 103707.8, 103684, 103645.1, 
    103596.1,
  102961, 103093.1, 103176.3, 103283.4, 103360.5, 103445.2, 103520, 103582.2, 
    103629.4, 103663.4, 103686.1, 103696.9, 103692, 103668.9, 103630.3,
  102880.6, 103005.6, 103088.6, 103190.2, 103275.7, 103362.8, 103440.8, 
    103516.5, 103575.5, 103620, 103650.3, 103669.8, 103677.7, 103669.8, 
    103641.9,
  102808.4, 102913.1, 103002.7, 103097.4, 103186.5, 103275.4, 103354.9, 
    103427.5, 103502.6, 103557.7, 103601, 103629.5, 103646.6, 103649.2, 
    103634.9,
  102753.4, 102822.9, 102908.7, 102998.7, 103085, 103177.4, 103261.7, 
    103337.6, 103405.7, 103475.9, 103529.5, 103571.6, 103595.6, 103607.9, 
    103608.3,
  102712.9, 102761.2, 102825.6, 102901.3, 102981.5, 103064.4, 103148, 
    103229.8, 103307.1, 103380.3, 103444.9, 103494.2, 103531.7, 103554, 
    103565.5,
  101971.1, 102088, 102196.7, 102314.2, 102435.9, 102553.9, 102675.3, 
    102787.9, 102892.1, 102979.1, 103041.5, 103098.3, 103143.4, 103179.1, 
    103213.1,
  102002.2, 102120.1, 102226.9, 102345.9, 102459.8, 102577.6, 102692.6, 
    102804.7, 102909.9, 103003.5, 103076.2, 103133.1, 103182.2, 103225.5, 
    103255.8,
  102021.9, 102135.1, 102244.1, 102362.2, 102475.6, 102590, 102707.4, 
    102819.4, 102925.2, 103021.8, 103099.9, 103160.7, 103213.4, 103258.1, 
    103289.2,
  102039.4, 102147.1, 102252.4, 102363.5, 102477.1, 102591.4, 102705.1, 
    102818, 102924.8, 103022.6, 103106.5, 103174.4, 103233.4, 103285.9, 
    103318.9,
  102049.6, 102148.9, 102247.7, 102354, 102469.2, 102581.9, 102695.5, 
    102806.1, 102913.5, 103013.1, 103101.9, 103176.8, 103240.7, 103298.9, 
    103343.1,
  102058.9, 102144.9, 102237.7, 102334.7, 102445.5, 102558.5, 102673.3, 
    102783.3, 102891.3, 102994.1, 103086.6, 103166.7, 103235.9, 103296.7, 
    103345.5,
  102064.1, 102138.2, 102225.5, 102310.9, 102416, 102528.6, 102645.3, 
    102754.3, 102862.3, 102967, 103063.4, 103146.6, 103218.9, 103280.9, 
    103330.8,
  102073.8, 102133.9, 102211.5, 102287, 102379.4, 102484.8, 102611.4, 102719, 
    102824.9, 102930.1, 103031.4, 103118.6, 103194, 103257.3, 103315.8,
  102087, 102140, 102206, 102269.2, 102354.3, 102450.9, 102562.1, 102677.1, 
    102785.6, 102885.8, 102991.5, 103080.9, 103158.3, 103223.5, 103284.9,
  102101.9, 102146.6, 102204, 102254.6, 102325.4, 102409.5, 102508.6, 
    102615.1, 102735.2, 102839.4, 102938.3, 103034.3, 103117.9, 103185.4, 
    103247.4,
  101691.2, 101666.3, 101651.6, 101643.1, 101646.4, 101658.1, 101681.5, 
    101718.7, 101766.3, 101816.9, 101872.1, 101925.5, 101983.3, 102042.5, 
    102104.9,
  101767.7, 101747.4, 101743.7, 101742.1, 101748.2, 101762.8, 101782.7, 
    101816.2, 101862.9, 101912.5, 101965.7, 102019.4, 102080.8, 102144.7, 
    102211.1,
  101839.6, 101832.7, 101835.8, 101833.7, 101841.5, 101852.5, 101871.9, 
    101901.9, 101947, 101996, 102054.4, 102115.7, 102177.5, 102244.1, 102315.1,
  101883.4, 101876.5, 101883.6, 101889, 101904.9, 101921.8, 101946.7, 
    101980.5, 102022.7, 102074.9, 102133.8, 102198.3, 102263, 102337.3, 
    102409.9,
  101885.6, 101901.1, 101918.3, 101936.1, 101954, 101975.1, 102005.4, 
    102043.5, 102091.5, 102147.8, 102208.8, 102277.4, 102346.7, 102419.3, 
    102495.5,
  101871.7, 101908.6, 101927.6, 101950.3, 101985, 102016.8, 102057.8, 
    102099.5, 102148.3, 102203.5, 102268.8, 102338.2, 102408.1, 102483.9, 
    102558.8,
  101877, 101917.1, 101946.1, 101978.4, 102020.9, 102055, 102095.3, 102140.7, 
    102198.6, 102251.4, 102317.8, 102389.6, 102463.8, 102536.2, 102614.4,
  101917.9, 101933, 101980.6, 102008.3, 102049.8, 102084.4, 102132.6, 
    102178.3, 102233.8, 102292.9, 102363.3, 102437.8, 102511.5, 102586.5, 
    102661.2,
  101966.6, 101966.1, 102008.5, 102042, 102085.5, 102119.7, 102162.4, 102207, 
    102267.2, 102328.2, 102393.9, 102468.9, 102546.9, 102622.1, 102699.4,
  101999.5, 101994, 102043.9, 102077.3, 102115.8, 102141.4, 102186.5, 
    102224.3, 102276.6, 102345.4, 102414, 102485.5, 102566.7, 102645.6, 
    102725.3,
  101205, 101271.7, 101346.6, 101403.8, 101467.1, 101526.7, 101586.4, 
    101641.2, 101697.9, 101742.2, 101782.4, 101819, 101847.8, 101863.3, 
    101871.7,
  101221.1, 101290.6, 101359.7, 101416.9, 101486.4, 101555.9, 101616.9, 
    101684.9, 101742.3, 101795.2, 101840.1, 101876.9, 101912.4, 101941.5, 
    101960.1,
  101237.4, 101309.9, 101382.6, 101439.2, 101512.3, 101580.6, 101655.9, 
    101729.5, 101796.4, 101855.7, 101905.8, 101946.7, 101984.4, 102012.9, 
    102036.4,
  101248, 101314.4, 101393.2, 101448.5, 101520.9, 101590.6, 101674.2, 
    101756.4, 101833.7, 101899.4, 101952.5, 101995.7, 102040.1, 102075.1, 
    102104.5,
  101256, 101335.3, 101419.4, 101462.4, 101537.9, 101606.6, 101692.3, 
    101777.9, 101862.6, 101935.6, 101996.8, 102046.6, 102091.8, 102132.6, 
    102168.9,
  101279.6, 101349.6, 101434.5, 101482.9, 101560.8, 101621.4, 101700.2, 
    101792.5, 101884, 101959.9, 102024.5, 102079.9, 102133.1, 102182.2, 
    102220.4,
  101306.8, 101386.8, 101463.7, 101508.6, 101582.6, 101649.4, 101728.1, 
    101810.9, 101900.6, 101978.5, 102048.9, 102110.7, 102172.6, 102227, 
    102275.3,
  101345.1, 101415.2, 101478.7, 101532.2, 101605.2, 101665.5, 101746.7, 
    101827.8, 101908.5, 101986.6, 102061.7, 102130.4, 102199, 102261.3, 
    102323.7,
  101389, 101441.3, 101495.5, 101557.6, 101628.5, 101706, 101777.3, 101852.9, 
    101927.2, 101996.9, 102074.7, 102146.2, 102217.7, 102283.8, 102362.2,
  101421.8, 101466.8, 101521.5, 101597.2, 101655.1, 101727.4, 101796.7, 
    101873.5, 101939.7, 102009.6, 102082.5, 102153.6, 102229.9, 102303.7, 
    102386.6,
  100465, 100437.2, 100413, 100391.5, 100410.3, 100399.2, 100482, 100522.6, 
    100618.7, 100706.5, 100810.8, 100953.8, 101099.5, 101230.4, 101354.7,
  100559.1, 100534.1, 100507.2, 100493.7, 100489.3, 100498.1, 100564.9, 
    100566.1, 100672.6, 100751.6, 100873.5, 101013.3, 101158, 101297.6, 
    101426.6,
  100661.6, 100632.4, 100607, 100589.9, 100567.9, 100606.5, 100604.5, 
    100659.9, 100744.5, 100827.3, 100956.4, 101088.1, 101224.3, 101361.1, 
    101487.6,
  100752.2, 100723.7, 100704.4, 100685.3, 100683, 100691.7, 100688.6, 
    100752.1, 100816.7, 100915.4, 101040.5, 101162.8, 101295.4, 101426.7, 
    101553.6,
  100831, 100802, 100792.8, 100773.6, 100770.7, 100769.5, 100793.7, 100842.8, 
    100915, 101035.1, 101139.5, 101246, 101371.2, 101497.9, 101623.7,
  100900.7, 100877.4, 100875, 100854, 100863.6, 100875.3, 100891.6, 100947.4, 
    101022.6, 101131.3, 101220, 101326.7, 101443.9, 101568.9, 101694.9,
  100944.2, 100942.2, 100946, 100949.1, 100960.3, 100959.8, 100986.3, 
    101031.6, 101121.7, 101217.3, 101294.2, 101402.3, 101516.3, 101640.7, 
    101760.5,
  101010.5, 101028.6, 101042.6, 101036.6, 101029.8, 101037.5, 101066.4, 
    101128.7, 101219.4, 101279.8, 101371.3, 101480.7, 101591.4, 101709.4, 
    101829.4,
  101063, 101059, 101077.1, 101079.5, 101108.7, 101123.8, 101160.6, 101231.6, 
    101284.1, 101355, 101453.3, 101551.2, 101666.1, 101779.4, 101891.3,
  101090.7, 101075.3, 101115.6, 101126.9, 101158.1, 101193.6, 101245.6, 
    101308.4, 101371.8, 101445.6, 101534.8, 101633.3, 101743.1, 101842.6, 
    101947.5,
  101445.3, 101327.9, 101245.5, 101159.6, 101080.5, 101012.9, 100955.8, 
    100905.8, 100855.4, 100808.1, 100769, 100722.6, 100711.9, 100738.8, 
    100790.8,
  101583.7, 101479.6, 101396.6, 101314.2, 101241.4, 101178, 101125.4, 
    101075.4, 101035.2, 100985.6, 100948.5, 100914, 100910.5, 100931.8, 
    100967.8,
  101738, 101637.6, 101556.1, 101472.4, 101402.2, 101338.5, 101288.5, 
    101239.8, 101203.2, 101160, 101131.7, 101100, 101092.9, 101098.3, 101124.4,
  101876, 101783.1, 101706.5, 101627.1, 101560.4, 101499.5, 101451.3, 
    101403.4, 101371.5, 101327.4, 101299.2, 101268.2, 101258.6, 101259.1, 
    101274.6,
  101992.1, 101911.1, 101844.1, 101772, 101708.2, 101650.4, 101603.2, 
    101559.2, 101524.9, 101478.9, 101454.1, 101435.1, 101417.2, 101407.2, 
    101409.8,
  102078, 102009.1, 101957.8, 101895.3, 101839.4, 101785.6, 101738.1, 
    101698.1, 101655.1, 101614.1, 101599.3, 101580.3, 101554.9, 101539.4, 
    101529.3,
  102137.9, 102079.5, 102039.3, 101983.8, 101936.9, 101888.5, 101845.9, 
    101806.5, 101756.2, 101733.1, 101719.1, 101688.6, 101661.7, 101639.9, 
    101625,
  102163.8, 102122.9, 102092.5, 102047.7, 102007.3, 101963.1, 101928, 
    101882.3, 101847.5, 101836.6, 101806.8, 101773.1, 101748.3, 101724.7, 
    101710.4,
  102158.1, 102128, 102111.1, 102075.4, 102043.2, 102004.5, 101968.4, 
    101929.9, 101915.4, 101893.2, 101863.8, 101840.3, 101807.4, 101782.6, 
    101769.5,
  102136.7, 102114.3, 102106.3, 102076.8, 102050.9, 102022.6, 101986.2, 
    101963.1, 101947.1, 101926.3, 101905.8, 101869.4, 101846.7, 101838.4, 
    101832.8,
  102672.7, 102584, 102479.4, 102380.9, 102273.1, 102171.7, 102063.2, 101955, 
    101854.8, 101746.4, 101636, 101527.7, 101420.9, 101323.4, 101230.2,
  102733.8, 102647.1, 102552, 102463.2, 102363.2, 102266.7, 102166.1, 
    102062.6, 101960.3, 101859.1, 101758, 101656.1, 101558.1, 101462.1, 
    101368.6,
  102805.8, 102733.1, 102646.8, 102556.9, 102458.4, 102354.5, 102249.4, 
    102146.1, 102043.5, 101943.2, 101846.1, 101751.8, 101661.3, 101573.8, 
    101491.9,
  102850.7, 102788.8, 102714.8, 102633.8, 102545.9, 102451.5, 102351.6, 
    102250.9, 102150.4, 102050.9, 101953.6, 101862.5, 101774.2, 101692.7, 
    101615,
  102893, 102839.7, 102778.8, 102710.4, 102629.1, 102540.6, 102445.7, 102348, 
    102249.8, 102154.9, 102060.2, 101971.1, 101884, 101803.6, 101730.8,
  102922.5, 102878.2, 102827.1, 102764.6, 102695.5, 102618.7, 102534.3, 
    102447.5, 102355.8, 102265.4, 102177.1, 102091, 102007.5, 101929, 101858.5,
  102940.3, 102903.5, 102865.5, 102812.9, 102752.2, 102686.4, 102611.2, 
    102533, 102449.6, 102365.4, 102281.6, 102201.9, 102123.7, 102049.5, 
    101980.4,
  102945.4, 102914.7, 102887.1, 102843.1, 102791.6, 102732.5, 102670.2, 
    102602.4, 102531.3, 102456.8, 102380.2, 102305.8, 102234.4, 102163.6, 
    102098,
  102928.8, 102910.3, 102893.7, 102855.7, 102819, 102767.5, 102716.9, 
    102656.6, 102594.4, 102528.1, 102460.8, 102391.6, 102326.6, 102261.8, 
    102199.9,
  102902.2, 102887.1, 102880.9, 102851.9, 102821.9, 102779.3, 102737.3, 
    102686.4, 102633.2, 102577.8, 102520, 102459.2, 102397.8, 102337.3, 
    102281.5 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
