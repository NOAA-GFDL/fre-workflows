netcdf atmos_daily.00010101-00010701.pr.tile5 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pr(time, grid_yt, grid_xt) ;
		pr:_FillValue = 1.e+20f ;
		pr:missing_value = 1.e+20f ;
		pr:units = "kg m-2 s-1" ;
		pr:long_name = "Precipitation" ;
		pr:cell_methods = "time: mean" ;
		pr:cell_measures = "area: area" ;
		pr:time_avg_info = "average_T1,average_T2,average_DT" ;
		pr:standard_name = "precipitation_flux" ;
		pr:interp_method = "conserve_order1" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:07 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile5.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile5.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pr =
  9.816134e-07, 1.678621e-06, 4.664818e-06, 5.187032e-06, 6.45335e-06, 
    1.436801e-05, 9.249137e-05, 0.0002974612, 0.0004440914, 0.0006232968, 
    0.0006139279, 0.0005943866, 0.0005973899, 0.0004980752, 0.0004329419,
  1.342153e-06, 1.244869e-06, 4.364524e-06, 5.237423e-06, 1.021241e-05, 
    9.908824e-06, 1.606805e-05, 4.661181e-05, 0.000255598, 0.0004670013, 
    0.0005305826, 0.0005464047, 0.0005463288, 0.00053419, 0.0005214045,
  4.149194e-06, 3.951347e-06, 7.572557e-06, 8.574475e-06, 1.191147e-05, 
    1.298931e-05, 1.261761e-05, 1.91915e-05, 1.927366e-05, 5.047521e-05, 
    0.0001087789, 0.0001994395, 0.0002809276, 0.0002875269, 0.0003180819,
  3.730499e-06, 5.301087e-06, 7.369629e-06, 9.423007e-06, 1.10741e-05, 
    1.032675e-05, 1.461238e-05, 1.408202e-05, 1.471724e-05, 1.386566e-05, 
    1.723638e-05, 2.063542e-05, 3.972662e-05, 7.077558e-05, 7.257869e-05,
  8.213956e-07, 1.125492e-06, 2.428405e-06, 5.623193e-06, 8.189284e-06, 
    9.226043e-06, 8.934613e-06, 1.096894e-05, 1.218274e-05, 1.194948e-05, 
    1.162731e-05, 1.193942e-05, 1.111983e-05, 1.132013e-05, 1.075345e-05,
  2.461473e-07, 2.810955e-07, 7.482278e-07, 1.740635e-06, 2.828449e-06, 
    4.089924e-06, 7.019775e-06, 8.175767e-06, 1.023437e-05, 8.886452e-06, 
    9.279584e-06, 1.044499e-05, 1.092655e-05, 1.149805e-05, 9.168725e-06,
  1.900247e-08, 2.340537e-08, 1.107269e-07, 4.613718e-07, 8.906667e-07, 
    1.891735e-06, 3.178534e-06, 4.743949e-06, 5.581455e-06, 8.108123e-06, 
    9.85758e-06, 8.978041e-06, 8.45136e-06, 8.020977e-06, 9.977368e-06,
  1.049792e-08, 1.620063e-08, 1.913641e-08, 2.016969e-08, 1.504261e-07, 
    6.698936e-07, 6.695241e-07, 1.311427e-06, 1.111788e-06, 3.696996e-06, 
    1.139981e-05, 1.392145e-05, 1.075757e-05, 7.968109e-06, 7.725235e-06,
  6.739029e-09, 1.885673e-08, 2.099205e-08, 2.724794e-08, 1.643163e-08, 
    2.779518e-08, 8.870781e-08, 2.771864e-07, 1.69453e-07, 6.592106e-07, 
    1.715277e-06, 5.517925e-06, 9.106365e-06, 1.052975e-05, 1.157994e-05,
  1.138184e-08, 2.787475e-08, 2.486239e-08, 3.414269e-08, 2.564846e-08, 
    1.595849e-08, 3.180646e-08, 1.973124e-08, 7.260748e-08, 1.817047e-07, 
    6.076303e-07, 2.656671e-07, 2.311957e-06, 5.754497e-06, 3.242404e-06,
  7.549204e-06, 3.676303e-06, 1.62896e-06, 2.002317e-06, 1.095254e-05, 
    6.389808e-05, 0.0002532421, 0.0004840804, 0.0003106322, 4.643913e-05, 
    1.147746e-06, 1.184216e-07, 2.86096e-09, 4.171934e-08, 9.736064e-08,
  3.804175e-06, 8.250333e-06, 7.384311e-06, 4.238464e-06, 3.174274e-06, 
    1.563601e-05, 0.0001454505, 0.0004402697, 0.0004312041, 0.0002713233, 
    0.0001087297, 3.156917e-05, 8.868562e-06, 8.810732e-06, 1.691935e-05,
  1.359188e-06, 2.345093e-06, 1.043366e-06, 6.425136e-06, 6.804601e-06, 
    4.794366e-06, 1.239947e-05, 0.0001113696, 0.0003684231, 0.0006182038, 
    0.0004816876, 0.0004200024, 0.000310826, 0.0002171754, 0.0001826872,
  3.344847e-08, 7.13961e-07, 8.176593e-07, 4.619095e-07, 7.790726e-06, 
    6.833717e-06, 3.267565e-06, 4.74526e-06, 5.684411e-05, 0.0001692911, 
    0.0004388771, 0.0005510947, 0.0004679296, 0.0004793778, 0.0004334079,
  5.616161e-09, 2.12503e-07, 7.60638e-07, 5.928585e-07, 9.48932e-07, 
    8.7446e-06, 9.220436e-06, 2.772863e-06, 2.754132e-06, 3.987319e-05, 
    0.000266341, 0.0006325027, 0.0007824808, 0.0007468842, 0.0006814072,
  3.59089e-08, 6.573611e-09, 3.204522e-07, 2.863408e-07, 6.92799e-07, 
    1.131817e-06, 2.64701e-06, 1.194974e-05, 6.323191e-06, 6.810787e-06, 
    0.0001581684, 0.000506701, 0.000765133, 0.0008545257, 0.0008897842,
  8.987658e-11, 1.299788e-08, 1.10741e-08, 1.106638e-07, 3.011801e-07, 
    5.500824e-07, 8.629647e-07, 2.138695e-06, 1.052677e-05, 9.084261e-06, 
    7.361569e-06, 6.087793e-05, 0.0002450753, 0.0003066156, 0.0003224103,
  2.007041e-11, 1.709854e-11, 3.312144e-11, 1.74652e-09, 1.593375e-07, 
    3.45961e-07, 2.565964e-07, 1.124385e-06, 2.697923e-06, 8.235074e-06, 
    1.218372e-05, 7.286063e-06, 7.335989e-06, 1.09279e-05, 2.840479e-05,
  1.773342e-11, 1.988452e-11, 7.811223e-10, 1.226537e-08, 9.768286e-08, 
    3.625573e-07, 4.742317e-07, 3.042837e-07, 9.246147e-07, 5.693372e-06, 
    5.691831e-06, 1.076094e-05, 1.229553e-05, 1.107108e-05, 1.032948e-05,
  3.947613e-12, 3.599153e-11, 1.283244e-09, 4.197928e-09, 3.847293e-09, 
    1.537378e-07, 2.157045e-06, 2.576327e-07, 1.403566e-07, 1.948922e-06, 
    6.415413e-06, 8.263378e-06, 1.370508e-05, 1.184706e-05, 8.941262e-06,
  5.987833e-06, 1.141438e-05, 5.203109e-05, 0.0001505357, 0.0002479537, 
    0.0002823778, 0.0002180825, 0.0001726369, 5.635803e-05, 3.335845e-05, 
    3.445533e-05, 3.973018e-05, 1.158924e-05, 6.182162e-06, 2.092764e-06,
  8.998321e-06, 9.450682e-06, 3.317531e-05, 0.0001223996, 0.0001943434, 
    0.0001660656, 0.0002238201, 0.0001614521, 6.937414e-05, 4.436401e-05, 
    1.957697e-05, 1.414828e-05, 8.605127e-06, 1.168731e-05, 6.517014e-06,
  7.465994e-06, 7.987186e-06, 7.283953e-06, 5.793935e-05, 0.0001160456, 
    0.0001579999, 0.0001423677, 0.0001282701, 0.0001202814, 6.330668e-05, 
    3.991165e-05, 7.914253e-06, 9.924595e-06, 7.978889e-06, 1.659789e-05,
  8.498169e-06, 7.758971e-06, 8.127276e-06, 8.940779e-06, 4.370936e-05, 
    7.135179e-05, 8.396726e-05, 0.0001174797, 0.0001297605, 4.832611e-05, 
    2.636068e-05, 1.215333e-05, 4.010494e-06, 3.659726e-06, 9.42439e-06,
  5.285582e-06, 3.993496e-06, 7.061921e-06, 5.629269e-06, 8.562504e-06, 
    3.611987e-05, 7.933665e-05, 0.0001172735, 0.0001321515, 0.0001849549, 
    0.0001380709, 9.743615e-05, 1.327673e-05, 1.452401e-06, 1.998037e-05,
  6.558617e-06, 6.752793e-06, 6.753097e-06, 7.180104e-06, 4.754672e-06, 
    1.314069e-05, 7.478076e-05, 0.0001796834, 0.000248282, 0.0003036138, 
    0.0004512341, 0.0004254962, 0.0002262042, 0.0001455821, 0.000132443,
  6.803414e-06, 8.303216e-06, 3.758218e-06, 5.698e-06, 9.147038e-06, 
    8.648484e-06, 2.334066e-05, 0.0001653496, 0.0004239844, 0.0005127026, 
    0.0005651346, 0.0006678681, 0.0007048014, 0.0007650791, 0.0007477964,
  6.998542e-06, 1.082507e-05, 5.949746e-06, 3.952795e-06, 5.539945e-06, 
    9.41183e-06, 7.707787e-06, 1.91272e-05, 0.0001797602, 0.0004309531, 
    0.0005499368, 0.0005992433, 0.000679689, 0.0006951465, 0.0008112748,
  6.888699e-06, 1.143514e-05, 9.382572e-06, 6.67499e-06, 6.598601e-06, 
    6.368321e-06, 5.703817e-06, 6.424023e-06, 1.18848e-05, 7.485037e-05, 
    0.0002449958, 0.0003672162, 0.0004202836, 0.0004367389, 0.0004077028,
  1.03204e-05, 6.481123e-06, 1.024948e-05, 8.615227e-06, 8.757415e-06, 
    4.962574e-06, 2.720867e-06, 5.32999e-06, 7.121768e-06, 6.010314e-06, 
    3.095069e-05, 7.985725e-05, 0.0001699955, 0.0002393835, 0.000328021,
  7.160423e-06, 1.282444e-05, 4.03897e-05, 4.347091e-05, 3.146256e-05, 
    1.623416e-05, 3.205046e-05, 6.679442e-05, 7.547323e-05, 5.391117e-05, 
    2.011359e-05, 5.182607e-06, 7.227922e-07, 9.169744e-07, 4.229701e-06,
  1.009066e-05, 1.1584e-05, 2.625236e-05, 5.90217e-05, 4.866534e-05, 
    4.002508e-05, 2.124426e-05, 1.355624e-05, 2.419563e-05, 1.253698e-05, 
    4.255098e-06, 1.158436e-06, 9.51219e-07, 1.784676e-07, 9.703397e-06,
  8.341204e-06, 7.934524e-06, 1.714095e-05, 4.542346e-05, 5.674582e-05, 
    8.217758e-05, 7.005973e-05, 1.650161e-05, 4.464369e-06, 6.851144e-06, 
    3.467749e-06, 7.63736e-07, 3.363763e-06, 7.900503e-07, 8.806839e-07,
  7.630107e-06, 5.566529e-06, 7.357937e-06, 2.471972e-05, 5.260135e-05, 
    6.180877e-05, 8.64195e-05, 5.945321e-05, 1.483066e-05, 4.931568e-06, 
    1.922245e-06, 1.070704e-06, 5.56727e-06, 6.985766e-06, 8.354023e-06,
  7.441765e-06, 6.752685e-06, 7.293525e-06, 1.526487e-05, 4.998449e-05, 
    9.103371e-05, 8.57258e-05, 9.448044e-05, 5.067239e-05, 6.434491e-06, 
    8.73448e-07, 1.413242e-06, 1.446378e-05, 5.804182e-06, 1.463642e-05,
  7.798787e-06, 6.989105e-06, 6.652671e-06, 6.91414e-06, 4.752977e-05, 
    0.000166765, 0.0002212076, 0.0002404319, 7.934034e-05, 2.620712e-05, 
    1.130342e-06, 4.872758e-06, 6.492839e-06, 1.632054e-05, 3.224265e-05,
  7.470073e-06, 9.605387e-06, 8.802257e-06, 5.71074e-06, 3.017353e-05, 
    0.0001563894, 0.000331021, 0.0003835563, 0.000211091, 6.563804e-05, 
    2.258903e-05, 4.479903e-06, 1.231065e-05, 5.433594e-05, 2.676538e-05,
  8.400827e-06, 7.929285e-06, 8.623795e-06, 6.944282e-06, 7.924838e-06, 
    8.121072e-05, 0.0002217965, 0.0003394336, 0.0003495867, 0.0001991294, 
    5.65074e-05, 4.969993e-05, 2.485363e-05, 8.807175e-05, 3.272027e-05,
  7.380931e-06, 1.093864e-05, 9.116041e-06, 8.569677e-06, 7.762063e-06, 
    2.848545e-05, 0.0001354617, 0.0002164032, 0.0003279708, 0.0003768666, 
    0.0003089284, 0.0002497489, 0.0002793109, 0.0003103236, 0.0001104685,
  8.137376e-06, 8.705456e-06, 1.017351e-05, 9.657867e-06, 7.310205e-06, 
    9.431848e-06, 7.409101e-05, 0.0001720563, 0.0002249832, 0.0003576269, 
    0.0004388054, 0.0004719223, 0.0004368157, 0.0003229475, 0.0002276451,
  0.0001330435, 0.0001781969, 0.0001662677, 0.0001599493, 0.0001629849, 
    0.0001697526, 0.0001666436, 0.0001401416, 0.0001056219, 6.896532e-05, 
    4.354501e-05, 3.616558e-05, 5.367217e-05, 0.0001463464, 0.000191438,
  0.000123297, 0.0001564702, 0.0001646729, 0.0001657891, 0.0001718454, 
    0.0001711427, 0.0001830518, 0.0001826416, 0.0001481199, 9.230619e-05, 
    4.151309e-05, 1.952162e-05, 5.592639e-05, 0.0001420622, 0.0002260805,
  0.000138277, 0.0001502489, 0.0001742839, 0.0001850796, 0.0001902875, 
    0.0001895735, 0.000175749, 0.0001611864, 0.0001247679, 7.366089e-05, 
    2.869341e-05, 2.253205e-05, 6.183505e-05, 0.0001283092, 0.0002946478,
  0.000118936, 0.0001646285, 0.0001850693, 0.0002080615, 0.000209297, 
    0.0001932359, 0.0001609203, 0.0001265456, 8.725305e-05, 5.02744e-05, 
    2.555413e-05, 1.686085e-05, 5.675351e-05, 8.558777e-05, 4.769176e-05,
  0.000105515, 0.000145942, 0.0001876737, 0.0002299158, 0.0002226526, 
    0.0002002605, 0.0001581514, 0.0001119359, 6.872604e-05, 3.94079e-05, 
    1.929308e-05, 2.244953e-05, 4.892893e-05, 4.219249e-05, 4.509541e-05,
  8.694766e-05, 0.0001192892, 0.0001726461, 0.0002146005, 0.0002303749, 
    0.0002187553, 0.0001689932, 0.0001236278, 5.837313e-05, 2.831656e-05, 
    1.528363e-05, 1.664252e-05, 2.547314e-05, 3.014567e-05, 8.104395e-06,
  4.445936e-05, 7.072368e-05, 0.0001190698, 0.0001845894, 0.0002227366, 
    0.0002298131, 0.0001821427, 0.0001382823, 7.180409e-05, 2.17153e-05, 
    1.586195e-05, 1.235122e-05, 1.978363e-05, 1.78434e-05, 8.330086e-06,
  1.017953e-05, 2.398793e-05, 6.890832e-05, 0.0001251766, 0.0001851796, 
    0.0002261639, 0.0002180697, 0.0001646308, 0.0001055847, 3.695092e-05, 
    1.75549e-05, 1.525536e-05, 1.127844e-05, 2.019978e-05, 1.219914e-05,
  4.118099e-06, 5.64449e-06, 1.92776e-05, 6.752738e-05, 0.0001437408, 
    0.000204308, 0.0002443217, 0.0002079956, 0.0001362489, 7.437291e-05, 
    2.886897e-05, 1.745172e-05, 1.004811e-05, 1.657222e-05, 1.787812e-06,
  3.759966e-06, 2.531353e-06, 4.951872e-06, 1.844811e-05, 8.09337e-05, 
    0.0001652454, 0.0002305239, 0.0002687516, 0.0001860005, 0.0001144008, 
    5.037947e-05, 3.069769e-05, 1.560356e-05, 1.478249e-05, 1.923453e-06,
  0.0002164863, 0.0002660363, 0.0003733526, 0.0003285779, 0.0001708998, 
    4.666859e-05, 6.372838e-06, 6.721956e-06, 9.154349e-06, 1.010325e-05, 
    6.426739e-06, 2.249938e-06, 4.413589e-06, 4.483601e-07, 1.514539e-06,
  0.0002632197, 0.0003105392, 0.000301477, 0.0002413806, 0.0001422676, 
    2.640955e-05, 7.76352e-06, 1.062813e-05, 1.629655e-05, 1.357225e-05, 
    1.055329e-05, 1.056025e-05, 3.991381e-06, 1.45329e-06, 1.311676e-06,
  0.0003165699, 0.0003110161, 0.0002774079, 0.0002073807, 0.0001120666, 
    2.836193e-05, 1.331587e-05, 1.897645e-05, 2.064502e-05, 1.411579e-05, 
    1.761295e-05, 9.021548e-06, 3.91654e-06, 4.923293e-06, 1.186528e-06,
  0.0003185079, 0.0002925575, 0.0002656341, 0.0002228255, 0.0001104603, 
    2.282357e-05, 1.85825e-05, 2.128581e-05, 2.379892e-05, 1.658884e-05, 
    1.139033e-05, 1.32504e-05, 5.671355e-06, 9.821288e-07, 6.110362e-07,
  0.0002543695, 0.0002341126, 0.0002199116, 0.0001900633, 9.897808e-05, 
    3.081916e-05, 2.357486e-05, 2.034311e-05, 2.195849e-05, 1.641181e-05, 
    1.126138e-05, 1.155623e-05, 3.018704e-06, 8.557084e-06, 1.114082e-05,
  0.0001836734, 0.0001662924, 0.0001799762, 0.0001729167, 9.580164e-05, 
    3.794911e-05, 3.232504e-05, 2.41779e-05, 1.562106e-05, 1.459044e-05, 
    9.254239e-06, 1.486798e-05, 5.31156e-06, 3.411005e-06, 1.711562e-05,
  0.0001842237, 0.0001365865, 0.0001266136, 0.0001215966, 9.403275e-05, 
    5.402862e-05, 3.110544e-05, 2.03582e-05, 1.12531e-05, 1.02249e-05, 
    7.098259e-06, 3.927981e-06, 8.419825e-06, 6.524139e-06, 5.465503e-07,
  0.000194462, 0.000166387, 0.0001288642, 9.26609e-05, 7.880016e-05, 
    6.348691e-05, 4.712666e-05, 1.885848e-05, 6.320423e-06, 4.937716e-06, 
    5.285521e-06, 3.780931e-06, 1.276079e-05, 1.101134e-05, 2.451538e-07,
  0.0001773712, 0.0001581216, 0.0001329294, 9.052997e-05, 6.248846e-05, 
    5.668536e-05, 3.923753e-05, 1.887749e-05, 7.16611e-06, 6.973174e-06, 
    6.081622e-06, 2.664207e-06, 1.710466e-05, 1.740274e-05, 1.134766e-07,
  0.0001249873, 0.0001376718, 0.000134803, 0.0001263195, 8.396176e-05, 
    5.920891e-05, 3.865149e-05, 1.708064e-05, 9.130833e-06, 9.787142e-06, 
    5.002247e-06, 1.133162e-06, 2.469395e-05, 3.379749e-05, 9.110248e-07,
  0.0002035361, 0.0001836317, 0.0001182715, 7.087482e-05, 0.0001099351, 
    0.0001391404, 0.0001897888, 0.0002393942, 0.0003573897, 0.0001858153, 
    6.346656e-06, 1.536223e-07, 2.342856e-08, 9.693554e-10, 6.816175e-10,
  0.0001698147, 0.0001771853, 0.0001407895, 7.388436e-05, 0.0001629711, 
    0.0002096974, 0.0002514934, 0.0003513692, 0.0004338666, 0.0001329022, 
    1.844811e-07, 1.821539e-08, 3.446688e-09, 1.374096e-09, 1.103784e-09,
  0.0001229053, 0.0001592995, 0.0001420257, 9.293894e-05, 0.0002237436, 
    0.0002926929, 0.0002951804, 0.0004898699, 0.0004821536, 4.854976e-05, 
    4.053348e-08, 1.335615e-08, 4.356935e-09, 1.519846e-08, 1.551485e-07,
  0.0001418638, 0.000128124, 0.0001126746, 0.0001150842, 0.0002490305, 
    0.0003363819, 0.0003439387, 0.0006170676, 0.0004789122, 7.940158e-07, 
    1.723708e-08, 1.134884e-07, 7.919854e-07, 1.058603e-06, 6.887991e-07,
  0.000214088, 0.0001539356, 0.0001017506, 0.0001411646, 0.0002604678, 
    0.0003343821, 0.0004056973, 0.0007156742, 0.0004135642, 1.018998e-07, 
    2.80661e-07, 1.81856e-06, 2.401528e-06, 1.265559e-06, 7.337178e-07,
  0.0003360385, 0.0002479809, 0.0001588423, 0.0002060115, 0.0002630922, 
    0.0002961594, 0.0004471956, 0.0007617818, 0.0003392736, 1.494896e-07, 
    2.270257e-06, 5.097611e-06, 2.638e-06, 9.149622e-07, 4.496326e-07,
  0.0004422426, 0.0003567273, 0.0002366443, 0.0002809477, 0.0002448443, 
    0.0002744525, 0.000425786, 0.0007646133, 0.0003234102, 1.978996e-06, 
    7.562101e-06, 7.421022e-06, 1.718714e-06, 6.698023e-07, 3.887565e-07,
  0.0005268729, 0.0004613682, 0.0003437709, 0.000338236, 0.0002539047, 
    0.0002789413, 0.0004342499, 0.0007366806, 0.0003043429, 6.229953e-06, 
    1.053541e-05, 5.610238e-06, 6.817054e-07, 2.957013e-07, 5.751179e-08,
  0.0006150464, 0.0005726008, 0.0004633265, 0.0003827014, 0.000274025, 
    0.0003015491, 0.0004452898, 0.000676797, 0.0002694354, 1.104257e-05, 
    8.299009e-06, 2.02419e-06, 1.101226e-07, 4.145402e-08, 7.900648e-09,
  0.0006553804, 0.0006419963, 0.0005230969, 0.000436242, 0.0002959319, 
    0.0003264221, 0.0004640701, 0.0006288987, 0.0002482853, 1.050001e-05, 
    2.554032e-06, 2.88624e-07, 3.032536e-08, 1.464788e-08, 3.463053e-09,
  0.0001602743, 0.0002051515, 0.0001960823, 0.0001554569, 0.0002054958, 
    0.0001394345, 0.0001293678, 0.0001253133, 1.955754e-05, 1.819443e-07, 
    5.561891e-08, 5.194599e-08, 6.750238e-08, 7.166314e-08, 2.452777e-07,
  0.0001482164, 0.0002173814, 0.0002560925, 0.0001898947, 0.0002207739, 
    0.000166636, 0.0001517019, 0.0001234488, 6.454979e-07, 5.628794e-08, 
    4.355504e-08, 4.118023e-08, 6.433817e-08, 1.779013e-07, 1.576382e-07,
  0.0001371637, 0.0002270713, 0.0003089045, 0.0002315518, 0.0002484633, 
    0.0001752171, 0.0001693739, 0.0001038902, 2.546819e-07, 3.071725e-08, 
    1.935593e-08, 7.706388e-09, 2.570847e-08, 9.88477e-08, 1.551306e-07,
  0.0001275749, 0.0002024877, 0.0003355179, 0.0002712158, 0.0002595109, 
    0.0001660047, 0.0001565525, 6.875656e-05, 7.602315e-08, 2.098657e-08, 
    4.687065e-08, 9.573109e-08, 1.894922e-07, 7.590939e-07, 4.270787e-07,
  0.0001277294, 0.0001760161, 0.0003335052, 0.0002964769, 0.0002708515, 
    0.0001672298, 0.0001370496, 3.947217e-05, 5.952836e-08, 2.29524e-08, 
    2.767504e-08, 4.370224e-08, 1.153514e-07, 1.641514e-07, 8.27807e-08,
  0.0001412738, 0.0001592247, 0.0003250724, 0.0003402981, 0.0002646991, 
    0.0001820292, 0.0001420822, 2.470995e-05, 7.590521e-08, 1.572989e-08, 
    7.590613e-09, 4.056906e-08, 2.031546e-07, 8.331412e-07, 9.994488e-07,
  0.0001499893, 0.000141496, 0.0003124226, 0.000386984, 0.0002568111, 
    0.0002060164, 0.0001519753, 2.431274e-05, 1.027798e-07, 3.04155e-08, 
    9.147429e-08, 2.150646e-07, 2.118978e-07, 1.234411e-07, 1.278311e-07,
  0.0001611629, 0.0001392642, 0.0002897171, 0.000404063, 0.0002275997, 
    0.0002106163, 0.0001598406, 4.378625e-05, 2.529642e-07, 2.643711e-08, 
    7.431616e-08, 1.988253e-07, 6.245017e-08, 9.724025e-09, 4.929423e-08,
  0.0001577016, 0.0001289595, 0.0002399524, 0.0003693871, 0.0002184116, 
    0.0002210321, 0.0001676936, 7.596714e-05, 2.753595e-06, 2.680135e-08, 
    2.616085e-08, 1.931212e-08, 2.415272e-08, 4.286357e-10, 6.571781e-10,
  0.0001411426, 0.0001148554, 0.0001812713, 0.0002848546, 0.0002324075, 
    0.0002218017, 0.000162488, 0.0001223102, 2.441758e-05, 3.637241e-08, 
    1.353463e-08, 8.790214e-10, 2.606704e-09, 3.189994e-09, 9.80461e-09,
  0.0002025868, 0.0002379446, 0.0002774377, 0.0002584809, 0.0002709883, 
    0.000212418, 9.120243e-05, 2.004092e-05, 3.927641e-06, 4.59641e-06, 
    5.372838e-06, 5.29678e-06, 4.452644e-06, 5.475374e-06, 3.098776e-06,
  0.0001900659, 0.0002505851, 0.0002834327, 0.000275095, 0.0002885812, 
    0.0002683126, 9.105074e-05, 2.353535e-05, 5.090265e-06, 5.331367e-06, 
    5.478559e-06, 4.668318e-06, 5.155973e-06, 5.694165e-06, 5.313874e-06,
  0.0002055302, 0.0002977776, 0.0003042692, 0.0003150297, 0.0003149604, 
    0.000339811, 8.768479e-05, 2.218848e-05, 6.055849e-06, 5.575906e-06, 
    4.393577e-06, 3.789467e-06, 2.989447e-06, 3.976024e-06, 3.506383e-06,
  0.0002307787, 0.0003252221, 0.0003338525, 0.0003333132, 0.0002982197, 
    0.0003546177, 7.237844e-05, 1.632845e-05, 5.76195e-06, 4.379329e-06, 
    4.632223e-06, 5.828618e-06, 4.675509e-06, 5.152559e-06, 3.313069e-06,
  0.0002560056, 0.0003484296, 0.0003724444, 0.0003404417, 0.0002760804, 
    0.0003447534, 6.508519e-05, 7.953149e-06, 5.023813e-06, 3.691619e-06, 
    4.016419e-06, 4.13283e-06, 3.004878e-06, 1.59275e-06, 9.835823e-07,
  0.0002736135, 0.0003410903, 0.0004045482, 0.0003527493, 0.000294112, 
    0.0003363839, 6.763791e-05, 4.819972e-06, 3.199756e-06, 3.455231e-06, 
    3.622415e-06, 4.454624e-06, 3.218371e-06, 5.090175e-06, 2.429368e-06,
  0.0002790776, 0.0003348191, 0.000414923, 0.0003752552, 0.0003284042, 
    0.000324199, 7.469647e-05, 3.90593e-06, 3.131238e-06, 2.903658e-06, 
    3.765351e-06, 5.399486e-06, 7.307196e-06, 4.599009e-06, 2.951214e-06,
  0.0002639198, 0.0003115978, 0.0004142919, 0.000423135, 0.0003923722, 
    0.0003106892, 0.0001039018, 3.809251e-06, 3.525966e-06, 3.378894e-06, 
    4.379359e-06, 5.646611e-06, 4.960445e-06, 2.05017e-06, 2.040946e-06,
  0.0002302218, 0.0003003455, 0.0004301443, 0.0005039603, 0.0004543084, 
    0.0003007578, 0.0001627168, 6.936541e-06, 3.611641e-06, 3.666904e-06, 
    4.536309e-06, 5.273397e-06, 2.62036e-06, 6.369425e-07, 1.006182e-06,
  0.0002079489, 0.0002921235, 0.0004347294, 0.0006255637, 0.0005377406, 
    0.0003042251, 0.0002038661, 1.559019e-05, 3.229301e-06, 2.344314e-06, 
    3.259958e-06, 4.858563e-06, 3.616775e-06, 1.396982e-06, 2.09698e-06,
  7.823324e-05, 0.0001179271, 0.0001311762, 0.0001042063, 0.0001336032, 
    0.0002000427, 0.0001860226, 0.0001224383, 5.843872e-05, 1.047976e-05, 
    4.348488e-06, 2.299476e-06, 2.855557e-06, 2.36392e-06, 6.181544e-06,
  6.259478e-05, 0.0001014232, 0.0001461938, 0.0001029068, 9.654028e-05, 
    0.000170934, 0.0001989634, 0.0001472828, 9.699705e-05, 1.89967e-05, 
    3.507085e-06, 2.050778e-06, 3.375174e-06, 1.928423e-06, 4.446111e-06,
  4.056821e-05, 8.115821e-05, 0.0001390385, 0.0001274423, 8.934829e-05, 
    0.0001662136, 0.0002480431, 0.0001979333, 0.0001317059, 4.381876e-05, 
    7.926391e-06, 6.714348e-06, 2.065711e-06, 1.54739e-06, 3.85956e-06,
  3.07761e-05, 5.077252e-05, 0.000108864, 0.0001391895, 0.0001019696, 
    0.0001672315, 0.0003058109, 0.0002317008, 0.0001381938, 7.146178e-05, 
    1.688694e-05, 7.97519e-06, 3.051795e-06, 8.317283e-07, 5.143836e-06,
  3.251891e-05, 3.917046e-05, 7.69709e-05, 0.0001182913, 0.0001150245, 
    0.000162386, 0.0003196637, 0.0002509566, 0.0001255793, 8.257922e-05, 
    2.748313e-05, 9.243029e-06, 6.163822e-06, 1.519408e-06, 4.136724e-06,
  2.673201e-05, 2.656927e-05, 5.29397e-05, 8.919155e-05, 0.0001075389, 
    0.0001510175, 0.0002812474, 0.0003030052, 0.0001299944, 7.812541e-05, 
    3.577039e-05, 9.884755e-06, 7.269382e-06, 1.422644e-06, 2.692953e-06,
  2.58815e-05, 2.174263e-05, 2.272803e-05, 5.011646e-05, 8.808174e-05, 
    0.0001388959, 0.0002487952, 0.0003500376, 0.000145449, 8.316718e-05, 
    4.933591e-05, 1.376437e-05, 8.712223e-06, 4.688524e-06, 3.421124e-06,
  3.994939e-05, 2.31202e-05, 1.737371e-05, 2.265269e-05, 5.935437e-05, 
    0.0001282008, 0.000211228, 0.000351834, 0.0001642323, 8.108485e-05, 
    5.905105e-05, 1.719089e-05, 6.528519e-06, 2.152052e-06, 4.217997e-06,
  5.679967e-05, 2.934273e-05, 1.907012e-05, 1.60096e-05, 2.509352e-05, 
    0.0001033018, 0.000182053, 0.0003203854, 0.0002088455, 8.825526e-05, 
    6.37234e-05, 2.466582e-05, 6.734121e-06, 1.39619e-06, 4.293174e-06,
  7.687388e-05, 3.796057e-05, 2.3658e-05, 1.889747e-05, 1.292083e-05, 
    7.220639e-05, 0.0001635105, 0.0002746596, 0.0002598441, 0.0001012361, 
    6.882069e-05, 3.346846e-05, 8.408228e-06, 2.354818e-06, 5.211977e-06,
  4.232287e-05, 5.246201e-05, 7.067039e-05, 9.221231e-05, 0.000176873, 
    0.0001796208, 6.224716e-05, 2.302866e-05, 1.109061e-05, 1.159325e-05, 
    1.517092e-05, 1.660098e-05, 1.011568e-05, 3.983139e-06, 3.278617e-06,
  6.803855e-05, 4.798883e-05, 6.753614e-05, 9.306415e-05, 0.0001980591, 
    0.0002134568, 7.953242e-05, 2.350887e-05, 1.22142e-05, 1.105996e-05, 
    1.751524e-05, 1.770297e-05, 4.519189e-06, 2.080448e-06, 3.149662e-06,
  5.681026e-05, 6.208495e-05, 4.936741e-05, 9.830129e-05, 0.0002171848, 
    0.0002592988, 0.0001023273, 3.04257e-05, 1.58053e-05, 1.166917e-05, 
    2.235785e-05, 2.266858e-05, 7.475065e-06, 2.102825e-06, 3.74687e-06,
  6.641197e-05, 5.40249e-05, 5.267364e-05, 9.685452e-05, 0.0002223929, 
    0.0003031377, 0.0001394081, 3.506051e-05, 2.114654e-05, 1.401905e-05, 
    2.816343e-05, 2.318541e-05, 6.992599e-06, 2.581855e-06, 3.645034e-06,
  5.200447e-05, 4.425896e-05, 6.944682e-05, 0.0001130302, 0.0002398299, 
    0.0003545887, 0.0001789123, 4.512849e-05, 2.84894e-05, 1.541166e-05, 
    2.897795e-05, 2.098368e-05, 6.967087e-06, 1.393479e-06, 4.093495e-06,
  5.785954e-05, 7.5699e-05, 6.7615e-05, 0.0001198151, 0.0002628676, 
    0.0004369901, 0.0002267637, 4.850979e-05, 3.411638e-05, 1.382684e-05, 
    2.394036e-05, 1.453642e-05, 5.917847e-06, 3.748002e-06, 2.623407e-06,
  0.0001036163, 5.65593e-05, 9.767958e-05, 0.0001363539, 0.0002868572, 
    0.000492986, 0.0002871639, 5.83507e-05, 3.107762e-05, 1.241194e-05, 
    1.640685e-05, 9.888739e-06, 6.352648e-06, 3.183151e-06, 2.468253e-06,
  0.0001099643, 9.368237e-05, 8.6835e-05, 0.0001414568, 0.000288597, 
    0.0005500732, 0.0003584248, 6.71722e-05, 3.884537e-05, 1.127544e-05, 
    9.836409e-06, 6.051594e-06, 5.566558e-06, 3.14308e-06, 6.352212e-06,
  0.0001113448, 7.613748e-05, 0.0001021964, 0.0001253803, 0.000300789, 
    0.0006091017, 0.0004441959, 8.223789e-05, 4.486648e-05, 8.699919e-06, 
    6.159898e-06, 6.159943e-06, 6.032896e-06, 4.285553e-06, 7.309071e-06,
  0.0001018116, 7.909483e-05, 8.649217e-05, 0.0001247119, 0.0002771636, 
    0.0006153019, 0.0005195605, 0.0001438242, 5.54359e-05, 9.488147e-06, 
    4.903463e-06, 6.29674e-06, 4.872961e-06, 3.892e-06, 4.187397e-06,
  3.01934e-05, 1.684482e-05, 9.796016e-06, 7.458898e-06, 5.845785e-06, 
    4.306709e-06, 4.696269e-06, 3.443509e-06, 2.957466e-06, 2.298791e-06, 
    3.850708e-06, 7.597981e-06, 2.327374e-05, 3.897088e-05, 1.15639e-05,
  3.598016e-05, 1.318555e-05, 8.446729e-06, 5.378674e-06, 4.713374e-06, 
    3.378924e-06, 4.076895e-06, 3.593174e-06, 3.422342e-06, 2.537514e-06, 
    4.873096e-06, 5.412088e-06, 3.334575e-05, 4.720098e-05, 1.325137e-05,
  3.362948e-05, 1.73643e-05, 1.023982e-05, 7.325931e-06, 4.218384e-06, 
    3.334114e-06, 4.3122e-06, 5.791193e-06, 3.577171e-06, 3.126007e-06, 
    4.598584e-06, 9.498447e-06, 4.036507e-05, 4.889035e-05, 1.014443e-05,
  3.034702e-05, 1.945362e-05, 1.361236e-05, 6.603711e-06, 4.617474e-06, 
    5.10239e-06, 5.454942e-06, 7.36177e-06, 4.615962e-06, 4.455846e-06, 
    5.095006e-06, 8.191449e-06, 3.69213e-05, 4.946114e-05, 6.745971e-06,
  3.52138e-05, 2.444034e-05, 1.631509e-05, 8.398363e-06, 5.120162e-06, 
    6.010009e-06, 7.292037e-06, 8.012166e-06, 6.389161e-06, 5.317848e-06, 
    6.545661e-06, 8.921989e-06, 3.407944e-05, 3.658811e-05, 4.778844e-06,
  3.706065e-05, 2.300384e-05, 1.567791e-05, 9.310441e-06, 6.297098e-06, 
    5.132452e-06, 7.937863e-06, 8.138746e-06, 5.47279e-06, 4.790102e-06, 
    8.17169e-06, 1.500808e-05, 3.118858e-05, 3.629268e-05, 1.403839e-06,
  4.054091e-05, 2.605297e-05, 1.400871e-05, 9.225349e-06, 6.83066e-06, 
    6.184478e-06, 1.124741e-05, 1.042592e-05, 7.119225e-06, 4.920111e-06, 
    1.326291e-05, 1.972669e-05, 4.435135e-05, 2.393563e-05, 3.104748e-06,
  4.251154e-05, 2.908829e-05, 1.730773e-05, 9.373035e-06, 7.564555e-06, 
    5.878001e-06, 1.057897e-05, 8.168883e-06, 8.264849e-06, 7.375865e-06, 
    1.974242e-05, 2.476793e-05, 4.048633e-05, 3.123418e-05, 3.326541e-06,
  4.678101e-05, 3.539232e-05, 1.623249e-05, 1.089721e-05, 7.076894e-06, 
    1.004747e-05, 8.406633e-06, 7.926703e-06, 5.76304e-06, 8.984612e-06, 
    2.678586e-05, 2.484402e-05, 6.105081e-05, 2.923772e-05, 3.759233e-06,
  5.391629e-05, 3.547612e-05, 1.794372e-05, 1.093897e-05, 1.065426e-05, 
    8.010664e-06, 5.190405e-06, 7.457254e-06, 8.207146e-06, 8.542428e-06, 
    2.269251e-05, 2.697431e-05, 7.424562e-05, 2.383829e-05, 4.066481e-06,
  3.913341e-06, 2.876525e-06, 2.155659e-06, 6.501011e-07, 1.860648e-07, 
    8.800763e-08, 2.482952e-08, 2.037285e-09, 4.242831e-12, 3.458219e-09, 
    5.618795e-09, 2.283062e-07, 1.811274e-06, 1.818515e-05, 3.102758e-05,
  5.100441e-06, 2.961895e-06, 1.655451e-06, 4.786688e-07, 1.156179e-07, 
    1.669018e-07, 3.885672e-08, 1.519247e-11, 2.249681e-12, 2.946127e-11, 
    2.509973e-08, 1.137749e-07, 3.470247e-07, 1.027866e-05, 3.70364e-05,
  8.096091e-06, 4.368972e-06, 2.001909e-06, 8.980084e-07, 3.831159e-07, 
    1.857305e-07, 2.094743e-07, 3.890459e-08, 3.693395e-08, 5.616647e-09, 
    2.241071e-08, 8.799054e-09, 5.747883e-07, 1.183923e-05, 3.20933e-05,
  1.038552e-05, 5.670366e-06, 3.482649e-06, 1.943067e-06, 7.203216e-07, 
    4.16837e-07, 3.546753e-07, 2.352143e-07, 1.206533e-07, 1.565729e-10, 
    6.762676e-08, 4.345851e-09, 9.183283e-07, 1.224944e-05, 2.22769e-05,
  1.268012e-05, 6.620533e-06, 6.852934e-06, 1.939898e-06, 6.838059e-07, 
    5.93174e-07, 4.820186e-07, 2.990159e-07, 2.431271e-07, 7.17256e-10, 
    2.356733e-08, 1.530739e-09, 1.414052e-06, 1.331399e-05, 2.302675e-05,
  1.308844e-05, 9.894668e-06, 1.02013e-05, 3.311954e-06, 1.125861e-06, 
    7.402885e-07, 6.765728e-07, 4.315204e-07, 3.282941e-07, 3.432082e-10, 
    1.194333e-07, 2.286903e-08, 1.542959e-06, 1.667538e-05, 1.742018e-05,
  1.881795e-05, 1.328371e-05, 9.670329e-06, 5.974536e-06, 1.419073e-06, 
    9.945129e-07, 1.12178e-06, 6.870558e-07, 4.036949e-07, 1.639703e-09, 
    1.758521e-07, 1.843666e-08, 6.013128e-07, 8.120752e-06, 1.770664e-05,
  3.043619e-05, 1.785302e-05, 1.273948e-05, 8.419777e-06, 2.920471e-06, 
    1.597345e-06, 1.018811e-06, 8.464515e-07, 5.87497e-07, 3.114448e-08, 
    1.997407e-07, 3.888791e-08, 5.003642e-07, 1.004248e-05, 1.55705e-05,
  3.673227e-05, 1.947576e-05, 1.459093e-05, 1.016172e-05, 4.639741e-06, 
    2.692671e-06, 2.152169e-06, 7.253028e-07, 6.167118e-07, 2.22701e-08, 
    7.292694e-08, 1.199681e-07, 8.904869e-07, 1.705423e-05, 1.265134e-05,
  3.698395e-05, 2.481439e-05, 2.043734e-05, 1.177368e-05, 7.033856e-06, 
    3.97099e-06, 1.731792e-06, 8.834904e-07, 6.759489e-07, 4.625316e-08, 
    4.232879e-07, 2.02288e-07, 7.040459e-06, 2.494504e-05, 1.225556e-05,
  2.469872e-05, 1.70902e-05, 1.331377e-05, 1.221596e-05, 6.965086e-06, 
    1.916761e-06, 1.122407e-06, 9.78402e-07, 1.788457e-06, 3.356422e-06, 
    3.78413e-06, 5.440566e-06, 1.060827e-05, 1.407424e-05, 1.035124e-05,
  1.768855e-05, 7.512541e-06, 1.379273e-05, 1.032893e-05, 8.555102e-06, 
    2.846893e-06, 1.720162e-06, 1.228516e-06, 1.405847e-06, 3.007624e-06, 
    3.032567e-06, 3.938465e-06, 7.891006e-06, 8.825473e-06, 1.095627e-05,
  1.576095e-05, 5.482208e-06, 1.0875e-05, 1.009337e-05, 6.265625e-06, 
    4.185404e-06, 1.197221e-06, 1.501063e-06, 1.524204e-06, 2.091551e-06, 
    3.318731e-06, 1.868442e-06, 4.829915e-06, 6.842405e-06, 1.580693e-05,
  1.324499e-05, 4.714188e-06, 8.71855e-06, 7.519893e-06, 5.415393e-06, 
    3.727793e-06, 1.837381e-06, 1.526773e-06, 1.385852e-06, 1.426588e-06, 
    9.611293e-07, 2.038746e-06, 2.517964e-06, 9.892447e-06, 9.036518e-06,
  1.113464e-05, 4.607463e-06, 2.813578e-06, 4.659195e-06, 3.857977e-06, 
    3.077068e-06, 2.036622e-06, 1.897186e-06, 1.048412e-07, 4.85857e-07, 
    9.057169e-07, 1.171993e-06, 1.439357e-06, 3.699003e-06, 9.715995e-06,
  1.522718e-05, 3.488383e-06, 1.762224e-06, 3.267619e-06, 4.341292e-06, 
    3.517093e-06, 1.813896e-06, 1.045036e-06, 8.28346e-08, 5.634602e-08, 
    6.206936e-08, 1.687498e-07, 3.234874e-07, 1.91322e-07, 1.712315e-06,
  4.627217e-05, 5.891476e-06, 2.360388e-06, 1.213083e-06, 2.18303e-06, 
    3.144641e-06, 2.324682e-06, 1.195169e-06, 6.853031e-07, 6.048379e-08, 
    7.328966e-09, 2.589501e-09, 3.919104e-10, 7.963893e-10, 8.967559e-08,
  0.0001030481, 2.678175e-05, 2.076517e-06, 1.129819e-06, 1.506497e-06, 
    2.10493e-06, 2.36364e-06, 1.15568e-06, 3.81258e-07, 1.328865e-07, 
    3.039866e-08, 6.849376e-08, 3.906533e-10, 2.359879e-09, 4.066247e-08,
  0.0001276813, 4.587341e-05, 4.092829e-06, 1.25282e-06, 1.655495e-06, 
    2.005035e-06, 1.733593e-06, 1.399948e-06, 9.163831e-08, 4.472927e-08, 
    3.493512e-08, 1.738355e-08, 1.542967e-08, 7.498133e-08, 2.536365e-07,
  0.0001207882, 6.179791e-05, 1.058796e-05, 2.249078e-06, 1.606873e-06, 
    1.389811e-06, 7.333087e-07, 8.387236e-07, 3.88363e-07, 1.765054e-07, 
    3.032949e-07, 7.326575e-08, 2.189784e-07, 6.402434e-08, 2.435773e-07,
  0.0001330839, 0.0002298933, 0.0002568801, 0.0002331414, 0.0002383229, 
    0.0003033633, 0.0002426684, 0.0001304698, 4.776713e-05, 4.470186e-06, 
    4.169877e-06, 5.520399e-06, 8.049345e-06, 3.091676e-06, 3.973302e-06,
  0.0001961006, 0.0003030916, 0.0003320946, 0.0003090854, 0.0003079298, 
    0.0002469109, 0.0001405254, 3.163748e-05, 4.524616e-06, 3.476595e-06, 
    7.534961e-06, 8.211965e-06, 8.699147e-06, 8.447309e-06, 3.822349e-06,
  0.0002768636, 0.0003661541, 0.0003868903, 0.0003470375, 0.0002766602, 
    0.0001536038, 4.370548e-05, 1.829479e-05, 7.006046e-06, 7.871099e-06, 
    8.240774e-06, 1.076626e-05, 9.825855e-06, 1.156391e-05, 7.436249e-06,
  0.0003780321, 0.0004009924, 0.0003643328, 0.0002593454, 0.0001379029, 
    3.833601e-05, 8.803046e-06, 5.396583e-06, 6.025335e-06, 5.919848e-06, 
    1.053076e-05, 1.222375e-05, 1.068702e-05, 1.03347e-05, 1.200972e-05,
  0.0004884398, 0.00036646, 0.0002688672, 0.0001333579, 3.299184e-05, 
    1.214662e-05, 9.650611e-06, 5.99375e-06, 4.731275e-06, 4.106474e-06, 
    6.050481e-06, 7.826163e-06, 9.531671e-06, 1.071659e-05, 8.65727e-06,
  0.0005266049, 0.0002694488, 0.0001643882, 4.702356e-05, 8.773792e-06, 
    9.205071e-06, 9.192893e-06, 6.525359e-06, 7.837173e-06, 7.400602e-06, 
    6.34801e-06, 5.557054e-06, 7.592677e-06, 8.247646e-06, 8.08849e-06,
  0.0004689186, 0.0001921652, 8.616867e-05, 1.639371e-05, 6.092866e-06, 
    6.558293e-06, 7.524392e-06, 4.143106e-06, 5.88763e-06, 5.518112e-06, 
    4.295249e-06, 5.348734e-06, 8.700526e-06, 7.27242e-06, 5.824782e-06,
  0.0003412446, 0.0001491821, 4.893474e-05, 7.996468e-06, 4.189783e-06, 
    4.824524e-06, 2.230094e-06, 3.097828e-06, 3.791164e-06, 4.044224e-06, 
    5.254526e-06, 5.908225e-06, 6.005443e-06, 6.651154e-06, 4.805622e-06,
  0.0002629551, 0.0001271596, 2.332291e-05, 4.575466e-06, 2.662653e-06, 
    3.135224e-06, 4.078517e-06, 4.033605e-06, 7.502865e-06, 9.35187e-06, 
    6.524075e-06, 6.435283e-06, 7.946964e-06, 6.558184e-06, 6.260068e-06,
  0.0002253618, 8.61257e-05, 1.552817e-05, 3.017284e-06, 1.28988e-06, 
    3.239503e-06, 4.758821e-06, 6.853201e-06, 9.79534e-06, 1.135477e-05, 
    9.030638e-06, 1.38829e-05, 1.005293e-05, 6.866875e-06, 7.526304e-06,
  4.978263e-05, 5.793299e-05, 5.057565e-05, 4.056957e-05, 3.241839e-05, 
    2.622136e-05, 4.982572e-05, 0.0001010002, 0.0001254734, 0.0001201101, 
    0.0001157657, 7.845498e-05, 2.097996e-05, 4.055201e-05, 2.072727e-05,
  5.852794e-05, 6.309001e-05, 5.58768e-05, 4.771836e-05, 3.749465e-05, 
    8.236188e-05, 0.0001386695, 0.0001958995, 0.0001718053, 0.0001210156, 
    8.313705e-05, 8.619587e-05, 3.896406e-05, 2.859763e-05, 2.483937e-05,
  4.885459e-05, 6.352967e-05, 4.813752e-05, 4.954184e-05, 0.00011864, 
    0.0001658197, 0.0001999338, 0.0001980316, 0.0001674504, 0.0001243438, 
    9.959532e-05, 6.679662e-05, 4.214812e-05, 5.326709e-05, 2.756197e-05,
  5.898836e-05, 6.076858e-05, 4.723397e-05, 0.0001081119, 0.0001987766, 
    0.000256083, 0.0002306821, 0.0002208551, 0.0001649113, 0.0001291338, 
    0.0001041682, 6.424722e-05, 4.994241e-05, 3.31756e-05, 2.535505e-05,
  4.523831e-05, 4.664441e-05, 0.0001217612, 0.0002307018, 0.0002711712, 
    0.0002441483, 0.0002939619, 0.0002270398, 0.0001657852, 0.0001388632, 
    0.0001063651, 7.443963e-05, 5.364861e-05, 4.174003e-05, 3.16625e-05,
  3.658607e-05, 0.0001056771, 0.0002414863, 0.0002816185, 0.0002533937, 
    0.000244915, 0.0002516168, 0.0002026681, 0.000181543, 0.0001521052, 
    0.0001101402, 8.111099e-05, 6.014231e-05, 4.335525e-05, 3.456232e-05,
  0.0001080252, 0.0002191152, 0.0003326388, 0.0002929223, 0.0002592802, 
    0.0002572332, 0.0002294788, 0.0002099941, 0.0001903311, 0.0001627491, 
    0.0001195123, 8.300554e-05, 6.021734e-05, 4.784295e-05, 3.588812e-05,
  0.0002601884, 0.0003409827, 0.0003788182, 0.000282067, 0.0002741577, 
    0.0002596018, 0.0002262966, 0.0002263803, 0.0002268734, 0.0001703502, 
    0.0001113757, 8.773088e-05, 5.863215e-05, 4.188344e-05, 3.13155e-05,
  0.0004067356, 0.0004341132, 0.00038917, 0.0002944366, 0.0002692166, 
    0.0002286292, 0.0002476706, 0.0002655695, 0.0002276323, 0.0001613196, 
    0.0001103254, 7.577897e-05, 5.688343e-05, 3.759778e-05, 2.767887e-05,
  0.0005382871, 0.0004880058, 0.0003605293, 0.0002849569, 0.0002634711, 
    0.0002615176, 0.0002714116, 0.0002614237, 0.0002067585, 0.0001403819, 
    0.0001044667, 7.229325e-05, 4.190851e-05, 3.503437e-05, 1.631824e-05,
  4.832299e-06, 5.506708e-06, 3.550608e-06, 1.850232e-06, 1.254382e-06, 
    1.549153e-06, 1.828548e-06, 2.000508e-06, 3.512361e-06, 4.878311e-06, 
    4.408826e-06, 8.009238e-06, 8.114022e-06, 7.420983e-06, 1.400009e-06,
  7.559684e-06, 5.423049e-06, 3.354306e-06, 2.240286e-06, 1.503284e-06, 
    1.472347e-06, 1.119715e-06, 2.124882e-06, 3.696958e-06, 5.095561e-06, 
    5.972548e-06, 7.779766e-06, 7.976631e-06, 4.342632e-06, 4.595747e-07,
  1.094094e-05, 9.074268e-06, 7.020744e-06, 3.378706e-06, 2.692665e-06, 
    2.641737e-06, 1.519612e-06, 2.202315e-06, 3.670847e-06, 5.144089e-06, 
    5.930538e-06, 5.898267e-06, 6.177859e-06, 3.716538e-06, 6.487142e-07,
  1.922057e-05, 1.050069e-05, 8.874112e-06, 5.915978e-06, 4.454455e-06, 
    3.236252e-06, 2.082795e-06, 1.602989e-06, 2.311529e-06, 3.176637e-06, 
    2.517315e-06, 3.659753e-06, 4.645777e-06, 3.476473e-06, 1.91133e-07,
  2.361804e-05, 1.858829e-05, 1.051514e-05, 8.240146e-06, 4.481069e-06, 
    4.482842e-06, 2.202416e-06, 2.320366e-06, 9.769665e-07, 2.057296e-06, 
    3.702502e-06, 4.241546e-06, 4.827439e-06, 4.586128e-06, 4.40117e-07,
  2.821465e-05, 2.016546e-05, 1.396666e-05, 1.27851e-05, 6.663147e-06, 
    4.702926e-06, 3.235872e-06, 1.605932e-06, 1.271984e-06, 6.959925e-07, 
    1.449609e-06, 4.362939e-06, 4.799089e-06, 4.088548e-06, 4.381462e-07,
  4.433183e-05, 2.675092e-05, 1.737008e-05, 1.149913e-05, 9.09183e-06, 
    6.739293e-06, 4.020415e-06, 3.178335e-06, 1.437366e-06, 3.464511e-07, 
    6.090151e-07, 1.627349e-06, 3.399322e-06, 4.197625e-06, 2.694999e-07,
  5.006395e-05, 3.120757e-05, 2.172333e-05, 1.540415e-05, 1.470274e-05, 
    7.216266e-06, 4.452103e-06, 2.650146e-06, 1.725322e-06, 7.150501e-07, 
    6.835923e-08, 5.667299e-07, 1.433495e-06, 1.577786e-06, 4.962712e-07,
  6.219729e-05, 3.976497e-05, 2.96251e-05, 2.067228e-05, 1.368121e-05, 
    7.894573e-06, 5.311785e-06, 2.808346e-06, 1.932213e-06, 1.056595e-06, 
    6.422509e-07, 1.056248e-07, 7.176735e-07, 4.831713e-07, 1.712075e-06,
  6.767263e-05, 5.624747e-05, 4.085768e-05, 2.975576e-05, 1.555454e-05, 
    1.202211e-05, 6.144917e-06, 3.368137e-06, 1.622438e-06, 9.363092e-07, 
    1.091617e-06, 4.15156e-07, 3.514861e-07, 1.376904e-06, 7.462318e-06,
  1.12527e-06, 2.736688e-06, 6.861357e-06, 3.539709e-06, 6.704088e-06, 
    1.02213e-05, 8.88755e-06, 9.620009e-06, 6.31404e-06, 9.726521e-06, 
    1.483693e-05, 1.029249e-05, 8.559943e-06, 4.412899e-06, 5.119362e-06,
  1.606418e-06, 4.082716e-06, 2.514841e-06, 3.080674e-06, 5.20947e-06, 
    7.532764e-06, 6.047489e-06, 9.22506e-06, 9.349284e-06, 9.57126e-06, 
    8.772784e-06, 1.109169e-05, 1.091434e-05, 4.740314e-06, 4.563523e-06,
  1.249254e-06, 2.437283e-06, 3.474875e-06, 2.278897e-06, 3.611255e-06, 
    7.125169e-06, 6.644048e-06, 1.044681e-05, 9.762037e-06, 1.017622e-05, 
    6.011435e-06, 1.031695e-05, 1.022714e-05, 7.878806e-06, 1.222503e-06,
  1.029544e-06, 1.656143e-06, 2.875224e-06, 1.402685e-06, 3.968003e-06, 
    4.169756e-06, 1.026107e-05, 7.873429e-06, 8.736014e-06, 9.091938e-06, 
    8.492467e-06, 1.10487e-05, 7.951138e-06, 1.444912e-05, 3.938263e-07,
  5.908609e-07, 8.764323e-07, 1.459115e-06, 1.088032e-06, 1.627803e-06, 
    1.949538e-06, 5.480257e-06, 1.335884e-05, 8.800223e-06, 9.93791e-06, 
    1.066262e-05, 8.513659e-06, 8.61273e-06, 9.219603e-06, 2.478438e-06,
  1.209531e-06, 1.766875e-06, 1.243957e-06, 1.040309e-06, 1.233793e-06, 
    9.722424e-07, 3.594744e-06, 9.684029e-06, 1.238971e-05, 1.115322e-05, 
    1.064351e-05, 1.22174e-05, 1.006196e-05, 8.400698e-06, 4.977878e-06,
  1.331774e-06, 2.017229e-06, 1.629334e-06, 2.536793e-06, 2.140311e-06, 
    8.62556e-07, 3.32452e-06, 3.922707e-06, 1.323424e-05, 1.20068e-05, 
    1.135026e-05, 1.313022e-05, 1.221781e-05, 1.338942e-05, 6.05556e-06,
  2.734754e-06, 2.828291e-06, 1.975895e-06, 3.614185e-06, 2.392569e-06, 
    3.494035e-06, 3.934731e-06, 5.972372e-06, 7.857478e-06, 1.164044e-05, 
    1.426189e-05, 1.335542e-05, 1.042697e-05, 1.177158e-05, 9.529385e-06,
  4.603368e-06, 3.812865e-06, 1.708123e-06, 3.771157e-06, 3.268303e-06, 
    5.477962e-06, 4.458561e-06, 4.258489e-06, 7.179773e-06, 1.187188e-05, 
    1.372209e-05, 1.549175e-05, 1.183879e-05, 9.342054e-06, 1.026096e-05,
  3.182624e-06, 4.274292e-06, 5.830482e-06, 4.059521e-06, 3.96379e-06, 
    5.107763e-06, 5.113148e-06, 4.959285e-06, 7.867655e-06, 8.412093e-06, 
    1.330934e-05, 1.590724e-05, 1.573623e-05, 1.028418e-05, 1.163036e-05,
  5.091337e-06, 4.633163e-06, 6.333094e-06, 7.946169e-06, 6.825219e-06, 
    8.411457e-06, 1.033496e-05, 9.800367e-06, 1.162169e-05, 1.31049e-05, 
    1.442258e-05, 1.127004e-05, 7.231034e-06, 5.914118e-06, 2.41681e-06,
  4.613993e-06, 6.217047e-06, 9.17047e-06, 9.241e-06, 6.590471e-06, 
    8.481938e-06, 9.037049e-06, 9.501186e-06, 1.124246e-05, 1.319189e-05, 
    1.372919e-05, 1.303761e-05, 1.052177e-05, 8.808911e-06, 2.120178e-06,
  5.387714e-06, 5.45388e-06, 9.22859e-06, 7.354116e-06, 9.540522e-06, 
    6.625236e-06, 8.249675e-06, 9.563112e-06, 1.051349e-05, 1.149252e-05, 
    1.326904e-05, 1.317994e-05, 1.360129e-05, 9.541449e-06, 4.807746e-06,
  5.768744e-06, 6.078891e-06, 8.793194e-06, 8.438044e-06, 8.537474e-06, 
    7.221451e-06, 7.238262e-06, 9.752566e-06, 8.387081e-06, 1.045082e-05, 
    1.287608e-05, 1.446507e-05, 1.543051e-05, 1.197606e-05, 8.312092e-06,
  5.069018e-06, 7.710294e-06, 8.139681e-06, 8.350948e-06, 4.161281e-06, 
    7.618176e-06, 5.889396e-06, 7.65444e-06, 1.030251e-05, 1.218088e-05, 
    1.151515e-05, 1.26467e-05, 1.49598e-05, 1.354678e-05, 9.772936e-06,
  1.594665e-06, 4.730173e-06, 4.982361e-06, 4.768554e-06, 5.733431e-06, 
    6.404815e-06, 4.015536e-06, 7.102389e-06, 1.257762e-05, 1.047962e-05, 
    9.406745e-06, 1.171568e-05, 1.360913e-05, 1.540005e-05, 1.104782e-05,
  1.708556e-06, 2.287811e-06, 2.842988e-06, 4.281398e-06, 4.018737e-06, 
    3.256607e-06, 6.408956e-06, 7.334715e-06, 1.108506e-05, 9.493889e-06, 
    1.0601e-05, 1.148386e-05, 1.127067e-05, 1.356487e-05, 1.287239e-05,
  1.593295e-06, 9.701005e-07, 3.39041e-06, 5.70553e-06, 3.505976e-06, 
    4.809076e-06, 6.939965e-06, 1.066228e-05, 1.137114e-05, 8.404903e-06, 
    1.035318e-05, 1.206546e-05, 1.239051e-05, 1.304585e-05, 1.395476e-05,
  1.256431e-06, 1.165344e-06, 2.568863e-06, 4.518165e-06, 4.937777e-06, 
    4.023311e-06, 4.174798e-06, 4.148573e-06, 6.414136e-06, 8.335524e-06, 
    7.831822e-06, 8.307511e-06, 1.140793e-05, 1.101256e-05, 1.284371e-05,
  3.41946e-06, 3.179647e-06, 2.716887e-06, 5.724769e-06, 8.214079e-06, 
    3.909905e-06, 5.243242e-06, 4.105958e-06, 3.376553e-06, 4.687633e-06, 
    6.986664e-06, 6.308326e-06, 9.701876e-06, 1.129812e-05, 1.412227e-05,
  2.850223e-06, 4.240215e-06, 4.251544e-06, 5.360039e-06, 6.833114e-06, 
    6.789116e-06, 7.571369e-06, 9.00989e-06, 1.040617e-05, 1.519866e-05, 
    1.856688e-05, 2.00347e-05, 1.519071e-05, 9.068895e-06, 5.610239e-06,
  4.47618e-06, 4.032649e-06, 5.391175e-06, 5.772105e-06, 6.062509e-06, 
    7.549689e-06, 7.986492e-06, 8.104189e-06, 8.579538e-06, 1.239348e-05, 
    1.729561e-05, 2.25628e-05, 1.996332e-05, 1.45913e-05, 8.778645e-06,
  4.307271e-06, 4.043658e-06, 4.653354e-06, 4.470043e-06, 6.77329e-06, 
    9.950388e-06, 1.004076e-05, 8.483094e-06, 9.719263e-06, 1.014525e-05, 
    1.42421e-05, 1.912423e-05, 2.001113e-05, 1.772523e-05, 1.04925e-05,
  5.035601e-06, 3.569042e-06, 2.45597e-06, 3.288749e-06, 6.835633e-06, 
    8.041553e-06, 1.017585e-05, 1.090616e-05, 1.05186e-05, 9.472272e-06, 
    1.102627e-05, 1.505346e-05, 2.168946e-05, 2.007816e-05, 1.544068e-05,
  3.722562e-06, 2.773848e-06, 3.170785e-06, 3.734011e-06, 7.175773e-06, 
    7.935762e-06, 1.024982e-05, 1.002434e-05, 1.094952e-05, 9.853308e-06, 
    9.411218e-06, 1.286997e-05, 1.812615e-05, 2.036511e-05, 1.767507e-05,
  4.037272e-06, 5.834693e-06, 2.725472e-06, 5.429676e-06, 5.378864e-06, 
    7.35396e-06, 8.277221e-06, 9.48773e-06, 1.065695e-05, 1.065267e-05, 
    1.15539e-05, 1.238782e-05, 1.501562e-05, 1.971261e-05, 2.007994e-05,
  3.817801e-06, 5.130134e-06, 6.509381e-06, 5.491637e-06, 4.655291e-06, 
    5.740438e-06, 6.068137e-06, 8.174956e-06, 9.601242e-06, 1.095462e-05, 
    1.132699e-05, 1.040713e-05, 1.368412e-05, 1.753306e-05, 1.905455e-05,
  4.122692e-06, 2.424869e-06, 4.36128e-06, 4.234476e-06, 4.868967e-06, 
    4.91179e-06, 5.595781e-06, 8.558253e-06, 9.226148e-06, 9.519087e-06, 
    1.069737e-05, 1.225051e-05, 1.316251e-05, 1.464429e-05, 1.737186e-05,
  2.272327e-06, 1.385716e-06, 3.40515e-06, 4.346774e-06, 5.326955e-06, 
    5.099152e-06, 6.279796e-06, 9.279072e-06, 9.597737e-06, 9.22082e-06, 
    9.307949e-06, 1.161134e-05, 1.251274e-05, 1.444475e-05, 1.725528e-05,
  2.321178e-06, 8.706181e-07, 3.498715e-06, 4.916132e-06, 6.60736e-06, 
    3.440384e-06, 6.181675e-06, 1.107406e-05, 6.946656e-06, 7.621867e-06, 
    9.148425e-06, 9.515179e-06, 1.085337e-05, 1.263847e-05, 1.533797e-05,
  2.137718e-06, 3.627186e-06, 7.201594e-06, 6.88618e-06, 8.501618e-06, 
    7.464015e-06, 7.57394e-06, 7.551128e-06, 8.63251e-06, 9.31763e-06, 
    1.343945e-05, 1.745263e-05, 1.562797e-05, 1.524921e-05, 1.762245e-05,
  2.269807e-06, 5.049286e-06, 7.509487e-06, 5.766928e-06, 6.937251e-06, 
    6.717454e-06, 8.40247e-06, 8.626665e-06, 8.13203e-06, 9.60194e-06, 
    1.270569e-05, 1.46539e-05, 1.521178e-05, 1.648446e-05, 1.605423e-05,
  2.507697e-06, 3.84634e-06, 5.786589e-06, 6.358918e-06, 6.789431e-06, 
    7.188829e-06, 8.971667e-06, 9.133402e-06, 1.212119e-05, 1.145561e-05, 
    1.198652e-05, 1.237148e-05, 1.599061e-05, 1.69596e-05, 1.695713e-05,
  2.792379e-06, 4.419718e-06, 5.545212e-06, 5.436694e-06, 6.252948e-06, 
    8.749607e-06, 9.366036e-06, 9.540385e-06, 1.151126e-05, 1.17468e-05, 
    1.148587e-05, 1.396415e-05, 1.526021e-05, 1.788957e-05, 2.03503e-05,
  2.364246e-06, 4.557518e-06, 4.00078e-06, 5.031836e-06, 5.916685e-06, 
    6.943788e-06, 8.24688e-06, 9.66107e-06, 1.059824e-05, 1.197204e-05, 
    1.188518e-05, 1.300044e-05, 1.543548e-05, 1.884997e-05, 2.055749e-05,
  2.870595e-06, 4.601384e-06, 4.787616e-06, 6.69361e-06, 5.238648e-06, 
    5.704065e-06, 8.291266e-06, 9.624513e-06, 1.071801e-05, 1.123034e-05, 
    1.139487e-05, 1.320459e-05, 1.582988e-05, 1.72463e-05, 2.196731e-05,
  1.887358e-06, 5.154116e-06, 4.864802e-06, 5.877657e-06, 5.129519e-06, 
    6.666609e-06, 7.167705e-06, 8.526824e-06, 8.344033e-06, 9.955436e-06, 
    1.218901e-05, 1.252258e-05, 1.443497e-05, 1.709665e-05, 2.145603e-05,
  3.081341e-06, 4.386242e-06, 5.592238e-06, 7.301347e-06, 5.604019e-06, 
    7.083243e-06, 7.827965e-06, 9.215393e-06, 8.284722e-06, 9.131761e-06, 
    9.844871e-06, 1.217138e-05, 1.252995e-05, 1.711497e-05, 1.957826e-05,
  1.850671e-06, 3.374073e-06, 5.382274e-06, 6.007338e-06, 7.335226e-06, 
    7.80533e-06, 7.641334e-06, 9.767271e-06, 9.408122e-06, 1.042397e-05, 
    9.431629e-06, 9.82346e-06, 1.275631e-05, 1.214234e-05, 1.892631e-05,
  1.72596e-06, 4.575058e-07, 4.019092e-06, 6.494033e-06, 6.268526e-06, 
    6.791076e-06, 7.7054e-06, 1.122245e-05, 1.046231e-05, 1.008293e-05, 
    9.995464e-06, 9.367258e-06, 1.0937e-05, 1.281297e-05, 1.566289e-05,
  3.660766e-06, 4.836072e-06, 9.759614e-06, 8.793343e-06, 8.446419e-06, 
    9.294424e-06, 9.612792e-06, 7.308841e-06, 7.209871e-06, 7.357787e-06, 
    1.065412e-05, 1.466294e-05, 1.616267e-05, 1.738976e-05, 1.600381e-05,
  3.530879e-06, 5.575889e-06, 8.090263e-06, 6.852445e-06, 8.657515e-06, 
    7.890008e-06, 8.784598e-06, 8.537364e-06, 8.046432e-06, 6.864097e-06, 
    9.237982e-06, 1.125798e-05, 1.456985e-05, 1.777899e-05, 2.014312e-05,
  4.143609e-06, 4.585496e-06, 6.688891e-06, 5.976999e-06, 7.923674e-06, 
    7.628583e-06, 8.747296e-06, 8.663907e-06, 8.807624e-06, 8.655524e-06, 
    7.718457e-06, 9.011348e-06, 1.369982e-05, 1.649293e-05, 2.046815e-05,
  5.039775e-06, 3.864044e-06, 5.536084e-06, 5.900529e-06, 7.669183e-06, 
    7.296704e-06, 8.453309e-06, 9.466165e-06, 8.928301e-06, 9.589034e-06, 
    1.013961e-05, 8.743678e-06, 1.14614e-05, 1.555374e-05, 1.877981e-05,
  5.668503e-06, 4.461715e-06, 4.706661e-06, 6.801331e-06, 7.61237e-06, 
    8.828556e-06, 8.196528e-06, 8.831867e-06, 1.000507e-05, 1.293285e-05, 
    1.032192e-05, 9.696796e-06, 9.233423e-06, 1.235493e-05, 1.751672e-05,
  4.983542e-06, 5.096502e-06, 4.774061e-06, 6.97556e-06, 8.093875e-06, 
    8.783474e-06, 8.390423e-06, 9.532701e-06, 1.066039e-05, 1.238697e-05, 
    1.154353e-05, 1.158599e-05, 9.673295e-06, 1.358925e-05, 1.639072e-05,
  4.860999e-06, 5.208103e-06, 7.302763e-06, 6.701595e-06, 7.397126e-06, 
    9.283676e-06, 1.107961e-05, 1.153477e-05, 1.145557e-05, 1.217496e-05, 
    1.307236e-05, 1.073886e-05, 1.01833e-05, 1.162151e-05, 1.615633e-05,
  4.346884e-06, 6.096207e-06, 7.679537e-06, 6.867152e-06, 6.456878e-06, 
    7.729749e-06, 1.097904e-05, 1.285081e-05, 1.156472e-05, 1.195914e-05, 
    1.332211e-05, 1.210828e-05, 1.189413e-05, 1.1346e-05, 1.401343e-05,
  8.638397e-06, 9.060572e-06, 5.807189e-06, 7.289521e-06, 9.224957e-06, 
    8.126162e-06, 1.056382e-05, 1.293708e-05, 1.280216e-05, 1.222978e-05, 
    1.531891e-05, 1.512128e-05, 1.24076e-05, 1.16363e-05, 1.498586e-05,
  7.995787e-06, 4.027126e-06, 6.671825e-06, 7.449436e-06, 8.138898e-06, 
    8.801247e-06, 9.218644e-06, 1.044539e-05, 1.264111e-05, 1.395081e-05, 
    1.369558e-05, 1.285227e-05, 1.477697e-05, 1.256506e-05, 1.347791e-05,
  9.215971e-06, 9.643222e-06, 1.861545e-05, 1.605282e-05, 2.035088e-05, 
    2.05714e-05, 2.32943e-05, 4.786989e-05, 8.743708e-05, 0.0001837415, 
    0.0002440446, 0.0002848, 0.0003231655, 0.0003421951, 0.0003574862,
  9.120804e-06, 1.091427e-05, 1.454756e-05, 1.421486e-05, 1.882678e-05, 
    1.618734e-05, 1.771924e-05, 2.008776e-05, 2.752435e-05, 5.140209e-05, 
    9.963936e-05, 0.0001482536, 0.0002094565, 0.0002112946, 0.0001871467,
  8.418856e-06, 8.824506e-06, 1.090442e-05, 1.392389e-05, 1.721617e-05, 
    1.899669e-05, 2.014425e-05, 1.797543e-05, 1.676365e-05, 2.208294e-05, 
    3.451417e-05, 5.002166e-05, 7.384459e-05, 0.0001035322, 8.141304e-05,
  1.114697e-05, 9.071358e-06, 8.694421e-06, 1.201951e-05, 1.32465e-05, 
    1.89994e-05, 1.962801e-05, 1.994426e-05, 1.790117e-05, 1.726678e-05, 
    1.906113e-05, 2.140629e-05, 2.844458e-05, 2.891632e-05, 3.00616e-05,
  1.399627e-05, 9.744048e-06, 1.108051e-05, 1.02969e-05, 9.810068e-06, 
    1.221532e-05, 2.120803e-05, 2.538643e-05, 2.642693e-05, 1.730887e-05, 
    1.574526e-05, 1.794209e-05, 1.733341e-05, 2.229152e-05, 2.429285e-05,
  1.593023e-05, 1.412263e-05, 1.465752e-05, 1.185204e-05, 9.830912e-06, 
    1.086546e-05, 1.465537e-05, 2.055359e-05, 2.149692e-05, 2.11254e-05, 
    1.82424e-05, 1.696837e-05, 1.632428e-05, 1.399938e-05, 1.744028e-05,
  1.391706e-05, 1.74949e-05, 1.709738e-05, 1.585231e-05, 1.377989e-05, 
    1.089806e-05, 1.095343e-05, 1.273081e-05, 1.834457e-05, 2.567403e-05, 
    2.206869e-05, 1.666019e-05, 1.442596e-05, 1.500031e-05, 1.414303e-05,
  1.345437e-05, 1.929383e-05, 1.749797e-05, 1.617351e-05, 1.495069e-05, 
    1.251858e-05, 1.094522e-05, 8.828397e-06, 1.215015e-05, 1.873748e-05, 
    2.048395e-05, 2.033384e-05, 1.644058e-05, 1.563672e-05, 1.54884e-05,
  1.303795e-05, 1.39703e-05, 1.687288e-05, 1.452797e-05, 1.559302e-05, 
    1.480545e-05, 1.399165e-05, 9.102174e-06, 7.027495e-06, 1.211996e-05, 
    1.664002e-05, 1.916748e-05, 1.718209e-05, 1.632204e-05, 1.621491e-05,
  1.40884e-05, 1.288867e-05, 1.376662e-05, 1.486776e-05, 1.714265e-05, 
    1.622062e-05, 1.490584e-05, 1.075164e-05, 8.279685e-06, 6.779946e-06, 
    1.051502e-05, 1.529959e-05, 1.662699e-05, 1.822797e-05, 1.728501e-05,
  0.0002286083, 0.00031248, 0.0002955293, 0.0003157223, 0.0003314877, 
    0.0003479241, 0.0003267572, 0.0003649189, 0.0002952267, 0.0002356783, 
    0.0001606725, 0.000136394, 0.000128883, 0.0001232585, 0.0001367978,
  0.0002218199, 0.0002835973, 0.0002932392, 0.0002932399, 0.0002910713, 
    0.0002940784, 0.0002851311, 0.0002749746, 0.0002735283, 0.0003006186, 
    0.0002924571, 0.0002987692, 0.0002695334, 0.0002444475, 0.0003401113,
  0.0002365474, 0.0003093196, 0.0003241688, 0.0002806162, 0.0002838406, 
    0.0002690434, 0.0002736507, 0.0002538778, 0.0002451825, 0.0002882364, 
    0.0003570367, 0.0003995092, 0.0004354947, 0.0004318234, 0.0005234266,
  0.0001941919, 0.0002598878, 0.0003171297, 0.000294192, 0.0002626778, 
    0.0002473881, 0.0002531706, 0.0002458599, 0.0002577964, 0.0002879637, 
    0.0003925323, 0.0004633621, 0.0005329982, 0.0005771384, 0.0005975975,
  0.000103201, 0.0001852779, 0.0002418823, 0.0002618889, 0.0002606891, 
    0.0002199719, 0.0002004409, 0.0002197698, 0.0002484887, 0.0003114434, 
    0.000406792, 0.0004577937, 0.0006637796, 0.0005798627, 0.0006065883,
  3.828252e-05, 8.827165e-05, 0.0001430326, 0.0001789364, 0.0002050008, 
    0.0001980863, 0.0001812155, 0.0001765443, 0.0002332915, 0.0002410235, 
    0.0004531586, 0.0005126416, 0.0006462337, 0.0006233741, 0.0005030942,
  1.107725e-05, 2.587899e-05, 5.744473e-05, 8.322445e-05, 0.0001149525, 
    0.0001369885, 0.0001709176, 0.0001856954, 0.0002224044, 0.0002677385, 
    0.0003905832, 0.0005548181, 0.0005502063, 0.0005737125, 0.000502634,
  3.729123e-06, 8.497205e-06, 2.288586e-05, 3.334753e-05, 4.874858e-05, 
    7.417094e-05, 0.0001251185, 0.0001663269, 0.0002043066, 0.0002339757, 
    0.0003485102, 0.0004539674, 0.0005135523, 0.0005001266, 0.000467208,
  4.206397e-06, 4.144131e-06, 7.629539e-06, 1.96062e-05, 2.44295e-05, 
    3.428765e-05, 5.533216e-05, 0.0001006586, 0.0001628953, 0.0002453535, 
    0.0003547698, 0.0004124734, 0.0004890424, 0.0004708774, 0.0005042201,
  6.914957e-06, 5.755498e-06, 6.068849e-06, 6.83059e-06, 1.420682e-05, 
    1.958729e-05, 2.643506e-05, 4.961556e-05, 0.000128395, 0.000222548, 
    0.0003364791, 0.0004240647, 0.0004323424, 0.0004296442, 0.0004412858,
  9.083901e-05, 0.0001460161, 0.0002288299, 0.0001868375, 0.0001665177, 
    0.0001225898, 0.0001435225, 0.0001595954, 0.0001424868, 0.0001699898, 
    0.0001917517, 0.0001902015, 0.0001471453, 0.0001779164, 7.852636e-05,
  3.815741e-05, 0.0001347399, 0.0001399135, 0.0001597743, 0.0001798891, 
    0.000189617, 9.453482e-05, 0.0001023918, 0.0001043801, 0.0001849732, 
    0.0001304611, 0.0001362162, 0.0001148756, 0.0001259905, 7.672387e-05,
  3.789566e-05, 4.242315e-05, 0.0001359007, 0.0001237748, 0.0001129955, 
    0.000129837, 0.0001823932, 0.0001327982, 8.133631e-05, 0.0001058899, 
    0.0001227924, 0.0001273284, 0.0001181925, 0.0001025185, 4.468171e-05,
  5.165399e-05, 5.254542e-05, 4.000814e-05, 0.0001194096, 9.740844e-05, 
    0.0001144035, 0.000108163, 0.0001110596, 0.0001183267, 7.649083e-05, 
    0.0001115432, 9.490539e-05, 0.0001177832, 0.0001087036, 4.319169e-05,
  0.0001563767, 7.129631e-05, 3.618955e-05, 3.883778e-05, 6.253341e-05, 
    9.180733e-05, 0.0001306254, 0.0001045651, 0.0001016084, 0.000102315, 
    7.583224e-05, 0.0001098469, 0.0001195933, 0.0001148583, 9.604358e-05,
  0.0002256896, 0.0001876071, 0.0001359932, 5.886286e-05, 4.306852e-05, 
    4.505147e-05, 9.111575e-05, 9.23559e-05, 0.0001042369, 7.081936e-05, 
    8.813539e-05, 0.0001278678, 0.0001064051, 9.131434e-05, 7.952305e-05,
  0.000262918, 0.0002494996, 0.0002164443, 0.0001652993, 8.214554e-05, 
    5.586646e-05, 3.656305e-05, 7.160915e-05, 7.243253e-05, 4.195435e-05, 
    4.904266e-05, 4.207439e-05, 3.992099e-05, 2.745472e-05, 1.396245e-05,
  0.0002654508, 0.0002702343, 0.0002300779, 0.0001885627, 0.0001549733, 
    8.729192e-05, 5.097192e-05, 1.267622e-05, 1.395518e-05, 2.189664e-05, 
    2.493117e-05, 1.517454e-05, 1.40676e-05, 9.113738e-06, 1.127002e-05,
  0.0002530309, 0.0002551192, 0.0002240386, 0.0001616765, 0.0001419825, 
    0.0001138806, 7.766187e-05, 5.758093e-05, 2.366082e-05, 2.922167e-06, 
    2.258065e-06, 2.641933e-06, 3.687561e-06, 5.932975e-06, 1.066521e-05,
  0.0002385724, 0.0002376121, 0.0002192544, 0.0001731948, 0.0001391647, 
    0.0001120585, 9.760615e-05, 9.942328e-05, 7.771848e-05, 4.304269e-05, 
    5.546321e-06, 3.234296e-06, 6.839159e-06, 1.786281e-05, 3.475909e-05,
  9.56441e-05, 0.0001347844, 8.243595e-05, 5.074771e-05, 4.305038e-05, 
    5.923555e-05, 6.743694e-05, 6.613816e-05, 4.098372e-05, 2.654202e-05, 
    1.254424e-05, 2.913595e-05, 1.705142e-05, 1.716459e-05, 2.30647e-05,
  7.193883e-05, 6.755989e-05, 7.846589e-05, 5.52678e-05, 6.493685e-05, 
    4.854328e-05, 5.345869e-05, 5.992059e-05, 5.527556e-05, 3.732795e-05, 
    2.087966e-05, 1.162155e-05, 1.026675e-05, 1.672279e-05, 3.254218e-05,
  3.898134e-05, 3.1254e-05, 6.367965e-05, 7.722015e-05, 5.971575e-05, 
    5.181198e-05, 5.233792e-05, 4.405319e-05, 5.012227e-05, 3.402801e-05, 
    2.181577e-05, 2.353743e-05, 2.048877e-05, 1.485223e-05, 3.972416e-05,
  1.941337e-05, 2.389024e-05, 4.349222e-05, 6.016149e-05, 5.885509e-05, 
    6.39534e-05, 4.61333e-05, 4.516886e-05, 4.100857e-05, 3.5424e-05, 
    1.962406e-05, 2.667167e-05, 1.457796e-05, 2.094817e-05, 2.515183e-05,
  3.132482e-05, 2.159395e-05, 1.817019e-05, 3.791076e-05, 5.46708e-05, 
    5.720088e-05, 5.276874e-05, 6.067509e-05, 6.121067e-05, 3.284321e-05, 
    1.732697e-05, 2.024042e-05, 1.999571e-05, 3.339825e-05, 8.781085e-05,
  1.714402e-05, 1.610428e-05, 1.695809e-05, 5.064829e-05, 4.048505e-05, 
    2.947157e-05, 5.722619e-05, 7.975064e-05, 9.156871e-05, 6.842912e-05, 
    4.621713e-05, 4.544496e-05, 8.547996e-05, 8.92129e-05, 0.0001085494,
  1.857758e-05, 1.594745e-05, 7.021819e-06, 2.274754e-05, 3.342989e-05, 
    5.886506e-05, 5.11521e-05, 6.573628e-05, 0.000144917, 0.0001223298, 
    9.619659e-05, 0.0001306428, 0.0001274197, 0.0001000602, 8.683975e-05,
  8.483713e-06, 1.638913e-05, 2.459975e-05, 1.275522e-05, 9.195345e-06, 
    8.05529e-05, 8.11445e-05, 0.0001360676, 0.0001605981, 8.607106e-05, 
    8.862063e-05, 7.658617e-05, 9.545284e-05, 8.813846e-05, 8.549706e-05,
  2.893699e-06, 9.648982e-06, 2.349112e-05, 2.166875e-05, 7.522517e-05, 
    5.951952e-05, 0.0001047312, 0.0001029328, 0.0001804594, 0.0001319723, 
    3.906948e-05, 3.768906e-05, 6.609273e-05, 5.42436e-05, 5.846133e-05,
  3.783362e-06, 6.972684e-06, 6.225953e-06, 1.458638e-06, 9.486059e-06, 
    2.841805e-05, 9.755366e-05, 7.483282e-05, 9.456915e-05, 0.0001140025, 
    5.414697e-05, 4.271508e-05, 3.851064e-05, 4.136429e-05, 6.582613e-05,
  2.536753e-05, 2.914542e-05, 6.739173e-05, 7.41954e-05, 8.980886e-05, 
    8.855135e-05, 7.333204e-05, 2.73668e-05, 1.519548e-05, 1.491622e-05, 
    1.368997e-05, 1.033537e-05, 9.2142e-06, 1.120243e-05, 1.034873e-05,
  1.817272e-05, 1.96048e-05, 3.380707e-05, 3.515555e-05, 3.977259e-05, 
    6.732322e-05, 4.498075e-05, 5.569166e-05, 2.990056e-05, 1.519999e-05, 
    1.061745e-05, 9.647542e-06, 8.076691e-06, 7.630815e-06, 8.718686e-06,
  1.628736e-05, 2.394748e-05, 1.992443e-05, 2.779495e-05, 2.821639e-05, 
    3.674056e-05, 2.515517e-05, 5.692061e-05, 5.70928e-05, 3.30639e-05, 
    1.407718e-05, 6.682962e-06, 1.970862e-05, 6.541416e-06, 7.514986e-06,
  2.135223e-05, 2.222939e-05, 1.802254e-05, 2.223314e-05, 2.213091e-05, 
    1.637753e-05, 1.310574e-05, 3.023402e-05, 0.0001034988, 9.537652e-05, 
    3.075621e-05, 1.0169e-05, 5.299724e-06, 6.49634e-06, 5.821897e-06,
  2.462976e-05, 1.887309e-05, 2.229594e-05, 2.078154e-05, 2.012384e-05, 
    1.817657e-05, 1.47399e-05, 1.68696e-05, 6.22712e-05, 6.427284e-05, 
    6.52753e-05, 1.824639e-05, 5.946757e-06, 3.969037e-06, 3.296469e-06,
  2.70752e-05, 1.829636e-05, 2.389677e-05, 2.412472e-05, 2.353773e-05, 
    2.642997e-05, 1.644114e-05, 1.569765e-05, 3.018185e-05, 6.240269e-05, 
    0.0001649857, 3.893885e-05, 1.129309e-05, 4.971598e-06, 3.728014e-06,
  4.452128e-05, 3.412697e-05, 3.598558e-05, 2.441819e-05, 2.031272e-05, 
    2.686521e-05, 2.181293e-05, 2.766639e-05, 2.048227e-05, 8.036503e-05, 
    0.0001558944, 0.0001247318, 2.914087e-05, 8.044286e-06, 6.519998e-06,
  3.828368e-05, 3.914563e-05, 4.035398e-05, 3.861103e-05, 3.042734e-05, 
    3.557157e-05, 3.120207e-05, 3.789515e-05, 2.532526e-05, 7.770486e-05, 
    0.0001365054, 0.0001508129, 3.89078e-05, 1.3549e-05, 6.345803e-06,
  3.571738e-05, 3.475324e-05, 3.226726e-05, 3.541974e-05, 4.164899e-05, 
    2.849613e-05, 2.359033e-05, 2.403517e-05, 3.363149e-05, 6.834399e-05, 
    0.0001236806, 0.0001145667, 7.137264e-05, 2.906372e-05, 1.674243e-05,
  3.003626e-05, 3.293823e-05, 3.335036e-05, 6.322615e-05, 5.525895e-05, 
    6.066287e-05, 4.857002e-05, 3.01348e-05, 5.757523e-05, 7.300126e-05, 
    0.0001516406, 0.0001190558, 8.454379e-05, 3.101919e-05, 1.511934e-05,
  0.000300183, 0.0001867896, 0.0001123427, 0.0001884899, 0.00026987, 
    0.0001885167, 0.0001798407, 8.076058e-05, 7.596547e-05, 6.351497e-05, 
    3.548398e-05, 2.107905e-05, 1.447577e-05, 9.946749e-06, 5.190641e-06,
  0.0002942368, 0.0002505953, 0.000160997, 0.0002469709, 0.0002935653, 
    0.0003447738, 0.0002511231, 0.0001330296, 0.000121673, 9.493137e-05, 
    6.014032e-05, 3.198453e-05, 1.702333e-05, 9.502893e-06, 4.970962e-06,
  0.0001919098, 0.0002594985, 0.0002520287, 0.0002198645, 0.00028292, 
    0.0004203696, 0.0002383707, 0.0001692115, 0.0001066872, 7.391139e-05, 
    5.136639e-05, 4.603581e-05, 2.464562e-05, 1.347062e-05, 8.928007e-06,
  0.0001397707, 0.0002496416, 0.0002813951, 0.0002498124, 0.0002692875, 
    0.0003677709, 0.0004286672, 0.0002331013, 8.447422e-05, 0.0001174257, 
    0.0001018664, 5.569063e-05, 3.84899e-05, 1.975903e-05, 1.266993e-05,
  0.0001784552, 0.0002464842, 0.0002762098, 0.0002719545, 0.0002655842, 
    0.0002563117, 0.0003529934, 0.0003113103, 0.0001806951, 9.186447e-05, 
    8.323301e-05, 6.741212e-05, 5.190289e-05, 3.14173e-05, 1.710028e-05,
  0.0002170212, 0.0002732646, 0.0003251505, 0.000259777, 0.0002574587, 
    0.0002411142, 0.0003195496, 0.0002871064, 0.0002179422, 0.0001397766, 
    8.479953e-05, 7.011064e-05, 6.320776e-05, 4.630649e-05, 2.101085e-05,
  0.000194338, 0.0002704065, 0.0002325278, 0.0002454781, 0.0002303803, 
    0.0002209772, 0.0002503772, 0.0002944321, 0.0001467472, 0.0001668414, 
    0.0001017955, 5.695964e-05, 5.031359e-05, 4.651565e-05, 2.766557e-05,
  0.0002018744, 0.000176825, 0.0002010421, 0.0002314607, 0.0002242288, 
    0.0002120018, 0.000237072, 0.0002530549, 0.0002193624, 0.0001717986, 
    8.977072e-05, 9.999777e-05, 6.218679e-05, 5.278602e-05, 4.024168e-05,
  0.0001362785, 0.0001703793, 0.0002039183, 0.0002026063, 0.0002130885, 
    0.0002222305, 0.0002134705, 0.0002119426, 0.0002121603, 0.0001145601, 
    0.0001466134, 6.416316e-05, 5.151602e-05, 3.273715e-05, 6.189648e-05,
  0.0001125854, 0.0001586903, 0.0001752021, 0.0001859881, 0.0002026732, 
    0.0001925661, 0.0001993896, 0.0002127609, 0.0002573156, 0.0001634781, 
    0.0001349733, 4.268549e-05, 5.131748e-05, 3.857606e-05, 4.628939e-05,
  3.115412e-05, 4.31642e-05, 3.924185e-05, 3.04098e-05, 1.015473e-05, 
    9.504767e-06, 1.777868e-05, 1.649149e-05, 1.384175e-05, 1.007821e-05, 
    8.33715e-06, 3.016386e-06, 1.177278e-06, 4.130818e-07, 1.422603e-07,
  4.632782e-05, 5.446652e-05, 6.560206e-05, 3.766074e-05, 2.724181e-05, 
    1.025335e-05, 1.184451e-05, 1.341639e-05, 1.208924e-05, 1.004714e-05, 
    7.491855e-06, 3.430225e-06, 1.559536e-06, 4.459011e-07, 2.350078e-07,
  5.114462e-05, 6.209606e-05, 8.843934e-05, 6.749056e-05, 4.719921e-05, 
    2.70095e-05, 1.444552e-05, 1.64536e-05, 1.581273e-05, 1.376933e-05, 
    8.613488e-06, 7.940123e-06, 3.862486e-06, 2.586394e-06, 1.567336e-07,
  5.405054e-05, 7.769786e-05, 7.821251e-05, 9.068751e-05, 5.467099e-05, 
    4.606151e-05, 2.471106e-05, 1.998126e-05, 1.672499e-05, 1.483372e-05, 
    1.290632e-05, 8.788281e-06, 7.319231e-06, 2.958409e-06, 3.026775e-06,
  4.429093e-05, 6.976114e-05, 0.0001006691, 9.684654e-05, 9.066224e-05, 
    6.017926e-05, 4.236144e-05, 2.702788e-05, 2.050334e-05, 1.434158e-05, 
    1.421105e-05, 1.145818e-05, 8.728993e-06, 5.196092e-06, 2.576881e-06,
  6.128845e-05, 7.433997e-05, 7.935733e-05, 9.862768e-05, 0.0001332745, 
    7.748965e-05, 5.931271e-05, 3.673641e-05, 2.645876e-05, 1.846958e-05, 
    1.487937e-05, 1.351114e-05, 1.107311e-05, 8.163256e-06, 4.531194e-06,
  5.653868e-05, 7.538418e-05, 8.270717e-05, 9.068405e-05, 0.0001193297, 
    8.853051e-05, 7.969957e-05, 5.25234e-05, 4.411352e-05, 2.578146e-05, 
    1.680106e-05, 1.377532e-05, 1.429338e-05, 1.010346e-05, 6.693359e-06,
  3.958611e-05, 5.43797e-05, 8.465769e-05, 9.821677e-05, 0.0001173481, 
    0.0001190252, 9.474839e-05, 6.029168e-05, 5.902186e-05, 3.32001e-05, 
    2.252885e-05, 1.899375e-05, 1.586305e-05, 1.346565e-05, 7.817011e-06,
  4.788934e-05, 4.183911e-05, 0.0001036353, 0.0001296067, 0.0001035799, 
    0.0001053262, 8.519302e-05, 6.715898e-05, 7.372628e-05, 5.208482e-05, 
    2.760412e-05, 1.978371e-05, 1.630383e-05, 1.48918e-05, 6.801156e-06,
  6.486342e-05, 5.753946e-05, 8.710969e-05, 0.0001140614, 0.0001043393, 
    9.815339e-05, 0.0001293135, 6.277795e-05, 8.840644e-05, 7.670793e-05, 
    3.553626e-05, 2.486413e-05, 1.9916e-05, 1.258352e-05, 8.765614e-06,
  5.841607e-05, 3.430436e-05, 6.982792e-05, 0.0001054091, 8.457274e-05, 
    2.809352e-05, 1.904331e-06, 2.308894e-06, 2.020346e-06, 2.616911e-06, 
    3.047065e-06, 2.354835e-06, 2.151701e-06, 1.836546e-06, 8.331713e-07,
  6.663952e-05, 3.362348e-05, 5.994827e-05, 0.0001109209, 8.580855e-05, 
    2.302471e-05, 1.414539e-06, 1.802935e-06, 3.313125e-06, 2.626986e-06, 
    3.505004e-06, 2.95097e-06, 1.976839e-06, 2.355413e-06, 1.486421e-06,
  7.819248e-05, 4.065371e-05, 6.44871e-05, 0.000105011, 6.744518e-05, 
    9.459254e-06, 1.752196e-06, 2.346815e-06, 2.627595e-06, 3.335699e-06, 
    3.563664e-06, 4.161408e-06, 4.469487e-06, 5.557603e-06, 2.419708e-06,
  9.627073e-05, 5.719387e-05, 7.211505e-05, 8.859563e-05, 4.193175e-05, 
    2.399885e-06, 2.088714e-06, 2.322352e-06, 2.778907e-06, 2.764286e-06, 
    3.38787e-06, 3.251251e-06, 3.256967e-06, 4.037247e-06, 2.10664e-06,
  0.0001499364, 8.168282e-05, 6.098414e-05, 5.33908e-05, 1.501856e-05, 
    8.157631e-07, 1.553993e-06, 1.995878e-06, 2.147969e-06, 2.103769e-06, 
    3.249923e-06, 2.341684e-06, 3.389661e-06, 2.903085e-06, 3.186583e-06,
  0.0002327226, 0.0001226903, 4.81657e-05, 2.823904e-05, 6.754208e-06, 
    1.520122e-06, 1.014056e-06, 1.621856e-06, 1.922241e-06, 2.289137e-06, 
    2.594928e-06, 3.019699e-06, 2.830694e-06, 1.999928e-06, 2.010886e-06,
  0.0002661218, 0.0001619117, 3.64704e-05, 1.499309e-05, 4.977534e-06, 
    2.117393e-06, 1.480969e-06, 7.970214e-07, 1.35915e-06, 2.010082e-06, 
    2.952421e-06, 2.760263e-06, 2.461252e-06, 1.942394e-06, 2.564713e-06,
  0.0002623609, 0.0001873475, 6.193347e-05, 1.044759e-05, 4.830605e-06, 
    5.185342e-06, 2.060425e-06, 1.285516e-06, 1.163664e-06, 1.422847e-06, 
    1.630891e-06, 2.050335e-06, 3.065856e-06, 2.530938e-06, 2.693827e-06,
  0.0002216522, 0.0001967766, 9.395862e-05, 7.716308e-06, 6.230945e-06, 
    5.800091e-06, 4.237943e-06, 2.299832e-06, 1.500189e-06, 1.300228e-06, 
    1.257856e-06, 1.402255e-06, 2.35712e-06, 2.660445e-06, 2.114403e-06,
  0.0001804714, 0.0001958717, 0.0001147225, 9.992828e-06, 6.332857e-06, 
    6.696792e-06, 4.350257e-06, 4.308316e-06, 2.834945e-06, 1.209539e-06, 
    1.140891e-06, 1.374478e-06, 1.479958e-06, 2.562655e-06, 2.800392e-06,
  3.893749e-06, 2.009372e-06, 9.944293e-07, 1.633499e-06, 1.685281e-05, 
    5.405984e-05, 6.465695e-05, 8.912947e-05, 3.029725e-05, 1.902689e-07, 
    1.977674e-08, 3.202215e-05, 2.080922e-05, 1.185685e-05, 1.24852e-05,
  3.581463e-06, 1.502109e-06, 1.458019e-06, 5.162729e-06, 2.917529e-05, 
    6.555669e-05, 6.895271e-05, 5.955317e-05, 4.950873e-05, 5.330959e-07, 
    1.881531e-07, 1.441936e-05, 4.1991e-05, 1.190375e-05, 1.571307e-05,
  4.975005e-06, 3.245745e-06, 4.101822e-06, 2.091246e-05, 5.536301e-05, 
    8.803535e-05, 8.388808e-05, 8.327948e-05, 7.931698e-05, 9.172802e-06, 
    3.616525e-07, 2.044915e-05, 4.276932e-05, 1.179578e-05, 1.043038e-05,
  7.851732e-06, 6.567512e-06, 2.172602e-05, 6.357814e-05, 9.816636e-05, 
    0.0001052417, 0.0001010372, 8.599564e-05, 9.36949e-05, 2.375585e-05, 
    1.935963e-07, 5.581693e-07, 2.559879e-05, 9.255102e-06, 4.012464e-06,
  7.131559e-06, 1.807857e-05, 6.154744e-05, 0.0001294242, 0.0001387789, 
    0.0001210294, 0.0001074595, 8.962434e-05, 8.919456e-05, 4.119725e-05, 
    2.590986e-07, 9.672322e-07, 7.69147e-06, 6.945951e-06, 2.46801e-06,
  5.361368e-06, 3.302679e-05, 0.0001057976, 0.0001823433, 0.0001786351, 
    0.0001350677, 0.0001206644, 9.499984e-05, 7.125303e-05, 5.512236e-05, 
    1.73443e-06, 5.072167e-07, 5.119905e-07, 1.425468e-06, 1.768742e-06,
  8.627771e-06, 4.558032e-05, 0.0001305246, 0.0002136832, 0.000186593, 
    0.0001590059, 0.0001441151, 0.0001036032, 6.464281e-05, 5.873459e-05, 
    7.085773e-06, 3.386358e-07, 4.106403e-07, 1.643367e-06, 2.578798e-06,
  1.133837e-05, 6.314e-05, 0.0001642941, 0.0002368557, 0.000207597, 
    0.000170343, 0.0001656619, 0.0001147604, 6.820475e-05, 5.543193e-05, 
    1.279147e-05, 3.836101e-07, 6.412033e-07, 1.212805e-06, 1.966073e-06,
  1.551334e-05, 7.803155e-05, 0.0001923326, 0.0002495762, 0.0002205184, 
    0.0001881925, 0.0001838376, 0.0001283803, 7.698491e-05, 5.864674e-05, 
    2.383472e-05, 9.77334e-07, 6.024275e-07, 1.770536e-06, 1.103998e-06,
  2.921246e-05, 9.348673e-05, 0.0001993767, 0.0002724309, 0.0002296847, 
    0.0001942726, 0.00019328, 0.0001522433, 9.105545e-05, 6.572992e-05, 
    3.594674e-05, 4.981741e-06, 1.404293e-06, 1.122004e-06, 1.038552e-06,
  0.0001015506, 5.75559e-05, 5.68773e-05, 9.188877e-05, 9.678226e-05, 
    5.937919e-05, 2.721154e-05, 1.046281e-05, 3.713836e-06, 5.158784e-07, 
    4.856892e-06, 3.0002e-06, 4.786185e-06, 6.833855e-06, 1.110383e-05,
  8.346646e-05, 7.811367e-05, 8.19975e-05, 0.000137128, 0.0001399197, 
    6.51371e-05, 1.915198e-05, 1.896863e-05, 3.694978e-06, 8.091026e-07, 
    5.630816e-06, 5.766244e-06, 6.501245e-06, 9.767258e-06, 1.339627e-05,
  6.831848e-05, 9.182291e-05, 0.0001288279, 0.0001882097, 0.0001830548, 
    7.732691e-05, 1.351043e-05, 2.371632e-05, 7.480857e-06, 7.915052e-07, 
    1.188035e-06, 7.820549e-06, 1.138086e-05, 1.12243e-05, 1.226609e-05,
  6.066487e-05, 0.0001057026, 0.0001595797, 0.0002235169, 0.0002165624, 
    8.023855e-05, 1.178191e-05, 1.772657e-05, 4.047036e-06, 6.61138e-07, 
    9.008131e-06, 2.539546e-05, 2.386994e-05, 1.272183e-05, 8.673069e-06,
  5.685887e-05, 0.0001226824, 0.0001935843, 0.0002434973, 0.0001883732, 
    5.974195e-05, 1.298252e-05, 1.01698e-05, 8.507665e-06, 2.340421e-07, 
    1.294667e-06, 2.648465e-05, 3.302403e-05, 8.653704e-06, 4.118693e-06,
  5.576628e-05, 0.0001139515, 0.0001476376, 0.0001658694, 0.0001018817, 
    2.900488e-05, 1.056428e-05, 5.594642e-06, 1.377829e-05, 6.401681e-07, 
    8.092604e-06, 1.696275e-05, 5.373675e-06, 3.775804e-06, 1.836601e-06,
  1.772119e-05, 4.929824e-05, 5.970715e-05, 6.792039e-05, 4.060261e-05, 
    2.824095e-05, 1.458746e-05, 3.779604e-06, 1.410515e-05, 3.982663e-06, 
    7.055402e-07, 1.612918e-05, 6.26182e-06, 8.794368e-07, 9.488454e-07,
  2.639031e-06, 6.619405e-06, 1.110197e-05, 2.145444e-05, 3.865786e-05, 
    3.579654e-05, 1.724862e-05, 3.254166e-06, 9.863042e-06, 7.849823e-06, 
    1.983536e-05, 7.865431e-07, 4.21918e-07, 1.110837e-06, 7.476926e-07,
  1.420064e-06, 4.061221e-06, 1.227294e-05, 3.468366e-05, 4.513669e-05, 
    3.711201e-05, 1.562095e-05, 3.354898e-06, 6.916314e-06, 1.071714e-05, 
    5.672663e-06, 6.380512e-07, 5.758458e-07, 1.267919e-06, 9.373572e-07,
  9.788253e-07, 3.462274e-06, 1.27341e-05, 3.229005e-05, 4.887098e-05, 
    4.164088e-05, 1.701944e-05, 3.709941e-06, 4.527836e-06, 8.885959e-06, 
    1.1104e-05, 4.356801e-06, 2.433567e-06, 8.031564e-07, 8.367122e-07,
  1.790045e-06, 8.92286e-05, 0.0002366983, 0.0002547914, 0.0001104426, 
    1.281434e-05, 4.710979e-07, 5.769873e-08, 2.751612e-07, 8.542894e-08, 
    4.257197e-06, 1.003573e-05, 7.492234e-06, 6.771651e-06, 4.569392e-06,
  5.749648e-07, 5.905403e-05, 0.000249393, 0.0002817529, 0.0001136057, 
    7.257625e-06, 2.070704e-07, 1.183788e-07, 1.199546e-07, 4.016996e-07, 
    4.691274e-06, 6.204511e-06, 3.997068e-06, 3.799188e-06, 3.90418e-06,
  2.128658e-07, 4.619133e-05, 0.000275688, 0.0003439252, 0.0001337714, 
    1.153125e-05, 2.73262e-07, 1.758655e-07, 1.226303e-07, 8.918833e-07, 
    3.379763e-06, 3.119872e-06, 2.553212e-06, 3.130759e-06, 4.241901e-06,
  1.071749e-06, 6.635105e-05, 0.0003154309, 0.0004366899, 0.000212623, 
    4.148518e-05, 6.108139e-07, 1.705985e-07, 3.751863e-07, 2.353536e-07, 
    9.735866e-07, 2.304485e-06, 4.253429e-06, 5.2583e-06, 3.58439e-06,
  3.672896e-06, 9.84746e-05, 0.0003516149, 0.0005279111, 0.0004137809, 
    0.000128789, 9.174726e-07, 1.551955e-07, 1.850871e-07, 5.328811e-07, 
    1.320849e-06, 2.601804e-06, 4.565184e-06, 5.726211e-06, 5.002964e-06,
  2.083008e-05, 0.0002051402, 0.0004552443, 0.000690805, 0.000648286, 
    0.0002283398, 2.485732e-06, 6.499838e-07, 3.408092e-07, 3.892052e-07, 
    1.485563e-06, 2.955302e-06, 4.578656e-06, 5.363197e-06, 4.769651e-06,
  8.665726e-05, 0.0002721161, 0.0004893399, 0.0008039978, 0.0008872079, 
    0.0003214265, 1.517962e-05, 1.336006e-06, 4.667209e-07, 2.064035e-07, 
    2.602711e-06, 3.978815e-06, 3.376655e-06, 4.355597e-06, 5.352508e-06,
  8.715471e-05, 0.0002362629, 0.0004215274, 0.000844743, 0.0009722456, 
    0.0003676326, 2.357938e-05, 8.058781e-07, 5.694196e-07, 3.403964e-07, 
    1.622839e-06, 3.48684e-06, 3.490263e-06, 4.290396e-06, 3.584397e-06,
  9.405199e-05, 0.0001803584, 0.0003677606, 0.0008715853, 0.001030722, 
    0.0004054109, 4.145837e-05, 5.243634e-07, 2.153288e-07, 3.580596e-07, 
    2.742863e-06, 4.699237e-06, 3.202002e-06, 3.759926e-06, 4.03067e-06,
  0.000101484, 0.0001652454, 0.0003792903, 0.0008635886, 0.001062668, 
    0.0004511212, 5.259475e-05, 3.248828e-07, 1.127814e-07, 8.13531e-07, 
    2.497879e-06, 3.432181e-06, 3.695684e-06, 4.380496e-06, 4.111282e-06,
  2.967928e-05, 1.969386e-05, 6.044479e-05, 7.04237e-05, 7.181416e-05, 
    4.345272e-05, 4.627537e-05, 5.020772e-05, 4.330769e-05, 3.973441e-05, 
    3.076555e-05, 1.52265e-05, 2.481526e-06, 2.208167e-06, 1.145039e-06,
  1.770146e-05, 3.779911e-05, 6.792929e-05, 0.0001098408, 6.612745e-05, 
    4.047645e-05, 6.708767e-05, 7.438236e-05, 5.503384e-05, 8.942114e-05, 
    2.393138e-05, 1.02688e-05, 2.726776e-06, 1.90477e-06, 1.492092e-06,
  1.136388e-05, 5.754186e-05, 0.0001259472, 0.0001450825, 7.597856e-05, 
    5.253833e-05, 9.115396e-05, 9.835567e-05, 7.294043e-05, 4.108011e-05, 
    6.543202e-05, 1.108668e-05, 3.733309e-06, 2.620789e-06, 1.741542e-06,
  7.287118e-06, 7.524479e-05, 0.0001745439, 0.0001861434, 8.002632e-05, 
    6.898632e-05, 0.0001174914, 0.0001304572, 9.416397e-05, 5.458268e-05, 
    6.345574e-05, 9.303488e-06, 2.461864e-06, 3.917937e-06, 2.985066e-06,
  6.78085e-06, 0.0001183944, 0.0002438695, 0.0002156798, 8.036981e-05, 
    8.896479e-05, 0.0001659582, 0.0001669882, 0.0001123184, 6.253942e-05, 
    6.136679e-05, 8.153919e-06, 3.206368e-06, 3.313426e-06, 3.729783e-06,
  3.575555e-05, 0.0001799856, 0.0003462739, 0.0002415322, 8.766785e-05, 
    0.0001074771, 0.0002161527, 0.0002068232, 0.0001293641, 7.065223e-05, 
    3.051399e-05, 3.107126e-06, 3.135589e-06, 3.512515e-06, 2.775548e-06,
  9.705983e-05, 0.0002809525, 0.0004845023, 0.0002706441, 9.528968e-05, 
    0.0001456623, 0.0002757238, 0.0002451338, 0.0001336485, 8.159772e-05, 
    3.838616e-05, 2.690826e-07, 1.563227e-06, 1.900001e-06, 3.107339e-06,
  0.000214473, 0.0004647318, 0.0006536518, 0.0003123426, 0.0001148897, 
    0.0001943666, 0.0003439947, 0.0002579447, 0.0001330453, 9.13768e-05, 
    3.51881e-05, 1.100783e-06, 1.222429e-06, 2.846079e-06, 2.199445e-06,
  0.0003090466, 0.000645726, 0.0007757772, 0.0003814903, 0.0001423241, 
    0.0002830009, 0.000383743, 0.0002987241, 0.0001583216, 9.635938e-05, 
    2.540986e-05, 2.904604e-06, 1.533937e-06, 3.086964e-06, 2.219418e-06,
  0.0003619734, 0.0007345101, 0.0008637785, 0.0004310191, 0.0001559695, 
    0.0003518338, 0.0004073314, 0.000309964, 0.000192755, 8.631692e-05, 
    1.740956e-05, 3.791047e-06, 1.588453e-06, 2.214025e-06, 3.237036e-06,
  0.0002286639, 8.544714e-05, 4.668119e-06, 1.235961e-06, 1.341703e-06, 
    5.542891e-07, 3.252567e-07, 7.79524e-08, 2.670364e-07, 2.292095e-06, 
    9.852183e-06, 1.260627e-05, 4.449545e-06, 4.067488e-06, 4.550801e-06,
  0.0002190452, 9.216911e-05, 9.069822e-06, 8.7764e-06, 8.08618e-06, 
    3.535758e-06, 4.559171e-07, 8.357156e-08, 2.606757e-07, 3.283807e-06, 
    8.76979e-06, 1.479252e-05, 6.462848e-06, 2.316348e-06, 2.333594e-06,
  0.0002032233, 9.491744e-05, 2.36585e-05, 2.008293e-05, 2.059338e-05, 
    1.581075e-05, 6.612444e-06, 1.108171e-06, 1.24157e-06, 1.675527e-06, 
    4.833041e-06, 2.494078e-05, 6.960873e-06, 2.058041e-06, 3.082474e-06,
  0.0001317751, 6.462471e-05, 2.296475e-05, 1.965505e-05, 1.969867e-05, 
    1.333918e-05, 7.586587e-06, 1.693218e-06, 6.167172e-07, 1.689885e-07, 
    1.02663e-05, 3.16925e-05, 8.319672e-06, 1.889123e-06, 1.844258e-06,
  6.42407e-05, 2.951116e-05, 9.724833e-06, 7.406969e-06, 5.628214e-06, 
    2.690977e-06, 1.389342e-06, 5.796519e-07, 1.04349e-07, 1.869743e-06, 
    4.551019e-06, 2.905919e-05, 1.164738e-05, 6.485501e-06, 2.164566e-06,
  3.655275e-05, 1.489984e-05, 3.407888e-06, 1.540292e-06, 1.459856e-07, 
    1.562302e-08, 1.7691e-08, 5.430772e-08, 1.151019e-08, 3.150928e-07, 
    4.068115e-06, 3.560481e-05, 2.137928e-05, 7.795186e-06, 2.740733e-06,
  3.393865e-05, 1.559264e-05, 1.475639e-06, 1.756956e-07, 4.353539e-08, 
    9.466385e-08, 2.79128e-07, 1.628657e-07, 1.096474e-08, 1.018549e-07, 
    6.961784e-06, 3.290588e-05, 2.608969e-05, 1.028755e-05, 4.67233e-06,
  2.959673e-05, 1.502941e-05, 1.778801e-06, 1.138178e-07, 6.911865e-08, 
    2.714953e-07, 1.095829e-06, 5.256695e-07, 2.583937e-08, 5.075133e-07, 
    1.584483e-05, 4.060436e-05, 3.139341e-05, 1.318167e-05, 3.295243e-06,
  1.685956e-05, 1.104009e-05, 4.391643e-06, 1.014667e-06, 2.156073e-06, 
    2.576325e-06, 2.043775e-06, 3.739898e-07, 1.60006e-07, 5.172035e-06, 
    2.451086e-05, 3.052687e-05, 2.729346e-05, 1.444358e-05, 2.199351e-06,
  2.697844e-06, 8.13933e-06, 4.601827e-06, 1.856241e-06, 9.59387e-06, 
    2.872691e-06, 2.973174e-06, 2.628673e-07, 8.420591e-07, 1.706707e-05, 
    4.492937e-05, 4.304769e-05, 3.972283e-05, 1.4716e-05, 1.513084e-06,
  0.0001269286, 0.0002747605, 0.0002196852, 3.193095e-05, 3.445072e-05, 
    7.891779e-05, 9.056904e-05, 3.555514e-05, 1.311074e-06, 1.73043e-06, 
    2.509431e-06, 1.908627e-06, 4.434025e-06, 7.385846e-06, 9.518237e-06,
  0.0001519986, 0.0004065735, 0.0003018069, 6.497658e-05, 3.488996e-05, 
    7.721226e-05, 0.0001050377, 4.111357e-05, 8.806965e-07, 1.239554e-06, 
    2.758252e-06, 3.599746e-06, 4.807921e-06, 7.359014e-06, 1.117581e-05,
  0.0001922215, 0.0004422415, 0.0004118036, 9.259942e-05, 3.914705e-05, 
    9.570409e-05, 0.0001323329, 5.262559e-05, 3.877054e-06, 1.651263e-06, 
    3.197287e-06, 6.357507e-06, 6.426581e-06, 7.061442e-06, 8.016006e-06,
  0.0002317496, 0.0004229347, 0.0004496254, 0.0001485594, 5.652706e-05, 
    0.0001358526, 0.000165392, 5.897583e-05, 5.556275e-06, 4.432044e-06, 
    2.625313e-06, 4.48279e-06, 6.618813e-06, 4.868065e-06, 5.90388e-06,
  0.0002496199, 0.0003735151, 0.0004478486, 0.0002138743, 7.242523e-05, 
    0.0001580601, 0.0001935344, 5.626749e-05, 2.880407e-06, 3.075409e-06, 
    6.042076e-06, 3.658988e-06, 4.719312e-06, 4.855631e-06, 5.84667e-06,
  0.0002433643, 0.0003228482, 0.0003905667, 0.0002272372, 8.204372e-05, 
    0.0001649519, 0.0001839192, 3.566077e-05, 2.587971e-06, 3.539562e-06, 
    6.23309e-06, 6.926967e-06, 5.92611e-06, 5.353163e-06, 3.89059e-06,
  0.0002370394, 0.0003237582, 0.0003597101, 0.0002080873, 9.41829e-05, 
    0.0001767714, 0.0001757271, 2.728286e-05, 4.661021e-06, 1.632002e-06, 
    4.634885e-06, 4.889725e-06, 8.290963e-06, 6.498807e-06, 5.345164e-06,
  0.0002443077, 0.0003240092, 0.0003475024, 0.0001912914, 0.0001072243, 
    0.0001982891, 0.0001704264, 2.991044e-05, 4.143847e-06, 7.60378e-07, 
    4.084958e-06, 4.873036e-06, 1.205678e-05, 7.995448e-06, 4.127328e-06,
  0.0002664929, 0.0002919534, 0.0002666855, 0.0001871138, 0.000122068, 
    0.0001890261, 0.0001659314, 4.700428e-05, 4.318696e-06, 3.218422e-07, 
    4.566232e-06, 8.050153e-06, 8.085291e-06, 8.357164e-06, 5.494252e-06,
  0.000259468, 0.0002632565, 0.0002266434, 0.0001716518, 0.00012411, 
    0.0001518502, 0.0001418342, 6.277537e-05, 5.61273e-06, 2.037681e-06, 
    5.96641e-06, 8.112403e-06, 9.581199e-06, 8.293626e-06, 6.731994e-06,
  9.214679e-05, 3.784741e-05, 9.893839e-06, 1.945317e-05, 3.108833e-05, 
    0.0001143929, 0.0001519326, 9.98598e-05, 6.991999e-05, 5.000012e-05, 
    5.093166e-05, 7.255293e-05, 4.214883e-05, 6.015803e-06, 2.93395e-06,
  6.865151e-05, 3.1278e-05, 4.69803e-07, 1.693212e-06, 1.466336e-05, 
    0.0001354912, 0.0002224403, 0.000121202, 6.774962e-05, 3.68805e-05, 
    4.399132e-05, 5.160891e-05, 2.577116e-05, 3.987735e-06, 2.848455e-06,
  4.320308e-05, 3.587165e-05, 1.043457e-05, 1.304787e-06, 2.561882e-06, 
    0.0001774728, 0.0003120782, 0.0001636665, 6.615814e-05, 4.537099e-05, 
    4.501609e-05, 2.173717e-05, 1.627549e-05, 5.895978e-06, 3.503225e-06,
  3.624917e-05, 5.766545e-05, 4.793779e-05, 8.34865e-06, 1.484897e-06, 
    0.0002140927, 0.0004346326, 0.000241346, 6.90319e-05, 5.804947e-05, 
    2.915691e-05, 4.030253e-05, 7.941737e-06, 6.008117e-06, 4.993276e-06,
  5.192848e-05, 7.739178e-05, 8.340465e-05, 8.610963e-06, 1.974339e-06, 
    0.0002003521, 0.0005073977, 0.0003242609, 8.669386e-05, 7.44389e-05, 
    4.325607e-05, 1.025715e-05, 1.547052e-06, 5.137671e-06, 6.399362e-06,
  6.106954e-05, 7.770201e-05, 4.729537e-05, 8.960181e-06, 2.252916e-06, 
    0.0001922852, 0.0005557737, 0.00047717, 0.0001268594, 9.210117e-05, 
    5.052089e-05, 1.493186e-06, 2.289239e-06, 5.110972e-06, 5.777103e-06,
  3.7966e-05, 5.715503e-05, 3.041748e-05, 7.499656e-07, 4.113155e-06, 
    0.0001886435, 0.0006504738, 0.0005819235, 0.0001815463, 0.0001055416, 
    7.16261e-05, 2.494248e-06, 3.816755e-06, 5.219549e-06, 6.263126e-06,
  2.569669e-05, 5.325169e-05, 1.297054e-05, 1.189539e-06, 3.069178e-06, 
    0.0001426774, 0.0007472942, 0.0007207366, 0.0002366394, 0.0001312782, 
    0.0001248333, 7.830683e-06, 3.573791e-06, 4.779833e-06, 5.907138e-06,
  2.734473e-05, 2.364012e-05, 9.801101e-06, 5.072811e-07, 2.992479e-06, 
    0.0001183998, 0.00071604, 0.0007699664, 0.0003081832, 0.0001546169, 
    0.0001621171, 2.913755e-05, 3.764418e-06, 4.035377e-06, 5.704858e-06,
  1.750657e-05, 3.048545e-05, 1.268904e-05, 4.599902e-06, 6.024767e-06, 
    0.0001568183, 0.0007531829, 0.0008366015, 0.0003858824, 0.0001540237, 
    0.0001446138, 4.230172e-05, 8.289207e-06, 5.088549e-06, 6.027164e-06,
  5.656622e-05, 8.792368e-05, 0.0001786455, 0.0001129188, 2.645045e-05, 
    1.185277e-05, 8.720825e-06, 5.417633e-06, 2.281801e-06, 5.699506e-06, 
    3.006198e-07, 2.457186e-06, 3.038983e-05, 5.064529e-05, 4.112059e-05,
  2.226179e-05, 0.0001076753, 0.0001966187, 0.0001382468, 3.556978e-05, 
    1.184436e-05, 1.139348e-05, 4.640789e-06, 6.774428e-07, 2.169017e-06, 
    1.550535e-05, 4.717273e-06, 1.502378e-05, 4.274943e-05, 3.629069e-05,
  2.254344e-05, 0.0001242084, 0.0001419948, 8.347388e-05, 3.234639e-05, 
    4.206138e-06, 8.490174e-06, 4.786112e-06, 5.023794e-07, 3.577265e-06, 
    3.374726e-06, 1.340505e-05, 4.767625e-05, 5.170621e-05, 7.343363e-05,
  2.768284e-05, 0.0001727112, 0.0001444983, 6.67569e-05, 5.027938e-05, 
    3.024022e-05, 1.274765e-05, 2.814369e-06, 1.124952e-06, 3.263962e-07, 
    7.376432e-07, 1.770419e-05, 2.788618e-05, 7.225944e-05, 7.989046e-05,
  5.97297e-05, 0.0001107562, 0.000184699, 7.329044e-05, 2.752725e-05, 
    1.196403e-05, 9.175312e-06, 3.571698e-06, 1.339153e-06, 1.184889e-06, 
    8.479396e-06, 1.397794e-05, 3.22918e-05, 4.565635e-05, 8.687576e-05,
  0.0001592923, 0.0002016633, 7.416117e-05, 4.753692e-05, 3.440752e-05, 
    2.319001e-05, 4.396744e-06, 5.193628e-06, 2.685991e-06, 6.193126e-06, 
    1.788816e-05, 2.927881e-05, 2.888265e-05, 4.659376e-05, 6.214681e-05,
  0.0001920304, 0.000125636, 5.53134e-05, 4.638262e-05, 3.507868e-05, 
    5.255853e-06, 1.882688e-06, 2.753892e-06, 4.441729e-06, 9.675918e-06, 
    2.593941e-05, 2.288284e-05, 1.491878e-05, 7.370747e-05, 5.917762e-05,
  0.0001788393, 8.544124e-05, 3.567666e-05, 3.49164e-05, 3.117751e-05, 
    1.497661e-05, 1.172206e-05, 1.084954e-06, 7.360278e-07, 9.235433e-06, 
    3.576662e-05, 3.157907e-05, 2.385325e-05, 3.152626e-05, 4.574632e-05,
  0.0001095852, 4.542256e-05, 2.267739e-05, 3.18044e-05, 2.131795e-05, 
    8.965913e-06, 3.687306e-06, 2.357291e-07, 2.318553e-07, 1.036082e-05, 
    6.107774e-05, 4.465716e-05, 2.188819e-05, 2.955349e-05, 3.742284e-05,
  8.596935e-05, 5.480119e-05, 3.547117e-05, 2.637946e-05, 1.368483e-05, 
    2.029395e-06, 8.108756e-08, 4.049884e-09, 1.705477e-07, 2.382236e-05, 
    0.0001209094, 7.51535e-05, 2.127608e-05, 1.708601e-05, 2.081445e-05,
  0.000156149, 0.0001154775, 8.337976e-05, 0.000118622, 0.0001665253, 
    0.0001294239, 1.953039e-05, 6.658506e-06, 9.67282e-06, 3.437167e-05, 
    2.340834e-05, 1.164864e-05, 1.278734e-05, 4.833292e-06, 5.966328e-06,
  0.0001818389, 0.0001179257, 7.185939e-05, 8.474337e-05, 0.0002170002, 
    0.0001524781, 8.010275e-06, 7.275379e-06, 1.036414e-05, 1.139371e-05, 
    8.522689e-06, 9.677884e-08, 1.217307e-05, 6.728409e-06, 6.469913e-06,
  0.0001784677, 0.0001181904, 7.813306e-05, 0.0001048902, 0.0002644394, 
    0.0001770243, 4.053984e-06, 6.229374e-06, 1.365632e-05, 1.63614e-05, 
    5.36002e-06, 1.426559e-07, 1.674387e-05, 7.391454e-06, 7.588707e-06,
  0.0001466745, 0.0001305565, 9.808628e-05, 0.0001416465, 0.0003478809, 
    0.0002082832, 2.448981e-06, 5.249976e-06, 2.161933e-05, 2.763939e-05, 
    9.520075e-06, 1.698624e-07, 1.552063e-05, 1.553544e-05, 5.764921e-06,
  0.0001305217, 0.0001142891, 0.0001064047, 0.0002060839, 0.0004352071, 
    0.0002521067, 1.99844e-06, 3.802505e-06, 3.675566e-05, 4.234672e-05, 
    9.339149e-06, 1.825007e-07, 7.731459e-06, 1.896932e-05, 5.977457e-06,
  0.0001256403, 0.0001238808, 0.0001173627, 0.0002606792, 0.0005399993, 
    0.0002732815, 2.341153e-06, 8.6817e-06, 5.163988e-05, 5.285265e-05, 
    7.140279e-06, 4.144654e-07, 9.009681e-06, 6.276207e-06, 7.926234e-06,
  0.0001460462, 0.0001292251, 0.0001332345, 0.0002769181, 0.0005813272, 
    0.0002839884, 1.907223e-06, 1.718339e-05, 7.088893e-05, 6.03032e-05, 
    4.619092e-06, 1.674247e-06, 7.757963e-06, 1.210262e-05, 8.936597e-06,
  0.0001568822, 0.0001328453, 0.0001203463, 0.0002794768, 0.0005956039, 
    0.0002779626, 2.728332e-06, 3.098935e-05, 9.06964e-05, 5.526619e-05, 
    5.773883e-06, 5.790489e-06, 4.645147e-06, 1.172704e-05, 8.781114e-06,
  0.0001605959, 0.0001176042, 0.0001167947, 0.0003064813, 0.0005975129, 
    0.0002549776, 5.739927e-06, 5.43793e-05, 0.0001058588, 3.353539e-05, 
    7.911141e-06, 8.923443e-06, 2.371118e-06, 8.636596e-07, 3.892886e-06,
  0.0001775129, 0.000120667, 0.0001237141, 0.0003375942, 0.000545752, 
    0.0002469762, 2.862391e-05, 8.143387e-05, 9.974711e-05, 5.40796e-06, 
    8.722615e-06, 7.885136e-06, 2.895579e-06, 2.845909e-06, 1.153515e-05,
  8.742758e-05, 4.849659e-05, 4.626867e-05, 2.767508e-05, 2.646235e-05, 
    4.943082e-05, 9.020407e-05, 6.68374e-05, 4.970065e-05, 2.704021e-05, 
    4.172103e-05, 4.660102e-05, 6.206289e-05, 5.839946e-05, 4.920709e-05,
  6.322417e-05, 5.216222e-05, 4.173614e-05, 3.118451e-05, 3.887617e-05, 
    8.01433e-05, 0.0001082539, 8.351948e-05, 7.564442e-05, 4.622938e-05, 
    5.658626e-05, 5.422651e-05, 6.841749e-05, 7.741522e-05, 5.161156e-05,
  4.67172e-05, 3.893731e-05, 3.256199e-05, 4.722669e-05, 7.784432e-05, 
    0.0001274691, 0.00014237, 0.0001013973, 7.159139e-05, 5.890168e-05, 
    6.149067e-05, 4.485266e-05, 6.763657e-05, 4.756551e-05, 4.956606e-05,
  3.343345e-05, 2.482483e-05, 4.635085e-05, 7.869752e-05, 0.0001238049, 
    0.0001583276, 0.0001514912, 0.000104563, 7.858553e-05, 7.022211e-05, 
    5.388161e-05, 6.740744e-05, 7.35733e-05, 6.65024e-05, 3.859106e-05,
  2.163652e-05, 3.825908e-05, 9.718061e-05, 0.0001408818, 0.0001536199, 
    0.0001710606, 0.0001380235, 9.657402e-05, 7.81385e-05, 8.1077e-05, 
    8.904613e-05, 6.204135e-05, 3.843318e-05, 3.549999e-05, 3.673277e-05,
  1.393681e-05, 8.074298e-05, 0.0001683258, 0.0002024093, 0.0001791206, 
    0.0001743674, 0.0001388471, 9.297047e-05, 0.0001091021, 8.834913e-05, 
    7.416723e-05, 4.041779e-05, 8.428032e-06, 2.601764e-05, 1.669092e-05,
  5.040009e-05, 0.0001604131, 0.0002365666, 0.0002324528, 0.0002109082, 
    0.0001667063, 0.0001334825, 9.60172e-05, 0.0001040426, 0.0001061013, 
    0.0001361321, 3.000433e-05, 5.599236e-06, 1.687411e-05, 3.207781e-06,
  0.0001607575, 0.000250314, 0.0002894586, 0.0002077187, 0.0001821442, 
    0.0001421796, 8.760028e-05, 8.135059e-05, 0.0001065273, 0.0001342007, 
    9.169926e-05, 1.166052e-05, 2.042653e-07, 5.531875e-07, 2.797093e-06,
  0.0002750945, 0.0003242825, 0.0003016269, 0.0001975875, 0.0001486947, 
    0.0001098802, 5.254033e-05, 0.0001025287, 0.000140777, 0.0001802242, 
    7.56649e-05, 1.517627e-06, 1.242684e-08, 5.10736e-07, 1.734542e-06,
  0.0003615708, 0.0003521577, 0.0002569425, 0.0001551607, 0.0001433638, 
    8.444803e-05, 6.849259e-05, 0.0001564539, 0.0002424203, 0.0001659642, 
    1.623839e-05, 1.548399e-07, 2.956772e-07, 9.117114e-07, 1.818088e-06,
  5.404057e-06, 1.601375e-05, 2.883555e-05, 3.497296e-05, 2.80152e-05, 
    2.154307e-05, 1.626217e-05, 7.967724e-06, 3.54544e-06, 9.807439e-07, 
    6.878803e-07, 1.734075e-07, 8.163862e-08, 1.447865e-09, 4.419399e-07,
  8.754011e-06, 1.950135e-05, 2.509651e-05, 3.515621e-05, 3.02734e-05, 
    2.384387e-05, 1.532619e-05, 1.08121e-05, 3.304935e-06, 2.144047e-06, 
    1.766341e-06, 8.399645e-07, 4.981973e-07, 4.783701e-07, 5.303793e-07,
  1.212608e-05, 2.066823e-05, 3.153286e-05, 3.271373e-05, 3.366378e-05, 
    2.392862e-05, 1.684952e-05, 8.980955e-06, 3.473498e-06, 3.491023e-06, 
    3.154785e-06, 1.692436e-06, 1.03493e-06, 1.098703e-06, 1.366302e-06,
  1.925364e-05, 3.008356e-05, 5.129642e-05, 3.763632e-05, 3.613262e-05, 
    2.53453e-05, 1.874173e-05, 1.070867e-05, 3.781766e-06, 2.997336e-06, 
    4.659249e-06, 1.931549e-06, 1.600547e-06, 1.060219e-06, 9.885753e-06,
  2.596652e-05, 3.310139e-05, 5.136625e-05, 3.928488e-05, 3.241146e-05, 
    2.809886e-05, 1.991661e-05, 9.658234e-06, 4.147165e-06, 3.36658e-06, 
    5.67593e-06, 3.763708e-06, 2.169813e-06, 2.199417e-06, 2.904485e-05,
  1.77869e-05, 2.703046e-05, 7.226779e-05, 4.639756e-05, 3.833229e-05, 
    3.164327e-05, 2.022882e-05, 1.006809e-05, 4.31871e-06, 6.230384e-06, 
    6.689232e-06, 5.8428e-06, 1.18466e-05, 1.343345e-05, 3.418635e-05,
  2.578959e-05, 2.289047e-05, 7.474328e-05, 5.153398e-05, 4.910923e-05, 
    4.226552e-05, 2.651022e-05, 1.792345e-05, 9.65965e-06, 1.261827e-05, 
    1.216144e-05, 7.114461e-06, 3.782524e-06, 1.826629e-05, 4.422899e-05,
  1.877549e-05, 2.457404e-05, 6.897571e-05, 5.870506e-05, 6.51198e-05, 
    6.660165e-05, 4.635226e-05, 2.852745e-05, 2.577693e-05, 1.159392e-05, 
    8.966538e-06, 1.955666e-05, 1.647521e-05, 2.909593e-05, 5.43798e-05,
  1.501559e-05, 2.47976e-05, 6.948817e-05, 6.17603e-05, 8.182912e-05, 
    7.592198e-05, 5.062394e-05, 3.762541e-05, 2.892137e-05, 1.612244e-05, 
    2.915118e-05, 1.620334e-05, 1.35852e-05, 2.385885e-05, 3.410563e-05,
  1.583088e-05, 2.120489e-05, 5.238637e-05, 7.097763e-05, 8.046407e-05, 
    7.109471e-05, 3.840945e-05, 1.487934e-05, 2.846728e-05, 2.184277e-05, 
    3.101819e-05, 2.402392e-05, 2.582769e-05, 5.691551e-05, 4.344297e-05,
  2.474624e-07, 3.090445e-07, 2.096915e-07, 2.533175e-08, 1.354745e-09, 
    9.954202e-10, 6.439989e-09, 8.846657e-09, 7.552134e-08, 3.86145e-07, 
    3.430455e-07, 3.712974e-07, 9.723146e-07, 1.938894e-06, 4.853521e-06,
  1.467408e-06, 2.925089e-07, 1.450792e-07, 5.229603e-08, 8.255074e-10, 
    3.439187e-09, 3.474442e-08, 1.155804e-09, 3.666062e-10, 2.286329e-09, 
    1.936689e-07, 7.438234e-07, 2.12183e-06, 3.04789e-06, 4.568235e-06,
  1.006475e-06, 8.470322e-07, 1.971561e-07, 8.884557e-08, 1.300819e-07, 
    1.236051e-08, 1.585287e-08, 9.815438e-08, 8.289384e-11, 1.339383e-09, 
    8.195444e-08, 2.124612e-07, 3.921592e-06, 2.977945e-06, 4.764087e-06,
  1.391466e-06, 1.101569e-06, 3.804254e-07, 1.699855e-07, 3.146077e-07, 
    1.00106e-07, 1.638862e-07, 7.026511e-08, 7.52563e-10, 1.983256e-09, 
    5.705247e-08, 3.546589e-07, 8.385596e-07, 3.015134e-06, 5.545717e-06,
  9.650181e-07, 8.728008e-07, 3.881592e-07, 5.837998e-08, 4.141594e-07, 
    2.366546e-07, 4.958823e-08, 8.929868e-09, 5.916125e-10, 1.814569e-09, 
    2.79431e-08, 1.199707e-07, 3.749968e-07, 2.061387e-06, 3.931258e-06,
  1.07303e-06, 1.063254e-06, 2.248128e-07, 2.00666e-07, 4.697793e-08, 
    1.004878e-08, 2.114699e-09, 1.294832e-08, 2.745206e-11, 1.471166e-10, 
    1.005029e-09, 3.840304e-08, 1.416324e-07, 2.39422e-06, 5.580519e-06,
  1.291874e-06, 8.439366e-07, 4.384634e-07, 7.024862e-08, 6.036178e-08, 
    7.258441e-09, 1.903784e-11, 3.974667e-11, 2.708745e-10, 2.365801e-11, 
    1.488886e-09, 1.307735e-10, 8.847458e-09, 1.114225e-06, 3.647799e-06,
  7.752074e-07, 4.900642e-07, 4.463705e-07, 2.934744e-07, 1.65605e-08, 
    1.231211e-08, 1.075269e-11, 1.480801e-12, 8.572086e-12, 5.065327e-11, 
    5.214201e-09, 4.336016e-10, 3.043136e-09, 9.103513e-09, 1.41551e-06,
  8.224611e-07, 6.165841e-07, 6.995734e-07, 1.999566e-07, 7.441124e-08, 
    1.986503e-08, 7.81337e-10, 2.532403e-12, 3.851594e-11, 7.507521e-12, 
    1.694177e-10, 9.3499e-10, 2.685913e-09, 1.318558e-08, 1.397785e-06,
  9.257093e-07, 8.592216e-07, 1.101248e-06, 2.737173e-07, 4.12496e-08, 
    2.449292e-09, 9.903997e-11, 1.239044e-11, 1.448136e-11, 2.044069e-10, 
    6.690014e-10, 1.379422e-09, 2.532684e-09, 2.661316e-07, 1.396528e-06,
  2.835847e-06, 7.672362e-08, 5.191303e-09, 1.193967e-06, 4.036307e-06, 
    3.581627e-06, 2.323972e-06, 2.84467e-06, 4.750671e-06, 5.864622e-06, 
    3.984185e-06, 3.140156e-06, 3.359102e-06, 4.919787e-06, 3.517243e-06,
  4.545248e-06, 2.025952e-07, 2.514254e-10, 7.926498e-07, 4.23718e-06, 
    1.553258e-06, 1.688816e-06, 4.725182e-06, 5.3024e-06, 4.256585e-06, 
    3.423014e-06, 3.339554e-06, 4.178958e-06, 5.927817e-06, 3.427367e-06,
  5.271501e-06, 1.129701e-07, 3.337565e-09, 7.459414e-07, 1.692258e-06, 
    1.089141e-06, 2.380332e-06, 5.15892e-06, 5.424048e-06, 5.18994e-06, 
    5.060719e-06, 6.372716e-06, 4.0296e-06, 4.419404e-06, 4.204948e-06,
  4.46219e-06, 4.598176e-08, 1.722508e-09, 8.520114e-08, 6.441072e-07, 
    1.402263e-06, 2.416651e-06, 4.309304e-06, 5.863786e-06, 3.921145e-06, 
    4.560131e-06, 7.493171e-06, 3.025738e-06, 4.881178e-06, 4.72631e-06,
  6.377255e-06, 8.660895e-08, 1.374555e-09, 1.595397e-07, 7.164593e-07, 
    1.102941e-06, 3.114161e-06, 3.312222e-06, 5.29539e-06, 5.076655e-06, 
    5.985251e-06, 4.129077e-06, 2.760315e-06, 5.004138e-06, 5.391128e-06,
  6.053463e-06, 4.346473e-07, 1.19124e-08, 1.022669e-08, 1.888343e-06, 
    2.095509e-06, 1.084533e-06, 2.764889e-06, 3.469835e-06, 3.755946e-06, 
    5.815904e-06, 4.991995e-06, 4.626563e-06, 2.631297e-06, 5.06234e-06,
  7.525123e-06, 2.241766e-06, 6.832586e-08, 9.517177e-09, 1.339291e-06, 
    2.790857e-06, 9.442845e-07, 2.178635e-06, 2.635114e-06, 2.095527e-06, 
    2.405537e-06, 3.884487e-06, 4.007442e-06, 3.994605e-06, 4.992611e-06,
  9.328831e-06, 4.313789e-06, 5.857567e-07, 6.441978e-09, 6.250023e-07, 
    2.418112e-06, 7.700528e-07, 1.05854e-06, 6.792172e-07, 1.23277e-07, 
    1.238046e-06, 3.896058e-06, 3.864891e-06, 5.598044e-06, 4.510574e-06,
  9.277303e-06, 5.271844e-06, 3.781215e-06, 6.550025e-08, 7.632232e-07, 
    5.627163e-07, 5.53401e-07, 8.967062e-07, 1.483525e-07, 4.5172e-08, 
    1.619416e-06, 2.138194e-06, 2.25195e-06, 2.200176e-06, 3.388102e-06,
  9.928546e-06, 4.635051e-06, 4.064149e-06, 1.092394e-07, 4.842583e-07, 
    2.622739e-06, 3.309565e-07, 7.773406e-08, 1.540717e-08, 1.957644e-10, 
    2.890995e-09, 6.328433e-07, 2.505753e-06, 2.865245e-06, 2.849123e-06,
  1.398999e-05, 1.18448e-05, 1.23266e-05, 1.360628e-05, 6.798928e-06, 
    6.878698e-07, 3.100989e-06, 3.93727e-06, 2.499771e-06, 2.288416e-06, 
    2.752966e-06, 2.409018e-06, 2.886625e-06, 5.536202e-06, 7.469707e-06,
  1.624693e-05, 1.780838e-05, 1.342941e-05, 1.495567e-05, 1.15984e-05, 
    3.780384e-06, 1.095664e-05, 9.873122e-06, 5.525194e-06, 4.057344e-06, 
    2.43563e-06, 2.498725e-06, 3.333417e-06, 3.07363e-06, 9.285657e-06,
  1.616931e-05, 2.12997e-05, 1.509588e-05, 9.87371e-06, 9.033195e-06, 
    7.284965e-06, 1.365773e-05, 9.756276e-06, 6.523515e-06, 5.083787e-06, 
    4.524404e-06, 2.245384e-06, 2.482934e-06, 3.919556e-06, 9.274302e-06,
  1.444275e-05, 2.234694e-05, 9.850404e-06, 9.630575e-06, 9.49408e-06, 
    1.058604e-05, 1.172399e-05, 9.651745e-06, 1.260177e-05, 1.099935e-05, 
    4.981945e-06, 4.71583e-06, 4.334087e-06, 5.451726e-06, 5.901424e-06,
  1.208321e-05, 1.744574e-05, 9.398424e-06, 3.897389e-06, 4.096077e-06, 
    9.375925e-06, 1.313581e-05, 1.012425e-05, 4.843235e-06, 5.430933e-06, 
    6.49632e-06, 7.414868e-06, 7.051738e-06, 1.048961e-05, 3.021119e-06,
  8.335859e-06, 1.426132e-05, 1.369489e-05, 3.935338e-06, 3.862529e-06, 
    7.584295e-06, 1.055487e-05, 1.032045e-05, 5.618898e-06, 4.188266e-06, 
    3.536097e-06, 5.024462e-06, 7.762129e-06, 9.368158e-06, 8.396524e-06,
  7.803072e-06, 1.139515e-05, 1.373869e-05, 6.841515e-06, 7.757833e-06, 
    7.770466e-06, 1.059012e-05, 1.113768e-05, 2.707433e-06, 1.577774e-06, 
    3.527306e-07, 1.441154e-06, 6.10606e-06, 7.097383e-06, 1.288007e-05,
  7.977893e-06, 6.216413e-06, 1.172406e-05, 8.724642e-06, 6.911341e-06, 
    9.157426e-06, 9.205959e-06, 6.566323e-06, 3.401104e-06, 1.083828e-06, 
    3.978873e-08, 2.65234e-07, 1.046736e-06, 3.373832e-06, 9.673156e-06,
  7.730551e-06, 7.210977e-06, 1.115766e-05, 9.868439e-06, 9.165388e-06, 
    8.593724e-06, 1.151767e-05, 5.546063e-06, 1.492718e-06, 3.77921e-08, 
    1.958926e-09, 2.350468e-09, 4.388886e-08, 1.345484e-07, 2.274452e-06,
  7.42704e-06, 6.146258e-06, 1.053582e-05, 1.162419e-05, 9.85809e-06, 
    9.606882e-06, 1.039495e-05, 4.489142e-06, 1.408563e-06, 4.614103e-08, 
    2.365831e-09, 4.459289e-10, 8.232475e-10, 1.040005e-08, 3.501322e-07,
  1.488635e-05, 6.67736e-06, 9.552504e-06, 1.219266e-05, 1.41035e-05, 
    9.204973e-06, 4.782217e-06, 3.215663e-06, 2.51066e-06, 2.176846e-06, 
    4.310008e-06, 7.78754e-06, 8.65741e-06, 1.045631e-05, 9.882054e-06,
  1.455624e-05, 8.437742e-06, 1.093036e-05, 1.082705e-05, 1.286237e-05, 
    1.007854e-05, 2.963653e-06, 2.600854e-06, 2.859581e-06, 2.717212e-06, 
    3.890549e-06, 6.057141e-06, 8.015045e-06, 1.239557e-05, 1.300943e-05,
  1.291489e-05, 7.645303e-06, 9.611612e-06, 1.190406e-05, 1.320325e-05, 
    8.775115e-06, 1.700686e-06, 4.40525e-06, 6.757546e-06, 1.43253e-06, 
    3.920414e-06, 5.888909e-06, 7.976449e-06, 1.042545e-05, 1.388416e-05,
  1.375048e-05, 9.812226e-06, 8.792464e-06, 1.155109e-05, 1.084197e-05, 
    8.128231e-06, 2.791329e-06, 4.06083e-06, 7.768882e-06, 4.301683e-06, 
    4.165382e-06, 9.869123e-06, 1.07612e-05, 1.073567e-05, 1.08213e-05,
  1.217585e-05, 9.453554e-06, 6.921463e-06, 1.029481e-05, 3.470309e-06, 
    2.677599e-06, 5.820343e-06, 4.028333e-06, 1.227178e-05, 9.845649e-06, 
    6.827932e-06, 9.145246e-06, 8.296571e-06, 9.652153e-06, 8.490485e-06,
  1.351188e-05, 1.1383e-05, 6.160647e-06, 7.596681e-06, 3.21744e-06, 
    3.91406e-06, 6.681077e-06, 4.577882e-06, 1.405112e-05, 8.564818e-06, 
    9.650704e-06, 7.240457e-06, 7.785146e-06, 3.578174e-06, 6.257276e-06,
  1.36476e-05, 1.27475e-05, 7.850836e-06, 8.153264e-06, 4.341047e-06, 
    3.313321e-06, 6.439093e-06, 5.706299e-06, 1.328572e-05, 7.91274e-06, 
    7.521847e-06, 1.015085e-05, 7.611677e-06, 6.290808e-06, 3.927758e-06,
  8.189731e-06, 1.385414e-05, 8.220174e-06, 5.4825e-06, 4.74225e-06, 
    2.517664e-06, 6.657641e-06, 6.635655e-06, 1.042417e-05, 7.2236e-06, 
    6.178672e-06, 6.88377e-06, 1.23267e-05, 9.114164e-06, 3.72963e-06,
  5.391933e-06, 1.283617e-05, 1.371824e-05, 6.818243e-06, 4.069819e-06, 
    1.137489e-06, 6.685837e-06, 8.473536e-06, 8.353534e-06, 6.313095e-06, 
    3.921058e-06, 3.773728e-06, 4.154304e-06, 6.922778e-06, 2.332639e-06,
  4.679682e-06, 1.321858e-05, 1.368887e-05, 8.144193e-06, 3.750857e-06, 
    2.750758e-06, 8.030385e-06, 9.827385e-06, 8.988573e-06, 6.02599e-06, 
    2.073017e-06, 1.585267e-06, 1.251049e-06, 5.524788e-06, 5.473085e-06,
  6.528147e-06, 8.083179e-06, 1.12392e-05, 1.094423e-05, 5.764093e-06, 
    3.093542e-06, 4.213274e-06, 2.416934e-06, 3.555052e-06, 6.502836e-06, 
    6.40298e-06, 4.360729e-06, 5.766363e-06, 7.563208e-06, 7.262409e-06,
  5.720429e-06, 7.577152e-06, 1.172298e-05, 9.928051e-06, 6.125718e-06, 
    6.73257e-06, 3.360115e-06, 4.16755e-06, 3.694164e-06, 4.123516e-06, 
    2.918949e-06, 4.654129e-06, 5.812366e-06, 7.914221e-06, 7.394309e-06,
  4.289634e-06, 7.21299e-06, 9.327468e-06, 9.020257e-06, 6.85359e-06, 
    7.547518e-06, 1.067739e-05, 4.868378e-06, 3.676301e-06, 5.213649e-06, 
    2.361853e-06, 4.249433e-06, 4.951225e-06, 6.266208e-06, 6.792607e-06,
  4.261374e-06, 6.809475e-06, 9.740765e-06, 1.194879e-05, 7.818358e-06, 
    2.090381e-06, 3.516769e-06, 3.165404e-06, 2.963991e-06, 4.733627e-06, 
    6.213947e-06, 5.678095e-06, 7.232767e-06, 7.329461e-06, 6.753194e-06,
  4.645766e-06, 8.49281e-06, 5.92747e-06, 4.607467e-06, 4.834608e-06, 
    2.892381e-06, 3.072872e-06, 4.445062e-06, 5.804584e-06, 6.633897e-06, 
    7.063725e-06, 8.747887e-06, 9.6337e-06, 7.362677e-06, 5.845088e-06,
  5.085195e-06, 7.985877e-06, 8.263043e-06, 4.476422e-06, 9.171213e-07, 
    2.235653e-06, 1.916814e-06, 5.5834e-06, 8.684635e-06, 6.55934e-06, 
    6.977383e-06, 9.506066e-06, 7.045199e-06, 4.952391e-06, 6.958625e-06,
  4.096535e-06, 5.253804e-06, 9.148523e-06, 4.381003e-06, 1.470863e-06, 
    9.869602e-07, 3.296314e-06, 5.74e-06, 8.234696e-06, 7.204973e-06, 
    5.742173e-06, 6.620867e-06, 7.493461e-06, 7.060814e-06, 4.716608e-06,
  3.809565e-06, 5.61641e-06, 8.325849e-06, 5.085259e-06, 3.69421e-06, 
    5.894897e-06, 6.014605e-06, 3.612155e-06, 8.869742e-06, 1.024649e-05, 
    1.241964e-05, 1.494529e-05, 1.54684e-05, 2.980045e-06, 2.36688e-06,
  3.908673e-06, 3.614443e-06, 2.390596e-06, 2.957757e-06, 4.889625e-06, 
    1.125194e-05, 1.327307e-05, 8.149515e-06, 1.165457e-05, 1.63236e-05, 
    1.420852e-05, 7.699284e-06, 1.767184e-06, 4.880001e-07, 1.368703e-06,
  4.106303e-06, 3.765327e-06, 2.017649e-06, 3.875014e-06, 3.842391e-06, 
    7.672096e-06, 1.324511e-05, 8.651731e-06, 7.505001e-06, 7.807178e-06, 
    9.185699e-06, 6.156557e-06, 8.787155e-07, 2.08186e-07, 1.42776e-07,
  7.3418e-05, 8.816768e-05, 9.633345e-05, 0.000106033, 0.0001181816, 
    6.297516e-05, 2.863143e-06, 4.039667e-07, 2.026274e-06, 4.97788e-06, 
    5.439862e-06, 5.843163e-06, 5.116454e-06, 4.639111e-06, 5.580989e-06,
  7.789371e-05, 0.0001064824, 0.0001052831, 0.0001066892, 0.0001240056, 
    4.62849e-05, 1.375386e-06, 4.96778e-08, 2.452402e-06, 5.641034e-06, 
    5.058572e-06, 6.014587e-06, 4.604917e-06, 5.913865e-06, 6.436318e-06,
  9.196495e-05, 0.0001157043, 0.0001142281, 0.0001122034, 0.0001254451, 
    3.725933e-05, 2.662617e-07, 7.832295e-07, 2.827774e-06, 3.420834e-06, 
    5.514121e-06, 6.670861e-06, 4.468503e-06, 5.480063e-06, 6.208685e-06,
  9.456131e-05, 0.0001089032, 0.0001162821, 0.0001170583, 0.0001110393, 
    2.231325e-05, 5.558857e-07, 1.986415e-06, 2.706587e-06, 5.102389e-06, 
    4.810052e-06, 3.765745e-06, 4.459634e-06, 4.908657e-06, 4.594477e-06,
  9.70254e-05, 0.0001135177, 0.0001080225, 0.0001140334, 8.001027e-05, 
    7.199602e-06, 2.114828e-06, 1.982092e-06, 2.372591e-06, 2.485667e-06, 
    3.851885e-06, 3.650038e-06, 3.290404e-06, 3.514476e-06, 3.934372e-06,
  9.025803e-05, 9.460292e-05, 9.589839e-05, 0.0001020094, 4.754369e-05, 
    5.250946e-06, 1.777284e-06, 2.588054e-06, 3.408705e-06, 4.242079e-06, 
    4.245821e-06, 5.156342e-06, 4.103968e-06, 5.123853e-06, 4.595594e-06,
  7.867974e-05, 8.476731e-05, 8.196157e-05, 6.987886e-05, 2.174185e-05, 
    4.446527e-06, 4.033267e-06, 3.551389e-06, 4.130219e-06, 4.968323e-06, 
    6.548148e-06, 1.042291e-05, 1.229901e-05, 7.996554e-06, 7.210814e-06,
  6.63688e-05, 6.713768e-05, 6.159216e-05, 4.023746e-05, 1.025831e-05, 
    8.544711e-06, 9.314675e-06, 5.502215e-06, 3.636241e-06, 5.106519e-06, 
    7.140513e-06, 9.355347e-06, 1.485861e-05, 1.098689e-05, 1.240186e-05,
  5.430214e-05, 5.102605e-05, 3.937758e-05, 1.79655e-05, 1.041028e-05, 
    5.185891e-06, 6.901349e-06, 8.789237e-06, 9.605386e-06, 5.847141e-06, 
    5.778822e-06, 8.575685e-06, 1.27381e-05, 1.879221e-05, 1.883951e-05,
  4.412766e-05, 3.102534e-05, 1.890072e-05, 9.822177e-06, 8.018528e-06, 
    8.107862e-06, 9.176376e-06, 8.628339e-06, 6.668673e-06, 8.068165e-06, 
    8.338576e-06, 1.107093e-05, 1.886872e-05, 1.701008e-05, 2.082818e-05,
  3.10858e-06, 4.885593e-07, 3.861021e-07, 1.54345e-05, 0.0001224689, 
    0.0001714446, 4.221251e-05, 4.044187e-07, 2.163698e-07, 2.164474e-06, 
    3.844172e-06, 5.787675e-06, 4.361858e-06, 4.538917e-06, 4.951157e-06,
  3.579259e-07, 2.740732e-07, 3.85675e-07, 1.16924e-05, 0.0001657841, 
    0.0002485673, 3.159593e-05, 9.113331e-08, 2.980519e-07, 2.044723e-06, 
    4.496261e-06, 4.135153e-06, 3.191356e-06, 3.60794e-06, 3.224015e-06,
  7.840137e-09, 9.652345e-09, 1.875318e-07, 9.167788e-06, 0.000226496, 
    0.0003220853, 4.195944e-05, 2.77724e-07, 1.050151e-06, 3.767889e-06, 
    6.606193e-06, 2.945983e-06, 3.145268e-06, 3.063518e-06, 3.254631e-06,
  1.349995e-09, 7.443695e-08, 6.060292e-07, 1.919721e-05, 0.0002619219, 
    0.0003774189, 4.29824e-05, 4.494125e-08, 2.157907e-06, 2.912326e-06, 
    3.052075e-06, 2.624945e-06, 2.614264e-06, 2.982604e-06, 2.022916e-06,
  3.804831e-09, 1.8254e-07, 2.717774e-06, 3.926604e-05, 0.0002923362, 
    0.0004031783, 4.181432e-05, 2.681153e-08, 2.235301e-06, 1.427102e-06, 
    2.699162e-06, 1.949094e-06, 2.220976e-06, 2.338442e-06, 2.526726e-06,
  4.275164e-08, 5.342919e-07, 1.184722e-05, 7.531299e-05, 0.0003214523, 
    0.0003730337, 3.279758e-05, 2.93152e-07, 1.648632e-06, 1.584503e-06, 
    2.542556e-06, 2.34875e-06, 2.710817e-06, 3.586103e-06, 2.857256e-06,
  1.793248e-07, 7.381365e-07, 1.334743e-05, 9.029858e-05, 0.0003133701, 
    0.0003216609, 3.633516e-05, 6.656872e-07, 2.1217e-06, 1.923406e-06, 
    2.620651e-06, 3.748005e-06, 4.886921e-06, 7.622792e-06, 6.386387e-06,
  3.886969e-07, 1.685186e-06, 6.084129e-06, 6.340126e-05, 0.0002625847, 
    0.0002757148, 3.292463e-05, 4.075698e-07, 2.349741e-06, 2.559085e-06, 
    2.802948e-06, 3.249007e-06, 4.281978e-06, 7.355872e-06, 1.45685e-05,
  3.207163e-07, 1.82078e-06, 1.873239e-05, 6.44405e-05, 0.0002236388, 
    0.0002267386, 1.896891e-05, 1.246022e-06, 2.82454e-06, 8.172023e-06, 
    6.923664e-06, 7.582806e-06, 6.485401e-06, 8.661168e-06, 1.298999e-05,
  2.941121e-06, 1.291744e-05, 3.799144e-05, 8.446813e-05, 0.000191051, 
    0.0001406, 6.961886e-06, 5.154692e-06, 8.762639e-06, 1.475089e-05, 
    1.416969e-05, 1.05533e-05, 7.180989e-06, 1.321824e-05, 1.705906e-05,
  0.0006349849, 0.0006872684, 0.0003589807, 5.088945e-05, 2.081059e-07, 
    4.495057e-08, 1.415115e-07, 2.018876e-06, 3.807533e-06, 4.735771e-06, 
    5.366583e-06, 6.194374e-06, 5.104509e-06, 6.912955e-06, 6.579295e-06,
  0.0006973158, 0.000720147, 0.0003516509, 4.147723e-05, 6.028314e-07, 
    6.702517e-07, 5.458597e-08, 1.406131e-06, 4.766884e-06, 4.225826e-06, 
    5.143798e-06, 4.941727e-06, 4.808216e-06, 6.202768e-06, 6.382812e-06,
  0.0007100504, 0.0007479245, 0.0004002708, 4.204918e-05, 2.192593e-06, 
    1.092302e-06, 6.324512e-08, 1.424718e-06, 4.936974e-06, 2.42211e-06, 
    3.294719e-06, 4.542493e-06, 4.904e-06, 5.571067e-06, 6.367222e-06,
  0.000645159, 0.0007607678, 0.0004681894, 4.959609e-05, 4.449786e-06, 
    3.573536e-06, 3.982493e-07, 4.59592e-07, 2.358985e-06, 2.778415e-06, 
    4.284316e-06, 4.11817e-06, 4.691545e-06, 6.926629e-06, 9.207559e-06,
  0.0005980263, 0.000747395, 0.0004992841, 6.906233e-05, 6.83115e-06, 
    9.740456e-06, 1.57923e-06, 4.315526e-07, 1.748558e-06, 1.502304e-06, 
    3.078604e-06, 4.297437e-06, 5.460684e-06, 7.918321e-06, 1.192793e-05,
  0.0005736243, 0.0007167218, 0.0004699468, 8.41287e-05, 1.367031e-05, 
    1.857196e-05, 4.909341e-06, 1.075707e-06, 2.167873e-06, 2.636814e-06, 
    5.151422e-06, 7.404644e-06, 1.218789e-05, 9.595431e-06, 8.518108e-06,
  0.0005718837, 0.0006704427, 0.0004293232, 0.0001068681, 3.22552e-05, 
    3.026628e-05, 7.243856e-06, 8.821189e-07, 1.399077e-06, 1.966015e-06, 
    4.461859e-06, 7.975737e-06, 8.700121e-06, 1.130776e-05, 5.873848e-06,
  0.0005423292, 0.000582532, 0.0003839933, 0.000130611, 7.134113e-05, 
    3.678848e-05, 5.407284e-06, 8.832327e-07, 1.862958e-06, 1.516691e-06, 
    5.086186e-06, 7.640793e-06, 9.249777e-06, 1.116529e-05, 7.88765e-06,
  0.0004819561, 0.0004753116, 0.0003026968, 0.0001294184, 9.010884e-05, 
    3.056685e-05, 3.846954e-06, 8.336589e-07, 2.180373e-06, 2.15309e-06, 
    2.990952e-06, 6.133585e-06, 9.011947e-06, 6.589831e-06, 1.064066e-05,
  0.0004060546, 0.0003383318, 0.0002350245, 0.0001237369, 9.540033e-05, 
    3.156328e-05, 1.8465e-06, 1.137493e-06, 2.790404e-06, 3.980352e-06, 
    5.832135e-06, 7.212238e-06, 7.804741e-06, 7.207516e-06, 1.30929e-05,
  0.0003136354, 0.0003276306, 0.0002102765, 0.0001596038, 0.0001551518, 
    0.0001371433, 8.383317e-05, 2.756416e-05, 7.537987e-06, 2.187783e-05, 
    2.120073e-05, 1.870261e-05, 1.974148e-05, 1.235473e-05, 5.751386e-06,
  0.0004207227, 0.0004050531, 0.0002418298, 0.0001932905, 0.0001858869, 
    0.0001633802, 9.570859e-05, 3.223004e-05, 8.703759e-06, 1.82001e-05, 
    1.658806e-05, 2.119255e-05, 2.353936e-05, 1.138796e-05, 6.107644e-06,
  0.0004797037, 0.0004786836, 0.0002763443, 0.0002243917, 0.0002263616, 
    0.0001738034, 9.859855e-05, 4.092445e-05, 1.219011e-05, 7.093459e-06, 
    1.536852e-05, 2.152348e-05, 2.504953e-05, 1.139559e-05, 6.278549e-06,
  0.0005343069, 0.0004747326, 0.0002675158, 0.0002219768, 0.0002367361, 
    0.0001833596, 0.0001096436, 4.858681e-05, 1.402706e-05, 1.136719e-05, 
    6.817771e-06, 1.684582e-05, 3.607993e-05, 9.099877e-06, 4.969735e-06,
  0.0005981853, 0.0004363985, 0.0002460715, 0.0002164836, 0.0002534376, 
    0.0002063928, 0.0001197286, 5.888419e-05, 1.662132e-05, 7.134748e-06, 
    1.025179e-05, 2.47333e-05, 2.501482e-05, 5.986018e-06, 3.210667e-06,
  0.0005539108, 0.0003582757, 0.0002182691, 0.0001872947, 0.0002707335, 
    0.0002134604, 0.0001256937, 6.397157e-05, 2.130942e-05, 6.452327e-06, 
    5.192164e-06, 1.719798e-05, 1.160631e-05, 6.219309e-06, 5.497243e-06,
  0.0004948204, 0.0002099793, 0.0001182885, 0.0001696306, 0.0002732, 
    0.0002487779, 0.0001358074, 6.584367e-05, 2.52554e-05, 7.223374e-06, 
    4.942541e-06, 1.541831e-05, 5.357497e-06, 4.306672e-06, 4.108855e-06,
  0.0004299275, 0.0002190284, 8.993799e-05, 0.0001565042, 0.0002618572, 
    0.0002531719, 0.0001520694, 8.099653e-05, 2.661923e-05, 7.162568e-06, 
    6.388773e-06, 1.111138e-05, 1.627478e-06, 4.466873e-06, 3.176759e-06,
  0.0003662192, 0.0001802535, 9.185448e-05, 0.0001511607, 0.00024159, 
    0.0002509659, 0.0001664325, 9.306081e-05, 3.832702e-05, 1.032604e-05, 
    9.474842e-06, 9.070563e-06, 5.796499e-06, 5.784421e-06, 5.869239e-06,
  0.000310935, 0.0001852462, 0.0001111291, 0.0001594173, 0.0002149161, 
    0.0002303843, 0.0001873653, 0.000118997, 4.990483e-05, 1.463146e-05, 
    8.759144e-06, 3.669481e-06, 5.281521e-06, 7.508477e-06, 7.139721e-06,
  3.11322e-06, 1.624744e-06, 9.227186e-07, 1.354976e-06, 1.380753e-06, 
    7.751498e-07, 1.373859e-06, 1.371443e-06, 9.367592e-07, 9.712784e-07, 
    2.446678e-06, 2.728014e-06, 1.349617e-05, 3.181447e-05, 4.011695e-05,
  3.330124e-06, 2.016138e-06, 1.631155e-06, 6.359578e-07, 4.675247e-07, 
    5.642669e-07, 4.050899e-07, 3.48955e-07, 7.23387e-09, 6.96115e-10, 
    1.320823e-06, 4.607108e-06, 5.582777e-06, 3.659556e-05, 3.900457e-05,
  5.688116e-06, 3.292162e-06, 1.777987e-06, 1.180855e-06, 1.58284e-08, 
    1.130507e-08, 2.029954e-07, 1.763029e-08, 7.251496e-11, 1.486665e-10, 
    8.336542e-07, 8.431538e-07, 1.168934e-05, 3.498664e-05, 4.836836e-05,
  1.37261e-05, 8.197388e-06, 3.209722e-06, 1.468541e-06, 6.269517e-07, 
    1.463583e-07, 1.107661e-07, 8.877127e-10, 8.249547e-13, 1.484004e-11, 
    1.297753e-10, 1.001088e-07, 1.039245e-05, 3.889414e-05, 4.225919e-05,
  2.328447e-05, 1.573068e-05, 6.824976e-06, 2.687212e-06, 1.902226e-06, 
    4.632829e-07, 1.055632e-07, 4.637106e-16, 2.643903e-13, 6.502509e-12, 
    1.312413e-11, 7.593206e-08, 1.100017e-05, 3.969581e-05, 4.288396e-05,
  2.423417e-05, 2.216338e-05, 1.672317e-05, 6.719936e-06, 2.946477e-06, 
    1.111415e-06, 2.271727e-07, 4.435092e-08, 6.242495e-18, 6.040558e-12, 
    7.85209e-11, 2.821834e-06, 1.611887e-05, 2.835146e-05, 4.848529e-05,
  4.134371e-05, 3.267474e-05, 2.606814e-05, 1.491367e-05, 5.778605e-06, 
    2.047339e-06, 4.797077e-07, 7.642389e-08, 3.314378e-08, 6.993901e-11, 
    2.680561e-08, 1.734301e-06, 2.093018e-05, 4.381519e-05, 4.773513e-05,
  3.798104e-05, 3.497366e-05, 3.316854e-05, 1.99552e-05, 1.023414e-05, 
    2.779973e-06, 6.336848e-07, 1.954049e-07, 1.129304e-07, 1.513678e-10, 
    2.917501e-07, 7.002415e-06, 2.21776e-05, 4.764121e-05, 3.504962e-05,
  6.919415e-05, 6.345801e-05, 4.506442e-05, 2.346111e-05, 1.105983e-05, 
    3.495614e-06, 1.1155e-06, 2.148133e-07, 1.101188e-07, 2.108846e-08, 
    1.171786e-07, 4.817125e-06, 3.053667e-05, 3.789629e-05, 3.064216e-05,
  6.739223e-05, 7.255386e-05, 5.551332e-05, 3.075738e-05, 1.39595e-05, 
    4.53697e-06, 1.13381e-06, 2.835766e-07, 1.053762e-07, 3.057031e-07, 
    2.237795e-06, 9.533548e-06, 1.990523e-05, 4.347939e-05, 3.358977e-05,
  7.380318e-05, 8.464616e-05, 8.410747e-05, 7.452946e-05, 6.827847e-05, 
    6.830655e-05, 9.615051e-05, 0.0001378711, 0.0001432255, 0.0001162084, 
    0.0001034523, 8.445464e-05, 6.384329e-05, 4.76358e-05, 3.150916e-05,
  9.160793e-05, 0.0001021677, 0.00010613, 8.891121e-05, 8.440122e-05, 
    9.355443e-05, 0.0001077479, 0.0001174884, 0.0001257807, 0.0001297429, 
    0.0001330017, 8.916645e-05, 6.55436e-05, 4.825493e-05, 3.447208e-05,
  0.0001133121, 0.0001159358, 0.0001098674, 9.97864e-05, 9.460234e-05, 
    0.0001045222, 0.000124357, 0.0001552673, 0.0001764089, 0.0001193803, 
    9.63101e-05, 8.779007e-05, 6.136148e-05, 4.727051e-05, 3.133366e-05,
  0.0001240507, 0.0001148775, 0.0001123125, 0.0001056142, 0.0001040529, 
    0.0001210264, 0.0001445197, 0.0001619697, 0.0001375225, 0.000117659, 
    8.36307e-05, 7.182816e-05, 5.155787e-05, 3.822015e-05, 2.858835e-05,
  0.0001264822, 0.0001159202, 0.0001125455, 0.0001150422, 0.0001211264, 
    0.0001276943, 0.0001566704, 0.0001582517, 0.0001421223, 9.877944e-05, 
    0.0001022629, 6.572983e-05, 5.083565e-05, 3.80075e-05, 2.213217e-05,
  0.0001276227, 0.0001068344, 0.0001123147, 0.0001184915, 0.000131509, 
    0.0001584339, 0.000159233, 0.0001609186, 0.0001330909, 0.000105479, 
    8.248278e-05, 6.128679e-05, 4.543262e-05, 3.800332e-05, 1.583988e-05,
  0.00012008, 0.000110332, 0.0001176837, 0.0001240021, 0.0001445146, 
    0.0001598731, 0.000166755, 0.0001618423, 0.0001264325, 0.0001041668, 
    7.9346e-05, 5.441956e-05, 4.864034e-05, 2.935601e-05, 1.124248e-05,
  0.000126173, 0.0001224389, 0.0001327449, 0.0001423416, 0.000160151, 
    0.0001742207, 0.0001636938, 0.0001507946, 0.0001268436, 0.0001069172, 
    7.757475e-05, 5.809838e-05, 3.552982e-05, 2.263667e-05, 1.005471e-05,
  0.000139699, 0.0001288069, 0.0001463492, 0.000167077, 0.0001729077, 
    0.0001763179, 0.0001655262, 0.0001434934, 0.0001251017, 9.376327e-05, 
    8.786427e-05, 4.811984e-05, 2.171871e-05, 1.493143e-05, 8.467052e-06,
  0.0001364796, 0.0001413463, 0.0001588936, 0.0001785703, 0.0001749146, 
    0.0001669708, 0.0001593091, 0.0001449954, 0.0001211008, 9.945681e-05, 
    7.160309e-05, 2.518639e-05, 1.04075e-05, 1.118984e-05, 7.896897e-06,
  6.34815e-05, 6.736643e-05, 0.0001021517, 7.530107e-05, 0.0001017664, 
    0.0001396068, 5.343205e-05, 3.432677e-05, 1.696282e-05, 6.867838e-06, 
    3.010534e-06, 1.587346e-06, 1.000073e-06, 1.169091e-06, 1.401405e-06,
  0.000114529, 9.820212e-05, 8.803985e-05, 0.0001012531, 9.573134e-05, 
    9.880408e-05, 6.341845e-05, 4.126137e-05, 2.991002e-05, 1.161817e-05, 
    4.735999e-06, 1.818123e-06, 6.083036e-07, 9.354828e-07, 3.481428e-06,
  9.863983e-05, 9.800872e-05, 8.083999e-05, 0.0001224703, 0.000123726, 
    0.0001594884, 8.155586e-05, 7.979507e-05, 2.682975e-05, 1.095498e-05, 
    4.166607e-06, 1.847994e-06, 1.021639e-06, 4.164877e-06, 7.55307e-06,
  0.0001292574, 0.0001051756, 0.0001138526, 0.0001037594, 0.0001007983, 
    0.0001110721, 7.773472e-05, 9.482223e-05, 4.413656e-05, 1.287119e-05, 
    4.871669e-06, 1.787455e-06, 2.28589e-06, 8.304803e-06, 1.712319e-05,
  0.0001309315, 0.0001095001, 0.0001015366, 0.0001028016, 9.453417e-05, 
    0.0001072965, 0.0001253688, 8.418599e-05, 4.730868e-05, 1.895021e-05, 
    4.942508e-06, 2.358729e-06, 4.159121e-06, 1.172204e-05, 2.585622e-05,
  0.0001440098, 0.0001195, 0.0001136025, 0.0001122227, 9.692794e-05, 
    7.719958e-05, 0.0001286551, 7.954138e-05, 4.270473e-05, 2.060164e-05, 
    7.119562e-06, 4.385729e-06, 6.799611e-06, 2.555399e-05, 3.487167e-05,
  0.0001520109, 0.0001410824, 0.0001242263, 0.0001171318, 0.000109709, 
    9.775562e-05, 8.674482e-05, 6.244263e-05, 5.988881e-05, 1.638159e-05, 
    9.123914e-06, 7.349792e-06, 2.182811e-05, 4.241874e-05, 3.908644e-05,
  0.0001551301, 0.0001412392, 0.0001200929, 0.000103172, 6.160256e-05, 
    6.397194e-05, 7.714589e-05, 7.065511e-05, 4.238005e-05, 3.881829e-05, 
    1.706107e-05, 2.555326e-05, 4.490574e-05, 5.174392e-05, 3.719179e-05,
  0.0001558443, 0.0001419882, 0.0001100281, 8.439821e-05, 8.19308e-05, 
    8.524382e-05, 6.47671e-05, 4.02185e-05, 3.259736e-05, 2.875064e-05, 
    2.816489e-05, 5.278646e-05, 6.769809e-05, 5.212357e-05, 3.355409e-05,
  0.0001374822, 0.0001263974, 0.0001030652, 0.0001063457, 8.853681e-05, 
    8.761938e-05, 7.511768e-05, 5.674865e-05, 6.078859e-05, 4.134449e-05, 
    6.481983e-05, 8.213102e-05, 8.215899e-05, 4.634035e-05, 3.043031e-05,
  2.198727e-05, 1.670074e-05, 1.883161e-05, 1.163321e-05, 9.843127e-06, 
    1.164773e-07, 1.14544e-07, 4.163371e-08, 2.550109e-08, 1.603657e-08, 
    4.589363e-08, 1.444405e-08, 3.935666e-07, 4.394146e-07, 5.594875e-07,
  2.517834e-05, 2.257e-05, 3.366009e-05, 1.773408e-05, 9.118844e-06, 
    1.078317e-07, 7.027204e-09, 2.180033e-09, 1.61617e-08, 8.812926e-09, 
    4.267029e-08, 1.220408e-08, 3.865746e-09, 1.274505e-08, 5.811553e-07,
  2.952307e-05, 1.933471e-05, 1.747742e-05, 1.976496e-05, 1.050992e-05, 
    4.639429e-07, 1.005023e-08, 1.708427e-08, 4.617038e-08, 2.229359e-08, 
    1.487022e-07, 5.277293e-09, 3.622518e-09, 1.579673e-07, 2.295713e-08,
  2.476936e-05, 2.03239e-05, 1.683596e-05, 1.697008e-05, 5.763516e-06, 
    3.015708e-06, 3.058411e-08, 6.33303e-08, 3.491505e-08, 1.724755e-07, 
    1.611478e-07, 8.797327e-10, 2.44035e-10, 2.680878e-08, 5.21933e-08,
  2.550882e-05, 2.327177e-05, 1.961239e-05, 1.1516e-05, 2.27916e-06, 
    2.807205e-06, 4.770135e-07, 8.127953e-08, 7.054988e-08, 2.096073e-07, 
    1.449869e-07, 1.633684e-09, 1.919001e-09, 3.085874e-10, 2.02712e-10,
  2.538074e-05, 3.111241e-05, 2.555994e-05, 1.71236e-05, 7.645292e-06, 
    5.649113e-06, 5.055811e-07, 1.643904e-07, 1.66981e-07, 3.487712e-07, 
    6.345994e-08, 4.666176e-08, 6.839437e-10, 1.014248e-09, 3.016474e-08,
  2.613236e-05, 3.919813e-05, 3.663128e-05, 2.583362e-05, 1.444622e-05, 
    2.184813e-06, 8.304575e-07, 3.662919e-07, 2.603341e-07, 3.310436e-07, 
    6.719392e-08, 6.232174e-09, 7.806275e-10, 2.975019e-10, 2.695648e-09,
  2.628313e-05, 4.204387e-05, 4.553997e-05, 3.583454e-05, 1.105292e-05, 
    2.367769e-06, 1.918608e-06, 4.324574e-07, 2.871066e-07, 4.654207e-07, 
    5.470499e-08, 9.225155e-09, 2.802948e-09, 2.711327e-09, 1.379822e-08,
  2.562748e-05, 4.714395e-05, 5.102801e-05, 3.834725e-05, 1.07689e-05, 
    3.696828e-06, 2.254767e-06, 7.743573e-07, 3.805628e-07, 8.735239e-07, 
    3.536854e-07, 1.045031e-08, 1.578038e-08, 3.613563e-08, 2.63215e-08,
  2.844604e-05, 5.042183e-05, 5.451541e-05, 3.376994e-05, 9.617293e-06, 
    4.064654e-06, 2.77953e-06, 1.780685e-06, 1.16922e-06, 1.235119e-06, 
    2.971414e-07, 4.744165e-07, 3.329193e-07, 5.428029e-09, 1.281737e-08,
  0.0002100548, 0.0002552332, 0.0002556801, 0.0001691671, 5.182603e-05, 
    1.385582e-06, 1.686056e-06, 3.039612e-06, 2.985706e-06, 4.225804e-06, 
    4.160469e-06, 4.111662e-06, 3.785788e-06, 6.956374e-06, 6.605576e-06,
  0.0002303244, 0.0002700033, 0.0002625532, 0.0001544504, 3.438107e-05, 
    6.523786e-07, 5.666595e-07, 3.625427e-06, 2.983117e-06, 4.286944e-06, 
    5.61607e-06, 7.13955e-06, 4.993336e-06, 7.166488e-06, 8.543596e-06,
  0.0002478654, 0.0002506522, 0.0002536268, 0.0001271384, 2.614878e-05, 
    2.993345e-06, 7.240043e-07, 6.071291e-06, 7.736232e-06, 8.247307e-06, 
    8.174632e-06, 5.353229e-06, 6.090679e-06, 6.806261e-06, 7.329314e-06,
  0.000254774, 0.0002492479, 0.000213796, 8.674465e-05, 1.457147e-05, 
    8.667897e-06, 2.1469e-06, 5.223667e-06, 7.916235e-06, 4.945693e-06, 
    3.829984e-06, 3.438238e-06, 4.899608e-06, 5.631643e-06, 6.950464e-06,
  0.0002494491, 0.0002275148, 0.0001606868, 7.913904e-05, 3.271314e-05, 
    1.696885e-05, 1.425752e-06, 5.146536e-06, 6.544965e-06, 4.757478e-06, 
    4.283786e-06, 2.725704e-06, 3.023183e-06, 4.667634e-06, 4.970661e-06,
  0.0002365003, 0.000174933, 0.000104715, 2.517541e-05, 4.189484e-05, 
    2.191203e-05, 2.836546e-06, 6.096131e-06, 7.990845e-06, 4.429347e-06, 
    4.943883e-06, 4.230338e-06, 2.88643e-06, 3.670392e-06, 3.419537e-06,
  0.0001831558, 0.0001030287, 2.481685e-05, 2.423696e-05, 2.229781e-05, 
    4.621347e-05, 1.354063e-05, 6.42207e-06, 1.001033e-05, 1.072403e-05, 
    8.36002e-06, 5.463319e-06, 2.399341e-06, 4.598495e-06, 3.328599e-06,
  9.485002e-05, 3.093155e-05, 1.32917e-05, 1.087835e-05, 2.397993e-05, 
    1.555059e-05, 5.789441e-06, 4.971105e-06, 6.211889e-06, 8.744007e-06, 
    7.148903e-06, 5.267083e-06, 3.88176e-06, 5.550731e-06, 3.515551e-06,
  1.744398e-05, 1.881532e-05, 1.310391e-05, 1.714989e-05, 2.80271e-05, 
    1.460151e-05, 1.48673e-06, 4.163053e-06, 3.894549e-06, 6.932952e-06, 
    5.561927e-06, 6.315785e-06, 6.45269e-06, 2.753756e-06, 7.036307e-06,
  1.655114e-05, 1.737205e-05, 1.748684e-05, 2.517534e-05, 3.863381e-05, 
    1.311886e-05, 1.554461e-06, 9.304638e-07, 3.150416e-06, 5.218887e-06, 
    4.116427e-06, 5.522244e-06, 5.866803e-06, 6.44424e-06, 4.130439e-06,
  1.058778e-05, 5.175309e-05, 0.0001627509, 0.0002982442, 0.0003127486, 
    0.0002417679, 0.0002903953, 0.0002774417, 0.0001977854, 0.0001547897, 
    0.0001350326, 0.0001085621, 5.100346e-05, 2.605495e-05, 7.670177e-06,
  1.263304e-05, 6.835445e-05, 0.0002151908, 0.0004377651, 0.0004106202, 
    0.0002615649, 0.0003424073, 0.0003067884, 0.000229105, 0.0001932639, 
    0.0001738036, 0.0001388013, 3.760941e-05, 7.477152e-06, 7.262294e-06,
  1.894452e-05, 0.0001201216, 0.0003031128, 0.000577151, 0.0004605736, 
    0.0003113528, 0.0003815595, 0.0003316369, 0.0002522393, 0.0002262063, 
    0.0001928899, 9.928314e-05, 1.601347e-05, 5.167647e-06, 7.560502e-06,
  4.883506e-05, 0.0001754393, 0.0003849913, 0.0006818669, 0.0004381794, 
    0.0003546315, 0.0003917856, 0.0003221114, 0.0002605732, 0.0002323477, 
    0.0001826, 5.610046e-05, 5.248455e-06, 5.027035e-06, 7.987634e-06,
  0.0001001454, 0.0002493798, 0.0005116647, 0.0007519273, 0.0004201872, 
    0.0004024621, 0.0004120548, 0.0003175299, 0.0002506094, 0.0002127284, 
    0.0001322112, 1.573437e-05, 2.32618e-06, 4.456968e-06, 8.463078e-06,
  0.000169718, 0.0003844876, 0.0006720802, 0.0007830602, 0.0004243582, 
    0.0004488001, 0.0004157285, 0.0003116269, 0.0002402511, 0.0001801398, 
    7.125841e-05, 1.883733e-07, 9.02062e-07, 4.593366e-06, 1.067873e-05,
  0.0002745276, 0.0005287311, 0.000820356, 0.0007558942, 0.0004365268, 
    0.0004890182, 0.0004193973, 0.0002865349, 0.0002047244, 0.0001266311, 
    1.39913e-05, 7.158049e-08, 1.176721e-06, 6.256828e-06, 8.57376e-06,
  0.0003796178, 0.0006680085, 0.000887882, 0.0006641797, 0.0004948, 
    0.0005009605, 0.0003931003, 0.0002502865, 0.0001508906, 5.680155e-05, 
    2.733762e-08, 3.648084e-07, 1.29845e-06, 5.24282e-06, 7.208207e-06,
  0.0005098426, 0.0007430332, 0.0008560172, 0.000484571, 0.0005232873, 
    0.000486742, 0.0003437201, 0.0001910079, 8.625233e-05, 3.561207e-06, 
    4.315402e-09, 7.557244e-07, 1.180638e-06, 3.619827e-06, 7.452602e-06,
  0.0005573583, 0.0007550335, 0.0007739308, 0.0004899165, 0.0005324666, 
    0.0004314439, 0.0002629166, 0.0001057278, 1.956986e-05, 3.754637e-08, 
    6.854811e-09, 4.835209e-07, 2.008871e-06, 4.015588e-06, 6.038414e-06,
  3.483054e-05, 4.191745e-05, 5.228359e-05, 5.818881e-05, 6.82687e-05, 
    8.115522e-05, 8.699088e-05, 7.940026e-05, 6.400846e-05, 4.995393e-05, 
    3.681307e-05, 3.960668e-05, 6.56776e-05, 8.504985e-05, 5.947825e-05,
  2.798994e-05, 3.734521e-05, 4.71914e-05, 6.635983e-05, 8.408331e-05, 
    8.899804e-05, 9.896994e-05, 9.605212e-05, 9.203175e-05, 6.480033e-05, 
    4.789648e-05, 6.262676e-05, 0.0001142583, 0.0001234459, 7.533305e-05,
  2.701891e-05, 3.224032e-05, 4.36552e-05, 6.460474e-05, 8.784088e-05, 
    8.823808e-05, 8.853614e-05, 8.378419e-05, 9.361786e-05, 8.295979e-05, 
    7.109481e-05, 0.0001110956, 0.0001651247, 0.0001344307, 8.037983e-05,
  2.584255e-05, 3.329704e-05, 4.354951e-05, 6.122737e-05, 6.709342e-05, 
    7.668264e-05, 0.0001188094, 0.0001235058, 0.0001014237, 0.0001156468, 
    0.000106877, 0.0001699257, 0.000175609, 0.0001304227, 6.904826e-05,
  2.487725e-05, 3.127858e-05, 4.481186e-05, 7.284914e-05, 8.054202e-05, 
    0.0001011837, 0.0001181184, 0.0001444459, 0.0001426908, 0.000145373, 
    0.0001707553, 0.0002178491, 0.0001890676, 0.0001366749, 9.222485e-05,
  2.05985e-05, 2.715544e-05, 3.372719e-05, 6.811306e-05, 9.425871e-05, 
    0.0001386171, 0.0001576499, 0.0001747285, 0.0001856485, 0.000196791, 
    0.0002679835, 0.0002469386, 0.0002016758, 0.0001441243, 7.929804e-05,
  1.221952e-05, 1.786038e-05, 3.086633e-05, 6.478256e-05, 0.0001198131, 
    0.0001711983, 0.0002091771, 0.0002018213, 0.0002047465, 0.0003140127, 
    0.0003142706, 0.0002579289, 0.0002158787, 0.000145377, 9.043797e-05,
  1.026563e-05, 1.791259e-05, 3.910452e-05, 7.916444e-05, 0.0001630072, 
    0.0002378487, 0.0002457204, 0.0002139031, 0.0002542516, 0.0003413472, 
    0.0003284925, 0.0002651699, 0.0002158252, 0.0001476318, 8.923593e-05,
  1.913017e-05, 2.050865e-05, 5.104264e-05, 0.000133305, 0.0002582, 
    0.0003104809, 0.0002783117, 0.0002395109, 0.0003084155, 0.0003838753, 
    0.0003394767, 0.0002729406, 0.000206352, 0.0001521248, 9.344452e-05,
  3.369946e-05, 3.877785e-05, 0.0001044808, 0.0002244485, 0.0003609194, 
    0.0003564737, 0.0002891614, 0.0002735648, 0.0003616509, 0.000386364, 
    0.000330278, 0.0002617599, 0.0002120288, 0.0001593808, 9.360656e-05,
  2.410932e-06, 1.975254e-06, 2.095377e-06, 1.727891e-06, 2.312117e-06, 
    1.163249e-06, 8.27646e-07, 1.727901e-07, 6.548005e-08, 1.399071e-07, 
    1.716934e-07, 1.088267e-07, 3.650727e-07, 4.758541e-07, 1.379655e-06,
  2.891198e-06, 2.239511e-06, 2.527956e-06, 2.094076e-06, 2.071114e-06, 
    4.766671e-07, 3.206843e-07, 1.005616e-07, 7.754091e-08, 8.715588e-08, 
    1.219407e-07, 6.098819e-09, 2.817614e-08, 2.348201e-07, 3.42112e-07,
  3.942266e-06, 3.046338e-06, 4.097842e-06, 2.670094e-06, 1.493473e-06, 
    7.168966e-07, 4.111359e-07, 5.468189e-07, 1.98552e-07, 1.553015e-09, 
    7.488532e-09, 3.722852e-08, 9.071059e-10, 1.465227e-08, 4.954018e-08,
  4.378208e-06, 3.812649e-06, 4.060305e-06, 4.384615e-06, 2.449597e-06, 
    1.41653e-06, 1.072165e-06, 1.109242e-06, 3.268032e-07, 1.099102e-07, 
    3.327373e-10, 5.844937e-10, 4.857348e-09, 8.520946e-10, 3.266497e-08,
  8.534882e-06, 5.334585e-06, 4.33182e-06, 5.24611e-06, 2.57317e-06, 
    2.47402e-06, 1.520998e-06, 1.075199e-06, 8.786338e-07, 2.043739e-07, 
    2.126477e-09, 1.88425e-10, 9.50795e-12, 2.854217e-11, 1.749015e-09,
  1.33943e-05, 1.143164e-05, 6.557479e-06, 4.034411e-06, 4.016269e-06, 
    3.597691e-06, 1.814825e-06, 1.338839e-06, 9.627627e-07, 4.83558e-07, 
    3.201738e-08, 2.634406e-09, 5.13365e-10, 3.964993e-10, 2.750804e-10,
  2.773032e-05, 2.002002e-05, 1.398947e-05, 7.171959e-06, 7.669706e-06, 
    4.977459e-06, 2.929033e-06, 1.880532e-06, 1.586235e-06, 6.124425e-07, 
    1.091262e-07, 6.394758e-09, 3.061244e-10, 1.241939e-08, 1.006686e-10,
  4.102349e-05, 3.269892e-05, 1.918383e-05, 1.354616e-05, 2.144748e-05, 
    7.632427e-06, 5.74574e-06, 3.336586e-06, 2.491797e-06, 9.284117e-07, 
    1.94785e-07, 4.852173e-09, 1.415952e-08, 6.599339e-08, 5.12058e-10,
  4.285635e-05, 3.264351e-05, 2.476528e-05, 2.412972e-05, 1.864171e-05, 
    1.303174e-05, 1.018646e-05, 5.66394e-06, 3.100922e-06, 1.726367e-06, 
    5.415919e-07, 1.047261e-07, 2.634353e-07, 5.530968e-08, 2.733781e-08,
  3.280914e-05, 3.432382e-05, 2.658705e-05, 2.883615e-05, 2.646389e-05, 
    2.810205e-05, 2.082887e-05, 1.213265e-05, 6.908946e-06, 3.51798e-06, 
    1.52745e-06, 7.17834e-07, 4.945321e-07, 1.565313e-07, 5.611491e-08,
  0.0003208292, 0.0002323227, 0.0001676517, 0.0001692352, 0.0001310275, 
    0.0001013466, 8.831172e-05, 7.706295e-05, 6.324195e-05, 7.201476e-05, 
    4.100167e-05, 3.261354e-05, 2.492848e-05, 1.909644e-05, 1.422116e-05,
  0.0003416398, 0.0002123334, 0.000195564, 0.000171866, 0.0001514006, 
    0.0001247973, 0.0001107669, 9.890104e-05, 7.547934e-05, 6.683514e-05, 
    6.060763e-05, 3.024027e-05, 2.963054e-05, 2.026091e-05, 1.538982e-05,
  0.0003498432, 0.0002309436, 0.0001960013, 0.0001921367, 0.0001453104, 
    0.0001296591, 0.0001183923, 0.0001037141, 9.232703e-05, 5.470789e-05, 
    6.951064e-05, 2.968176e-05, 3.469531e-05, 1.758975e-05, 1.707691e-05,
  0.0002952447, 0.0002113206, 0.000177026, 0.0001355031, 0.0001411224, 
    0.0001252675, 0.000117782, 0.000102144, 0.0001034028, 6.836046e-05, 
    6.832558e-05, 3.247985e-05, 2.377141e-05, 1.72485e-05, 1.738501e-05,
  0.0002590757, 0.0001890877, 0.000164465, 0.0001480524, 0.0001445535, 
    0.0001237772, 0.0001169154, 0.0001009085, 8.841342e-05, 8.063867e-05, 
    5.482798e-05, 2.91598e-05, 1.423142e-05, 1.528058e-05, 1.329664e-05,
  0.0001996083, 0.000161421, 0.0001466145, 0.0001463694, 0.0001382577, 
    0.000129521, 0.0001145963, 0.0001166115, 9.636261e-05, 8.099665e-05, 
    5.46564e-05, 2.080581e-05, 1.089683e-05, 1.240662e-05, 1.369458e-05,
  0.0001415811, 0.0001439632, 0.0001387396, 0.0001290845, 0.0001205792, 
    0.0001258969, 0.0001165288, 0.0001078071, 9.763656e-05, 6.779428e-05, 
    3.16935e-05, 1.221369e-05, 9.307176e-06, 1.106425e-05, 1.212694e-05,
  0.0001224555, 0.0001246035, 0.0001254561, 0.0001318309, 0.0001162433, 
    0.0001172421, 0.0001124854, 9.182029e-05, 6.502173e-05, 2.65539e-05, 
    1.121225e-05, 1.07131e-05, 9.376192e-06, 8.95879e-06, 9.607029e-06,
  8.438195e-05, 9.907796e-05, 0.0001067307, 0.0001028088, 9.277579e-05, 
    8.9801e-05, 6.673235e-05, 4.776548e-05, 2.337657e-05, 7.765912e-06, 
    8.468312e-06, 7.900567e-06, 9.344204e-06, 9.056829e-06, 8.557608e-06,
  4.059239e-05, 4.960505e-05, 5.334623e-05, 5.12671e-05, 4.42558e-05, 
    3.511424e-05, 2.101501e-05, 1.292005e-05, 7.731924e-06, 6.100212e-06, 
    7.642781e-06, 7.883454e-06, 8.289735e-06, 7.673872e-06, 8.151704e-06,
  8.779206e-07, 5.986411e-09, 1.681424e-09, 6.889723e-09, 4.127262e-09, 
    1.839715e-10, 1.339399e-11, 1.396261e-25, 1.549296e-26, 0, 0, 
    2.133206e-14, 2.513427e-08, 2.66642e-06, 3.805814e-06,
  1.23027e-06, 7.026564e-09, 5.623866e-09, 4.083954e-09, 7.790324e-09, 
    2.749292e-09, 5.171358e-10, 1.097152e-11, 5.46521e-26, 2.084306e-27, 0, 
    4.552361e-11, 9.464687e-07, 4.65741e-06, 4.860263e-06,
  6.634937e-07, 1.428548e-08, 1.07582e-08, 8.570803e-09, 8.443816e-09, 
    3.353423e-08, 2.940847e-09, 6.627415e-10, 4.908672e-12, 2.228712e-26, 
    1.955534e-27, 3.548085e-07, 2.955409e-06, 7.164786e-06, 6.656425e-06,
  9.424797e-08, 8.055147e-09, 1.33231e-08, 1.806836e-08, 9.895479e-09, 
    5.320787e-09, 2.082936e-08, 2.99636e-09, 2.357006e-10, 4.956798e-26, 
    2.153358e-08, 1.916631e-06, 8.09442e-06, 1.806718e-05, 9.778414e-06,
  1.868632e-08, 2.327507e-08, 2.183802e-08, 2.147116e-08, 1.090405e-08, 
    2.704626e-09, 3.771449e-09, 4.19675e-09, 1.336385e-09, 3.971423e-10, 
    1.160427e-06, 1.235624e-05, 1.509491e-05, 1.968959e-05, 1.23503e-05,
  2.077566e-08, 2.745069e-08, 3.721255e-08, 2.553998e-08, 1.602683e-08, 
    8.327347e-09, 3.257881e-09, 3.361674e-10, 6.715914e-09, 2.483761e-06, 
    1.553215e-05, 2.685031e-05, 2.325753e-05, 1.600525e-05, 1.918361e-05,
  2.860932e-08, 1.624148e-07, 4.158165e-08, 3.195649e-08, 1.003354e-07, 
    5.845135e-09, 1.215676e-07, 1.003897e-07, 3.018369e-06, 2.247478e-05, 
    4.324434e-05, 3.768025e-05, 2.39076e-05, 1.692454e-05, 2.16005e-05,
  4.718913e-07, 1.367355e-07, 6.251012e-07, 2.78658e-08, 1.103788e-06, 
    2.501943e-06, 6.983152e-06, 1.338314e-05, 3.993303e-05, 5.630627e-05, 
    5.97493e-05, 4.288779e-05, 2.66546e-05, 2.955403e-05, 1.629527e-05,
  1.369542e-05, 1.651598e-05, 1.797129e-05, 1.531285e-05, 1.913464e-05, 
    2.501469e-05, 3.914754e-05, 5.720729e-05, 6.519452e-05, 7.223528e-05, 
    5.943846e-05, 4.768218e-05, 3.752834e-05, 2.567008e-05, 1.586741e-05,
  6.168673e-05, 6.38511e-05, 6.339719e-05, 7.113405e-05, 7.099388e-05, 
    7.404818e-05, 8.397878e-05, 7.879678e-05, 8.415119e-05, 7.666013e-05, 
    6.208522e-05, 4.841473e-05, 3.199552e-05, 2.805713e-05, 1.738118e-05,
  1.945919e-06, 9.198934e-07, 9.603721e-08, 3.442632e-09, 1.55559e-09, 
    3.517657e-07, 2.329845e-07, 1.900027e-07, 1.486231e-07, 1.475462e-07, 
    2.555437e-09, 5.244285e-09, 7.163439e-10, 6.115702e-10, 1.216799e-09,
  4.028707e-07, 1.538135e-07, 1.986723e-08, 2.938897e-10, 3.013838e-10, 
    2.306763e-08, 3.600166e-08, 1.16916e-07, 1.719819e-08, 3.542487e-10, 
    2.062968e-10, 8.905934e-10, 6.360468e-11, 9.063091e-11, 8.081618e-10,
  2.924475e-07, 6.821238e-08, 1.649226e-09, 4.084719e-11, 7.068551e-08, 
    2.890898e-09, 1.04087e-08, 2.40995e-09, 3.213771e-08, 1.601325e-11, 
    1.173311e-11, 3.89363e-11, 4.158009e-11, 3.445546e-10, 1.115772e-10,
  1.788425e-07, 2.042498e-08, 2.45683e-11, 1.213703e-10, 7.528326e-09, 
    1.326594e-09, 2.822643e-09, 7.766637e-10, 1.315793e-10, 5.974851e-15, 
    2.115724e-15, 1.812449e-16, 6.87729e-14, 1.915616e-11, 1.574168e-10,
  9.237733e-08, 3.376424e-09, 1.97529e-10, 7.851232e-10, 1.312045e-09, 
    7.573901e-10, 2.706247e-09, 4.098543e-11, 1.959569e-11, 2.125384e-16, 
    5.456197e-16, 3.476746e-18, 3.812143e-17, 9.718616e-12, 1.235369e-10,
  9.740793e-09, 2.137475e-09, 1.094866e-09, 7.005543e-09, 6.081192e-09, 
    4.579393e-09, 1.557822e-09, 4.235171e-09, 9.734322e-11, 3.41674e-12, 
    2.652099e-12, 4.549422e-23, 3.087695e-23, 1.459163e-12, 5.037198e-12,
  9.788601e-09, 1.549493e-08, 2.096066e-08, 2.794284e-08, 2.336967e-08, 
    1.266275e-08, 3.444909e-09, 5.818336e-09, 6.713036e-09, 3.40706e-09, 
    6.130678e-11, 2.952762e-23, 1.82175e-23, 1.120872e-23, 3.204896e-24,
  2.011009e-08, 3.011419e-08, 4.851306e-08, 7.224347e-08, 5.734605e-08, 
    4.906649e-08, 2.465534e-08, 7.921937e-08, 1.52898e-08, 5.412723e-10, 
    7.813073e-10, 1.422816e-11, 1.385305e-23, 5.337144e-24, 1.264238e-24,
  3.578062e-08, 4.211993e-08, 8.404761e-08, 9.886885e-08, 7.185023e-08, 
    2.596669e-08, 2.019373e-08, 1.528301e-08, 7.565059e-09, 6.35248e-10, 
    8.384858e-10, 6.131329e-11, 2.124667e-11, 2.048351e-13, 2.891738e-24,
  4.730142e-08, 7.041365e-08, 1.259731e-07, 1.259969e-07, 8.076953e-08, 
    3.616738e-08, 2.19266e-08, 1.605697e-08, 7.628612e-09, 8.740406e-10, 
    1.129934e-09, 2.627337e-10, 3.742046e-10, 2.160325e-11, 1.127087e-12,
  0.0001123455, 0.0001548528, 0.0001989381, 0.0002182679, 0.0001808538, 
    0.0001200518, 9.986755e-05, 9.202537e-05, 7.352795e-05, 6.736146e-05, 
    5.859098e-05, 4.165094e-05, 2.687465e-05, 3.378875e-05, 2.892784e-05,
  0.0001211949, 0.0001648925, 0.0002106174, 0.0001916454, 0.0001499635, 
    0.0001112212, 0.0001730592, 0.000107247, 7.865003e-05, 8.143948e-05, 
    6.879192e-05, 5.254298e-05, 3.37611e-05, 3.183193e-05, 2.952664e-05,
  0.0001621099, 0.0002013068, 0.0002325964, 0.0001995682, 0.000188249, 
    0.0001555742, 9.651032e-05, 0.0001181228, 9.39708e-05, 9.047556e-05, 
    7.988816e-05, 7.765552e-05, 6.433221e-05, 4.728182e-05, 3.35903e-05,
  0.0002133801, 0.0002456246, 0.0002535696, 0.0002230637, 0.0002460296, 
    0.0001850589, 0.000147248, 0.0001425464, 0.0001085326, 0.0001067814, 
    8.12987e-05, 8.92464e-05, 7.779381e-05, 5.622312e-05, 2.080593e-05,
  0.0002663177, 0.0002683182, 0.0002676972, 0.0002239164, 0.0002124176, 
    0.0001968038, 0.0001576685, 9.161672e-05, 0.0001375956, 0.0001251308, 
    0.000107235, 9.174481e-05, 8.415205e-05, 4.10774e-05, 1.015272e-05,
  0.000293963, 0.0002919738, 0.0002951929, 0.0002408509, 0.0002273277, 
    0.00023043, 0.0001687098, 0.0001237315, 0.0001060622, 0.0001302661, 
    0.0001329654, 8.718474e-05, 6.808277e-05, 4.60217e-05, 5.470018e-06,
  0.0003057188, 0.0002976113, 0.000297174, 0.000260702, 0.0002676929, 
    0.000247728, 0.0001741608, 0.0001355285, 0.0001574954, 0.0001151381, 
    0.0001203543, 9.075163e-05, 4.585973e-05, 1.130234e-05, 5.144814e-06,
  0.0003024887, 0.0003075755, 0.000278979, 0.0002618042, 0.000274892, 
    0.000244113, 0.0001783722, 0.0001546869, 0.0001344631, 0.000139162, 
    0.0001363774, 6.48768e-05, 1.519623e-05, 4.046589e-06, 4.196548e-06,
  0.0003206203, 0.0002790074, 0.0002565534, 0.0002646348, 0.0002749107, 
    0.0002165333, 0.0001671757, 0.0001698921, 0.0001636326, 0.0001247479, 
    8.358435e-05, 2.728874e-05, 2.547866e-06, 3.052074e-06, 4.758511e-06,
  0.0002804184, 0.0002503725, 0.0002424989, 0.0002555607, 0.0002465429, 
    0.0001883639, 0.0001783899, 0.0001714013, 0.0001381847, 0.0001085832, 
    2.863156e-05, 3.915926e-06, 2.188378e-06, 3.101843e-06, 6.085475e-06,
  1.293021e-05, 1.227364e-05, 9.127548e-06, 6.750297e-06, 2.672248e-06, 
    2.618186e-06, 1.834347e-06, 1.302357e-06, 8.699967e-07, 3.446708e-07, 
    1.63422e-07, 2.333089e-11, 2.233774e-08, 3.099355e-07, 4.303987e-06,
  1.302202e-05, 1.182391e-05, 1.052743e-05, 6.34456e-06, 4.904772e-06, 
    4.218061e-06, 3.395463e-06, 2.442112e-06, 1.124273e-06, 3.720381e-07, 
    1.131994e-07, 1.849698e-10, 1.392263e-10, 6.558156e-07, 1.017138e-05,
  1.806777e-05, 1.508865e-05, 1.219701e-05, 9.995601e-06, 1.079991e-05, 
    7.263945e-06, 5.824851e-06, 3.896941e-06, 1.890707e-06, 6.618265e-07, 
    1.644037e-07, 5.841611e-10, 1.50455e-08, 3.85047e-06, 1.991418e-05,
  2.156437e-05, 1.797506e-05, 1.201686e-05, 1.210122e-05, 1.098753e-05, 
    1.101813e-05, 1.048449e-05, 6.357486e-06, 4.337264e-06, 1.430333e-06, 
    4.398158e-07, 7.0804e-08, 4.629921e-07, 1.084921e-05, 5.485912e-05,
  3.627894e-05, 1.823573e-05, 1.107516e-05, 9.951889e-06, 1.138504e-05, 
    2.872055e-05, 2.586821e-05, 1.191331e-05, 5.514238e-06, 2.955304e-06, 
    9.319307e-07, 3.884065e-07, 2.88036e-06, 2.638709e-05, 6.834231e-05,
  4.243181e-05, 2.126691e-05, 1.405325e-05, 9.388556e-06, 1.238642e-05, 
    2.677183e-05, 4.360617e-05, 1.693436e-05, 1.332333e-05, 4.519389e-06, 
    1.350968e-06, 1.027622e-06, 1.598265e-05, 4.525198e-05, 6.531423e-05,
  5.468079e-05, 2.722286e-05, 1.671054e-05, 1.107395e-05, 1.550354e-05, 
    4.477333e-05, 4.41576e-05, 3.363072e-05, 1.232059e-05, 5.499966e-06, 
    2.168923e-06, 7.854856e-06, 4.650494e-05, 7.075399e-05, 8.077628e-05,
  5.499714e-05, 3.884475e-05, 1.969811e-05, 1.387254e-05, 1.642336e-05, 
    4.939433e-05, 7.519831e-05, 4.609432e-05, 1.345286e-05, 4.913145e-06, 
    1.381886e-05, 3.920234e-05, 8.512677e-05, 9.429705e-05, 8.547336e-05,
  4.183064e-05, 4.773651e-05, 2.264145e-05, 1.80726e-05, 1.817746e-05, 
    7.460912e-05, 9.663392e-05, 7.911164e-05, 2.6565e-05, 3.197595e-05, 
    5.843583e-05, 9.086775e-05, 0.0001076947, 0.0001051552, 9.021574e-05,
  2.039109e-05, 2.949737e-05, 1.574366e-05, 1.233182e-05, 1.861175e-05, 
    4.539072e-05, 9.248009e-05, 8.592393e-05, 7.259345e-05, 8.134075e-05, 
    0.0001210238, 0.0001283002, 0.000118218, 0.0001077218, 0.000100339,
  3.36471e-05, 1.903509e-05, 3.416284e-05, 0.0001096471, 0.0001435768, 
    0.0001066523, 6.753797e-05, 4.754804e-05, 3.194415e-05, 1.966445e-05, 
    1.815754e-05, 1.81224e-05, 2.874014e-05, 3.524143e-05, 2.135865e-05,
  1.150156e-05, 5.060776e-05, 0.0001126744, 0.0001659745, 0.0001486135, 
    9.038251e-05, 4.616949e-05, 3.105549e-05, 1.981924e-05, 1.458654e-05, 
    2.311849e-05, 2.436879e-05, 2.404944e-05, 2.231369e-05, 1.796223e-05,
  1.416551e-05, 0.00010191, 0.0001470061, 0.0001553638, 0.0001014295, 
    4.395128e-05, 1.61078e-05, 9.324476e-06, 1.347192e-05, 2.028881e-05, 
    1.714486e-05, 2.833051e-05, 2.777526e-05, 2.620847e-05, 1.76412e-05,
  2.910979e-05, 8.765743e-05, 0.0001070658, 8.616095e-05, 3.378489e-05, 
    6.115024e-06, 5.193144e-06, 5.361356e-06, 5.482911e-06, 1.303014e-05, 
    1.857374e-05, 1.625774e-05, 1.482533e-05, 2.489785e-05, 1.793193e-05,
  1.284137e-05, 3.271407e-05, 3.669451e-05, 1.982338e-05, 4.11108e-06, 
    3.797752e-06, 5.092085e-06, 6.464739e-06, 4.701272e-06, 2.51149e-06, 
    5.20699e-06, 1.400325e-05, 1.168241e-05, 1.470769e-05, 1.435304e-05,
  1.018081e-06, 2.110057e-06, 4.236215e-06, 3.090116e-06, 2.612696e-06, 
    3.290085e-06, 3.780633e-06, 5.544408e-06, 4.612757e-06, 2.118592e-06, 
    2.675745e-06, 6.908394e-06, 5.769336e-06, 9.830052e-06, 7.701297e-06,
  3.413134e-07, 4.291091e-07, 1.174487e-06, 1.512331e-06, 1.632011e-06, 
    1.840034e-06, 3.572589e-06, 4.234172e-06, 2.723179e-06, 1.358888e-06, 
    1.207479e-06, 1.463588e-06, 2.731678e-06, 6.250389e-06, 3.657895e-06,
  4.079058e-07, 2.87896e-07, 5.625612e-07, 8.996527e-07, 1.649242e-06, 
    9.59544e-07, 3.358441e-06, 2.615237e-06, 2.036859e-06, 1.47798e-06, 
    1.121387e-06, 1.289178e-06, 8.237088e-07, 2.11658e-06, 1.40251e-06,
  2.018132e-07, 3.788068e-07, 3.656871e-07, 4.699425e-07, 9.483005e-07, 
    2.11039e-06, 1.102881e-06, 1.699331e-06, 1.127792e-06, 1.329419e-06, 
    1.834622e-06, 1.200601e-06, 2.486585e-07, 2.058977e-07, 8.439109e-07,
  2.743419e-07, 3.58595e-07, 2.726859e-07, 3.331342e-07, 5.873745e-07, 
    7.098753e-07, 4.641308e-07, 5.674353e-07, 9.298529e-07, 6.338943e-07, 
    9.898559e-07, 8.090539e-07, 4.976216e-08, 1.918594e-07, 5.808295e-07,
  1.216609e-05, 7.916062e-06, 1.186416e-05, 3.367983e-05, 4.163066e-05, 
    3.529699e-05, 6.761496e-05, 5.993843e-05, 9.75953e-05, 8.401737e-05, 
    5.330686e-05, 2.384572e-05, 7.248763e-05, 9.602492e-05, 6.133023e-05,
  1.776686e-05, 5.636575e-06, 2.178449e-05, 5.089519e-05, 5.731528e-05, 
    5.012231e-05, 7.561431e-05, 0.0001019786, 0.000100509, 8.332147e-05, 
    7.537689e-05, 1.398048e-05, 4.612745e-06, 4.279144e-05, 6.436726e-05,
  2.563172e-05, 3.895073e-05, 7.735132e-05, 0.000111405, 0.000112789, 
    0.0001053695, 0.0001381945, 0.0001562771, 0.0001187302, 0.0001049484, 
    0.0001877965, 1.310233e-05, 2.214006e-07, 2.817081e-05, 4.3023e-05,
  7.743345e-05, 0.0001224509, 0.0001787783, 0.0001828529, 0.0001699602, 
    0.0001621159, 0.0001938817, 0.0001958604, 0.0001694196, 0.0001545482, 
    9.874986e-05, 1.741723e-05, 4.802248e-06, 3.569046e-05, 3.43464e-05,
  0.0001524633, 0.0002214904, 0.0002554532, 0.0002417926, 0.0001889383, 
    0.0001823232, 0.0002199151, 0.0002332242, 0.0002019839, 0.0001752332, 
    0.0001456747, 1.814504e-05, 6.169769e-06, 2.778052e-05, 1.846198e-05,
  0.0002259995, 0.0002991703, 0.0002875572, 0.0002368605, 0.0001870137, 
    0.0001957007, 0.0002659927, 0.0002718129, 0.0002276711, 0.000200332, 
    0.00015508, 2.179909e-05, 1.436394e-05, 3.542291e-05, 2.344817e-05,
  0.0003022793, 0.0003302463, 0.0003192046, 0.0002301861, 0.0001937319, 
    0.000217736, 0.0002912358, 0.0002917056, 0.0002540892, 0.0002397989, 
    0.0001571459, 1.241771e-05, 3.357662e-05, 2.82188e-05, 1.718384e-05,
  0.0003423033, 0.0003652134, 0.0003479236, 0.000268922, 0.0002034888, 
    0.0002332402, 0.0003196655, 0.000290957, 0.0002751922, 0.0002750313, 
    0.0001414459, 6.475845e-06, 9.177677e-06, 2.187542e-05, 1.487784e-05,
  0.000339643, 0.0003561297, 0.0003595916, 0.0002908531, 0.0002399722, 
    0.0002657639, 0.0003043696, 0.000272694, 0.0002814451, 0.0003019477, 
    0.0001202469, 2.463719e-07, 1.194585e-05, 1.572277e-05, 1.101224e-05,
  0.0003187781, 0.0003430373, 0.0003517225, 0.0003113819, 0.0002730082, 
    0.0002996855, 0.0002979218, 0.00025353, 0.0003101348, 0.0002926696, 
    8.877416e-05, 4.664397e-07, 9.230494e-06, 1.348322e-05, 1.039625e-05,
  0.0001445197, 0.0001413376, 0.0001576437, 0.0001620745, 0.0001616171, 
    0.0001605894, 0.0001633134, 0.0001725445, 0.0001756752, 0.0001788973, 
    0.0001773981, 0.0001547368, 9.063727e-05, 3.19825e-05, 2.979429e-06,
  0.0001729968, 0.0001907327, 0.0002074262, 0.0002097027, 0.0001956446, 
    0.0001970621, 0.0002034205, 0.0002028715, 0.0002084524, 0.0002157277, 
    0.000210262, 0.000120916, 3.697695e-05, 1.20058e-05, 5.611539e-06,
  0.0002308076, 0.0002309893, 0.0002223664, 0.0002166956, 0.0002218067, 
    0.0002175123, 0.0002287798, 0.0002363987, 0.0002381513, 0.0002265324, 
    0.0001397015, 5.010216e-05, 1.041011e-05, 6.130941e-07, 7.066502e-06,
  0.0002362841, 0.0002292348, 0.0002089069, 0.0001978922, 0.0002114258, 
    0.0002136431, 0.0002171815, 0.0002296554, 0.0001967985, 0.0001142468, 
    3.652131e-05, 2.70135e-06, 7.671155e-07, 2.309604e-07, 4.343345e-06,
  0.0002199762, 0.0001967409, 0.0001890817, 0.0001908936, 0.000195456, 
    0.000218983, 0.0002127008, 0.0001570697, 8.137269e-05, 1.512255e-05, 
    6.759669e-06, 4.956919e-06, 5.54693e-07, 3.615452e-07, 4.884966e-06,
  0.0002065032, 0.0001789658, 0.0001880301, 0.0001733405, 0.0001810805, 
    0.0001561421, 0.0001196809, 5.085687e-05, 4.140735e-06, 2.229287e-06, 
    9.365803e-06, 7.489178e-06, 7.920405e-07, 4.118677e-07, 7.160573e-08,
  0.0001334583, 0.0001273459, 0.0001408445, 0.0001296225, 9.499118e-05, 
    5.650687e-05, 1.753485e-05, 3.903309e-06, 3.102383e-06, 2.812457e-06, 
    1.366546e-05, 1.200324e-05, 4.497439e-07, 3.496291e-07, 8.154234e-07,
  2.921642e-05, 3.727962e-05, 4.449835e-05, 3.288653e-05, 1.224701e-05, 
    3.464842e-06, 2.686412e-06, 4.075934e-06, 3.505889e-06, 3.75803e-06, 
    2.449054e-05, 1.802041e-05, 7.720207e-07, 4.530599e-07, 2.324051e-07,
  1.746239e-06, 2.442265e-06, 3.607453e-06, 3.095597e-06, 3.108432e-06, 
    4.216933e-06, 3.950323e-06, 3.709146e-06, 7.845807e-06, 1.40053e-05, 
    3.943165e-05, 2.124734e-05, 2.720452e-07, 2.042111e-07, 7.773244e-08,
  1.926633e-06, 1.724431e-06, 2.854775e-06, 3.552185e-06, 3.929346e-06, 
    4.32962e-06, 3.317858e-06, 3.065965e-06, 1.860126e-05, 4.710486e-05, 
    6.21576e-05, 2.308295e-05, 1.185896e-07, 5.629596e-08, 2.756238e-07,
  4.544241e-05, 4.378969e-05, 4.197023e-05, 3.799065e-05, 4.199429e-05, 
    2.73099e-05, 2.268661e-05, 9.908073e-06, 3.675192e-06, 2.37386e-06, 
    1.782897e-06, 1.22654e-05, 6.570104e-05, 0.0001023123, 0.0001039272,
  4.592523e-05, 4.899991e-05, 5.27801e-05, 6.141301e-05, 7.92205e-05, 
    5.642431e-05, 2.116337e-05, 1.257409e-05, 7.159588e-06, 4.618665e-06, 
    1.996451e-05, 7.809007e-05, 0.0001414734, 0.0001351286, 8.322797e-05,
  4.135817e-05, 3.937523e-05, 3.982074e-05, 8.466017e-05, 6.622002e-05, 
    4.063756e-05, 1.844741e-05, 1.182589e-05, 6.288073e-06, 2.290489e-05, 
    9.493165e-05, 0.0001704019, 0.0001849977, 0.0001416333, 9.321483e-05,
  3.738488e-05, 3.26217e-05, 5.858596e-05, 6.143231e-05, 6.309109e-05, 
    3.367645e-05, 1.868988e-05, 9.758031e-06, 4.166119e-05, 0.0001246633, 
    0.0002028199, 0.0002157849, 0.0001901579, 0.0001269749, 7.481897e-05,
  3.58448e-05, 3.532811e-05, 6.433126e-05, 0.0001063447, 5.291426e-05, 
    2.357515e-05, 2.087522e-05, 7.575299e-05, 0.0001646061, 0.000236115, 
    0.0002438588, 0.0002176257, 0.0001806678, 0.0001124098, 9.168994e-05,
  3.938746e-05, 3.343071e-05, 5.40227e-05, 7.017129e-05, 5.804269e-05, 
    5.799943e-05, 0.0001214212, 0.0001930279, 0.0002524822, 0.0002494247, 
    0.0002419735, 0.0002295995, 0.0001619945, 0.0001121098, 0.0001090037,
  0.0001310275, 7.667548e-05, 0.0001416148, 0.0001253321, 0.000123465, 
    0.0001662971, 0.0002214287, 0.0002587205, 0.0002607802, 0.0002589262, 
    0.0002603747, 0.0002239934, 0.0001574559, 0.0001241386, 0.0001337547,
  0.0002166971, 0.0002122369, 0.0002294541, 0.0001880204, 0.0002100518, 
    0.0002353131, 0.0002526893, 0.0002709336, 0.0002714718, 0.0002900846, 
    0.0002710077, 0.0002106421, 0.0001559581, 0.0001378188, 0.0001473398,
  0.0002812123, 0.0002576925, 0.0002244717, 0.0002303131, 0.0002492473, 
    0.0002828347, 0.0002984197, 0.0003040465, 0.0003118326, 0.0002989387, 
    0.0002498583, 0.0001964947, 0.0001541569, 0.0001462382, 0.0001624424,
  0.0003242897, 0.0002269715, 0.0002461741, 0.0002796576, 0.0003136975, 
    0.0003381891, 0.0003396261, 0.0003296373, 0.0003029596, 0.0002768471, 
    0.0002326209, 0.0001963074, 0.0001726994, 0.0001659739, 0.0002043407,
  0.000128735, 0.0001603148, 0.0001866328, 0.0001548491, 0.0001252607, 
    0.0001160924, 0.0001117728, 4.750106e-05, 3.8877e-05, 2.596818e-05, 
    1.644023e-05, 3.619791e-06, 8.161694e-06, 3.641235e-06, 9.324484e-06,
  0.000142595, 0.0002023728, 0.0001520407, 0.0001399539, 0.0001361062, 
    9.731652e-05, 5.955891e-05, 3.524976e-05, 2.123824e-05, 1.595911e-05, 
    8.572907e-06, 2.435727e-06, 4.145439e-06, 6.030969e-06, 1.760026e-06,
  0.0001242162, 0.0001670921, 0.000156299, 0.0001155568, 9.846775e-05, 
    6.712082e-05, 3.81677e-05, 1.981868e-05, 2.125826e-05, 1.594217e-05, 
    8.042823e-06, 3.419915e-06, 2.677526e-06, 6.080936e-06, 2.247791e-06,
  7.216573e-05, 7.640894e-05, 7.057426e-05, 6.22461e-05, 5.246144e-05, 
    3.885339e-05, 2.654883e-05, 1.783323e-05, 1.879809e-05, 1.541299e-05, 
    5.779101e-06, 3.565782e-06, 3.551012e-06, 1.276383e-05, 1.426658e-06,
  1.936886e-05, 2.232845e-05, 2.251053e-05, 1.639018e-05, 1.231085e-05, 
    1.120404e-05, 1.044255e-05, 1.136934e-05, 1.418674e-05, 1.135557e-05, 
    4.868788e-06, 2.77079e-06, 3.87486e-06, 4.750528e-06, 1.735354e-06,
  5.421145e-06, 2.54676e-06, 2.829844e-06, 3.573964e-06, 4.076186e-06, 
    5.077293e-06, 7.383108e-06, 8.635849e-06, 1.024375e-05, 8.680729e-06, 
    4.144038e-06, 2.927669e-06, 2.120139e-06, 1.237025e-06, 2.79669e-06,
  5.406645e-06, 3.198924e-06, 1.398037e-06, 2.190478e-06, 3.396383e-06, 
    5.810029e-06, 6.525219e-06, 8.513559e-06, 8.902231e-06, 7.808342e-06, 
    2.820125e-06, 1.975268e-06, 6.170227e-07, 3.307151e-07, 3.099361e-06,
  6.921871e-06, 3.343333e-06, 1.952415e-06, 2.051799e-06, 3.298555e-06, 
    5.202995e-06, 7.837752e-06, 8.190955e-06, 9.100627e-06, 7.034961e-06, 
    3.494395e-06, 5.591609e-07, 4.645358e-07, 1.520115e-07, 3.89051e-06,
  8.09127e-06, 4.317249e-06, 2.45618e-06, 2.316866e-06, 2.371551e-06, 
    3.893547e-06, 6.051647e-06, 7.690384e-06, 6.620427e-06, 5.564838e-06, 
    2.42028e-06, 6.066799e-07, 3.779625e-07, 1.882883e-07, 7.927165e-06,
  1.454851e-05, 7.531284e-06, 3.686323e-06, 2.556247e-06, 1.14033e-06, 
    1.933967e-06, 3.274892e-06, 5.682851e-06, 5.273815e-06, 3.884849e-06, 
    2.328986e-06, 5.493346e-07, 2.094087e-07, 1.068236e-06, 1.586586e-05,
  3.224473e-08, 1.498475e-08, 3.259399e-09, 3.401874e-09, 1.26935e-08, 
    1.286498e-05, 1.42466e-05, 2.645006e-05, 4.333918e-05, 7.734323e-05, 
    8.142099e-05, 5.776104e-05, 3.023689e-05, 1.830053e-05, 1.445979e-05,
  3.005345e-07, 1.610597e-07, 2.526447e-07, 4.476283e-06, 5.228118e-07, 
    1.91508e-05, 2.849668e-05, 5.356976e-05, 5.68255e-05, 6.017179e-05, 
    6.473478e-05, 4.421575e-05, 3.231002e-05, 5.015615e-06, 1.630757e-05,
  1.409292e-05, 2.096671e-05, 2.060064e-05, 2.646962e-05, 4.10463e-05, 
    5.107792e-05, 5.160283e-05, 5.796998e-05, 6.301443e-05, 4.767516e-05, 
    4.621881e-05, 4.715391e-05, 1.558917e-05, 2.00191e-05, 2.546482e-05,
  7.602395e-05, 8.275002e-05, 8.980091e-05, 8.060643e-05, 9.335362e-05, 
    0.000107253, 6.183292e-05, 7.334172e-05, 6.413607e-05, 4.391391e-05, 
    5.929951e-05, 4.087459e-05, 4.649363e-05, 5.31719e-05, 5.420092e-05,
  0.0001359857, 0.000143658, 0.0001300939, 0.0001122955, 9.659356e-05, 
    7.873818e-05, 0.0001137239, 8.953269e-05, 7.734129e-05, 5.847901e-05, 
    3.901937e-05, 8.722526e-05, 5.803327e-05, 6.071584e-05, 6.755813e-05,
  0.0001540722, 0.000172374, 0.0001591365, 0.0001231707, 9.485313e-05, 
    0.0001031812, 9.845091e-05, 9.784653e-05, 7.197436e-05, 5.730585e-05, 
    5.360056e-05, 6.825375e-05, 8.474341e-05, 7.231213e-05, 5.421673e-05,
  0.0001576728, 0.0001613367, 0.0001488689, 0.0001239089, 9.458313e-05, 
    8.862594e-05, 8.097103e-05, 9.802457e-05, 7.67723e-05, 6.724082e-05, 
    6.112731e-05, 0.0001190356, 0.0001178521, 8.26843e-05, 6.757955e-05,
  0.0001444603, 0.0001500674, 0.0001391859, 0.0001204638, 9.104926e-05, 
    7.564585e-05, 0.0001084519, 7.683766e-05, 0.0001063986, 8.202836e-05, 
    9.788132e-05, 0.0001075302, 0.0001137743, 9.579203e-05, 7.344539e-05,
  0.0001324683, 0.0001422764, 0.0001260233, 0.0001057653, 8.360662e-05, 
    7.649319e-05, 8.584918e-05, 0.0001016139, 0.000135117, 0.0001064559, 
    7.749521e-05, 9.316771e-05, 0.0001114596, 9.310116e-05, 5.912624e-05,
  0.0001295633, 0.0001395446, 0.0001168119, 9.670096e-05, 7.257899e-05, 
    6.183828e-05, 6.694182e-05, 0.0001021259, 0.0001209624, 8.403061e-05, 
    8.636684e-05, 9.50695e-05, 0.0001070511, 0.0001105901, 6.641203e-05,
  3.704117e-05, 3.828523e-05, 4.082955e-05, 4.238574e-05, 4.169584e-05, 
    4.385409e-05, 6.426147e-05, 3.816649e-05, 2.777944e-05, 3.43334e-05, 
    2.376819e-05, 1.285635e-05, 8.12276e-06, 6.786378e-06, 3.54436e-06,
  3.287597e-05, 3.001039e-05, 3.23254e-05, 3.197919e-05, 2.504677e-05, 
    2.418221e-05, 3.270133e-05, 3.849603e-05, 4.982336e-05, 3.028906e-05, 
    2.602223e-05, 1.481099e-05, 1.424932e-05, 7.102072e-06, 3.671226e-06,
  3.941502e-05, 3.830463e-05, 3.782458e-05, 3.699536e-05, 3.790098e-05, 
    4.020441e-05, 3.325906e-05, 3.763573e-05, 3.606594e-05, 5.144768e-05, 
    3.828069e-05, 3.717204e-05, 2.357813e-05, 1.289967e-05, 4.589113e-06,
  4.474304e-05, 4.448702e-05, 4.248153e-05, 4.735342e-05, 4.2876e-05, 
    4.17678e-05, 3.621854e-05, 3.569797e-05, 3.71389e-05, 5.383475e-05, 
    5.113264e-05, 3.900354e-05, 2.336628e-05, 9.583278e-06, 3.139207e-06,
  4.820126e-05, 5.302809e-05, 5.499935e-05, 5.139475e-05, 4.954983e-05, 
    4.076613e-05, 3.81017e-05, 3.163873e-05, 2.308618e-05, 1.868809e-05, 
    2.82911e-05, 3.168844e-05, 1.958464e-05, 1.107943e-05, 3.177713e-06,
  6.03542e-05, 6.066799e-05, 6.33442e-05, 5.806179e-05, 5.568436e-05, 
    4.436983e-05, 3.500551e-05, 3.180548e-05, 1.949008e-05, 1.420169e-05, 
    2.031588e-05, 3.638075e-05, 2.012591e-05, 7.58027e-06, 1.68231e-06,
  6.429786e-05, 6.44593e-05, 7.165404e-05, 6.784739e-05, 5.819868e-05, 
    4.926976e-05, 3.560476e-05, 2.730636e-05, 1.306063e-05, 2.94427e-06, 
    9.74341e-06, 1.097167e-05, 8.983067e-06, 3.910699e-06, 5.042174e-07,
  6.870868e-05, 7.259511e-05, 7.535695e-05, 8.17974e-05, 7.711342e-05, 
    5.829602e-05, 4.210329e-05, 2.693546e-05, 1.149172e-05, 1.802644e-06, 
    1.563939e-06, 3.498492e-06, 2.511383e-06, 1.68629e-06, 2.361629e-07,
  6.236034e-05, 6.414804e-05, 7.89343e-05, 8.712277e-05, 8.787106e-05, 
    7.00968e-05, 5.180009e-05, 3.175853e-05, 1.149451e-05, 1.391879e-06, 
    4.894742e-09, 8.35326e-07, 2.819505e-07, 3.262551e-07, 5.864413e-08,
  4.736514e-05, 5.517777e-05, 6.47882e-05, 7.575213e-05, 8.153851e-05, 
    7.776848e-05, 6.429333e-05, 4.161175e-05, 1.299289e-05, 5.939565e-07, 
    1.353205e-09, 3.745612e-10, 1.495037e-09, 2.511827e-09, 1.414965e-09,
  3.20713e-05, 3.898911e-05, 3.814795e-05, 2.384446e-05, 1.439825e-05, 
    5.957112e-05, 0.0001130814, 8.575232e-05, 4.850832e-05, 0.0001004723, 
    1.373041e-05, 5.943075e-06, 7.827726e-06, 8.531502e-06, 6.320638e-06,
  5.497697e-05, 3.969314e-05, 4.480322e-05, 3.030088e-05, 1.280725e-05, 
    2.255565e-05, 0.0001141891, 9.548373e-05, 4.353114e-05, 5.307375e-05, 
    1.139211e-05, 5.947266e-06, 1.177084e-05, 7.890163e-06, 6.522178e-06,
  7.992772e-05, 5.31797e-05, 5.189966e-05, 4.20497e-05, 1.843605e-05, 
    2.033344e-05, 9.688444e-05, 0.0001121765, 4.947732e-05, 4.061748e-05, 
    1.854119e-05, 1.690904e-05, 1.46582e-05, 1.056406e-05, 7.131279e-06,
  0.0001020317, 7.187043e-05, 6.912054e-05, 5.367752e-05, 3.178939e-05, 
    1.652086e-05, 8.63581e-05, 0.0001387971, 7.199917e-05, 3.174039e-05, 
    2.615374e-05, 1.106726e-05, 1.417237e-05, 1.302095e-05, 7.357947e-06,
  9.832153e-05, 8.415798e-05, 9.861544e-05, 6.671971e-05, 4.854742e-05, 
    2.126782e-05, 6.35774e-05, 0.0001556018, 9.269339e-05, 1.197462e-05, 
    1.612871e-05, 8.188971e-06, 1.410312e-05, 1.361108e-05, 9.904159e-06,
  8.092014e-05, 9.00996e-05, 0.0001006254, 8.02908e-05, 4.728034e-05, 
    1.767754e-05, 4.42801e-05, 0.0001571324, 0.0001158681, 2.183485e-05, 
    6.789343e-06, 1.121926e-05, 1.217898e-05, 1.030094e-05, 8.180678e-06,
  6.484969e-05, 8.739272e-05, 0.0001128351, 9.063395e-05, 5.196449e-05, 
    1.871583e-05, 2.430469e-05, 0.0001550305, 0.0001347457, 3.694161e-05, 
    7.611183e-06, 6.134528e-06, 1.49359e-05, 1.195093e-05, 1.154038e-05,
  4.392025e-05, 8.918036e-05, 0.0001160003, 0.0001115421, 6.283325e-05, 
    2.349191e-05, 3.808257e-05, 0.0001474669, 0.0001485868, 4.510643e-05, 
    9.241437e-06, 1.464634e-05, 9.720975e-06, 1.232099e-05, 1.21353e-05,
  3.720077e-05, 8.671916e-05, 0.000123375, 0.0001023131, 7.226757e-05, 
    2.866453e-05, 2.464648e-05, 0.0001386989, 0.0001602311, 6.135058e-05, 
    1.965262e-05, 7.661812e-06, 1.143164e-05, 1.138962e-05, 9.261019e-06,
  4.777631e-05, 7.417934e-05, 0.0001201303, 0.0001010252, 7.807215e-05, 
    4.051622e-05, 3.0247e-05, 0.0001354156, 0.000150846, 6.690482e-05, 
    2.340407e-05, 1.295053e-05, 8.473615e-06, 8.296657e-06, 6.746362e-06,
  0.0001274559, 0.0001433243, 0.0001418772, 9.434287e-05, 7.478757e-05, 
    7.099463e-05, 0.0001116017, 9.894716e-05, 7.159497e-05, 6.711702e-05, 
    7.18567e-05, 5.76454e-05, 4.138262e-05, 2.98154e-05, 2.175865e-05,
  0.0001633396, 0.0001069831, 0.0001304206, 0.0001065117, 7.687207e-05, 
    7.479422e-05, 7.881416e-05, 9.473314e-05, 7.839245e-05, 9.046645e-05, 
    5.406379e-05, 4.048297e-05, 3.222596e-05, 2.813678e-05, 1.794922e-05,
  0.0001294411, 0.0001228007, 0.0001502095, 0.0001240314, 7.750271e-05, 
    7.423828e-05, 8.972978e-05, 7.855168e-05, 9.062062e-05, 6.745038e-05, 
    5.053623e-05, 4.344918e-05, 2.889921e-05, 1.950301e-05, 3.992384e-05,
  0.0001348574, 0.0001203053, 0.0001378728, 0.0001120141, 7.050818e-05, 
    9.593068e-05, 0.0001288525, 0.0001145622, 0.0001307637, 0.0001485567, 
    9.571278e-05, 0.0001002052, 0.0001167021, 4.870169e-05, 1.618001e-05,
  0.0001211853, 0.0001167403, 0.0001394578, 0.0001074178, 7.446425e-05, 
    9.934112e-05, 0.0001366129, 0.0001299155, 9.558348e-05, 0.0001448314, 
    0.000135213, 8.914235e-05, 3.818002e-05, 4.504666e-05, 4.549709e-05,
  0.000149093, 0.0001320699, 0.0001263373, 9.351792e-05, 7.892301e-05, 
    0.0001140436, 0.0001528207, 0.0001594162, 0.0001370722, 0.0001607824, 
    0.0002029781, 6.723073e-05, 8.522701e-05, 3.735842e-05, 3.419889e-05,
  0.0002058717, 0.000155747, 0.0001217264, 6.945912e-05, 6.773634e-05, 
    0.0001229035, 0.0001992528, 0.0001692262, 0.0001581403, 0.0001372122, 
    0.0001642644, 9.52054e-05, 5.996306e-05, 4.41425e-05, 1.417047e-05,
  0.0002294895, 0.0001589111, 9.389332e-05, 5.004205e-05, 6.580166e-05, 
    0.0001647943, 0.0002098917, 0.0001750955, 0.0001298273, 0.0001672354, 
    0.0001282617, 0.0001466315, 7.522957e-05, 4.021744e-05, 2.197992e-05,
  0.0002307459, 0.0001566103, 7.11407e-05, 4.33657e-05, 7.73565e-05, 
    0.000182445, 0.0002321689, 0.0001753987, 0.0001409826, 0.0001586121, 
    0.0001782715, 0.00010958, 0.0001010135, 4.389736e-05, 2.780991e-05,
  0.0002007032, 0.0001253872, 5.836484e-05, 4.599538e-05, 0.0001118191, 
    0.0002497596, 0.0002549682, 0.0001654784, 0.0001561137, 0.0001725497, 
    0.0001326599, 0.0001122622, 8.936745e-05, 4.630252e-05, 4.318985e-05,
  0.0001522511, 0.0001128859, 0.0001155772, 0.0001076239, 6.403586e-05, 
    8.551228e-05, 0.0001813159, 0.0001056078, 1.77543e-05, 6.708281e-06, 
    2.18862e-06, 1.443852e-06, 8.457951e-07, 8.661085e-07, 1.034233e-06,
  0.0001342183, 0.0001318685, 0.0001324947, 0.0001660155, 0.0001119029, 
    0.0001443871, 5.870248e-05, 6.743784e-05, 1.510026e-05, 4.021058e-06, 
    1.225903e-06, 1.464062e-06, 5.480296e-07, 5.04887e-07, 6.900449e-07,
  0.0001525608, 0.0001111182, 0.0001059684, 0.0001037837, 0.0001090077, 
    0.000131373, 8.712249e-05, 1.900066e-05, 8.314953e-06, 4.249621e-06, 
    1.515763e-06, 1.061072e-06, 5.292961e-07, 4.649008e-07, 2.14214e-07,
  0.0001414438, 0.0001234323, 0.0001153786, 9.478939e-05, 9.927952e-05, 
    0.0001116558, 0.0001186621, 5.240806e-05, 1.129858e-05, 6.123481e-06, 
    2.454012e-06, 1.299803e-06, 4.806992e-07, 1.700937e-07, 7.321206e-08,
  0.0001557612, 0.0001413587, 0.0001526577, 0.000190469, 0.0001741881, 
    0.0001324746, 0.0001282348, 2.926759e-05, 1.347527e-05, 5.921123e-06, 
    3.394966e-06, 9.904553e-07, 5.460241e-07, 1.087544e-07, 5.861936e-08,
  0.0001552574, 0.0001658338, 0.0001515539, 0.0001338659, 0.0001644648, 
    0.0001388387, 9.576747e-05, 4.398072e-05, 1.490435e-05, 5.89913e-06, 
    3.21045e-06, 1.12215e-06, 6.029933e-07, 1.25411e-08, 7.088236e-09,
  0.0001423276, 0.0001557129, 0.000164898, 0.0001540317, 0.0001694219, 
    0.0001460944, 7.685695e-05, 3.109954e-05, 1.529511e-05, 6.435577e-06, 
    3.137743e-06, 1.453195e-06, 3.04032e-07, 1.950061e-10, 8.080271e-08,
  0.0001331112, 0.0001614506, 0.0002053174, 0.0001988227, 0.000169796, 
    0.0001329098, 6.73111e-05, 2.065558e-05, 1.768859e-05, 6.232448e-06, 
    3.159301e-06, 1.591741e-06, 9.519304e-08, 1.620368e-10, 2.324254e-10,
  0.000123633, 0.0001571532, 0.0001682699, 0.000186484, 0.0001841275, 
    0.0001161113, 4.680942e-05, 2.11917e-05, 1.577581e-05, 7.487559e-06, 
    3.847729e-06, 1.83862e-06, 3.75271e-07, 2.134623e-08, 1.165685e-07,
  0.0001280778, 0.0001511655, 0.0001689351, 0.0002091136, 0.000174955, 
    8.200342e-05, 3.918747e-05, 2.85463e-05, 1.535632e-05, 1.049967e-05, 
    4.546861e-06, 2.33338e-06, 7.44103e-07, 2.665394e-08, 3.224351e-07,
  0.0001107413, 8.001598e-05, 5.210025e-05, 7.239901e-05, 6.618902e-05, 
    5.535101e-05, 5.688153e-05, 4.210262e-05, 0.0001134313, 6.845739e-05, 
    6.358036e-05, 4.368134e-05, 1.727645e-05, 1.046377e-05, 6.889971e-06,
  0.0001463737, 8.756776e-05, 5.636842e-05, 7.241151e-05, 8.004992e-05, 
    4.337919e-05, 5.1057e-05, 5.44491e-05, 9.680774e-05, 6.368088e-05, 
    6.309296e-05, 3.972676e-05, 2.447379e-05, 1.000939e-05, 6.626827e-06,
  0.0001562287, 0.0001117707, 9.753589e-05, 8.943343e-05, 7.331243e-05, 
    6.440441e-05, 6.064853e-05, 6.51233e-05, 7.214423e-05, 7.29435e-05, 
    5.167873e-05, 3.513627e-05, 2.699977e-05, 1.224664e-05, 5.959519e-06,
  0.000169873, 0.0001635949, 0.0001137703, 4.950487e-05, 8.421783e-05, 
    8.834946e-05, 7.750392e-05, 0.0001281716, 7.720357e-05, 8.017113e-05, 
    4.845151e-05, 5.180727e-05, 3.078537e-05, 1.484956e-05, 7.036081e-06,
  0.0001746298, 0.0001790722, 0.0001204591, 6.30994e-05, 8.392804e-05, 
    8.274998e-05, 7.083092e-05, 0.0001726862, 0.0001344753, 5.9857e-05, 
    7.029466e-05, 4.211875e-05, 2.671615e-05, 2.000034e-05, 9.385579e-06,
  0.0001381669, 0.0001818928, 0.000138227, 0.0001099223, 4.548332e-05, 
    6.988712e-05, 0.0001260667, 0.0001590218, 0.0001577818, 0.0001079068, 
    9.064475e-05, 5.291652e-05, 3.05367e-05, 2.100004e-05, 1.300023e-05,
  0.0001077029, 0.0001558136, 0.0001760195, 0.000107323, 6.347225e-05, 
    9.1494e-05, 0.0001824285, 0.0001651127, 0.000175025, 0.000146309, 
    6.603867e-05, 5.69556e-05, 2.640956e-05, 1.60037e-05, 1.099691e-05,
  8.523452e-05, 0.0001475107, 0.0001684371, 0.0001309227, 9.242262e-05, 
    0.0001574405, 0.000208082, 0.000225155, 0.0001290593, 0.0001171549, 
    0.0001063637, 8.202476e-05, 2.821691e-05, 2.207136e-05, 1.117429e-05,
  8.773032e-05, 0.0001318265, 0.0001739032, 0.0001741349, 0.0001352545, 
    0.0002120976, 0.000194243, 0.0001792855, 0.0001724385, 0.0001187581, 
    7.286049e-05, 8.902195e-05, 3.210619e-05, 2.221295e-05, 5.508364e-06,
  7.883376e-05, 9.65413e-05, 0.0001505456, 0.0001370957, 0.0001518796, 
    0.0001903348, 0.0002537767, 0.0001595054, 0.0001356554, 0.0001283184, 
    0.0001170356, 5.352531e-05, 2.796703e-05, 2.690253e-05, 7.623909e-06,
  2.586339e-05, 5.95071e-05, 6.119989e-05, 4.845133e-05, 3.458594e-05, 
    2.577314e-05, 1.740097e-05, 1.076775e-05, 6.674501e-06, 7.109095e-06, 
    5.956462e-06, 3.218831e-06, 2.11468e-06, 1.225157e-06, 1.774836e-06,
  1.599613e-05, 2.746706e-05, 5.953393e-05, 6.289632e-05, 4.038763e-05, 
    3.087013e-05, 2.454731e-05, 1.54241e-05, 1.056984e-05, 9.267027e-06, 
    6.119291e-06, 4.484873e-06, 3.370604e-06, 2.353104e-06, 1.81956e-06,
  2.072222e-05, 1.472634e-05, 4.399075e-05, 7.436057e-05, 5.556926e-05, 
    3.467281e-05, 2.642036e-05, 1.808331e-05, 1.069457e-05, 1.186295e-05, 
    1.07204e-05, 7.650122e-06, 3.565125e-06, 3.458131e-06, 3.212849e-06,
  3.099352e-05, 1.557598e-05, 3.201808e-05, 6.097747e-05, 7.098947e-05, 
    4.659788e-05, 2.940838e-05, 2.084739e-05, 1.779369e-05, 1.396599e-05, 
    1.10801e-05, 7.765251e-06, 6.421505e-06, 5.240844e-06, 4.616592e-06,
  5.435021e-05, 3.194927e-05, 2.249254e-05, 3.903661e-05, 7.25012e-05, 
    5.939719e-05, 4.234291e-05, 2.812301e-05, 2.449085e-05, 2.009357e-05, 
    1.41305e-05, 1.003114e-05, 8.609384e-06, 6.411668e-06, 6.780252e-06,
  5.99799e-05, 5.87752e-05, 2.653655e-05, 2.887113e-05, 5.483227e-05, 
    7.667785e-05, 5.150288e-05, 3.456138e-05, 3.036949e-05, 3.076554e-05, 
    2.259052e-05, 1.342569e-05, 8.650917e-06, 1.009589e-05, 7.856363e-06,
  6.841794e-05, 8.214191e-05, 4.705388e-05, 2.451192e-05, 3.431532e-05, 
    6.851663e-05, 6.700215e-05, 4.405582e-05, 4.096332e-05, 3.901052e-05, 
    2.86322e-05, 2.021557e-05, 1.277675e-05, 1.057372e-05, 6.936556e-06,
  5.867844e-05, 8.104987e-05, 6.793516e-05, 2.689476e-05, 3.263324e-05, 
    5.134158e-05, 7.40214e-05, 5.40361e-05, 7.585956e-05, 6.38998e-05, 
    4.161169e-05, 3.128294e-05, 2.409451e-05, 1.105481e-05, 9.068413e-06,
  4.827305e-05, 9.116733e-05, 8.956114e-05, 3.512959e-05, 2.521127e-05, 
    3.552609e-05, 7.494825e-05, 0.0001059002, 9.097942e-05, 5.836341e-05, 
    5.634191e-05, 3.737981e-05, 1.938146e-05, 8.239966e-06, 1.123543e-05,
  5.081802e-05, 0.0001225823, 0.0001261932, 7.483784e-05, 2.810523e-05, 
    5.152063e-05, 9.830287e-05, 0.0001183601, 0.0001051491, 9.189707e-05, 
    3.945439e-05, 4.036427e-05, 2.740702e-05, 1.855417e-05, 1.418118e-05,
  6.148892e-05, 5.952718e-05, 5.880594e-05, 5.578269e-05, 4.770971e-05, 
    4.110526e-05, 4.133521e-05, 2.309653e-05, 1.311065e-05, 6.690313e-06, 
    6.626612e-06, 5.054387e-07, 2.810453e-07, 6.4333e-09, 5.559978e-10,
  5.264368e-05, 5.197255e-05, 5.732551e-05, 5.77443e-05, 5.526578e-05, 
    3.760701e-05, 2.918145e-05, 5.108505e-05, 1.469063e-05, 9.711516e-06, 
    7.781759e-06, 2.283458e-06, 1.287469e-07, 5.325498e-10, 7.259381e-11,
  6.87248e-05, 5.424613e-05, 6.248548e-05, 5.880284e-05, 5.163273e-05, 
    4.285478e-05, 2.471089e-05, 3.10512e-05, 1.107839e-05, 1.202323e-05, 
    8.117694e-06, 3.40437e-06, 3.479125e-07, 1.685365e-10, 3.998749e-10,
  7.409858e-05, 6.342911e-05, 5.921693e-05, 5.768071e-05, 5.320086e-05, 
    4.330366e-05, 3.334747e-05, 1.687499e-05, 3.127875e-05, 1.600666e-05, 
    7.838721e-06, 4.803073e-06, 4.780747e-07, 2.809412e-09, 2.964073e-11,
  7.026279e-05, 7.543304e-05, 7.510107e-05, 6.674659e-05, 5.809401e-05, 
    4.778122e-05, 3.844975e-05, 2.804282e-05, 1.387061e-05, 1.602461e-05, 
    9.239856e-06, 6.120641e-06, 5.856023e-07, 1.06233e-08, 1.463425e-11,
  6.857074e-05, 6.675803e-05, 5.787628e-05, 6.598532e-05, 5.791917e-05, 
    5.195758e-05, 3.832546e-05, 2.939528e-05, 1.966405e-05, 1.997942e-05, 
    9.1241e-06, 9.041152e-06, 1.885664e-06, 1.17147e-08, 3.903735e-12,
  6.522555e-05, 6.39037e-05, 7.23417e-05, 6.246488e-05, 6.851978e-05, 
    4.926375e-05, 4.04778e-05, 2.705434e-05, 2.232683e-05, 2.946242e-05, 
    7.44836e-06, 7.654452e-06, 2.354199e-06, 3.220085e-08, 5.78309e-13,
  6.102756e-05, 6.734391e-05, 6.32154e-05, 6.856432e-05, 6.172362e-05, 
    6.183994e-05, 4.466753e-05, 2.972562e-05, 2.357053e-05, 1.836941e-05, 
    2.031687e-05, 4.609957e-06, 1.767104e-06, 5.339002e-08, 2.935043e-14,
  8.120317e-05, 6.702371e-05, 7.216838e-05, 6.033631e-05, 6.133344e-05, 
    5.86696e-05, 4.066014e-05, 3.252925e-05, 2.200587e-05, 1.600282e-05, 
    9.676675e-06, 8.04963e-06, 2.76406e-06, 2.828737e-07, 9.646013e-10,
  8.659913e-05, 8.354722e-05, 7.525075e-05, 6.658517e-05, 5.991153e-05, 
    5.52612e-05, 4.73089e-05, 3.509727e-05, 2.396819e-05, 1.368312e-05, 
    7.695633e-06, 8.273291e-06, 2.902195e-06, 4.351596e-08, 1.457041e-10,
  7.434337e-06, 8.080727e-06, 4.534312e-06, 3.886504e-06, 1.694962e-06, 
    7.912129e-07, 3.45432e-08, 2.703361e-07, 8.193895e-07, 3.337304e-06, 
    8.892599e-06, 5.99584e-06, 2.391974e-06, 3.214953e-08, 6.998921e-09,
  1.191546e-05, 8.065012e-06, 6.839516e-06, 4.511053e-06, 2.31242e-06, 
    9.426304e-07, 1.081573e-07, 6.15773e-07, 9.505573e-07, 1.698429e-06, 
    8.400964e-06, 8.520767e-06, 3.657005e-06, 1.361746e-07, 4.323469e-09,
  1.406099e-05, 7.371699e-06, 6.407876e-06, 4.179823e-06, 3.181424e-06, 
    1.45973e-06, 6.26951e-07, 7.698523e-07, 1.01481e-06, 1.668305e-06, 
    7.506442e-06, 9.68119e-06, 5.057009e-06, 6.23499e-07, 1.394212e-08,
  1.719954e-05, 1.088506e-05, 7.531197e-06, 5.913232e-06, 3.39705e-06, 
    1.640178e-06, 1.486368e-06, 4.510908e-07, 1.23793e-06, 1.72986e-06, 
    5.35922e-06, 9.939849e-06, 6.310543e-06, 2.232419e-06, 3.381149e-08,
  3.155944e-05, 1.641426e-05, 8.961867e-06, 6.767063e-06, 3.710672e-06, 
    3.489418e-06, 1.234974e-06, 1.079265e-06, 1.060279e-06, 1.458973e-06, 
    4.838499e-06, 9.922236e-06, 6.242236e-06, 6.481301e-06, 1.120174e-07,
  3.712609e-05, 1.765434e-05, 1.222785e-05, 9.295517e-06, 6.142487e-06, 
    3.685989e-06, 1.899221e-06, 1.994488e-06, 1.366012e-06, 1.534539e-06, 
    3.046321e-06, 6.473444e-06, 9.11915e-06, 6.647916e-06, 8.285297e-07,
  5.5633e-05, 2.758128e-05, 1.41485e-05, 8.77903e-06, 6.459413e-06, 
    3.517025e-06, 3.127223e-06, 1.929117e-06, 1.777972e-06, 1.279626e-06, 
    3.485012e-06, 6.629015e-06, 1.14027e-05, 7.516953e-06, 1.263441e-06,
  8.323413e-05, 4.128511e-05, 2.45934e-05, 1.575134e-05, 7.522295e-06, 
    4.508673e-06, 3.718821e-06, 2.464664e-06, 1.744013e-06, 1.162191e-06, 
    2.976185e-06, 5.172102e-06, 1.214015e-05, 8.408193e-06, 1.982718e-06,
  7.400648e-05, 4.86782e-05, 3.215535e-05, 2.09788e-05, 1.049278e-05, 
    6.916221e-06, 5.074851e-06, 3.419085e-06, 2.386457e-06, 1.678938e-06, 
    1.685217e-06, 3.090438e-06, 8.611541e-06, 1.109393e-05, 5.717835e-06,
  8.327106e-05, 6.699112e-05, 4.452604e-05, 2.444703e-05, 1.64347e-05, 
    8.295446e-06, 4.989182e-06, 4.052437e-06, 3.372785e-06, 2.157289e-06, 
    1.53153e-06, 2.485679e-06, 1.107475e-05, 8.939045e-06, 6.289978e-06,
  6.348665e-08, 3.383226e-07, 4.308912e-07, 1.71685e-06, 1.250848e-06, 
    1.330822e-06, 2.319122e-06, 1.998932e-06, 4.780837e-06, 3.008445e-06, 
    4.528276e-06, 4.954269e-06, 3.601208e-06, 5.168788e-06, 4.895518e-06,
  4.760118e-08, 4.251049e-07, 3.90764e-07, 2.507677e-06, 1.447242e-06, 
    9.874173e-07, 1.008103e-06, 1.466675e-06, 1.633029e-06, 2.366595e-06, 
    3.087623e-06, 3.53915e-06, 3.584959e-06, 4.266066e-06, 7.022838e-06,
  6.689552e-08, 9.761621e-07, 1.209754e-06, 2.82811e-06, 3.999046e-06, 
    1.768494e-06, 1.056506e-06, 5.206853e-08, 1.006091e-06, 8.943956e-07, 
    1.541786e-06, 1.935832e-06, 2.389547e-06, 3.446149e-06, 6.473398e-06,
  9.278613e-08, 3.683704e-07, 7.671453e-07, 2.12771e-06, 5.318796e-06, 
    4.558828e-06, 1.914725e-06, 6.786505e-08, 6.01072e-10, 1.151168e-07, 
    2.663931e-07, 7.1502e-07, 1.844513e-06, 2.720575e-06, 3.557959e-06,
  1.061556e-07, 2.23938e-07, 1.314885e-06, 3.386304e-06, 4.098648e-06, 
    3.922364e-06, 3.64791e-06, 7.524512e-07, 1.620572e-08, 1.557979e-09, 
    2.598163e-10, 2.263151e-07, 5.445679e-07, 1.643182e-06, 2.540188e-06,
  3.668765e-08, 9.916831e-08, 1.026525e-06, 3.244916e-06, 3.740462e-06, 
    1.767e-06, 3.080221e-06, 2.925528e-06, 2.223425e-06, 9.782523e-07, 
    2.799597e-08, 2.97369e-09, 2.983335e-10, 1.596903e-06, 1.692392e-06,
  1.224097e-07, 1.834839e-07, 9.453084e-07, 2.26966e-06, 1.170247e-06, 
    1.349027e-06, 1.468778e-06, 2.284122e-06, 2.329862e-06, 1.80894e-06, 
    1.006569e-06, 6.468531e-08, 2.920346e-10, 4.16e-07, 1.562652e-06,
  3.646856e-07, 3.506857e-07, 2.904465e-07, 1.607314e-06, 5.451357e-07, 
    1.723891e-07, 3.930038e-07, 1.158441e-06, 4.865268e-07, 1.092785e-06, 
    4.337595e-07, 3.562069e-07, 5.487358e-08, 1.170418e-07, 5.755291e-07,
  5.37245e-07, 3.781759e-07, 2.762477e-07, 9.820504e-08, 7.335399e-08, 
    1.004701e-07, 2.38268e-07, 4.27744e-07, 7.635379e-07, 9.346046e-07, 
    1.571565e-06, 5.58043e-08, 2.574875e-07, 3.294379e-07, 2.891542e-07,
  7.083637e-07, 7.046753e-07, 5.219782e-07, 2.70821e-07, 1.987452e-07, 
    1.610322e-07, 1.063857e-07, 3.257253e-07, 2.815837e-07, 8.376301e-07, 
    1.105103e-06, 2.564178e-07, 2.049291e-07, 2.579133e-07, 7.472887e-07,
  0.0002658612, 0.0002294846, 0.0001969029, 0.0002226331, 0.0002319591, 
    0.0002133424, 0.000189581, 0.0002152736, 0.0002233247, 0.0001499606, 
    0.0001799482, 0.0001000129, 8.317372e-05, 5.069005e-05, 1.254797e-05,
  0.000279421, 0.0002402177, 0.0002243337, 0.0002462337, 0.0002617078, 
    0.00023917, 0.0002146193, 0.0002112202, 0.0001361083, 0.0002194064, 
    0.0001204548, 0.0001816494, 0.0001059223, 1.264817e-05, 6.016992e-06,
  0.0003136019, 0.0002670257, 0.0002822277, 0.0002832718, 0.0002906119, 
    0.0002635179, 0.0001955177, 0.0001369451, 0.0001065239, 0.000233071, 
    0.0001039058, 5.034363e-05, 1.453992e-05, 5.408006e-06, 6.480466e-06,
  0.0002788364, 0.0002653344, 0.0002955121, 0.0003166797, 0.0002630845, 
    0.0001988028, 0.0001557148, 0.0001478589, 0.0001433353, 0.0001271148, 
    9.616086e-05, 2.553459e-05, 8.301184e-06, 6.559149e-06, 7.526577e-06,
  0.0002322471, 0.0002824874, 0.0002896736, 0.0002873874, 0.0002474887, 
    0.0001956573, 0.0001184033, 0.0001289398, 0.0001108146, 5.40224e-05, 
    1.66161e-05, 1.0909e-05, 1.200441e-05, 1.177257e-05, 1.180672e-05,
  0.0001670365, 0.0002350289, 0.0002603738, 0.0002072743, 0.0001793312, 
    0.0001457779, 0.0001056118, 7.371913e-05, 3.282647e-05, 1.271316e-05, 
    3.30525e-06, 5.29098e-06, 6.501956e-06, 8.501179e-06, 1.077363e-05,
  9.088236e-05, 0.0001436945, 0.0001507394, 0.000120802, 9.407422e-05, 
    6.550689e-05, 3.507178e-05, 1.749699e-05, 5.026674e-06, 4.04837e-06, 
    1.904696e-06, 1.429914e-06, 4.322165e-06, 5.58069e-06, 4.333943e-06,
  1.719717e-05, 4.120659e-05, 4.742543e-05, 2.826065e-05, 1.19571e-05, 
    9.066538e-06, 4.837822e-06, 7.035679e-06, 1.029904e-05, 8.329425e-06, 
    2.801512e-06, 9.979047e-07, 5.889001e-07, 1.644713e-06, 2.81172e-06,
  3.903319e-07, 2.665907e-06, 2.463634e-06, 4.894675e-06, 3.841057e-06, 
    5.179937e-06, 6.921338e-06, 7.29239e-06, 6.952955e-06, 1.019022e-05, 
    5.173187e-06, 1.131678e-06, 3.904673e-07, 1.176809e-06, 2.266296e-06,
  2.02624e-06, 3.695803e-06, 4.730866e-06, 6.485926e-06, 5.243016e-06, 
    7.901996e-06, 3.213192e-06, 2.219632e-06, 3.259125e-06, 3.492548e-06, 
    3.332926e-06, 5.149366e-06, 7.571217e-06, 2.435644e-06, 9.939133e-07,
  5.602545e-06, 4.444014e-06, 1.650028e-06, 1.731565e-06, 8.971174e-07, 
    4.070756e-07, 3.46415e-08, 1.205404e-09, 2.739876e-10, 3.061939e-11, 
    1.179581e-10, 7.248681e-08, 9.224789e-06, 1.24681e-05, 5.08273e-05,
  4.237593e-06, 4.297866e-06, 2.637538e-06, 1.258804e-06, 7.774952e-07, 
    4.670188e-07, 6.680865e-08, 9.945452e-10, 3.193403e-10, 2.376095e-12, 
    2.959674e-09, 8.713736e-06, 6.589983e-05, 0.0001109506, 5.548555e-05,
  6.260546e-06, 6.63879e-06, 2.06028e-06, 1.915358e-06, 1.274628e-06, 
    6.629822e-07, 8.029962e-08, 1.730897e-08, 2.641276e-10, 3.112605e-09, 
    7.952984e-06, 0.0001019742, 5.528456e-05, 0.0001135728, 6.185419e-05,
  4.061574e-06, 3.199096e-06, 1.430833e-06, 1.221917e-06, 1.335982e-06, 
    2.886138e-07, 9.327844e-08, 2.223877e-08, 1.768057e-07, 7.233706e-06, 
    6.2965e-05, 9.015549e-05, 9.374551e-05, 0.0001056371, 0.0001033236,
  7.567964e-06, 3.740242e-06, 1.859251e-06, 9.472287e-07, 4.919901e-07, 
    4.272032e-07, 5.580607e-07, 2.43996e-06, 2.877329e-05, 6.581828e-05, 
    0.0001224179, 0.0001340559, 0.0001123228, 5.072644e-05, 7.625399e-05,
  3.350186e-05, 1.836621e-05, 8.365767e-06, 4.699683e-06, 8.765175e-06, 
    2.067121e-05, 4.179847e-05, 6.392875e-05, 9.829536e-05, 0.0001174344, 
    0.000151475, 0.0001409823, 0.0001040324, 7.443575e-05, 2.436118e-05,
  8.840564e-05, 7.171983e-05, 5.323487e-05, 4.864767e-05, 5.529971e-05, 
    7.802961e-05, 9.424282e-05, 0.0001125364, 0.0001415836, 0.0001310871, 
    0.00013639, 0.000133737, 0.0001130303, 7.663693e-05, 3.417225e-05,
  0.0001303964, 0.0001208617, 0.0001100095, 0.0001001126, 0.000102472, 
    0.0001038259, 0.0001153101, 0.0001311338, 0.0001288955, 0.0001277582, 
    0.0001325412, 0.0001296531, 0.0001114145, 7.908056e-05, 4.031205e-05,
  0.0001207237, 0.000125895, 0.0001234117, 0.0001144815, 0.0001198277, 
    0.0001285224, 0.0001339696, 0.0001411688, 0.0001277805, 0.0001031643, 
    0.0001128868, 0.0001109619, 9.738487e-05, 7.098319e-05, 4.173252e-05,
  0.0001147638, 0.0001212335, 0.0001221014, 0.0001214734, 0.0001259047, 
    0.0001312232, 0.0001507348, 0.0001431355, 0.0001261478, 0.000102746, 
    0.0001006607, 9.336192e-05, 7.971728e-05, 5.260448e-05, 3.727915e-05,
  0.0001849778, 0.0001997143, 0.000203325, 0.0002217434, 0.000178569, 
    0.0001332404, 6.604021e-05, 9.000243e-06, 4.123711e-06, 8.434928e-07, 
    1.460328e-05, 5.093482e-06, 5.71016e-06, 8.004547e-06, 8.264528e-06,
  0.0001966257, 0.0002369253, 0.0002193345, 0.0001854469, 0.0001495247, 
    6.72067e-05, 1.610185e-05, 9.732586e-06, 2.023814e-06, 6.564146e-07, 
    5.374897e-07, 2.307068e-06, 4.640158e-06, 1.054625e-05, 1.089546e-05,
  0.0002075445, 0.0002029904, 0.0001500067, 0.0001121043, 7.097374e-05, 
    2.643867e-05, 1.095343e-05, 8.418176e-06, 1.25722e-06, 9.875255e-07, 
    4.301449e-07, 3.538384e-06, 6.600337e-06, 6.190976e-06, 1.025083e-05,
  7.823102e-05, 6.642556e-05, 4.982813e-05, 3.526677e-05, 1.446136e-05, 
    5.074981e-06, 5.171492e-06, 3.29692e-06, 1.477284e-06, 5.658678e-07, 
    8.981116e-07, 1.130915e-06, 6.314872e-06, 7.727373e-06, 1.055095e-05,
  5.399462e-06, 8.998254e-06, 8.015627e-06, 9.64383e-06, 7.805405e-06, 
    3.254522e-06, 1.717046e-06, 1.734045e-06, 1.967323e-06, 1.019597e-06, 
    7.477827e-07, 8.915769e-07, 4.298252e-06, 6.021648e-06, 6.516972e-06,
  5.905266e-07, 6.856436e-07, 9.072343e-07, 1.792414e-06, 1.248321e-06, 
    5.79827e-07, 7.159848e-07, 2.321673e-06, 3.606644e-06, 8.977158e-07, 
    6.124836e-07, 1.052906e-06, 1.687749e-06, 4.075399e-06, 6.612602e-06,
  5.007112e-07, 5.770789e-07, 4.930536e-07, 1.267606e-06, 2.381355e-07, 
    1.268649e-07, 7.069332e-08, 4.149983e-07, 9.708887e-07, 9.617408e-08, 
    5.79002e-08, 9.369926e-07, 2.106072e-06, 4.187114e-06, 7.380534e-06,
  1.407284e-06, 7.802299e-07, 6.299227e-07, 1.006952e-06, 3.527065e-07, 
    5.885538e-08, 1.575163e-08, 2.887029e-08, 3.076297e-08, 1.490161e-08, 
    7.505796e-08, 2.171618e-06, 3.876991e-06, 4.114903e-06, 8.532342e-06,
  1.9349e-06, 1.727752e-06, 9.408687e-07, 7.841053e-07, 3.20901e-07, 
    2.427038e-08, 7.265306e-09, 4.36736e-08, 5.734318e-08, 1.990569e-08, 
    1.043858e-07, 1.130356e-06, 1.983784e-06, 3.640291e-06, 7.243455e-06,
  1.769665e-06, 1.261083e-06, 8.623904e-07, 6.729509e-07, 2.815448e-07, 
    4.296163e-08, 1.528235e-08, 4.826494e-08, 6.54079e-08, 2.350894e-08, 
    2.077565e-08, 4.963361e-07, 1.927897e-06, 4.331416e-06, 1.220132e-05,
  8.072853e-06, 4.311464e-06, 5.998209e-07, 3.893755e-07, 1.720017e-05, 
    7.406124e-05, 0.0001586607, 0.0001889217, 0.0001293968, 9.239157e-05, 
    5.028844e-05, 1.724716e-05, 6.269081e-05, 2.380934e-05, 2.005565e-05,
  1.765748e-05, 4.620011e-06, 1.445693e-05, 4.470299e-05, 8.263748e-05, 
    0.0001693459, 0.0002513049, 0.0002290142, 0.0001474412, 0.000108709, 
    7.175984e-05, 3.522312e-05, 6.064926e-05, 2.549795e-05, 1.843918e-05,
  7.07368e-05, 6.208281e-05, 9.763634e-05, 0.0001356924, 0.0001960181, 
    0.0002661112, 0.0002781213, 0.00023777, 0.0001724436, 0.0001245908, 
    9.289422e-05, 5.0132e-05, 8.910977e-05, 2.532806e-05, 2.476616e-05,
  0.000185832, 0.0001750845, 0.0002055576, 0.0002477194, 0.0002841082, 
    0.000315942, 0.0003024622, 0.0002259235, 0.0001875968, 0.0001418707, 
    0.0001053555, 5.570667e-05, 4.652228e-05, 4.150915e-05, 1.125266e-05,
  0.0002623315, 0.0002278703, 0.0002472042, 0.000281347, 0.000305349, 
    0.0003387787, 0.000298107, 0.0002554867, 0.0001876767, 0.0001442909, 
    0.0001115115, 6.17092e-05, 4.886813e-05, 1.998633e-05, 8.441857e-06,
  0.0002548083, 0.0002528028, 0.0002864913, 0.0003165836, 0.000346355, 
    0.0003388597, 0.0002873821, 0.0002460259, 0.0002028529, 0.0001419524, 
    0.0001148274, 6.74851e-05, 2.628237e-05, 1.979685e-05, 4.146309e-06,
  0.0002524777, 0.0002613737, 0.000301681, 0.000349309, 0.0003456941, 
    0.0003281059, 0.0003013362, 0.0002537156, 0.0002077816, 0.0001476933, 
    0.0001259772, 8.225704e-05, 4.275853e-05, 1.494643e-05, 4.876324e-06,
  0.0002620804, 0.0002964378, 0.0003217634, 0.0003521709, 0.000353018, 
    0.0003021009, 0.0002686084, 0.0002456198, 0.0002096415, 0.0001534249, 
    0.0001252954, 9.321063e-05, 5.46065e-05, 2.876321e-05, 4.284208e-06,
  0.0002857382, 0.0003097943, 0.0003224588, 0.0003230325, 0.0002902489, 
    0.0002591926, 0.000258673, 0.0002452904, 0.0001999245, 0.0001506152, 
    0.0001246876, 8.88112e-05, 5.613492e-05, 2.172858e-05, 3.942332e-06,
  0.000276173, 0.0002722363, 0.0002894644, 0.0002599739, 0.0002368414, 
    0.0001972004, 0.0001956498, 0.0002127014, 0.0002025529, 0.0001580509, 
    0.0001214104, 8.120462e-05, 4.926791e-05, 8.391731e-06, 1.651556e-06,
  1.778099e-05, 9.836923e-06, 5.927968e-06, 1.63368e-06, 4.012564e-07, 
    1.3134e-06, 5.954282e-07, 1.478762e-06, 6.575892e-06, 5.200106e-06, 
    2.165629e-06, 1.616951e-06, 1.94348e-05, 1.216191e-05, 5.446326e-06,
  1.274309e-05, 7.427909e-06, 1.589318e-06, 1.891361e-06, 7.709307e-07, 
    1.529137e-06, 8.004739e-07, 1.217665e-06, 3.620505e-06, 3.521223e-06, 
    1.873456e-06, 1.132728e-06, 1.148186e-05, 1.984928e-05, 7.229518e-06,
  6.13471e-06, 3.727459e-06, 6.15193e-07, 1.828041e-06, 1.394433e-06, 
    8.461261e-07, 4.844739e-07, 9.031754e-07, 1.42672e-06, 2.018019e-06, 
    3.341401e-06, 1.191095e-06, 1.624295e-05, 2.179533e-05, 7.082954e-06,
  5.756062e-07, 1.273265e-06, 5.635582e-07, 8.172312e-07, 8.188639e-07, 
    8.211073e-07, 6.95869e-08, 5.420675e-07, 3.027102e-07, 9.757744e-07, 
    2.954257e-06, 1.729756e-06, 1.45002e-05, 2.763405e-05, 1.199668e-05,
  2.502724e-07, 1.643491e-06, 5.883696e-07, 1.201696e-06, 8.739852e-07, 
    9.113315e-07, 4.619185e-07, 5.814207e-07, 3.094384e-07, 3.507651e-07, 
    1.613571e-06, 7.593345e-07, 8.993457e-06, 3.056894e-05, 1.789451e-05,
  1.049264e-06, 1.926484e-06, 3.585065e-07, 4.63265e-07, 4.214709e-07, 
    7.259603e-07, 3.070538e-07, 2.612774e-07, 4.524169e-07, 1.374094e-06, 
    2.893647e-07, 2.102591e-06, 1.580752e-05, 1.440854e-05, 1.166365e-05,
  3.923587e-06, 7.404076e-07, 1.370735e-07, 1.059475e-07, 2.285575e-08, 
    2.335913e-07, 3.397957e-07, 1.176152e-07, 1.331935e-06, 1.163779e-06, 
    9.597301e-08, 2.653395e-06, 1.5181e-05, 1.857978e-05, 6.000407e-06,
  4.300981e-06, 5.697464e-07, 5.553857e-08, 1.547601e-07, 6.879086e-09, 
    1.395162e-08, 2.497666e-08, 2.975672e-08, 3.46485e-07, 9.39957e-08, 
    1.152949e-08, 1.880147e-06, 1.913131e-05, 4.01663e-05, 5.349529e-06,
  2.110389e-06, 4.524315e-07, 8.455111e-09, 6.268963e-08, 3.249628e-08, 
    1.898857e-08, 9.487443e-09, 1.49718e-08, 2.598302e-08, 1.27438e-08, 
    3.181287e-09, 1.809371e-07, 2.176223e-05, 6.564464e-05, 1.51444e-05,
  1.597925e-06, 4.57087e-07, 4.312296e-07, 4.711335e-07, 1.345557e-07, 
    2.696602e-08, 1.258701e-08, 2.167947e-08, 1.084322e-08, 2.689265e-08, 
    3.537084e-08, 1.025478e-08, 1.812245e-05, 7.005545e-05, 1.613233e-05,
  1.676228e-05, 2.341362e-05, 4.048513e-05, 5.65298e-05, 8.721364e-05, 
    0.0001090321, 7.997425e-05, 3.849872e-05, 6.7086e-06, 8.354693e-07, 
    5.069458e-06, 7.611058e-06, 6.194814e-06, 2.510142e-06, 2.528396e-06,
  3.906627e-05, 3.687581e-05, 5.049258e-05, 6.447123e-05, 9.921637e-05, 
    0.0001352742, 0.0001074753, 6.420074e-05, 1.383904e-05, 3.073858e-06, 
    7.005428e-06, 2.077325e-06, 5.074477e-06, 2.624121e-06, 1.567132e-06,
  5.340792e-05, 5.553603e-05, 6.130303e-05, 6.936776e-05, 0.0001102662, 
    0.0001512932, 0.0001308394, 8.29592e-05, 2.192761e-05, 4.32626e-06, 
    1.683018e-06, 2.239347e-06, 6.57242e-06, 3.002679e-06, 1.969107e-06,
  5.908288e-05, 6.097649e-05, 6.265105e-05, 6.682306e-05, 0.0001001788, 
    0.0001375509, 0.0001288009, 8.481868e-05, 2.844213e-05, 5.32355e-06, 
    2.560601e-06, 9.630072e-07, 1.017585e-05, 4.261444e-06, 2.035964e-06,
  5.291986e-05, 6.317425e-05, 6.35726e-05, 6.405408e-05, 9.408892e-05, 
    0.0001293346, 0.0001260783, 9.802976e-05, 4.049944e-05, 8.507615e-06, 
    5.597919e-06, 6.035381e-06, 6.572238e-06, 4.321223e-06, 2.209744e-06,
  6.61831e-05, 7.458419e-05, 7.733807e-05, 6.986618e-05, 9.205766e-05, 
    0.0001355627, 0.0001491282, 0.0001121355, 5.867259e-05, 1.453693e-05, 
    4.624832e-06, 6.254307e-07, 4.747901e-07, 3.120131e-06, 1.874666e-06,
  8.374449e-05, 8.738769e-05, 8.658745e-05, 7.674639e-05, 8.753718e-05, 
    0.0001379319, 0.0001518719, 0.0001265184, 7.421385e-05, 3.059473e-05, 
    1.054948e-05, 1.570554e-06, 7.574308e-07, 4.901416e-06, 1.477032e-06,
  9.791915e-05, 0.0001130261, 0.0001027876, 9.119202e-05, 9.291406e-05, 
    0.0001288419, 0.0001372153, 0.0001230814, 7.569465e-05, 3.596964e-05, 
    1.179977e-05, 1.432617e-06, 7.966756e-07, 3.918639e-06, 5.076113e-06,
  0.0001146696, 0.0001265451, 0.000116421, 8.74225e-05, 9.292665e-05, 
    0.0001231198, 0.0001246995, 0.0001075806, 7.401464e-05, 3.667593e-05, 
    9.970196e-06, 1.163566e-06, 9.840289e-07, 4.778803e-06, 5.840982e-06,
  0.0001256476, 0.0001428874, 0.0001289872, 0.000104058, 9.706936e-05, 
    0.0001135654, 0.0001118667, 9.330162e-05, 6.833911e-05, 3.17942e-05, 
    9.992377e-06, 3.862311e-07, 2.763697e-06, 7.590316e-06, 3.242409e-06,
  1.184465e-06, 1.091491e-06, 4.270453e-07, 5.910846e-08, 2.191562e-06, 
    4.122545e-05, 6.717459e-05, 2.640852e-05, 4.965569e-06, 5.835062e-05, 
    8.057756e-05, 2.145038e-05, 2.09845e-06, 1.674903e-06, 2.372128e-06,
  2.318491e-06, 1.563942e-06, 7.237321e-07, 4.219949e-07, 1.324702e-07, 
    1.188746e-05, 4.605899e-05, 2.930141e-05, 1.444574e-06, 2.912656e-05, 
    7.976999e-05, 4.182344e-05, 3.338894e-06, 1.689758e-06, 2.473038e-06,
  1.482544e-06, 1.230029e-06, 1.210042e-06, 5.39879e-07, 6.346297e-08, 
    1.957892e-06, 1.424868e-05, 1.612971e-05, 1.228566e-06, 1.022905e-05, 
    8.437402e-05, 7.599215e-05, 5.586585e-06, 1.657246e-06, 2.18637e-06,
  2.174256e-06, 2.167935e-06, 1.179591e-06, 7.434433e-07, 2.848888e-07, 
    6.65033e-08, 1.166831e-06, 2.793946e-06, 6.024979e-07, 3.819477e-06, 
    6.779992e-05, 0.0001014212, 9.348253e-06, 2.739562e-06, 1.963327e-06,
  3.191998e-06, 3.924327e-06, 1.631483e-06, 1.123575e-06, 5.986327e-07, 
    2.500118e-07, 2.409554e-07, 1.575972e-07, 2.949731e-07, 1.410937e-06, 
    4.725438e-05, 7.874303e-05, 1.117989e-05, 3.490196e-06, 1.304108e-06,
  2.976358e-06, 5.754717e-06, 2.007362e-06, 1.489017e-06, 7.937282e-07, 
    1.170387e-08, 1.669944e-07, 1.32628e-07, 7.369949e-08, 2.6106e-06, 
    2.140193e-05, 6.540571e-05, 1.690832e-05, 1.807477e-06, 3.888827e-06,
  3.590513e-06, 3.224665e-06, 1.87377e-06, 1.374883e-06, 9.697558e-07, 
    3.912731e-07, 1.48363e-07, 4.900956e-08, 7.637201e-08, 5.165477e-06, 
    1.270338e-05, 8.015824e-05, 1.997027e-05, 9.86206e-07, 6.028403e-07,
  7.686424e-06, 4.092532e-06, 3.536281e-06, 1.797164e-06, 1.302611e-06, 
    4.716996e-07, 8.518709e-08, 7.338588e-08, 2.144073e-07, 5.527032e-06, 
    1.380586e-05, 7.880891e-05, 4.358481e-05, 2.211935e-06, 7.983559e-07,
  1.180719e-05, 6.840494e-06, 4.983509e-06, 2.653639e-06, 1.914966e-06, 
    7.319901e-07, 3.844167e-08, 2.607107e-07, 1.499044e-06, 8.071089e-06, 
    1.035741e-05, 1.249026e-05, 5.369379e-05, 5.333984e-06, 8.320496e-07,
  1.102708e-05, 8.484166e-06, 4.909726e-06, 2.310952e-06, 1.917712e-06, 
    5.195143e-07, 2.788062e-07, 3.986815e-07, 4.213245e-06, 1.093428e-05, 
    1.246886e-05, 1.597732e-05, 8.752979e-05, 7.591136e-06, 1.358438e-06,
  4.310664e-06, 7.058588e-06, 3.83022e-06, 2.926776e-05, 4.164891e-05, 
    2.833641e-05, 3.388926e-05, 2.073857e-05, 1.492996e-05, 1.603431e-05, 
    1.048224e-05, 5.71373e-07, 1.262855e-07, 5.260723e-07, 2.127816e-06,
  9.444055e-06, 8.900875e-06, 4.466159e-06, 1.123626e-05, 2.695074e-05, 
    5.133439e-05, 7.255042e-05, 5.131661e-05, 1.17207e-05, 1.404388e-05, 
    1.739231e-05, 1.715781e-06, 5.725324e-07, 6.70448e-07, 2.001236e-06,
  1.146616e-05, 5.263398e-06, 4.410397e-06, 5.781171e-06, 2.134717e-05, 
    5.054248e-05, 0.0001061411, 9.016519e-05, 1.807503e-05, 2.119706e-05, 
    2.005511e-05, 1.317926e-05, 5.291088e-07, 4.935453e-07, 2.541673e-06,
  9.999841e-06, 1.426892e-05, 3.206071e-06, 2.388399e-06, 1.688102e-05, 
    3.302042e-05, 0.0001061622, 0.0001164256, 3.07759e-05, 2.114079e-05, 
    2.687916e-05, 1.36275e-05, 1.654628e-06, 1.563219e-06, 1.802053e-06,
  1.376892e-05, 1.588019e-05, 2.32457e-07, 2.004448e-06, 1.461275e-05, 
    2.17723e-05, 8.220557e-05, 0.0001258919, 5.476868e-05, 1.659354e-05, 
    2.6101e-05, 2.188109e-05, 7.966923e-07, 1.906592e-06, 2.570355e-06,
  1.639197e-05, 5.934956e-06, 2.671446e-07, 2.357163e-06, 1.106836e-05, 
    1.426537e-05, 6.31579e-05, 0.0001258894, 7.71638e-05, 1.830861e-05, 
    6.218699e-06, 2.5877e-05, 1.409883e-06, 2.065662e-06, 1.739733e-06,
  1.491156e-05, 4.106796e-06, 4.049077e-07, 5.034876e-07, 7.219654e-06, 
    1.567171e-05, 5.618141e-05, 0.0001173476, 8.647388e-05, 1.91013e-05, 
    1.844799e-05, 1.638314e-05, 1.391048e-06, 2.557138e-06, 1.979502e-06,
  1.082571e-05, 6.704626e-07, 2.751715e-07, 5.242814e-07, 3.294102e-06, 
    1.316657e-05, 5.776585e-05, 0.0001026509, 7.482336e-05, 8.244276e-06, 
    1.103397e-05, 3.511313e-05, 1.47212e-06, 2.131917e-06, 1.200395e-06,
  3.806941e-06, 1.859271e-07, 4.926762e-07, 9.328303e-07, 1.384246e-06, 
    6.31486e-06, 5.53721e-05, 0.0001056592, 6.945914e-05, 3.687109e-06, 
    6.666474e-06, 3.457558e-05, 1.24077e-05, 7.909203e-07, 4.750651e-06,
  6.336087e-07, 1.224604e-07, 3.505473e-07, 3.790425e-07, 1.216535e-06, 
    6.076207e-06, 4.892408e-05, 0.0001172399, 8.305581e-05, 5.051981e-06, 
    4.465862e-06, 5.802106e-06, 2.914718e-05, 2.620473e-06, 4.028127e-06,
  8.307836e-07, 8.305568e-07, 4.545705e-06, 1.500123e-05, 2.804446e-05, 
    2.64521e-05, 1.439102e-05, 1.056456e-05, 1.322731e-05, 1.186194e-05, 
    6.112357e-06, 1.426047e-06, 7.607163e-08, 1.417558e-06, 3.836262e-06,
  7.080259e-07, 1.198696e-06, 6.178068e-06, 1.908386e-05, 2.847221e-05, 
    2.887631e-05, 1.736902e-05, 6.536738e-06, 2.141324e-05, 9.07908e-06, 
    3.922198e-06, 1.922393e-06, 2.663429e-09, 1.102167e-06, 3.579217e-06,
  1.983834e-07, 6.129296e-06, 1.086193e-05, 2.161137e-05, 3.202907e-05, 
    3.267657e-05, 1.877661e-05, 7.789754e-06, 9.172911e-06, 7.201719e-06, 
    3.60376e-06, 1.484661e-06, 8.051147e-08, 1.328602e-06, 3.345342e-06,
  1.30505e-07, 7.278025e-06, 1.099206e-05, 1.728766e-05, 3.179456e-05, 
    3.56562e-05, 2.084253e-05, 5.154935e-06, 3.428269e-06, 6.731421e-06, 
    8.115231e-06, 2.247223e-06, 6.380968e-07, 9.668979e-07, 1.820445e-06,
  3.171409e-06, 1.015105e-05, 1.54075e-05, 1.489761e-05, 2.794179e-05, 
    3.409458e-05, 2.424156e-05, 1.005669e-05, 1.484996e-06, 4.278781e-06, 
    8.50681e-06, 1.589009e-06, 9.793931e-07, 8.694806e-07, 2.3107e-06,
  2.973599e-06, 7.469828e-06, 1.016271e-05, 1.36687e-05, 2.520996e-05, 
    3.640429e-05, 2.126478e-05, 8.784737e-06, 2.6856e-06, 5.703934e-06, 
    1.29929e-05, 8.699298e-07, 3.876958e-07, 1.058327e-06, 3.058087e-06,
  1.194973e-05, 1.195777e-05, 1.552673e-05, 8.318518e-06, 1.915403e-05, 
    3.425825e-05, 1.883898e-05, 4.321877e-06, 2.682021e-06, 5.266818e-06, 
    1.217793e-05, 7.460662e-07, 7.433555e-08, 1.106865e-06, 4.816982e-06,
  2.510947e-05, 1.656742e-05, 1.98589e-05, 1.445254e-05, 1.557432e-05, 
    2.322727e-05, 1.372589e-05, 4.477099e-06, 3.24012e-06, 6.338389e-06, 
    1.350527e-05, 7.277953e-07, 2.10063e-08, 4.722613e-07, 5.57344e-06,
  3.546393e-05, 2.160038e-05, 1.280676e-05, 7.291211e-06, 1.376738e-05, 
    1.16824e-05, 8.197301e-06, 4.429199e-06, 2.487523e-06, 1.540204e-05, 
    1.02475e-05, 1.401461e-06, 1.043046e-07, 1.643913e-06, 8.343772e-06,
  4.994673e-05, 2.491229e-05, 8.940934e-06, 3.891196e-06, 4.027485e-06, 
    5.635051e-06, 2.847413e-06, 1.38877e-06, 2.542237e-06, 9.969741e-06, 
    1.528267e-05, 3.217589e-06, 6.215951e-07, 3.892984e-06, 9.754555e-06,
  1.867941e-06, 2.940144e-06, 5.194257e-06, 4.401484e-06, 1.842228e-05, 
    1.19091e-05, 1.159916e-05, 1.109091e-05, 6.382567e-06, 3.876968e-06, 
    1.557282e-05, 1.471039e-05, 2.128897e-05, 1.262317e-05, 7.858072e-06,
  2.336947e-06, 2.574139e-06, 5.516667e-06, 4.348918e-06, 1.549029e-05, 
    1.519098e-05, 5.58121e-06, 6.042112e-06, 3.193723e-06, 1.824861e-06, 
    1.166893e-05, 1.462828e-05, 2.341001e-05, 8.116163e-06, 6.365794e-06,
  3.27573e-06, 3.65438e-06, 4.882247e-06, 4.332444e-06, 1.602612e-05, 
    1.632162e-05, 7.747643e-06, 8.530117e-06, 2.540464e-06, 1.296053e-06, 
    3.360773e-06, 1.009446e-05, 9.01049e-06, 4.061222e-06, 4.033847e-06,
  2.880279e-06, 3.344698e-06, 4.748318e-06, 4.48425e-06, 1.330397e-05, 
    1.336709e-05, 1.098806e-05, 7.775402e-06, 5.972392e-06, 2.766669e-06, 
    4.150389e-06, 3.603054e-06, 6.432658e-06, 5.711057e-06, 4.128791e-06,
  3.687242e-06, 2.263424e-06, 3.991772e-06, 4.671058e-06, 1.068078e-05, 
    1.032926e-05, 1.235841e-05, 8.121466e-06, 4.213979e-06, 2.49976e-06, 
    2.569897e-06, 5.383152e-06, 6.538716e-06, 5.594489e-06, 5.360416e-06,
  3.82868e-06, 1.199745e-06, 3.113732e-06, 4.920169e-06, 1.163056e-05, 
    1.062235e-05, 1.127737e-05, 5.076378e-06, 4.674283e-06, 5.632356e-07, 
    4.592873e-06, 6.936952e-06, 7.005292e-06, 8.475813e-06, 4.114087e-06,
  4.930255e-06, 7.181347e-07, 2.420619e-06, 6.053504e-06, 1.411022e-05, 
    1.248836e-05, 9.981864e-06, 4.677232e-06, 6.776128e-06, 1.641505e-07, 
    6.029143e-06, 5.494544e-06, 1.343049e-05, 1.249297e-05, 6.569153e-06,
  2.871437e-06, 2.337839e-07, 1.871563e-06, 8.002909e-06, 1.715043e-05, 
    1.257861e-05, 4.960179e-06, 5.84915e-06, 8.156923e-06, 1.256139e-06, 
    4.201649e-06, 3.953249e-06, 3.142509e-06, 1.320639e-05, 8.264564e-06,
  4.334497e-06, 4.438672e-07, 1.950732e-06, 9.903685e-06, 2.372409e-05, 
    2.03083e-05, 5.943146e-06, 3.216841e-06, 7.706127e-06, 3.344857e-06, 
    4.598484e-06, 4.220044e-06, 1.030432e-05, 6.826833e-06, 7.703774e-06,
  6.063233e-06, 8.950689e-07, 4.416339e-06, 1.130774e-05, 2.617158e-05, 
    2.511029e-05, 1.140365e-05, 3.197223e-06, 1.020153e-05, 2.84182e-06, 
    4.606184e-06, 4.74624e-06, 2.967191e-06, 8.067035e-06, 6.399166e-06,
  4.799555e-06, 7.918893e-06, 5.113195e-06, 1.105978e-05, 7.834672e-06, 
    3.045579e-06, 4.443954e-06, 1.257368e-05, 2.563907e-05, 2.964504e-05, 
    1.848468e-05, 1.5759e-05, 9.993108e-06, 6.104337e-06, 4.882961e-06,
  4.958833e-06, 8.107031e-06, 5.928725e-06, 9.575318e-06, 1.099968e-05, 
    5.228987e-06, 3.245726e-06, 2.997328e-05, 2.566995e-05, 3.471398e-05, 
    3.009589e-05, 1.321763e-05, 7.626393e-06, 4.541503e-06, 4.916292e-06,
  4.159732e-06, 7.551958e-06, 6.524563e-06, 1.300278e-05, 1.531467e-05, 
    5.703396e-06, 5.807469e-06, 6.806172e-07, 4.376505e-05, 4.03047e-05, 
    2.961359e-05, 9.553513e-06, 8.978053e-06, 4.408912e-06, 5.284005e-06,
  4.353762e-06, 5.413959e-06, 5.557134e-06, 1.215902e-05, 1.542449e-05, 
    6.241521e-06, 6.258945e-06, 5.567207e-07, 1.994525e-05, 2.433453e-05, 
    2.133915e-05, 1.164614e-05, 8.357515e-06, 6.040945e-06, 6.900815e-06,
  3.181067e-06, 5.020484e-06, 5.931496e-06, 1.005784e-05, 1.295079e-05, 
    9.772542e-06, 2.936666e-06, 1.74262e-06, 6.686566e-07, 2.668887e-05, 
    2.37138e-05, 6.101517e-06, 5.807928e-06, 7.02682e-06, 6.273008e-06,
  2.13858e-06, 5.430144e-06, 5.893733e-06, 8.184606e-06, 1.056734e-05, 
    1.395152e-05, 2.217788e-06, 1.357709e-06, 3.82324e-06, 6.847283e-06, 
    3.063884e-05, 1.158409e-05, 1.456386e-05, 6.09334e-06, 6.689219e-06,
  2.061647e-06, 6.089555e-06, 4.846393e-06, 7.482168e-06, 1.490976e-05, 
    1.383728e-05, 2.858925e-06, 3.199493e-06, 6.422738e-06, 1.55966e-05, 
    3.475832e-05, 1.122813e-05, 6.710642e-06, 4.032295e-06, 5.350442e-06,
  3.737992e-06, 6.088127e-06, 4.670901e-06, 5.065543e-06, 1.384004e-05, 
    1.563647e-05, 2.740484e-06, 6.492884e-06, 1.035961e-05, 8.217071e-06, 
    6.852023e-06, 9.390987e-06, 3.371104e-06, 3.003066e-06, 2.832741e-06,
  6.98313e-06, 6.841043e-06, 4.360424e-06, 3.732292e-06, 9.526543e-06, 
    1.595618e-05, 3.699628e-06, 2.96721e-06, 6.451094e-06, 1.192745e-05, 
    8.489951e-06, 4.694738e-06, 3.525363e-06, 1.888258e-06, 2.834804e-06,
  9.004258e-06, 6.846165e-06, 5.263704e-06, 6.219647e-06, 8.72016e-06, 
    1.805507e-05, 4.948539e-06, 4.674922e-06, 8.974504e-06, 1.137548e-05, 
    1.135737e-05, 8.871851e-06, 4.10808e-06, 2.942934e-06, 5.020644e-06,
  2.11153e-06, 2.534448e-06, 1.378278e-05, 1.155568e-05, 5.987237e-06, 
    5.795352e-06, 4.556923e-06, 2.292049e-05, 3.433246e-05, 2.405028e-05, 
    1.513613e-05, 9.844161e-06, 6.372848e-06, 7.949578e-06, 1.110337e-05,
  2.36219e-06, 2.975037e-06, 1.649225e-05, 1.396793e-05, 5.56154e-06, 
    4.526422e-06, 1.473269e-05, 4.331482e-06, 2.137305e-05, 1.601158e-05, 
    1.15658e-05, 6.20719e-06, 5.19515e-06, 7.887059e-06, 1.029323e-05,
  1.364224e-06, 3.714671e-06, 1.468054e-05, 1.56563e-05, 6.005644e-06, 
    2.120817e-06, 1.765386e-06, 1.869745e-05, 1.016084e-05, 7.213964e-06, 
    4.752417e-06, 3.284711e-06, 3.924576e-06, 5.886227e-06, 7.856836e-06,
  8.450015e-07, 3.96478e-06, 1.39577e-05, 1.691869e-05, 8.757055e-06, 
    9.500906e-06, 5.889177e-06, 1.571206e-05, 1.319467e-05, 3.441624e-06, 
    1.773383e-06, 2.39549e-06, 3.400752e-06, 4.752882e-06, 7.317224e-06,
  9.474314e-07, 3.036356e-06, 1.364384e-05, 1.91714e-05, 8.532239e-06, 
    5.580291e-06, 7.391837e-06, 1.257462e-05, 3.814585e-06, 1.339495e-06, 
    1.143395e-06, 1.95643e-06, 2.381726e-06, 3.186736e-06, 6.122757e-06,
  1.716685e-06, 2.895074e-06, 1.090211e-05, 1.683259e-05, 8.325665e-06, 
    5.309507e-06, 9.996058e-06, 6.313773e-06, 6.40019e-06, 1.738217e-06, 
    2.699014e-06, 1.168607e-06, 3.231126e-06, 3.331807e-06, 4.331678e-06,
  3.191925e-06, 3.667962e-06, 8.654258e-06, 1.294655e-05, 6.551027e-06, 
    7.014291e-06, 1.107982e-05, 9.704119e-06, 9.108709e-06, 4.396832e-06, 
    3.729259e-06, 2.284335e-06, 3.785278e-06, 3.232199e-06, 3.517767e-06,
  3.430324e-06, 5.153947e-06, 7.483615e-06, 1.417061e-05, 8.280523e-06, 
    5.960106e-06, 8.122122e-06, 1.097933e-05, 6.326375e-06, 3.586175e-06, 
    2.654293e-06, 4.076658e-06, 1.759128e-06, 3.365582e-06, 3.545073e-06,
  4.262238e-06, 6.469057e-06, 9.049402e-06, 1.194312e-05, 1.093353e-05, 
    4.835191e-06, 6.505647e-06, 1.086336e-05, 4.540677e-06, 4.798132e-06, 
    4.259419e-06, 4.884943e-06, 3.951092e-06, 5.005416e-06, 3.478015e-06,
  4.226493e-06, 7.346669e-06, 8.453216e-06, 9.903953e-06, 9.408452e-06, 
    4.588687e-06, 3.754307e-06, 1.121604e-05, 7.501006e-06, 7.378256e-06, 
    9.331583e-06, 4.292222e-06, 3.035474e-06, 7.226655e-06, 4.556604e-06,
  2.315485e-06, 4.07508e-06, 1.119188e-05, 1.099323e-05, 1.096631e-05, 
    1.122114e-05, 2.084595e-06, 4.907018e-06, 3.46508e-06, 4.742989e-06, 
    2.637723e-06, 3.233973e-06, 4.416133e-06, 5.818833e-06, 6.191394e-06,
  3.229491e-06, 4.333102e-06, 1.121026e-05, 1.050973e-05, 1.274078e-05, 
    9.756818e-06, 3.209311e-06, 4.069917e-06, 3.325754e-06, 3.239502e-06, 
    3.040987e-06, 3.558253e-06, 4.907381e-06, 5.448453e-06, 5.24903e-06,
  5.171674e-06, 4.369068e-06, 7.533984e-06, 1.200047e-05, 9.996452e-06, 
    3.622704e-06, 3.088776e-06, 3.974398e-06, 2.925703e-06, 2.697639e-06, 
    2.310512e-06, 3.786745e-06, 4.087516e-06, 5.459907e-06, 5.478645e-06,
  5.78971e-06, 4.104485e-06, 5.282358e-06, 1.098061e-05, 7.648638e-06, 
    6.24311e-06, 5.093266e-06, 3.658359e-06, 3.079152e-06, 3.854747e-06, 
    3.256819e-06, 3.637246e-06, 3.200489e-06, 5.263235e-06, 4.700979e-06,
  6.25825e-06, 4.30752e-06, 5.752995e-06, 1.077598e-05, 5.651621e-06, 
    1.003799e-05, 8.145818e-06, 6.494526e-06, 2.875898e-06, 4.985074e-06, 
    3.802132e-06, 3.067315e-06, 4.478092e-06, 4.047675e-06, 4.773322e-06,
  7.224886e-06, 6.473931e-06, 4.474052e-06, 7.329073e-06, 8.859129e-06, 
    6.148865e-06, 8.812098e-06, 8.095426e-06, 4.306587e-06, 4.154299e-06, 
    3.501377e-06, 3.246302e-06, 5.17062e-06, 4.65762e-06, 5.253871e-06,
  4.991816e-06, 5.143817e-06, 1.296503e-06, 9.070868e-06, 1.099974e-05, 
    5.224479e-06, 9.747997e-06, 8.548537e-06, 7.699439e-06, 3.86204e-06, 
    5.862948e-06, 3.936982e-06, 3.72216e-06, 5.355871e-06, 5.056786e-06,
  6.788072e-06, 5.176611e-06, 8.317803e-07, 2.89436e-06, 1.036609e-05, 
    8.2123e-06, 8.89674e-06, 6.645336e-06, 4.88513e-06, 2.762392e-06, 
    5.048698e-06, 4.153829e-06, 4.495843e-06, 5.745168e-06, 5.635855e-06,
  4.031813e-06, 2.69361e-06, 4.492282e-07, 4.563969e-06, 3.794184e-06, 
    9.427985e-06, 1.06707e-05, 6.65062e-06, 6.412977e-06, 5.387269e-06, 
    4.90442e-06, 5.660341e-06, 5.631723e-06, 5.710629e-06, 6.393458e-06,
  4.080443e-06, 3.373933e-06, 4.405896e-07, 4.757949e-06, 3.80101e-06, 
    1.045018e-05, 1.024614e-05, 7.915829e-06, 5.425468e-06, 6.807e-06, 
    5.101244e-06, 5.71043e-06, 5.592482e-06, 6.468054e-06, 7.910491e-06,
  2.227851e-05, 1.053424e-05, 6.084405e-06, 1.109522e-05, 9.428773e-06, 
    4.313006e-06, 7.760783e-07, 1.27377e-06, 2.408106e-06, 3.129877e-06, 
    2.641346e-06, 3.442414e-06, 2.969934e-06, 5.122367e-06, 4.424182e-06,
  1.749738e-05, 1.264721e-05, 1.057849e-05, 7.377259e-06, 3.975992e-06, 
    9.984933e-07, 3.293161e-06, 1.56872e-06, 1.63817e-06, 2.67468e-06, 
    4.707599e-06, 4.594328e-06, 4.441781e-06, 6.032015e-06, 7.593056e-06,
  1.15599e-05, 1.20601e-05, 1.19939e-05, 1.034171e-05, 6.835722e-06, 
    1.177454e-06, 2.264974e-06, 1.547318e-06, 2.497118e-06, 3.897734e-06, 
    4.463415e-06, 5.420999e-06, 4.240006e-06, 6.716285e-06, 6.662487e-06,
  9.690594e-06, 1.254258e-05, 1.345298e-05, 7.423825e-06, 2.626632e-06, 
    7.590785e-07, 2.073828e-06, 2.926961e-06, 2.514202e-06, 3.74753e-06, 
    4.397628e-06, 5.25825e-06, 6.607948e-06, 7.556449e-06, 8.310473e-06,
  8.410419e-06, 1.115152e-05, 1.352804e-05, 5.681193e-06, 2.0624e-06, 
    3.331042e-06, 1.386398e-06, 3.468227e-06, 2.652765e-06, 3.984966e-06, 
    4.409431e-06, 4.941646e-06, 7.570407e-06, 8.489166e-06, 9.358712e-06,
  8.16501e-06, 1.088236e-05, 1.232945e-05, 6.441395e-06, 2.371154e-06, 
    5.529488e-06, 5.206696e-06, 5.191109e-06, 3.361625e-06, 3.954392e-06, 
    3.947887e-06, 5.835058e-06, 6.235294e-06, 7.224486e-06, 9.075174e-06,
  8.96061e-06, 9.284588e-06, 1.190471e-05, 8.436284e-06, 3.734297e-06, 
    7.09597e-06, 6.421504e-06, 3.622163e-06, 2.31067e-06, 4.382599e-06, 
    4.562084e-06, 4.971902e-06, 5.548091e-06, 6.755432e-06, 7.230694e-06,
  7.383341e-06, 8.593e-06, 1.095169e-05, 7.49202e-06, 3.384037e-06, 
    2.6216e-06, 5.744762e-06, 4.977214e-06, 4.909702e-06, 5.05934e-06, 
    5.612801e-06, 5.368439e-06, 7.010732e-06, 5.885193e-06, 6.961574e-06,
  5.664705e-06, 8.878949e-06, 9.340423e-06, 7.10797e-06, 5.296468e-06, 
    3.425853e-06, 3.549884e-06, 6.49921e-06, 4.598822e-06, 4.666744e-06, 
    7.456326e-06, 6.207132e-06, 4.759208e-06, 6.308874e-06, 6.559346e-06,
  3.716322e-06, 6.423396e-06, 8.440018e-06, 5.032819e-06, 4.643894e-06, 
    5.594242e-06, 3.616731e-06, 6.488817e-06, 5.781835e-06, 7.341714e-06, 
    5.472429e-06, 4.466514e-06, 4.375856e-06, 6.067268e-06, 6.012628e-06,
  3.69792e-05, 5.364393e-05, 6.363312e-05, 4.610444e-05, 3.488175e-05, 
    3.058956e-05, 4.88647e-05, 2.733411e-05, 2.574972e-05, 1.824559e-05, 
    4.721275e-06, 2.163763e-06, 2.639631e-06, 6.000249e-06, 7.461303e-06,
  5.801887e-05, 7.509623e-05, 8.461913e-05, 6.345032e-05, 3.636243e-05, 
    4.157528e-05, 5.064882e-05, 3.941768e-05, 4.19244e-05, 1.981251e-05, 
    5.35609e-06, 2.382304e-06, 4.053316e-06, 6.970624e-06, 8.836168e-06,
  7.121977e-05, 0.0001051522, 0.0001097461, 7.946455e-05, 5.066139e-05, 
    5.15726e-05, 5.143651e-05, 5.922244e-05, 3.354729e-05, 2.507507e-05, 
    5.505142e-06, 3.140177e-06, 4.533712e-06, 6.180581e-06, 7.087856e-06,
  0.0001014383, 0.0001348593, 0.0001321069, 8.88006e-05, 5.845294e-05, 
    4.956611e-05, 5.25847e-05, 4.234139e-05, 2.471842e-05, 1.288831e-05, 
    3.59822e-06, 2.253174e-06, 2.658718e-06, 4.042503e-06, 4.595822e-06,
  0.0001390858, 0.0001802703, 0.0001506542, 9.869094e-05, 5.512339e-05, 
    4.062815e-05, 3.259512e-05, 3.218291e-05, 2.223031e-05, 1.08373e-05, 
    3.432187e-06, 2.354099e-06, 2.452989e-06, 2.905824e-06, 5.298581e-06,
  0.0001853327, 0.0002155689, 0.0001766095, 0.0001022674, 6.487554e-05, 
    5.216242e-05, 3.413585e-05, 2.546859e-05, 1.69061e-05, 8.266829e-06, 
    3.662975e-06, 1.644887e-06, 1.75709e-06, 2.62261e-06, 3.413791e-06,
  0.0002189393, 0.0002191786, 0.0001846996, 0.0001018282, 6.655778e-05, 
    3.845397e-05, 3.803784e-05, 1.864122e-05, 1.332017e-05, 5.885387e-06, 
    2.279986e-06, 1.418944e-06, 2.038863e-06, 2.800618e-06, 3.395034e-06,
  0.0002406259, 0.0002281051, 0.0001801405, 0.0001081871, 6.691891e-05, 
    4.749715e-05, 2.748595e-05, 1.819886e-05, 1.042427e-05, 5.435995e-06, 
    1.373708e-06, 1.465729e-06, 1.691986e-06, 3.681421e-06, 3.032774e-06,
  0.0002473412, 0.0002151642, 0.000165303, 9.906952e-05, 6.353466e-05, 
    4.144532e-05, 2.325283e-05, 1.582302e-05, 1.543081e-05, 4.106553e-06, 
    1.207428e-06, 6.337004e-07, 1.501482e-06, 4.418371e-06, 4.277008e-06,
  0.0002456391, 0.0001926286, 0.0001393659, 8.812339e-05, 5.752403e-05, 
    3.049514e-05, 2.431108e-05, 1.66787e-05, 7.682683e-06, 2.36437e-06, 
    1.426979e-06, 1.552193e-06, 2.59789e-06, 4.170745e-06, 6.392504e-06,
  5.955416e-06, 4.259814e-06, 2.332389e-06, 1.30055e-06, 5.563368e-07, 
    1.286117e-07, 4.702267e-08, 5.445323e-07, 4.334153e-06, 1.041688e-05, 
    1.822052e-05, 1.613232e-05, 9.134514e-06, 2.91274e-06, 1.864892e-06,
  2.624534e-06, 1.55198e-06, 1.692281e-06, 1.169997e-06, 1.221147e-06, 
    3.621585e-07, 5.58692e-08, 2.686108e-07, 2.451691e-06, 7.617663e-06, 
    1.735688e-05, 2.236586e-05, 1.472757e-05, 5.796418e-06, 1.218196e-06,
  2.488311e-06, 1.313711e-06, 1.304376e-06, 1.349202e-06, 2.096189e-07, 
    1.364754e-07, 1.12528e-07, 1.205829e-08, 3.025363e-06, 6.847761e-06, 
    1.93097e-05, 2.501425e-05, 1.866917e-05, 4.135661e-06, 1.533944e-06,
  2.875806e-06, 1.006189e-06, 5.483995e-07, 1.742043e-07, 7.699051e-08, 
    9.970118e-08, 2.402969e-08, 1.529438e-07, 3.094138e-06, 5.321969e-06, 
    1.393314e-05, 2.387271e-05, 2.201516e-05, 9.655679e-06, 2.426125e-06,
  2.247437e-06, 4.404486e-07, 2.904918e-07, 1.810267e-07, 1.381506e-07, 
    1.115896e-07, 9.202293e-09, 4.883016e-07, 3.729905e-06, 8.986173e-06, 
    1.527078e-05, 2.832993e-05, 2.660496e-05, 1.256023e-05, 2.38501e-06,
  2.840567e-06, 1.111697e-06, 5.500345e-07, 1.166344e-07, 7.728629e-08, 
    4.020348e-07, 2.979171e-08, 9.560748e-07, 5.339423e-06, 1.165735e-05, 
    1.599745e-05, 2.820344e-05, 2.651239e-05, 1.382879e-05, 3.744226e-06,
  1.982897e-06, 2.150277e-06, 4.616876e-07, 2.449573e-07, 1.451525e-07, 
    6.559446e-08, 7.539123e-08, 2.531387e-06, 6.792193e-06, 1.624281e-05, 
    1.997539e-05, 2.925764e-05, 2.980404e-05, 1.372185e-05, 3.403434e-06,
  2.569252e-06, 1.995479e-06, 9.665615e-07, 7.985863e-07, 1.262055e-07, 
    1.549348e-07, 2.570183e-07, 3.78136e-06, 8.460531e-06, 1.881975e-05, 
    2.472193e-05, 3.506388e-05, 2.915346e-05, 1.889645e-05, 1.359323e-06,
  2.08798e-06, 2.07779e-06, 2.309223e-06, 1.025418e-06, 2.169568e-07, 
    2.018196e-07, 7.122392e-07, 3.560937e-06, 9.181826e-06, 2.287489e-05, 
    2.619745e-05, 2.240867e-05, 3.71054e-05, 1.336362e-05, 5.132252e-07,
  2.367298e-06, 3.381704e-06, 3.064838e-06, 1.53417e-06, 5.559153e-07, 
    6.750067e-07, 1.29166e-06, 3.538312e-06, 9.613386e-06, 2.10941e-05, 
    3.096678e-05, 4.279523e-05, 2.582494e-05, 6.85463e-06, 4.609101e-07,
  4.78202e-05, 6.247031e-05, 5.337826e-05, 2.707321e-05, 1.732172e-05, 
    1.2915e-05, 9.744884e-06, 7.397653e-06, 8.824813e-06, 6.830874e-06, 
    2.733875e-06, 3.640149e-06, 7.635318e-06, 9.656259e-06, 8.827969e-06,
  4.337114e-05, 4.067801e-05, 4.052357e-05, 2.875909e-05, 1.79914e-05, 
    1.29732e-05, 1.26168e-05, 6.320807e-06, 8.489856e-06, 7.867266e-06, 
    2.988059e-06, 2.399724e-06, 5.976985e-06, 1.140342e-05, 9.684822e-06,
  6.209989e-05, 4.983877e-05, 5.037548e-05, 3.992592e-05, 1.648327e-05, 
    1.794105e-05, 1.316749e-05, 1.12e-05, 9.72666e-06, 9.596311e-06, 
    7.044483e-06, 3.833105e-06, 6.46361e-06, 1.268696e-05, 1.307489e-05,
  7.034914e-05, 7.524412e-05, 6.667589e-05, 4.873395e-05, 3.307263e-05, 
    2.09121e-05, 1.531019e-05, 1.529721e-05, 1.152697e-05, 8.789478e-06, 
    7.012443e-06, 3.699669e-06, 4.78741e-06, 1.35269e-05, 1.414904e-05,
  9.109431e-05, 0.0001003364, 8.371739e-05, 6.13263e-05, 3.873006e-05, 
    2.679673e-05, 2.305996e-05, 1.869052e-05, 1.48935e-05, 9.179072e-06, 
    7.148888e-06, 5.003173e-06, 3.909665e-06, 1.233829e-05, 1.801785e-05,
  9.995892e-05, 0.0001025542, 9.71077e-05, 6.808404e-05, 5.173247e-05, 
    3.407771e-05, 1.862892e-05, 2.020239e-05, 1.586749e-05, 1.210836e-05, 
    1.00619e-05, 4.826031e-06, 4.482605e-06, 1.196653e-05, 1.690546e-05,
  0.0001182436, 0.0001101067, 0.0001010624, 7.627335e-05, 5.380854e-05, 
    3.605237e-05, 2.122233e-05, 1.94364e-05, 1.610538e-05, 1.265691e-05, 
    1.033805e-05, 5.54465e-06, 4.244738e-06, 1.28652e-05, 1.770111e-05,
  0.0001386086, 0.0001221015, 0.0001082856, 8.651197e-05, 6.604369e-05, 
    3.329148e-05, 2.354741e-05, 1.765985e-05, 2.005534e-05, 1.441896e-05, 
    7.788106e-06, 4.963186e-06, 5.705988e-06, 1.617764e-05, 1.66594e-05,
  0.000139617, 0.0001350264, 0.0001209784, 9.258914e-05, 6.759461e-05, 
    4.224234e-05, 2.921645e-05, 2.017705e-05, 2.386262e-05, 1.635455e-05, 
    5.325906e-06, 4.458979e-06, 7.53799e-06, 1.770769e-05, 1.841928e-05,
  0.0001292384, 0.0001260139, 0.000111267, 9.320409e-05, 7.419224e-05, 
    5.318684e-05, 3.339056e-05, 2.915477e-05, 2.680346e-05, 1.230289e-05, 
    4.602648e-06, 5.186276e-06, 9.427542e-06, 2.062978e-05, 2.189876e-05,
  7.512946e-06, 3.801545e-06, 1.997288e-07, 5.633991e-07, 6.715917e-07, 
    4.084361e-07, 3.572477e-07, 1.767316e-07, 3.158749e-06, 7.471193e-06, 
    7.278838e-06, 1.211588e-05, 7.27552e-06, 1.044441e-05, 9.384404e-06,
  6.863822e-06, 4.843601e-06, 2.83008e-06, 8.52805e-07, 2.862776e-07, 
    3.557463e-07, 4.943377e-07, 4.981571e-07, 6.976436e-07, 3.712999e-06, 
    8.492309e-06, 9.763255e-06, 1.140138e-05, 1.166806e-05, 9.462639e-06,
  8.508615e-06, 6.661769e-06, 6.686877e-06, 5.027577e-06, 2.84829e-06, 
    1.163874e-06, 2.392447e-06, 3.602087e-06, 8.258186e-07, 1.941178e-06, 
    3.932431e-06, 1.203968e-05, 1.572665e-05, 7.331143e-06, 1.209711e-05,
  1.069015e-05, 8.407412e-06, 7.863452e-06, 5.292284e-06, 4.341352e-06, 
    3.322802e-06, 3.968591e-06, 4.492953e-06, 2.746135e-06, 7.017509e-07, 
    4.116968e-06, 9.579036e-06, 1.75071e-05, 1.106592e-05, 1.152168e-05,
  1.165329e-05, 1.045753e-05, 1.011491e-05, 8.229687e-06, 5.331568e-06, 
    3.921716e-06, 2.070176e-06, 3.412246e-06, 3.287252e-06, 5.716406e-07, 
    4.8459e-06, 1.189193e-05, 1.504752e-05, 1.256743e-05, 1.260549e-05,
  1.334872e-05, 9.863677e-06, 1.027268e-05, 7.409521e-06, 5.885984e-06, 
    5.227252e-06, 2.266144e-06, 4.311607e-06, 5.753923e-06, 3.804302e-06, 
    5.784598e-06, 1.159408e-05, 1.60612e-05, 1.209314e-05, 1.171668e-05,
  1.516431e-05, 1.267191e-05, 1.182347e-05, 1.06111e-05, 8.012295e-06, 
    5.980053e-06, 5.547832e-06, 4.296452e-06, 6.681192e-06, 2.570825e-06, 
    8.252894e-06, 1.35804e-05, 1.707642e-05, 1.223595e-05, 1.264753e-05,
  1.628835e-05, 1.263765e-05, 1.282999e-05, 1.17677e-05, 9.558089e-06, 
    8.889058e-06, 7.882036e-06, 4.772554e-06, 4.010944e-06, 4.516195e-06, 
    1.109596e-05, 1.596647e-05, 1.623401e-05, 1.575753e-05, 1.583783e-05,
  1.801643e-05, 1.293986e-05, 1.245766e-05, 1.193203e-05, 9.528228e-06, 
    8.015253e-06, 7.104298e-06, 7.310795e-06, 5.990097e-06, 1.101614e-05, 
    1.807272e-05, 1.98076e-05, 1.891975e-05, 1.928053e-05, 1.509481e-05,
  1.835832e-05, 1.497242e-05, 1.42005e-05, 1.319584e-05, 8.959718e-06, 
    8.206262e-06, 6.498723e-06, 4.151174e-06, 9.174756e-06, 2.202753e-05, 
    2.747195e-05, 2.27774e-05, 2.730263e-05, 1.955843e-05, 1.751146e-05,
  5.66971e-06, 7.001236e-06, 6.962925e-06, 7.433517e-06, 5.327166e-06, 
    8.427165e-06, 6.158249e-06, 4.077979e-06, 2.512935e-06, 2.560479e-07, 
    1.885573e-06, 4.056129e-06, 9.030628e-06, 1.067933e-05, 7.890252e-06,
  5.929262e-06, 6.668656e-06, 7.99607e-06, 6.563781e-06, 1.046852e-05, 
    8.523316e-06, 5.567377e-06, 3.3449e-06, 1.462577e-06, 2.218398e-07, 
    2.091844e-07, 3.040476e-06, 7.030045e-06, 8.372458e-06, 4.696597e-06,
  7.828407e-06, 7.569044e-06, 9.626099e-06, 8.765901e-06, 9.702306e-06, 
    9.135282e-06, 5.235823e-06, 3.789637e-06, 1.193863e-06, 1.000267e-06, 
    3.528556e-07, 3.342525e-06, 6.13962e-06, 2.008713e-06, 2.304778e-06,
  9.264063e-06, 7.202448e-06, 1.106369e-05, 8.595533e-06, 9.45058e-06, 
    6.86901e-06, 4.650126e-06, 3.332073e-06, 1.484653e-06, 1.2676e-06, 
    1.143e-06, 1.321083e-06, 4.930639e-06, 1.312158e-06, 2.186177e-06,
  6.796983e-06, 8.480654e-06, 8.786948e-06, 8.730205e-06, 6.088045e-06, 
    3.797554e-06, 4.036459e-06, 3.63998e-06, 3.632643e-06, 1.621687e-06, 
    1.641224e-06, 1.250138e-06, 4.560813e-06, 6.444508e-07, 3.673668e-06,
  5.198385e-06, 6.136634e-06, 6.30164e-06, 7.049609e-06, 6.333796e-06, 
    3.166178e-06, 2.689724e-06, 1.657499e-06, 2.808782e-06, 1.125326e-06, 
    9.034091e-07, 1.521005e-06, 2.07488e-06, 7.530293e-07, 4.490778e-06,
  3.156138e-06, 5.290443e-06, 3.757404e-06, 4.489772e-06, 4.771188e-06, 
    2.941599e-06, 1.334946e-06, 2.109802e-06, 1.29641e-06, 7.48375e-07, 
    3.318671e-07, 7.927119e-07, 6.977275e-07, 9.323655e-07, 4.923029e-06,
  4.965281e-06, 4.413268e-06, 2.901879e-06, 2.944983e-06, 3.520555e-06, 
    2.064438e-06, 1.813336e-06, 1.277373e-06, 6.491649e-07, 1.595624e-07, 
    5.481006e-07, 1.28026e-07, 5.3554e-07, 2.565114e-06, 5.301536e-06,
  4.772386e-06, 3.503661e-06, 2.495098e-06, 3.159854e-06, 2.32124e-06, 
    1.545319e-06, 6.584189e-07, 8.599172e-07, 1.425778e-06, 1.436236e-06, 
    6.094746e-07, 1.683395e-07, 1.30851e-06, 6.353189e-06, 5.647587e-06,
  5.553532e-06, 3.07141e-06, 3.605877e-06, 2.701161e-06, 2.674761e-06, 
    1.833627e-06, 1.450912e-06, 1.019048e-06, 2.612545e-06, 1.011953e-06, 
    1.067677e-06, 4.811734e-07, 2.498062e-06, 6.928658e-06, 6.666002e-06,
  0.000183867, 4.463392e-05, 1.251042e-05, 4.819652e-06, 3.719937e-06, 
    5.29253e-06, 7.922284e-06, 6.612601e-06, 7.626489e-06, 6.405733e-06, 
    9.803353e-06, 8.7482e-06, 7.381691e-06, 7.746803e-06, 6.065303e-06,
  0.0001939921, 4.928066e-05, 1.231839e-05, 5.447971e-06, 4.984123e-06, 
    5.025979e-06, 5.86111e-06, 8.607174e-06, 6.76358e-06, 4.568045e-06, 
    6.152739e-06, 7.428062e-06, 8.182979e-06, 9.012346e-06, 5.958146e-06,
  0.0001890517, 4.477827e-05, 1.10393e-05, 5.706566e-06, 7.06264e-06, 
    4.725275e-06, 3.461015e-06, 8.789137e-06, 2.841243e-06, 6.113064e-06, 
    5.11541e-06, 7.822107e-06, 6.282067e-06, 9.270359e-06, 6.497665e-06,
  0.0001648242, 2.956495e-05, 9.846092e-06, 6.265993e-06, 6.539321e-06, 
    4.16881e-06, 6.296577e-06, 4.788913e-06, 5.035961e-06, 7.795879e-06, 
    5.295909e-06, 9.291268e-06, 7.228396e-06, 8.071385e-06, 6.702051e-06,
  0.0001350047, 1.33721e-05, 6.313114e-06, 5.213112e-06, 3.51423e-06, 
    5.516512e-06, 4.719698e-06, 8.108488e-06, 5.790539e-06, 5.29309e-06, 
    5.705936e-06, 4.74016e-06, 7.731292e-06, 6.817029e-06, 7.599989e-06,
  0.0001052508, 8.798694e-06, 6.726581e-06, 6.064128e-06, 5.015685e-06, 
    5.18094e-06, 5.937429e-06, 5.569587e-06, 7.39939e-06, 2.621328e-06, 
    2.825552e-06, 4.699123e-06, 6.45631e-06, 8.93893e-06, 8.918721e-06,
  7.319631e-05, 7.885214e-06, 5.816952e-06, 5.625622e-06, 7.279563e-06, 
    8.785059e-06, 4.068149e-06, 5.364586e-06, 6.442295e-06, 1.11278e-06, 
    3.536171e-06, 5.69884e-06, 6.795901e-06, 8.363379e-06, 7.908832e-06,
  4.18218e-05, 5.482226e-06, 5.855562e-06, 8.728891e-06, 8.182953e-06, 
    8.136178e-06, 1.675465e-06, 6.319378e-06, 4.923289e-06, 1.816722e-06, 
    2.065005e-06, 3.118402e-06, 6.361766e-06, 8.866494e-06, 8.945623e-06,
  1.604325e-05, 5.056673e-06, 7.348203e-06, 1.095355e-05, 1.163052e-05, 
    5.502473e-06, 4.272043e-06, 4.813031e-06, 1.597404e-06, 7.017588e-07, 
    1.025594e-06, 4.25993e-06, 5.745178e-06, 8.602377e-06, 8.688466e-06,
  7.173724e-06, 6.460202e-06, 9.483608e-06, 1.269053e-05, 1.015288e-05, 
    4.255556e-06, 4.935308e-06, 3.579495e-06, 1.178565e-06, 3.903058e-07, 
    1.07796e-06, 4.123442e-06, 6.089777e-06, 8.856832e-06, 1.233632e-05,
  4.18236e-06, 1.362873e-05, 1.234308e-05, 6.355377e-06, 1.1645e-05, 
    1.334229e-05, 9.278435e-06, 3.359924e-06, 3.038668e-06, 4.572561e-06, 
    8.14123e-06, 8.514108e-06, 7.463305e-06, 6.651568e-06, 5.960112e-06,
  1.550232e-05, 3.25255e-05, 3.314255e-05, 1.736755e-05, 1.795319e-05, 
    1.729863e-05, 6.778365e-06, 4.134079e-07, 1.139691e-06, 4.401317e-06, 
    6.893554e-06, 9.421494e-06, 8.578685e-06, 6.115541e-06, 5.440244e-06,
  2.965925e-05, 5.018189e-05, 4.828162e-05, 2.561501e-05, 2.089745e-05, 
    2.06405e-05, 5.278679e-06, 2.643693e-07, 5.708383e-06, 2.74273e-06, 
    1.052519e-05, 1.34371e-05, 8.788233e-06, 5.798851e-06, 3.509638e-06,
  5.394061e-05, 5.284213e-05, 4.673756e-05, 3.083011e-05, 2.192964e-05, 
    1.62131e-05, 6.246467e-06, 2.675795e-06, 3.070763e-06, 3.272212e-06, 
    7.571237e-06, 1.044263e-05, 9.970998e-06, 7.13172e-06, 7.950474e-06,
  8.415045e-05, 5.123459e-05, 3.96342e-05, 3.314126e-05, 1.963983e-05, 
    1.465736e-05, 2.622731e-06, 2.955358e-06, 2.918927e-06, 4.58196e-06, 
    8.887581e-06, 1.002239e-05, 1.068474e-05, 6.990836e-06, 6.189983e-06,
  0.0001040292, 4.129403e-05, 3.113253e-05, 3.409857e-05, 2.366352e-05, 
    8.508531e-06, 3.767052e-06, 1.792854e-06, 3.409083e-06, 3.467906e-06, 
    4.836884e-06, 7.041072e-06, 8.324689e-06, 6.366276e-06, 6.408809e-06,
  0.0001092104, 3.10007e-05, 2.748142e-05, 3.196099e-05, 2.499547e-05, 
    1.064504e-05, 4.585063e-06, 2.392949e-06, 1.955827e-06, 2.546979e-06, 
    2.886025e-06, 5.780419e-06, 6.366879e-06, 7.53652e-06, 7.665307e-06,
  0.0001072838, 2.41297e-05, 2.67813e-05, 2.83483e-05, 2.254524e-05, 
    1.162532e-05, 7.81654e-06, 2.40758e-06, 1.574962e-06, 2.020015e-06, 
    5.203718e-06, 5.868737e-06, 7.788921e-06, 8.684481e-06, 6.750957e-06,
  9.31093e-05, 1.995331e-05, 2.36539e-05, 2.361807e-05, 1.967634e-05, 
    9.403047e-06, 9.967131e-06, 2.83011e-06, 1.617053e-06, 2.309194e-06, 
    4.783425e-06, 5.674151e-06, 6.51732e-06, 7.986831e-06, 4.910575e-06,
  8.023202e-05, 1.612726e-05, 2.046763e-05, 1.920721e-05, 1.459153e-05, 
    1.178202e-05, 6.160279e-06, 4.301385e-06, 2.097746e-06, 5.683182e-06, 
    5.615307e-06, 4.479493e-06, 6.283486e-06, 5.502437e-06, 4.746162e-06,
  5.873326e-07, 1.561668e-06, 2.075759e-06, 1.215728e-06, 1.8145e-06, 
    1.709011e-06, 2.741754e-06, 4.896573e-06, 5.231873e-06, 6.96134e-06, 
    8.518832e-06, 6.659398e-06, 4.974656e-06, 4.440428e-06, 3.637003e-06,
  5.936569e-09, 1.262169e-08, 5.333116e-08, 4.715376e-07, 2.002689e-06, 
    1.87371e-06, 3.528447e-06, 3.519118e-06, 2.846614e-06, 4.487418e-06, 
    7.051138e-06, 7.902877e-06, 5.791984e-06, 5.72023e-06, 4.527756e-06,
  8.075669e-09, 2.97395e-08, 2.088203e-07, 3.839627e-07, 1.157022e-06, 
    5.361459e-06, 2.074574e-06, 3.368008e-06, 2.90315e-06, 3.96328e-06, 
    6.156817e-06, 7.09262e-06, 7.404219e-06, 6.604419e-06, 6.006318e-06,
  2.432431e-09, 3.862008e-09, 8.717089e-09, 4.092331e-08, 1.013152e-06, 
    4.592075e-06, 3.598405e-06, 3.308676e-06, 2.957255e-06, 5.018407e-06, 
    5.912863e-06, 7.407261e-06, 6.798549e-06, 7.426815e-06, 6.348796e-06,
  1.713469e-09, 3.095686e-09, 2.508808e-09, 2.818176e-08, 1.115456e-06, 
    2.011269e-06, 4.679422e-06, 3.707037e-06, 1.921221e-06, 3.168882e-06, 
    4.059371e-06, 6.125176e-06, 8.023228e-06, 9.054603e-06, 9.661476e-06,
  6.145195e-09, 1.170102e-09, 7.624601e-10, 6.743378e-09, 1.345663e-09, 
    6.457911e-07, 2.194671e-06, 5.630081e-06, 3.085614e-06, 3.866769e-06, 
    3.448847e-06, 7.321762e-06, 9.197398e-06, 1.218665e-05, 7.824946e-06,
  1.243976e-08, 6.95852e-10, 2.392114e-09, 8.918661e-09, 4.061359e-08, 
    2.813504e-07, 5.250584e-06, 4.633006e-06, 3.619695e-06, 3.406871e-06, 
    4.107762e-06, 7.156298e-06, 8.665319e-06, 8.000499e-06, 7.079494e-06,
  2.442145e-08, 1.466825e-09, 2.180757e-09, 2.281368e-09, 1.024401e-08, 
    1.161972e-07, 4.194345e-06, 5.434816e-06, 5.609152e-06, 3.605292e-06, 
    4.642359e-06, 7.045241e-06, 9.043083e-06, 9.160483e-06, 1.084076e-05,
  3.363298e-08, 1.929302e-09, 8.092498e-10, 6.484578e-09, 7.514949e-09, 
    6.782182e-08, 1.899551e-06, 1.01761e-05, 6.858897e-06, 3.926297e-06, 
    6.072421e-06, 5.594651e-06, 1.109734e-05, 1.254573e-05, 1.046997e-05,
  2.624265e-08, 4.091364e-09, 3.703914e-09, 6.247181e-09, 2.096801e-08, 
    1.200983e-08, 4.576881e-07, 7.416696e-06, 7.295585e-06, 6.920685e-06, 
    6.631798e-06, 6.628712e-06, 1.164429e-05, 1.235982e-05, 1.252472e-05,
  8.395669e-07, 3.275322e-07, 1.585006e-08, 1.82399e-08, 1.2727e-08, 
    1.047837e-08, 3.135864e-06, 5.62176e-06, 4.191538e-06, 4.912529e-06, 
    7.78233e-06, 7.916253e-06, 9.069357e-06, 8.58088e-06, 8.456581e-06,
  8.36041e-07, 1.48718e-06, 9.945891e-07, 1.798421e-07, 6.34798e-09, 
    3.692753e-07, 1.919746e-06, 3.519529e-06, 2.647575e-06, 3.280619e-06, 
    5.037247e-06, 7.312689e-06, 7.882288e-06, 1.145312e-05, 9.171368e-06,
  6.106457e-06, 8.515292e-06, 5.983559e-06, 1.469322e-06, 3.828604e-07, 
    1.066552e-06, 1.761889e-06, 2.744668e-06, 9.404868e-07, 3.859203e-06, 
    5.341511e-06, 6.800064e-06, 8.495374e-06, 8.622104e-06, 9.914622e-06,
  7.802225e-06, 7.218208e-06, 5.017194e-06, 1.769004e-06, 1.211561e-06, 
    2.92455e-07, 1.277233e-06, 2.185882e-06, 2.820938e-06, 4.049199e-06, 
    5.72033e-06, 6.120561e-06, 6.293906e-06, 7.807476e-06, 9.304081e-06,
  2.338873e-06, 4.775079e-07, 5.586121e-08, 2.207088e-08, 1.18533e-06, 
    1.802022e-06, 3.953398e-06, 2.354282e-06, 3.403761e-06, 3.573405e-06, 
    4.778227e-06, 6.652809e-06, 7.308383e-06, 9.287877e-06, 1.082516e-05,
  1.022123e-08, 5.641587e-09, 4.72012e-09, 6.09614e-09, 4.021394e-07, 
    1.975848e-06, 1.270252e-06, 4.269684e-06, 2.936884e-06, 4.071108e-06, 
    6.375018e-06, 6.694198e-06, 5.248074e-06, 9.041328e-06, 7.71905e-06,
  2.235061e-08, 5.879927e-08, 2.790541e-07, 2.026211e-07, 3.613793e-07, 
    8.113727e-07, 2.099518e-06, 3.963006e-06, 6.649943e-06, 6.021583e-06, 
    7.023907e-06, 7.785134e-06, 7.193174e-06, 8.685327e-06, 9.437748e-06,
  3.630746e-08, 5.136142e-08, 6.506518e-07, 1.930016e-06, 2.552205e-06, 
    6.927261e-06, 4.621307e-06, 6.873805e-06, 9.012184e-06, 5.874106e-06, 
    6.454325e-06, 6.753889e-06, 7.677833e-06, 7.807766e-06, 1.096405e-05,
  9.994178e-08, 1.161624e-07, 2.249418e-07, 1.473786e-07, 1.987502e-07, 
    7.478884e-07, 3.892469e-06, 5.802059e-06, 5.833292e-06, 8.59187e-06, 
    1.067625e-05, 9.197895e-06, 8.270757e-06, 8.443988e-06, 1.267849e-05,
  1.858169e-08, 1.179891e-08, 1.683586e-08, 6.69825e-09, 6.823302e-09, 
    7.85564e-09, 4.074157e-08, 6.661638e-07, 9.484519e-06, 9.817856e-06, 
    8.207942e-06, 8.999252e-06, 7.820165e-06, 8.791956e-06, 1.073987e-05,
  0.0002011121, 0.0001740253, 0.0001730166, 0.0001606382, 0.0001468373, 
    0.000129475, 0.0001002238, 8.049484e-05, 5.943434e-05, 8.224008e-05, 
    7.270509e-05, 5.166122e-05, 2.943881e-05, 1.705524e-05, 9.246422e-06,
  0.0001396603, 0.0001478803, 0.0001533235, 0.0001393809, 0.0001214692, 
    9.58692e-05, 7.622794e-05, 5.96726e-05, 6.521709e-05, 5.65944e-05, 
    3.555021e-05, 2.643075e-05, 9.398922e-06, 7.877613e-06, 6.112429e-06,
  5.565632e-05, 6.602142e-05, 6.745518e-05, 6.404839e-05, 5.88405e-05, 
    4.634364e-05, 3.847137e-05, 3.085766e-05, 2.344466e-05, 1.507626e-05, 
    1.043775e-05, 6.893428e-06, 5.091656e-06, 7.096647e-06, 5.545686e-06,
  4.277953e-06, 5.092012e-06, 7.581382e-06, 1.071206e-05, 1.214742e-05, 
    8.521733e-06, 4.774451e-06, 2.816981e-06, 1.808462e-06, 3.196202e-06, 
    4.895712e-06, 6.399112e-06, 6.432883e-06, 6.364844e-06, 6.479397e-06,
  8.279669e-07, 6.670821e-07, 2.116537e-06, 3.728597e-06, 5.497706e-06, 
    7.171018e-06, 7.72613e-06, 8.179269e-06, 6.014798e-06, 3.314663e-06, 
    5.523399e-06, 7.376659e-06, 6.290927e-06, 6.198091e-06, 5.187005e-06,
  3.383433e-06, 2.680976e-06, 9.713351e-07, 3.32477e-07, 7.162698e-07, 
    2.441759e-06, 3.709078e-06, 6.099009e-06, 6.076727e-06, 5.199667e-06, 
    9.361828e-06, 7.190736e-06, 6.579359e-06, 7.328712e-06, 7.556209e-06,
  6.249603e-07, 1.614064e-06, 2.927792e-06, 3.178109e-06, 3.322894e-06, 
    4.487104e-06, 3.673895e-06, 3.112835e-06, 4.171541e-06, 5.388124e-06, 
    8.998706e-06, 8.989598e-06, 9.462156e-06, 1.029778e-05, 7.784407e-06,
  2.667292e-07, 7.893271e-07, 2.188591e-06, 3.700496e-06, 3.989729e-06, 
    9.830179e-06, 1.296007e-05, 8.127305e-06, 4.756573e-06, 5.823409e-06, 
    5.119585e-06, 7.142285e-06, 8.16514e-06, 7.974755e-06, 7.527094e-06,
  1.188912e-07, 5.311804e-07, 7.281586e-07, 1.718323e-06, 2.866665e-06, 
    2.96902e-06, 7.495457e-06, 1.294759e-05, 1.131938e-05, 7.525524e-06, 
    9.446172e-06, 8.494199e-06, 7.320733e-06, 7.012994e-06, 7.885138e-06,
  3.971458e-08, 3.465442e-08, 7.682166e-08, 2.508204e-07, 7.318291e-07, 
    1.917976e-06, 3.461614e-06, 8.048202e-06, 7.045867e-06, 9.728856e-06, 
    1.138198e-05, 1.032355e-05, 8.572001e-06, 4.688816e-06, 6.443535e-06,
  6.321228e-06, 3.909376e-06, 2.512881e-06, 1.176377e-06, 4.887283e-07, 
    2.991383e-07, 3.662121e-07, 2.249795e-07, 1.396156e-07, 1.850418e-08, 
    8.365618e-08, 1.807176e-06, 7.730036e-06, 1.320478e-05, 2.379178e-05,
  2.502491e-05, 3.070258e-06, 1.531156e-06, 2.071083e-07, 7.387211e-08, 
    6.715915e-09, 5.136599e-09, 8.330661e-09, 1.056428e-07, 2.486959e-06, 
    6.851595e-06, 1.579209e-05, 1.4524e-05, 2.47343e-05, 4.484709e-05,
  8.43754e-05, 4.388875e-05, 2.500086e-05, 1.219524e-05, 5.741117e-06, 
    2.957873e-06, 3.390765e-06, 6.705392e-06, 1.113326e-05, 1.674446e-05, 
    1.811837e-05, 1.547866e-05, 1.59253e-05, 2.884037e-05, 2.348918e-05,
  8.656506e-05, 6.955348e-05, 5.678256e-05, 4.283224e-05, 3.007674e-05, 
    2.463856e-05, 2.256109e-05, 2.043833e-05, 2.064168e-05, 1.840006e-05, 
    1.746762e-05, 1.2285e-05, 2.41838e-05, 3.338627e-05, 1.654011e-05,
  5.471898e-05, 4.958172e-05, 4.010445e-05, 3.190583e-05, 2.695265e-05, 
    2.328405e-05, 1.998875e-05, 1.588426e-05, 1.488374e-05, 1.347795e-05, 
    1.500449e-05, 1.802466e-05, 2.788341e-05, 2.471411e-05, 6.476783e-06,
  2.824118e-05, 2.990372e-05, 2.682983e-05, 2.061891e-05, 1.580013e-05, 
    1.338523e-05, 1.200275e-05, 1.092827e-05, 8.092195e-06, 1.221077e-05, 
    2.255848e-05, 2.966521e-05, 2.652209e-05, 1.009249e-05, 9.102786e-07,
  1.042212e-05, 1.286005e-05, 1.243092e-05, 1.101056e-05, 1.005238e-05, 
    7.881513e-06, 7.976181e-06, 8.637876e-06, 1.711559e-05, 2.925631e-05, 
    3.552094e-05, 3.12243e-05, 1.438583e-05, 2.722119e-06, 3.865725e-07,
  4.137238e-06, 5.23538e-06, 5.740528e-06, 6.737234e-06, 7.810635e-06, 
    1.418691e-05, 1.669279e-05, 2.346955e-05, 2.837377e-05, 3.402915e-05, 
    2.267629e-05, 8.975255e-06, 2.986275e-06, 7.064457e-08, 1.51051e-07,
  1.825236e-06, 2.236167e-06, 3.224087e-06, 5.379219e-06, 6.873948e-06, 
    1.326576e-05, 1.643636e-05, 1.609751e-05, 1.084575e-05, 6.367308e-06, 
    1.786795e-06, 5.422916e-08, 3.587492e-09, 1.149287e-06, 2.118303e-06,
  1.737604e-06, 1.604422e-06, 8.982273e-07, 2.725104e-06, 2.166434e-06, 
    5.456852e-06, 3.89838e-06, 3.023298e-06, 1.927491e-06, 1.888215e-06, 
    1.49748e-06, 4.179886e-07, 5.293888e-08, 9.877953e-07, 1.604369e-06,
  3.193884e-06, 6.882342e-06, 7.324075e-06, 8.479708e-06, 1.145733e-05, 
    9.276883e-06, 8.806138e-06, 8.741514e-06, 8.282925e-06, 6.919689e-06, 
    6.597159e-06, 4.355408e-06, 5.506048e-06, 2.58189e-05, 3.986959e-05,
  4.399677e-06, 4.37483e-06, 5.296388e-06, 8.674818e-06, 6.989223e-06, 
    8.530227e-06, 9.40796e-06, 8.112998e-06, 7.1974e-06, 3.600549e-06, 
    3.179321e-06, 6.353014e-07, 1.462311e-05, 4.964686e-05, 5.868442e-05,
  3.154048e-06, 3.273507e-06, 3.521211e-06, 5.927863e-06, 7.810389e-06, 
    9.518241e-06, 7.00565e-06, 5.099252e-06, 1.875351e-06, 2.670017e-06, 
    3.078902e-06, 3.501874e-06, 2.269541e-05, 5.88016e-05, 3.954433e-05,
  1.13124e-06, 1.319565e-06, 1.478317e-06, 4.196194e-06, 5.288977e-06, 
    3.259587e-06, 2.670868e-06, 1.597748e-06, 2.301131e-06, 3.151515e-06, 
    2.824816e-07, 3.784627e-06, 2.19916e-05, 5.556273e-05, 2.860818e-05,
  3.077998e-07, 5.770385e-07, 3.665285e-07, 1.223732e-06, 2.779492e-06, 
    1.786336e-06, 7.249817e-07, 2.325177e-06, 1.89741e-06, 2.122341e-06, 
    2.235789e-06, 5.725468e-06, 2.745059e-05, 4.952707e-05, 1.654909e-05,
  1.190329e-08, 1.20919e-07, 1.313887e-07, 5.599444e-07, 1.685594e-06, 
    2.21122e-06, 1.756647e-06, 3.277149e-06, 3.144432e-06, 4.219308e-06, 
    7.051267e-06, 2.063664e-05, 3.432684e-05, 1.772675e-05, 1.194373e-05,
  1.663415e-10, 2.473998e-09, 1.17238e-08, 2.129578e-07, 1.423222e-06, 
    2.448155e-06, 2.74174e-06, 1.240438e-06, 7.989232e-06, 1.64492e-05, 
    2.317057e-05, 3.189577e-05, 3.75856e-05, 1.506165e-05, 1.085818e-05,
  4.681098e-10, 2.356174e-09, 2.771748e-08, 3.133817e-07, 2.380661e-06, 
    3.859544e-06, 4.780698e-06, 5.090484e-06, 1.516553e-05, 2.794622e-05, 
    3.444603e-05, 3.834194e-05, 2.190404e-05, 1.349405e-05, 7.542551e-06,
  1.637665e-07, 3.570169e-07, 1.248559e-06, 1.057978e-06, 4.821462e-06, 
    5.782894e-06, 1.127091e-05, 1.273404e-05, 1.504178e-05, 2.462899e-05, 
    1.607898e-05, 1.259092e-05, 1.028025e-05, 5.19627e-06, 4.004585e-06,
  3.279202e-06, 3.794691e-06, 5.803098e-06, 9.269639e-06, 6.574445e-06, 
    8.401616e-06, 7.426241e-06, 1.181544e-05, 9.927917e-06, 6.901613e-06, 
    8.681765e-06, 5.013977e-06, 4.146665e-06, 2.757919e-06, 3.818286e-06,
  1.175314e-05, 9.611445e-06, 9.448619e-06, 7.656989e-06, 7.560441e-06, 
    7.652571e-06, 9.99889e-06, 9.921134e-06, 5.529618e-06, 4.939884e-06, 
    1.223713e-05, 2.829844e-05, 2.89782e-05, 2.128358e-05, 7.597512e-06,
  1.096917e-05, 1.311092e-05, 1.13145e-05, 7.649331e-06, 7.885171e-06, 
    6.370077e-06, 1.063419e-05, 1.025526e-05, 6.517265e-06, 2.379429e-06, 
    8.111723e-06, 2.062787e-05, 3.36232e-05, 2.009921e-05, 7.562061e-06,
  6.224189e-06, 1.068825e-05, 1.198399e-05, 6.353695e-06, 5.839051e-06, 
    8.459197e-06, 9.511928e-06, 9.264968e-06, 9.289945e-06, 6.002778e-06, 
    7.202438e-06, 1.59929e-05, 2.717158e-05, 2.00439e-05, 1.028827e-05,
  3.66457e-06, 4.398713e-06, 6.871854e-06, 6.340829e-06, 5.096477e-06, 
    7.531738e-06, 8.32451e-06, 8.830031e-06, 1.028553e-05, 8.163427e-06, 
    9.143239e-06, 1.795381e-05, 2.631414e-05, 1.926057e-05, 7.545244e-06,
  2.116196e-06, 8.725074e-07, 4.796969e-06, 4.301743e-06, 1.541914e-05, 
    1.20511e-05, 5.510065e-06, 7.413196e-06, 8.065963e-06, 9.230394e-06, 
    1.227652e-05, 1.942636e-05, 2.462792e-05, 1.677573e-05, 6.076662e-06,
  2.036176e-06, 6.831001e-06, 1.216415e-05, 5.070735e-06, 1.636582e-05, 
    1.58996e-05, 7.973288e-06, 7.764519e-06, 5.456787e-06, 1.115367e-05, 
    1.767059e-05, 2.021045e-05, 2.187752e-05, 1.237952e-05, 5.857097e-06,
  1.228533e-07, 5.175386e-07, 7.904064e-06, 1.160438e-05, 1.769314e-05, 
    1.61279e-05, 1.5252e-05, 6.930547e-06, 3.386261e-06, 3.927922e-06, 
    1.157667e-05, 2.012818e-05, 1.499927e-05, 5.882919e-06, 4.780794e-06,
  5.050028e-08, 2.182314e-07, 1.39686e-06, 9.045597e-06, 1.54397e-05, 
    1.880153e-05, 1.882558e-05, 8.566926e-06, 4.795304e-06, 4.45876e-06, 
    4.732477e-06, 1.12072e-05, 6.638816e-06, 4.564718e-06, 3.168535e-06,
  1.459028e-08, 1.079455e-07, 2.640349e-07, 3.612766e-06, 1.168534e-05, 
    1.414417e-05, 1.70486e-05, 1.470396e-05, 8.615939e-06, 3.183967e-06, 
    2.001724e-06, 1.585063e-06, 2.820396e-06, 4.577962e-06, 3.528358e-06,
  1.91666e-08, 4.27882e-07, 2.924876e-06, 4.022711e-06, 6.139332e-06, 
    9.027077e-06, 1.291824e-05, 1.262704e-05, 1.318626e-05, 7.540642e-06, 
    4.563738e-06, 2.182559e-06, 2.33051e-06, 5.684369e-06, 5.462859e-06,
  1.899606e-05, 1.47193e-05, 9.238831e-06, 4.196351e-06, 2.706464e-06, 
    1.419244e-06, 4.828743e-06, 3.109357e-05, 2.864655e-05, 1.724416e-05, 
    1.419647e-05, 8.791479e-06, 7.951729e-06, 8.183589e-06, 1.133258e-05,
  7.991078e-06, 4.974511e-06, 1.357387e-06, 1.508077e-07, 5.68084e-07, 
    3.947864e-06, 2.234714e-06, 1.087452e-05, 1.323815e-05, 2.157137e-05, 
    1.484084e-05, 9.811643e-06, 7.269944e-06, 8.711851e-06, 1.186465e-05,
  4.694128e-06, 4.795243e-06, 2.192211e-06, 5.609975e-07, 3.153865e-07, 
    3.095167e-07, 1.432663e-06, 1.608531e-06, 6.294543e-06, 1.083018e-05, 
    1.262948e-05, 1.10797e-05, 5.630192e-06, 6.882152e-06, 1.002878e-05,
  7.804416e-06, 5.590699e-06, 3.495178e-06, 2.473258e-06, 1.916724e-06, 
    5.049549e-07, 5.680762e-07, 8.857861e-08, 4.888991e-06, 5.378794e-06, 
    5.922532e-06, 6.706793e-06, 3.999675e-06, 5.306984e-06, 6.975788e-06,
  1.031973e-05, 1.074777e-05, 6.412222e-06, 6.008152e-06, 3.727413e-06, 
    2.770194e-06, 8.090597e-07, 1.895371e-07, 1.369809e-07, 6.92021e-07, 
    1.582619e-06, 3.563739e-06, 6.193048e-06, 6.612388e-06, 5.479099e-06,
  1.49734e-05, 1.199742e-05, 1.240095e-05, 1.147548e-05, 8.401572e-06, 
    7.104175e-06, 5.64249e-06, 4.350839e-06, 3.658256e-07, 4.027774e-06, 
    2.637609e-06, 3.721895e-06, 5.417359e-06, 3.533832e-06, 5.758104e-06,
  5.739616e-06, 9.162986e-06, 1.118763e-05, 1.205282e-05, 1.363156e-05, 
    1.048853e-05, 6.808458e-06, 7.833889e-06, 5.974082e-06, 3.160892e-06, 
    3.115223e-06, 5.217497e-06, 5.435655e-06, 5.110581e-06, 7.438065e-06,
  9.159295e-06, 1.290384e-05, 1.160959e-05, 1.114995e-05, 1.059556e-05, 
    9.179053e-06, 9.739894e-06, 9.715836e-06, 6.390102e-06, 6.412643e-06, 
    7.740951e-06, 6.812602e-06, 7.59551e-06, 5.342719e-06, 1.013443e-05,
  1.108026e-05, 1.378976e-05, 1.878388e-05, 1.958572e-05, 1.225019e-05, 
    6.875488e-06, 9.322762e-06, 8.708815e-06, 8.653272e-06, 9.068706e-06, 
    7.889594e-06, 4.943045e-06, 3.93292e-06, 6.509878e-06, 5.36421e-06,
  1.140677e-05, 1.79525e-05, 1.700295e-05, 1.396829e-05, 1.453765e-05, 
    1.443949e-05, 1.411346e-05, 5.513361e-06, 5.503333e-06, 1.148175e-05, 
    1.143032e-05, 1.155108e-05, 4.141828e-06, 3.74287e-06, 4.347466e-06,
  2.278475e-05, 2.252536e-05, 2.262603e-05, 2.497993e-05, 3.951549e-05, 
    5.351657e-05, 0.0001250757, 7.791191e-05, 6.557177e-05, 6.697563e-05, 
    3.504982e-05, 1.248365e-05, 3.350732e-05, 2.679449e-05, 1.700904e-05,
  3.746429e-05, 3.581526e-05, 3.25591e-05, 6.144738e-05, 7.950272e-05, 
    5.148894e-05, 5.982246e-06, 2.132981e-06, 1.421378e-05, 2.201685e-05, 
    1.381819e-05, 9.80491e-06, 8.027985e-06, 1.074814e-05, 1.246303e-05,
  3.305086e-05, 3.492645e-05, 6.921355e-05, 7.411157e-05, 2.677795e-05, 
    6.398896e-08, 1.299003e-08, 2.710247e-09, 2.682366e-07, 4.765742e-06, 
    8.381631e-06, 7.615661e-06, 5.160186e-06, 6.140875e-06, 8.073e-06,
  3.436532e-05, 5.210338e-05, 5.281708e-05, 1.179441e-05, 4.694268e-08, 
    1.06409e-08, 1.548418e-08, 3.229712e-08, 1.149662e-07, 1.683986e-06, 
    4.364586e-06, 6.24539e-06, 4.56901e-06, 4.884019e-06, 4.970046e-06,
  4.24303e-05, 2.438594e-05, 4.847391e-06, 1.184595e-07, 1.047955e-07, 
    5.534441e-07, 1.480071e-07, 1.360501e-07, 3.118969e-06, 1.57481e-06, 
    4.202271e-06, 4.064116e-06, 4.259065e-06, 4.353351e-06, 3.620287e-06,
  5.936532e-06, 9.885935e-07, 1.180434e-07, 5.718663e-08, 1.005212e-07, 
    3.871428e-07, 2.872117e-07, 2.240424e-06, 3.430856e-06, 2.084975e-06, 
    3.335901e-06, 4.243023e-06, 4.388822e-06, 5.404876e-06, 4.617675e-06,
  9.816609e-07, 1.218015e-06, 3.142861e-07, 7.432936e-07, 8.972011e-07, 
    2.51886e-06, 2.324699e-06, 4.253027e-06, 3.35557e-06, 3.500568e-06, 
    6.519791e-06, 6.469539e-06, 7.116086e-06, 5.668934e-06, 6.734654e-06,
  3.244148e-06, 4.019858e-06, 2.677893e-06, 2.614596e-06, 1.767802e-06, 
    1.848304e-06, 3.605392e-06, 4.983433e-06, 2.448062e-06, 2.582404e-06, 
    4.591397e-06, 5.697943e-06, 6.083143e-06, 6.964309e-06, 6.66026e-06,
  3.546979e-06, 2.333515e-06, 3.712574e-06, 2.949891e-06, 5.818307e-06, 
    2.550611e-06, 2.637115e-06, 3.441013e-06, 6.077415e-06, 3.613228e-06, 
    2.390349e-06, 2.544621e-06, 6.523997e-06, 6.708288e-06, 8.127327e-06,
  5.95197e-06, 5.385662e-06, 5.826043e-06, 5.490432e-06, 4.878018e-06, 
    3.748189e-06, 3.840967e-06, 5.07444e-06, 7.081226e-06, 5.371958e-06, 
    4.069469e-06, 6.357649e-06, 5.057931e-06, 7.085383e-06, 6.803537e-06,
  3.945888e-07, 1.776237e-06, 8.430041e-06, 5.289373e-05, 9.748861e-05, 
    7.979998e-05, 0.0001141591, 0.000165602, 0.0002655087, 0.0002216465, 
    0.0001886609, 7.537209e-05, 3.923358e-05, 1.458048e-05, 7.057511e-06,
  4.086287e-06, 4.099964e-05, 0.0001691031, 0.0002355627, 0.0002579349, 
    0.0002180685, 0.0002520174, 0.0002067471, 0.0002427926, 0.000131655, 
    7.519304e-05, 2.203956e-05, 1.004611e-05, 7.92966e-06, 8.332515e-06,
  0.0004415928, 0.000469855, 0.0004834857, 0.0003908461, 0.0002651549, 
    0.0001438618, 0.0001531844, 0.0001053461, 3.732929e-05, 1.886099e-05, 
    8.244971e-06, 4.950661e-06, 5.4725e-06, 6.693721e-06, 8.682192e-06,
  0.0004764225, 0.0004651276, 0.0003393514, 0.0001494229, 7.726644e-05, 
    4.734872e-05, 9.407792e-06, 3.375914e-06, 3.074235e-06, 5.664587e-06, 
    4.61037e-06, 5.22242e-06, 5.991535e-06, 9.476794e-06, 1.00914e-05,
  0.0001506671, 5.590574e-05, 1.906298e-05, 6.159548e-06, 3.358651e-07, 
    6.858487e-07, 3.116849e-06, 1.943226e-06, 1.683624e-06, 2.789919e-06, 
    5.55904e-06, 8.299723e-06, 1.003544e-05, 1.07919e-05, 9.288551e-06,
  1.94742e-05, 4.402143e-07, 1.412052e-07, 2.168081e-08, 7.05831e-09, 
    1.9222e-06, 3.339693e-06, 3.987577e-06, 3.964768e-06, 4.115825e-06, 
    5.987216e-06, 1.038359e-05, 9.881619e-06, 9.429928e-06, 8.444676e-06,
  1.405678e-06, 7.978936e-07, 1.352012e-07, 2.230425e-07, 8.533155e-07, 
    2.91847e-06, 3.794469e-06, 7.497616e-06, 6.506577e-06, 6.699202e-06, 
    8.909899e-06, 1.217604e-05, 1.207215e-05, 9.703153e-06, 1.169259e-05,
  1.975556e-06, 6.397484e-06, 2.699988e-06, 1.620103e-06, 1.316315e-06, 
    2.42252e-06, 1.494089e-06, 3.503614e-06, 6.874142e-06, 6.868129e-06, 
    9.284069e-06, 1.22666e-05, 1.128178e-05, 1.172946e-05, 1.094526e-05,
  1.238217e-06, 8.000673e-07, 1.652254e-06, 2.583358e-06, 2.202837e-06, 
    2.217585e-06, 3.490621e-06, 1.668056e-06, 2.933862e-06, 3.456643e-06, 
    8.428915e-06, 9.991092e-06, 1.008955e-05, 1.073223e-05, 1.074422e-05,
  2.900746e-06, 1.938645e-06, 4.286911e-06, 7.163605e-06, 6.636504e-06, 
    3.505983e-06, 4.160217e-06, 2.84683e-06, 5.66222e-06, 3.884935e-06, 
    3.763716e-06, 6.453794e-06, 6.980372e-06, 8.896955e-06, 8.158635e-06,
  2.207102e-05, 3.178971e-05, 3.494248e-05, 1.909417e-05, 1.200738e-05, 
    7.760116e-06, 5.598245e-06, 3.998175e-06, 4.213887e-06, 1.014506e-05, 
    2.54861e-05, 8.174564e-05, 0.0001081305, 9.060692e-05, 9.154713e-05,
  9.9672e-06, 1.0996e-05, 8.925728e-06, 1.28214e-05, 1.083003e-05, 
    6.133235e-06, 1.525447e-05, 3.093247e-05, 4.247984e-05, 5.103394e-05, 
    0.0001221447, 0.0001173914, 0.0001490999, 0.0001228762, 0.0001595484,
  4.394206e-05, 2.235758e-05, 2.519739e-05, 4.629999e-05, 8.437008e-05, 
    0.0001138945, 0.0001351355, 0.0001387536, 0.0002298884, 0.0002378595, 
    0.0002091851, 0.0001284402, 9.609499e-05, 0.0001332298, 0.00012683,
  0.0002139607, 0.0001792191, 0.0001990173, 0.0002416389, 0.0002692466, 
    0.0002635017, 0.0002449356, 0.000192603, 0.0002402836, 0.0001741776, 
    0.0001594787, 0.0001409882, 0.0001316512, 0.0001469418, 8.934076e-05,
  0.0002513287, 0.0002976531, 0.000325432, 0.0003360177, 0.0003156129, 
    0.0002620905, 0.0002013452, 0.0001555968, 0.0001671002, 0.0002303876, 
    0.0001987958, 0.0001717914, 0.000177475, 0.0001340745, 6.065014e-05,
  0.0003040253, 0.0002809603, 0.0002727091, 0.0002467739, 0.0002323177, 
    0.0002006437, 0.00016891, 0.0001462076, 0.0001982976, 0.000201258, 
    0.0002064902, 0.0002109596, 0.000191424, 9.723869e-05, 3.901051e-05,
  0.0003036798, 0.0003157992, 0.000278241, 0.0002198208, 0.0001730339, 
    0.0001515558, 0.0001409514, 0.0001505386, 0.0001936572, 0.0002090869, 
    0.0002353508, 0.0002299344, 0.0001681209, 6.83086e-05, 2.139303e-05,
  0.0001721701, 0.0002003047, 0.0001967009, 0.0001660347, 0.0001449619, 
    0.0001364438, 0.0001461527, 0.0001743565, 0.0002197351, 0.000263995, 
    0.0002772246, 0.0002170595, 9.381783e-05, 3.6299e-05, 1.314998e-05,
  9.480169e-05, 0.000133272, 0.0001434223, 0.0001409368, 0.0001498618, 
    0.0001630463, 0.0001970342, 0.0002376509, 0.0003057121, 0.0003031657, 
    0.000246373, 0.0001160442, 3.188847e-05, 1.083387e-05, 6.736983e-06,
  2.131816e-05, 5.448111e-05, 6.861702e-05, 7.323734e-05, 9.739678e-05, 
    0.0001462771, 0.000201682, 0.0002467272, 0.000237481, 0.0001864674, 
    9.163861e-05, 2.279514e-05, 8.515473e-06, 6.18314e-06, 5.163115e-06,
  0.0001129534, 7.586501e-05, 5.932876e-05, 2.869029e-05, 1.970211e-05, 
    1.771682e-05, 2.275043e-05, 2.258677e-05, 1.886249e-05, 1.149917e-05, 
    5.544886e-06, 2.897192e-06, 2.082318e-06, 4.005832e-06, 3.561971e-06,
  7.287742e-05, 6.402069e-05, 4.158731e-05, 2.914786e-05, 1.731207e-05, 
    1.561223e-05, 1.709741e-05, 1.612786e-05, 1.606153e-05, 1.232421e-05, 
    5.983205e-06, 3.156213e-06, 2.474242e-06, 6.223252e-06, 4.480527e-06,
  4.163593e-05, 7.838171e-05, 8.32708e-05, 3.448362e-05, 2.276974e-05, 
    2.064894e-05, 1.938385e-05, 2.022093e-05, 1.713563e-05, 1.185382e-05, 
    6.601274e-06, 5.502423e-06, 4.773931e-06, 6.337002e-06, 4.732728e-06,
  2.505198e-05, 5.069318e-05, 8.986098e-05, 4.966027e-05, 2.519108e-05, 
    2.221852e-05, 2.39861e-05, 2.20965e-05, 1.900032e-05, 1.10904e-05, 
    8.242958e-06, 7.544012e-06, 6.96487e-06, 7.770522e-06, 7.082182e-06,
  5.914596e-06, 2.440429e-05, 5.906589e-05, 0.0001011788, 3.554345e-05, 
    1.895006e-05, 1.935898e-05, 1.731009e-05, 1.40717e-05, 1.157823e-05, 
    1.021826e-05, 1.144119e-05, 8.490088e-06, 7.22808e-06, 2.423478e-05,
  5.472256e-06, 1.142545e-05, 1.577194e-05, 3.645212e-05, 3.783358e-05, 
    1.83893e-05, 1.56102e-05, 9.507597e-06, 1.193684e-05, 1.093712e-05, 
    1.363961e-05, 1.406658e-05, 9.24802e-06, 1.30605e-05, 6.439529e-05,
  7.267441e-07, 3.176979e-06, 3.204923e-06, 1.55552e-05, 1.589809e-05, 
    1.737934e-05, 1.29791e-05, 8.456754e-06, 7.569211e-06, 1.14205e-05, 
    1.500045e-05, 1.245695e-05, 1.134914e-05, 6.113212e-05, 0.0001052139,
  4.127235e-06, 1.067938e-06, 1.986262e-06, 7.370803e-06, 5.296537e-06, 
    6.230654e-06, 4.798368e-06, 3.784477e-06, 5.783674e-06, 9.640186e-06, 
    1.315503e-05, 2.244325e-05, 7.024281e-05, 0.0001266366, 0.0001266837,
  0.0001067089, 4.512455e-05, 1.871702e-05, 6.353068e-06, 2.479609e-06, 
    2.908783e-06, 2.27848e-06, 2.463667e-06, 7.199984e-06, 2.222689e-05, 
    5.776624e-05, 0.0001122827, 0.0001703104, 0.000179574, 0.0001494811,
  0.0002504373, 0.000202849, 0.0001405341, 8.415795e-05, 5.252254e-05, 
    3.206822e-05, 3.120335e-05, 5.661272e-05, 9.558498e-05, 0.0001384428, 
    0.0001887604, 0.00024391, 0.0002298714, 0.0001716229, 0.0001340151,
  9.218389e-06, 1.620413e-05, 1.030328e-05, 6.363569e-06, 9.286007e-06, 
    1.284127e-05, 1.189519e-05, 8.787343e-06, 6.268295e-06, 5.299099e-06, 
    3.340244e-06, 3.844724e-06, 5.502672e-06, 4.539073e-06, 2.775795e-06,
  9.296614e-06, 1.214111e-05, 1.038998e-05, 7.164683e-06, 7.648029e-06, 
    1.105219e-05, 1.195859e-05, 1.093119e-05, 7.887785e-06, 5.367947e-06, 
    3.517114e-06, 4.193584e-06, 5.005042e-06, 6.839592e-06, 2.810381e-06,
  4.284814e-06, 1.235126e-05, 1.152782e-05, 1.190958e-05, 9.332995e-06, 
    9.660203e-06, 1.176246e-05, 1.304567e-05, 1.004068e-05, 6.227414e-06, 
    4.159218e-06, 3.879576e-06, 5.401158e-06, 6.000117e-06, 2.033052e-06,
  7.147989e-06, 4.339028e-05, 1.193935e-05, 1.380857e-05, 1.2842e-05, 
    9.594977e-06, 1.047755e-05, 1.417704e-05, 1.015236e-05, 7.141107e-06, 
    5.156655e-06, 4.731584e-06, 5.453059e-06, 6.033691e-06, 2.166727e-06,
  1.76078e-05, 2.576401e-05, 2.80366e-05, 2.62465e-05, 1.885531e-05, 
    1.467636e-05, 1.030621e-05, 1.245924e-05, 1.175383e-05, 7.9018e-06, 
    5.850221e-06, 5.232267e-06, 5.826384e-06, 5.257565e-06, 1.904642e-06,
  3.215876e-05, 3.227901e-05, 2.301388e-05, 7.346809e-05, 4.786316e-05, 
    1.912123e-05, 9.879171e-06, 1.063343e-05, 1.023956e-05, 7.817539e-06, 
    6.443872e-06, 6.329977e-06, 5.561002e-06, 4.398132e-06, 1.654339e-06,
  2.414662e-05, 4.345897e-05, 4.379075e-05, 6.416268e-05, 0.0001122144, 
    4.41354e-05, 1.854038e-05, 1.45389e-05, 1.09397e-05, 8.542101e-06, 
    8.064674e-06, 7.167179e-06, 5.320922e-06, 2.897217e-06, 1.233732e-06,
  8.655417e-06, 3.202545e-05, 4.992524e-05, 6.713622e-05, 0.0001128129, 
    0.0001074616, 3.025478e-05, 1.692807e-05, 1.077347e-05, 8.324184e-06, 
    7.43002e-06, 7.645755e-06, 4.495021e-06, 2.701798e-06, 9.697808e-07,
  7.566044e-07, 1.25222e-05, 5.548628e-05, 7.892755e-05, 0.0001137538, 
    0.0001171958, 4.065713e-05, 1.634092e-05, 1.120603e-05, 8.23125e-06, 
    7.999238e-06, 5.371653e-06, 3.702484e-06, 2.66304e-06, 4.481053e-07,
  2.516443e-06, 8.12903e-06, 4.080068e-05, 8.344277e-05, 9.473615e-05, 
    9.832819e-05, 5.700121e-05, 1.979337e-05, 1.296146e-05, 9.141038e-06, 
    6.791571e-06, 4.166656e-06, 3.331507e-06, 1.688783e-06, 3.989273e-07,
  1.836121e-05, 3.945226e-06, 3.050466e-06, 1.872599e-06, 1.866241e-06, 
    2.576015e-06, 4.257985e-06, 4.240082e-06, 3.686325e-06, 4.474505e-06, 
    5.606134e-06, 5.391068e-06, 4.694417e-06, 5.133501e-06, 4.708434e-06,
  6.257103e-06, 2.681244e-06, 2.972062e-06, 1.860445e-06, 3.587861e-06, 
    3.855002e-06, 2.631397e-06, 3.078356e-06, 2.293619e-06, 4.735808e-06, 
    5.293938e-06, 4.353399e-06, 3.695837e-06, 3.802691e-06, 4.923788e-06,
  4.261551e-06, 2.153485e-06, 2.323629e-06, 3.274896e-06, 3.424717e-06, 
    2.268883e-06, 3.412216e-06, 3.257623e-06, 1.756753e-06, 2.593333e-06, 
    3.629782e-06, 5.933326e-06, 5.99435e-06, 2.669868e-06, 4.225118e-06,
  3.736711e-06, 2.546654e-06, 2.850585e-06, 1.333507e-06, 2.602253e-06, 
    2.060453e-06, 2.675044e-06, 1.537337e-06, 2.615641e-06, 1.929173e-06, 
    3.942508e-06, 5.218911e-06, 3.084469e-06, 3.10347e-06, 4.076969e-06,
  4.312831e-06, 2.551256e-06, 1.909978e-06, 2.20904e-06, 2.113271e-06, 
    2.669878e-06, 3.669623e-06, 2.003206e-06, 2.756347e-06, 1.552044e-06, 
    2.526192e-06, 4.069631e-06, 4.30236e-06, 3.089629e-06, 3.339795e-06,
  3.70573e-06, 2.690267e-06, 2.702479e-06, 1.715611e-06, 2.061658e-06, 
    2.904751e-06, 2.248984e-06, 3.365658e-06, 3.445076e-06, 2.657827e-06, 
    3.277301e-06, 6.812969e-06, 5.924616e-06, 3.9883e-06, 2.814578e-06,
  3.847797e-06, 2.356504e-06, 1.231508e-06, 1.907638e-06, 1.949069e-06, 
    1.717885e-06, 1.545931e-06, 2.036775e-06, 4.017408e-06, 2.805098e-06, 
    3.03698e-06, 3.883015e-06, 2.769759e-06, 2.136936e-06, 2.212759e-06,
  3.319174e-06, 1.273038e-06, 7.010013e-07, 1.851442e-06, 1.520115e-06, 
    2.197034e-06, 1.124841e-06, 1.319113e-06, 1.736506e-06, 3.316866e-06, 
    3.247844e-06, 2.628322e-06, 2.297497e-06, 1.568461e-06, 1.182653e-06,
  3.447279e-06, 2.8607e-06, 2.241893e-06, 1.305437e-06, 8.414623e-07, 
    1.315267e-06, 8.672354e-07, 6.83008e-07, 8.478967e-07, 2.871307e-06, 
    2.604248e-06, 2.542523e-06, 1.270203e-06, 6.299128e-07, 3.564698e-07,
  3.122664e-06, 3.567738e-06, 1.402996e-06, 1.549596e-06, 5.511866e-07, 
    6.949572e-07, 1.334071e-06, 3.042817e-07, 8.093133e-07, 1.497582e-06, 
    1.630111e-06, 1.578706e-06, 1.304979e-06, 8.85046e-07, 4.844322e-07,
  7.508647e-05, 6.13739e-05, 5.481519e-05, 5.63786e-05, 4.945249e-05, 
    3.903099e-05, 3.862721e-05, 0.0001089756, 0.0001024837, 0.0001067272, 
    8.39866e-05, 4.159372e-05, 6.310517e-05, 0.0001386344, 0.0001569391,
  9.058714e-05, 7.889883e-05, 6.993393e-05, 6.612458e-05, 6.224793e-05, 
    5.441446e-05, 5.141667e-05, 0.0001334965, 0.0001161625, 0.0001687196, 
    9.621694e-05, 8.354672e-05, 0.000125276, 0.0002030132, 0.0002713697,
  9.694175e-05, 8.559135e-05, 7.689679e-05, 6.755691e-05, 6.578425e-05, 
    6.995234e-05, 7.464017e-05, 7.192892e-05, 8.494307e-05, 6.963294e-05, 
    0.0001288978, 0.0001078223, 0.0001656097, 0.0003028206, 0.0004208878,
  8.972405e-05, 8.185884e-05, 7.321395e-05, 6.978685e-05, 7.950236e-05, 
    7.647274e-05, 6.628393e-05, 7.110294e-05, 9.068297e-05, 0.0001769326, 
    0.0002449438, 0.000319329, 0.0003258845, 0.0004385856, 0.0004166109,
  7.850827e-05, 7.939355e-05, 7.45927e-05, 7.606228e-05, 7.534245e-05, 
    7.524175e-05, 6.952668e-05, 7.959136e-05, 9.926802e-05, 0.0001268638, 
    0.0001457249, 0.0002359194, 0.0003102346, 0.000362723, 0.0003637917,
  5.608035e-05, 6.310413e-05, 6.77221e-05, 7.415112e-05, 7.623248e-05, 
    8.000568e-05, 9.067864e-05, 0.0001018266, 0.0001170165, 0.0001396438, 
    0.0002100252, 0.0003771289, 0.0004952879, 0.0004294685, 0.0002759349,
  5.162277e-05, 6.259159e-05, 7.47308e-05, 7.910871e-05, 8.263325e-05, 
    9.009399e-05, 0.000109211, 0.0001288231, 0.0001435438, 0.0002100218, 
    0.0002982407, 0.0003557734, 0.000355802, 0.0002967257, 0.0001580264,
  6.384101e-05, 7.288148e-05, 7.991106e-05, 8.289687e-05, 9.803034e-05, 
    0.0001236279, 0.0001533044, 0.0001853302, 0.0002531235, 0.0003010324, 
    0.000307391, 0.0002468427, 0.0001938887, 0.0001552426, 2.945471e-05,
  8.600976e-05, 9.006811e-05, 0.0001082131, 0.0001270431, 0.0001700344, 
    0.0002076879, 0.0002412558, 0.0003023946, 0.0003247593, 0.0002585542, 
    0.0001587245, 7.466729e-05, 6.986805e-05, 2.721814e-05, 1.123136e-05,
  0.000151443, 0.0001671171, 0.0001905035, 0.0002237395, 0.0002578838, 
    0.0002964634, 0.0003351462, 0.0003026675, 0.00021316, 9.846272e-05, 
    2.336233e-05, 1.505116e-05, 1.818487e-05, 1.274183e-05, 9.473775e-06,
  5.925734e-06, 5.125301e-06, 3.578285e-06, 2.999389e-06, 1.964425e-06, 
    1.468074e-06, 8.503772e-07, 2.173838e-07, 2.633086e-07, 4.22033e-07, 
    9.470154e-08, 1.112739e-06, 1.169605e-06, 6.219634e-07, 2.828288e-08,
  6.08966e-06, 5.517619e-06, 3.569427e-06, 3.759684e-06, 2.948458e-06, 
    1.859989e-06, 6.206587e-07, 8.610692e-08, 2.311256e-07, 5.329047e-07, 
    2.124205e-07, 9.840144e-07, 6.147743e-07, 2.778789e-07, 1.556416e-06,
  7.086543e-06, 6.205443e-06, 5.17367e-06, 3.845388e-06, 3.011102e-06, 
    1.936104e-06, 7.729616e-07, 3.451465e-07, 1.624559e-07, 7.432101e-07, 
    2.174844e-06, 1.240756e-06, 2.715653e-07, 2.367441e-07, 9.880803e-07,
  7.108797e-06, 5.881549e-06, 4.211545e-06, 2.936365e-06, 1.80204e-06, 
    1.123881e-06, 3.578237e-07, 1.573287e-07, 6.190232e-07, 7.730867e-07, 
    4.953014e-08, 1.424732e-06, 2.167128e-07, 5.882594e-08, 1.254902e-05,
  4.263287e-06, 3.093815e-06, 2.282672e-06, 9.291169e-07, 1.232276e-06, 
    6.234798e-07, 3.886055e-07, 8.174555e-07, 5.132974e-07, 6.037749e-07, 
    2.087092e-07, 1.415294e-07, 1.648504e-06, 6.716044e-07, 7.140979e-05,
  2.153564e-06, 2.494545e-06, 2.122952e-06, 1.174981e-06, 8.327067e-07, 
    9.540061e-07, 6.184913e-07, 1.119645e-07, 1.945205e-08, 1.19815e-08, 
    1.136065e-09, 5.247296e-08, 4.194107e-07, 5.181019e-05, 0.0002011419,
  2.350019e-06, 2.129397e-06, 1.517607e-06, 9.413423e-07, 5.161876e-07, 
    2.700825e-07, 1.977142e-07, 1.963362e-09, 1.511303e-08, 2.748688e-10, 
    1.013392e-07, 4.797149e-06, 6.698871e-05, 0.0002368656, 0.0003574727,
  2.573293e-06, 2.131185e-06, 1.567331e-06, 1.255737e-06, 2.671334e-07, 
    1.227151e-07, 1.135563e-08, 4.628885e-10, 1.353089e-08, 4.948804e-06, 
    2.702403e-05, 0.0001106414, 0.0002749718, 0.0004558339, 0.0004289625,
  9.741093e-07, 7.557764e-07, 6.534087e-07, 1.998947e-07, 1.756619e-07, 
    7.47586e-08, 1.710168e-08, 2.474337e-06, 2.193996e-05, 6.434072e-05, 
    0.0001547063, 0.0002970696, 0.0004367087, 0.0005330885, 0.0002951799,
  1.321528e-06, 4.586468e-07, 1.92561e-07, 1.054498e-07, 7.806194e-07, 
    7.452133e-06, 3.419679e-05, 8.520346e-05, 0.0001267348, 0.0001705139, 
    0.0002520676, 0.0003032273, 0.0003475828, 0.0001839665, 0.0001242515,
  1.636402e-05, 6.930608e-06, 9.88491e-07, 1.231417e-06, 8.260754e-07, 
    9.158671e-08, 1.324546e-08, 6.248914e-08, 7.45367e-08, 1.610495e-07, 
    2.406042e-07, 1.249379e-07, 1.650017e-07, 8.411585e-07, 1.57514e-06,
  1.224996e-05, 5.570823e-06, 6.254526e-07, 1.250833e-07, 9.210615e-07, 
    1.194742e-07, 9.487211e-08, 4.612682e-08, 6.907316e-07, 2.783442e-07, 
    3.520666e-07, 6.49959e-09, 4.623177e-09, 1.221422e-06, 1.889526e-06,
  7.29047e-06, 2.819673e-06, 5.153015e-07, 2.060572e-07, 1.018825e-06, 
    2.491109e-08, 1.368562e-08, 7.544491e-08, 5.629494e-07, 2.393301e-07, 
    3.023734e-07, 9.029068e-08, 1.99686e-08, 1.205504e-07, 1.988126e-06,
  6.56778e-06, 2.619532e-06, 5.367112e-07, 2.538535e-07, 1.543365e-07, 
    8.045031e-08, 7.870129e-08, 3.063746e-07, 3.67343e-07, 4.601316e-07, 
    4.530417e-07, 3.966465e-07, 1.639279e-07, 5.705318e-09, 5.038243e-07,
  5.522007e-06, 2.919565e-06, 9.37997e-07, 2.957018e-07, 8.193045e-07, 
    2.379561e-07, 4.504945e-07, 3.887447e-07, 7.40851e-07, 7.254202e-07, 
    9.443931e-07, 4.766614e-07, 2.578282e-07, 1.497408e-08, 2.965575e-07,
  2.59742e-06, 1.726436e-06, 1.226506e-06, 7.095247e-07, 5.74994e-07, 
    4.172904e-07, 3.108844e-07, 1.108589e-07, 3.426811e-07, 9.673299e-07, 
    6.727013e-07, 9.47048e-08, 1.324856e-08, 4.856151e-08, 3.808498e-07,
  5.409843e-07, 9.792062e-07, 8.625889e-07, 6.10414e-07, 5.957088e-07, 
    4.010181e-07, 2.956588e-07, 1.035097e-06, 7.361946e-07, 9.163788e-07, 
    4.982017e-07, 1.739263e-07, 7.768065e-09, 1.855342e-07, 7.740902e-07,
  4.040714e-07, 6.408322e-07, 9.416944e-07, 1.132101e-06, 5.087212e-07, 
    4.29869e-07, 7.358824e-07, 7.219474e-07, 2.108129e-07, 6.099871e-08, 
    2.13885e-07, 1.175051e-07, 1.983431e-08, 2.189984e-06, 3.355549e-06,
  2.301046e-06, 8.444299e-07, 1.258735e-06, 1.589034e-06, 1.25948e-06, 
    8.046758e-07, 6.944913e-08, 3.246423e-07, 6.668012e-08, 1.90477e-07, 
    1.984774e-07, 2.250557e-08, 1.211291e-06, 2.531844e-06, 1.625408e-05,
  2.095085e-06, 1.532655e-06, 1.182968e-06, 1.666559e-06, 9.966254e-07, 
    1.540731e-07, 5.049041e-08, 4.986307e-08, 2.808239e-08, 2.383851e-07, 
    9.743142e-08, 7.794724e-08, 6.389059e-07, 8.69469e-06, 2.432456e-05,
  1.039332e-05, 8.167901e-07, 9.228433e-08, 1.309606e-08, 7.18265e-08, 
    2.145423e-08, 1.598367e-07, 2.88031e-08, 2.788219e-09, 1.699551e-09, 
    8.418046e-10, 2.451245e-09, 1.142453e-08, 1.81376e-07, 4.237343e-07,
  4.90941e-07, 1.772464e-08, 1.318831e-08, 7.367077e-09, 1.634355e-08, 
    1.712755e-08, 1.634122e-07, 2.601049e-08, 2.485617e-09, 4.468983e-09, 
    8.134614e-09, 7.074905e-09, 1.321689e-07, 4.187698e-07, 1.392526e-06,
  2.794745e-08, 1.217788e-08, 8.120264e-09, 7.215402e-09, 8.250405e-09, 
    4.796569e-08, 3.058224e-08, 1.77606e-09, 3.403968e-10, 5.307805e-10, 
    7.609438e-09, 1.209239e-08, 1.462136e-07, 7.531081e-07, 2.072987e-06,
  3.381956e-07, 2.780167e-08, 6.870439e-09, 3.173228e-09, 5.983608e-09, 
    2.391428e-08, 3.768521e-09, 6.208538e-10, 2.774856e-10, 3.470764e-10, 
    3.916183e-08, 4.457135e-08, 2.687706e-07, 7.67583e-07, 4.648296e-07,
  3.452341e-06, 1.015343e-06, 5.128435e-08, 2.912249e-09, 2.251546e-08, 
    2.008159e-09, 1.436737e-09, 7.395646e-10, 2.753288e-10, 1.741245e-09, 
    1.540331e-08, 3.240847e-08, 3.608923e-07, 4.116359e-07, 9.265419e-07,
  1.029979e-05, 2.024688e-06, 1.942822e-07, 5.565598e-09, 3.778113e-09, 
    7.36425e-09, 2.251134e-09, 1.606343e-09, 5.889603e-10, 7.055659e-10, 
    5.873264e-08, 3.023338e-08, 6.044144e-08, 1.344988e-06, 3.063199e-06,
  1.63675e-05, 2.982768e-06, 3.478125e-07, 1.607645e-08, 1.52318e-09, 
    2.458864e-09, 1.90082e-09, 1.035719e-09, 9.668827e-10, 6.83696e-09, 
    1.94603e-08, 6.435932e-08, 3.238211e-07, 2.252567e-06, 4.863222e-06,
  1.688676e-05, 3.670221e-06, 2.009679e-07, 2.298804e-08, 2.92122e-08, 
    1.314911e-09, 5.696535e-10, 1.674746e-09, 3.499266e-08, 4.660521e-08, 
    5.641513e-09, 1.420326e-07, 5.242921e-08, 3.176757e-06, 8.399431e-06,
  2.015401e-05, 5.0925e-06, 5.431099e-07, 2.966213e-08, 6.694593e-08, 
    7.166318e-10, 5.402356e-10, 1.346672e-09, 1.038047e-07, 1.88082e-08, 
    1.87006e-08, 1.900661e-07, 2.683558e-07, 7.744419e-06, 1.294207e-05,
  2.48075e-05, 9.444523e-06, 1.099416e-06, 6.069472e-08, 1.25666e-07, 
    3.015647e-09, 1.478633e-09, 6.503489e-10, 1.288114e-08, 5.578314e-08, 
    2.649662e-08, 2.820316e-09, 3.416394e-07, 1.288445e-05, 3.042339e-05,
  8.684349e-05, 0.0001678022, 0.0002068861, 0.0001807118, 0.0001086574, 
    5.014721e-05, 4.692143e-05, 3.327916e-05, 1.298375e-05, 9.135822e-06, 
    8.706822e-06, 5.607085e-06, 4.017484e-06, 3.685469e-06, 3.148072e-06,
  9.398803e-05, 0.0001630312, 0.0002082549, 0.000176175, 0.0001113876, 
    5.745657e-05, 4.463606e-05, 2.875371e-05, 9.252502e-06, 9.340906e-06, 
    8.172382e-06, 4.700998e-06, 4.003658e-06, 1.986819e-06, 2.041881e-06,
  0.0001107452, 0.0001808027, 0.0002084368, 0.0001628669, 0.00010006, 
    6.477282e-05, 5.108212e-05, 3.877754e-05, 8.555415e-06, 6.042879e-06, 
    4.496003e-06, 3.018473e-06, 5.345257e-06, 3.33041e-06, 2.403267e-06,
  0.0001512471, 0.0001866442, 0.0001789162, 0.0001245952, 7.644565e-05, 
    5.597477e-05, 4.518618e-05, 4.162767e-05, 1.725732e-05, 4.47695e-06, 
    4.570466e-06, 5.153554e-06, 5.465721e-06, 4.35118e-06, 2.668916e-06,
  0.0001616512, 0.0001573127, 0.0001436769, 8.689589e-05, 4.92405e-05, 
    3.769347e-05, 3.012823e-05, 3.193302e-05, 1.71193e-05, 4.587933e-06, 
    2.00777e-06, 3.207731e-06, 2.684375e-06, 2.640026e-06, 2.239606e-06,
  0.000158803, 0.0001347872, 9.606437e-05, 6.52455e-05, 4.210702e-05, 
    3.061382e-05, 2.203211e-05, 2.164371e-05, 1.068203e-05, 4.547572e-06, 
    3.48693e-06, 2.914907e-06, 4.434779e-06, 4.656328e-06, 2.371953e-06,
  0.0001617767, 0.0001022425, 7.483087e-05, 5.571119e-05, 4.25044e-05, 
    1.993168e-05, 8.612612e-06, 8.568406e-06, 8.314546e-06, 3.724601e-06, 
    6.989003e-06, 5.837103e-06, 7.638584e-06, 6.618703e-06, 3.292556e-06,
  0.0001442536, 7.07135e-05, 6.100914e-05, 5.062131e-05, 2.806793e-05, 
    7.78819e-06, 3.218669e-06, 5.866679e-06, 4.572706e-06, 4.819074e-06, 
    7.868388e-06, 7.106301e-06, 9.515943e-06, 1.075866e-05, 5.798721e-06,
  9.548199e-05, 4.481453e-05, 5.196871e-05, 3.37538e-05, 9.618171e-06, 
    2.162307e-06, 1.61216e-06, 2.917132e-06, 2.788104e-06, 1.793571e-06, 
    2.551052e-06, 3.265591e-06, 7.905967e-06, 9.12938e-06, 6.221266e-06,
  4.870227e-05, 3.3723e-05, 3.717537e-05, 1.799472e-05, 2.638495e-06, 
    1.376801e-06, 1.877139e-06, 1.643681e-06, 2.163258e-06, 2.036025e-06, 
    1.26631e-06, 2.362868e-06, 3.334301e-06, 2.878449e-06, 4.964982e-06,
  1.987029e-06, 6.877114e-07, 4.120373e-07, 1.911697e-07, 1.789378e-07, 
    2.32514e-08, 2.019501e-08, 9.734524e-08, 9.336597e-06, 3.248552e-05, 
    3.967853e-05, 1.292201e-05, 5.596773e-06, 2.396787e-06, 5.703755e-06,
  2.520717e-06, 1.790683e-06, 6.080813e-07, 3.364804e-07, 1.307033e-07, 
    6.258676e-08, 2.00963e-08, 9.357849e-07, 1.626755e-05, 3.709449e-05, 
    5.029206e-05, 1.15598e-05, 4.174193e-06, 1.878627e-06, 4.781302e-06,
  3.924012e-06, 3.157861e-06, 6.995527e-07, 3.27552e-07, 1.286971e-07, 
    7.256883e-08, 5.830623e-08, 3.421356e-06, 2.192618e-05, 3.963169e-05, 
    4.951404e-05, 1.597823e-05, 3.486213e-06, 2.140776e-06, 2.884681e-06,
  3.620857e-06, 2.431839e-06, 1.01501e-06, 1.407733e-07, 1.598364e-07, 
    1.837527e-08, 6.231625e-08, 5.861651e-06, 2.090016e-05, 3.062224e-05, 
    4.009593e-05, 1.694652e-05, 3.874295e-06, 5.141589e-06, 2.954375e-06,
  3.348645e-06, 2.935087e-06, 1.376729e-06, 2.717941e-07, 2.472177e-07, 
    2.967925e-08, 8.414107e-07, 9.469062e-06, 2.334103e-05, 2.370221e-05, 
    3.339105e-05, 1.559171e-05, 5.394508e-06, 5.728262e-06, 1.442873e-06,
  3.310153e-06, 2.469894e-06, 1.49921e-06, 2.287584e-07, 1.419645e-07, 
    6.044332e-07, 6.423617e-06, 1.837222e-05, 2.957485e-05, 2.152981e-05, 
    2.36796e-05, 1.078039e-05, 4.81076e-06, 4.296723e-06, 1.117444e-06,
  2.83039e-06, 2.536547e-06, 8.564956e-07, 4.282662e-07, 2.658448e-07, 
    6.593439e-06, 1.402004e-05, 2.339177e-05, 3.217023e-05, 1.974889e-05, 
    1.355362e-05, 1.118765e-05, 6.319583e-06, 6.86366e-06, 1.183386e-06,
  2.810533e-06, 2.338056e-06, 1.56094e-06, 4.745989e-07, 4.675876e-06, 
    1.397083e-05, 1.570281e-05, 2.201791e-05, 2.781626e-05, 1.583653e-05, 
    8.024123e-06, 1.378625e-05, 1.094959e-05, 9.029697e-06, 2.959402e-06,
  3.585853e-06, 2.018784e-06, 1.545172e-06, 4.0916e-06, 1.619285e-05, 
    1.611069e-05, 1.707806e-05, 1.756637e-05, 2.139149e-05, 1.709166e-05, 
    1.453169e-05, 1.616695e-05, 1.306863e-05, 9.831239e-06, 3.54943e-06,
  3.153444e-06, 1.759224e-06, 7.932188e-06, 1.647896e-05, 2.024302e-05, 
    1.640318e-05, 1.695521e-05, 1.78199e-05, 1.682729e-05, 1.855601e-05, 
    1.52459e-05, 1.369148e-05, 8.241834e-06, 5.424416e-06, 1.373726e-06,
  1.636097e-05, 1.056284e-05, 3.496599e-06, 5.009622e-08, 5.417499e-09, 
    9.878223e-09, 6.924692e-09, 1.116006e-08, 4.23209e-07, 4.144183e-06, 
    1.707472e-05, 1.136307e-05, 6.97836e-07, 6.381764e-07, 3.598789e-06,
  1.537584e-05, 1.059857e-05, 5.257568e-06, 1.380509e-07, 5.504848e-09, 
    6.106128e-09, 7.681976e-09, 6.974253e-09, 4.578158e-08, 6.479319e-07, 
    2.550453e-05, 2.210679e-05, 8.932489e-07, 1.950288e-07, 1.908704e-06,
  1.09877e-05, 7.770383e-06, 4.311863e-06, 3.463514e-07, 1.452778e-07, 
    1.691237e-09, 4.40541e-09, 3.024818e-09, 4.783935e-09, 3.73828e-08, 
    3.172614e-05, 3.839976e-05, 2.120275e-06, 1.806938e-07, 1.546528e-06,
  4.587834e-06, 4.808482e-06, 1.437262e-06, 2.430727e-07, 3.810994e-07, 
    5.151318e-08, 1.27142e-09, 1.0633e-09, 2.403814e-09, 2.529081e-08, 
    1.739164e-05, 3.907266e-05, 1.299029e-06, 1.028298e-07, 1.220379e-06,
  4.418612e-06, 3.9436e-06, 1.397867e-06, 7.738641e-07, 5.306911e-07, 
    1.479757e-07, 4.102587e-10, 1.637393e-09, 7.704462e-10, 5.936124e-09, 
    5.571323e-06, 4.89581e-05, 5.679013e-06, 1.094497e-07, 7.11763e-07,
  3.457003e-06, 3.258261e-06, 2.442669e-06, 1.639092e-06, 8.064613e-07, 
    1.519931e-07, 6.821736e-08, 2.528145e-09, 1.480368e-09, 9.955153e-10, 
    4.986255e-07, 4.587476e-05, 1.764171e-05, 1.012516e-06, 1.048378e-06,
  1.201389e-06, 1.88524e-06, 2.672995e-06, 2.025897e-06, 1.643892e-06, 
    7.828637e-08, 1.259905e-07, 1.940718e-09, 3.989198e-09, 1.952459e-09, 
    9.497937e-08, 4.501147e-05, 3.4045e-05, 5.669434e-06, 1.714487e-06,
  6.08828e-07, 1.083218e-06, 1.370033e-06, 3.385634e-06, 1.841535e-06, 
    1.512824e-06, 5.341727e-08, 1.597095e-09, 2.007294e-09, 6.346557e-10, 
    3.614824e-08, 4.228677e-05, 3.641479e-05, 1.18296e-05, 4.658494e-06,
  1.910105e-07, 7.419472e-07, 8.077199e-07, 2.446227e-06, 2.050172e-06, 
    1.238054e-06, 1.059849e-07, 1.301967e-10, 8.456007e-09, 2.283531e-09, 
    3.775618e-08, 3.782272e-05, 4.082541e-05, 1.408523e-05, 4.067316e-06,
  1.112394e-07, 4.791994e-07, 8.929235e-07, 1.958565e-06, 1.979406e-06, 
    1.219832e-06, 3.599512e-09, 7.300598e-09, 1.197178e-09, 8.704826e-10, 
    1.76137e-07, 3.055482e-05, 3.091875e-05, 1.470319e-05, 1.557469e-06,
  0.000158563, 0.0001435957, 0.0001433816, 0.0001343449, 0.000120916, 
    9.23136e-05, 6.225219e-05, 4.737713e-05, 4.50777e-05, 2.992878e-05, 
    1.927151e-05, 6.695215e-06, 1.897289e-06, 2.757606e-06, 2.00634e-06,
  0.0001827551, 0.0001733507, 0.0001794324, 0.0001689134, 0.0001523216, 
    0.0001165646, 8.759912e-05, 4.246425e-05, 4.750645e-05, 2.178329e-05, 
    1.835946e-05, 1.524604e-05, 2.203141e-06, 2.083548e-06, 1.850129e-06,
  0.0002057522, 0.0002150918, 0.0002138877, 0.0002046736, 0.0001788362, 
    0.0001434245, 0.000103408, 6.076683e-05, 4.683909e-05, 4.437476e-05, 
    1.587538e-05, 1.6582e-05, 3.604479e-07, 2.041817e-06, 1.431696e-06,
  0.0002156639, 0.0002411402, 0.0002383577, 0.0002184446, 0.0001920173, 
    0.0001540876, 0.0001169986, 7.214294e-05, 3.880003e-05, 1.957976e-05, 
    1.528913e-05, 1.625296e-05, 6.269354e-06, 2.220721e-06, 1.68737e-06,
  0.0002036692, 0.0002071928, 0.0002270673, 0.0002290744, 0.0002060975, 
    0.0001567154, 0.0001140513, 7.891656e-05, 4.562661e-05, 1.30094e-05, 
    9.682441e-06, 1.999837e-05, 1.317415e-05, 2.761589e-06, 2.005676e-06,
  0.0001754266, 0.0001927579, 0.0002071648, 0.0002176458, 0.0002173293, 
    0.0001641977, 0.0001106525, 8.008311e-05, 4.739456e-05, 2.3252e-05, 
    1.417508e-05, 1.716323e-05, 2.483359e-05, 9.915833e-06, 4.334172e-06,
  0.0001467758, 0.0001640407, 0.0001923791, 0.0002254926, 0.0002127785, 
    0.0001676559, 0.0001104215, 7.922434e-05, 5.244403e-05, 6.609881e-06, 
    2.428697e-06, 8.25074e-06, 2.471579e-05, 2.037278e-05, 5.53056e-06,
  0.0001332342, 0.0001473796, 0.000170243, 0.000211505, 0.0002131114, 
    0.0001706686, 0.0001124333, 7.570413e-05, 3.911006e-05, 2.908601e-06, 
    3.490382e-08, 5.125308e-06, 3.099296e-05, 3.382792e-05, 3.965312e-06,
  0.0001364114, 0.0001375639, 0.0001497634, 0.0001897881, 0.0002009238, 
    0.000157442, 0.0001079646, 7.327808e-05, 2.415391e-05, 5.444698e-07, 
    2.17706e-06, 9.468962e-06, 4.863807e-05, 3.826179e-05, 5.943798e-06,
  0.0001470324, 0.0001382018, 0.0001411017, 0.0001676307, 0.0001844886, 
    0.0001563714, 0.0001156812, 5.597895e-05, 7.708871e-06, 2.844756e-07, 
    3.353024e-07, 2.8076e-05, 6.825201e-05, 2.623416e-05, 2.382922e-06,
  2.098927e-06, 2.109467e-06, 1.638838e-06, 2.200457e-06, 1.1456e-06, 
    7.759102e-07, 4.815002e-07, 3.955059e-07, 6.568868e-07, 5.88656e-06, 
    1.522032e-05, 1.801825e-05, 1.651604e-05, 8.813086e-06, 3.944028e-06,
  2.248543e-06, 2.661149e-06, 1.97185e-06, 2.34152e-06, 2.02507e-06, 
    1.204455e-06, 1.062262e-06, 1.266242e-06, 3.418347e-07, 6.909257e-06, 
    1.438584e-05, 2.252842e-05, 2.309382e-05, 1.424951e-05, 5.078005e-06,
  3.123193e-06, 3.903173e-06, 3.625851e-06, 3.087813e-06, 2.281189e-06, 
    2.667447e-06, 7.724799e-07, 1.492e-06, 7.351442e-07, 6.955129e-06, 
    1.807551e-05, 2.586925e-05, 2.634177e-05, 1.3545e-05, 1.837159e-06,
  4.85165e-06, 3.800526e-06, 3.609166e-06, 3.09142e-06, 3.855923e-06, 
    2.220043e-06, 2.908644e-06, 1.138934e-06, 1.150849e-06, 8.621505e-06, 
    1.651946e-05, 2.145954e-05, 3.089452e-05, 1.54807e-05, 3.202087e-06,
  5.878339e-06, 3.529027e-06, 3.28175e-06, 2.887897e-06, 2.884174e-06, 
    1.995231e-06, 1.712231e-06, 1.949109e-07, 6.127337e-07, 9.185875e-06, 
    7.513323e-06, 2.424308e-05, 3.302192e-05, 2.324455e-05, 3.322733e-06,
  5.969021e-06, 5.257066e-06, 3.817347e-06, 3.348926e-06, 2.275815e-06, 
    1.376893e-06, 1.596997e-06, 4.877701e-07, 1.11126e-06, 7.324327e-06, 
    1.598246e-05, 1.929612e-05, 3.208618e-05, 2.944196e-05, 8.719227e-06,
  5.543277e-06, 5.24237e-06, 3.319269e-06, 3.421035e-06, 3.216808e-06, 
    1.33572e-06, 4.202808e-07, 4.293456e-07, 2.177442e-06, 1.133804e-05, 
    8.602666e-06, 1.950581e-05, 3.228878e-05, 2.884154e-05, 1.962905e-05,
  5.450912e-06, 2.582581e-06, 3.553673e-06, 2.85744e-06, 3.016553e-06, 
    1.052344e-06, 1.047932e-06, 1.317721e-07, 5.087818e-06, 1.228912e-05, 
    7.650887e-06, 1.230614e-05, 1.596239e-05, 3.452669e-05, 1.796008e-05,
  2.419475e-06, 2.639971e-06, 1.95316e-06, 1.640787e-06, 2.534603e-06, 
    2.68292e-06, 6.955922e-07, 1.107133e-06, 1.351439e-05, 1.573263e-05, 
    6.243424e-06, 1.605843e-05, 3.251954e-05, 3.411776e-05, 2.216887e-05,
  3.200576e-06, 1.783308e-06, 2.187508e-06, 3.004593e-06, 2.351883e-06, 
    1.494947e-06, 1.522887e-06, 1.281977e-05, 2.613239e-05, 5.890412e-06, 
    7.597901e-06, 2.515476e-05, 2.268144e-05, 3.953772e-05, 2.564174e-05,
  1.084443e-05, 5.306845e-06, 2.444661e-06, 9.591309e-07, 1.967523e-06, 
    9.606545e-07, 4.748823e-07, 3.678387e-08, 4.133855e-09, 3.464251e-10, 
    6.819455e-09, 2.33012e-07, 3.693429e-06, 6.752331e-06, 9.960985e-06,
  1.475975e-05, 7.948956e-06, 4.591848e-06, 2.257962e-06, 1.859941e-06, 
    1.734327e-06, 4.69186e-07, 7.883636e-08, 4.64487e-08, 1.420108e-08, 
    1.153293e-08, 5.096996e-08, 3.016065e-06, 7.970085e-06, 1.085905e-05,
  2.039211e-05, 1.455714e-05, 8.475653e-06, 3.475569e-06, 2.181056e-06, 
    1.829317e-06, 1.024012e-06, 2.289972e-07, 1.160574e-08, 2.899588e-07, 
    9.878823e-10, 1.530135e-08, 3.362303e-06, 7.875731e-06, 1.120658e-05,
  2.467028e-05, 1.928305e-05, 1.036269e-05, 4.772893e-06, 1.945538e-06, 
    2.024198e-06, 8.862257e-07, 6.79056e-07, 8.783591e-08, 2.825267e-08, 
    6.213586e-08, 1.870506e-07, 4.752112e-06, 9.557307e-06, 1.282279e-05,
  2.385081e-05, 2.199585e-05, 1.257635e-05, 6.247169e-06, 3.062145e-06, 
    2.555253e-06, 1.487281e-06, 1.036983e-06, 1.670679e-08, 1.901076e-08, 
    2.843301e-07, 1.520306e-06, 2.167631e-06, 7.506066e-06, 1.730422e-05,
  2.668481e-05, 2.599492e-05, 1.445408e-05, 6.168678e-06, 2.76065e-06, 
    2.822715e-06, 1.437921e-06, 1.952335e-06, 9.506384e-07, 1.226937e-07, 
    1.103048e-06, 1.162389e-06, 1.997034e-06, 7.748436e-06, 1.391975e-05,
  2.770818e-05, 2.321004e-05, 1.584905e-05, 8.27515e-06, 5.97132e-06, 
    4.578822e-06, 3.5173e-06, 1.820219e-06, 4.888263e-07, 9.480535e-07, 
    2.374371e-06, 1.18836e-06, 1.476003e-06, 5.433079e-06, 1.600884e-05,
  2.055975e-05, 1.968352e-05, 1.473631e-05, 1.24257e-05, 8.203718e-06, 
    6.25378e-06, 5.00942e-06, 1.900856e-06, 1.209826e-06, 1.455792e-06, 
    1.398493e-06, 7.880595e-07, 1.411745e-06, 3.926207e-06, 1.910073e-05,
  1.175382e-05, 1.174736e-05, 1.220046e-05, 1.033889e-05, 1.010829e-05, 
    6.685646e-06, 4.2471e-06, 2.141167e-06, 1.242102e-06, 8.677241e-07, 
    7.601668e-07, 1.391551e-06, 3.968415e-07, 3.260477e-06, 2.140402e-05,
  6.678602e-06, 7.857625e-06, 7.995792e-06, 8.430942e-06, 8.888327e-06, 
    5.586982e-06, 3.343611e-06, 2.319469e-06, 8.744274e-07, 7.078849e-07, 
    1.332261e-06, 2.395582e-06, 2.06152e-06, 1.20915e-06, 1.517273e-05,
  5.210305e-06, 4.855273e-06, 3.974358e-06, 2.148386e-06, 1.553191e-06, 
    1.491029e-06, 2.738579e-06, 1.716641e-06, 1.33351e-06, 2.489917e-06, 
    3.891619e-06, 3.587445e-06, 2.138114e-06, 4.053723e-07, 3.689564e-06,
  4.166208e-06, 4.054481e-06, 6.300227e-06, 3.87771e-06, 2.233982e-06, 
    2.883789e-06, 2.852747e-06, 3.832455e-06, 3.043775e-06, 3.355047e-06, 
    4.178971e-06, 4.375498e-06, 3.373753e-06, 1.213545e-06, 9.344263e-07,
  5.586924e-06, 4.329365e-06, 5.964034e-06, 4.968692e-06, 3.847758e-06, 
    2.801121e-06, 3.699505e-06, 4.186364e-06, 2.798924e-06, 3.526839e-06, 
    4.795229e-06, 3.268266e-06, 3.52646e-06, 1.24022e-06, 8.049802e-07,
  6.401763e-06, 2.676785e-06, 3.841656e-06, 5.55469e-06, 4.834602e-06, 
    4.528484e-06, 3.101083e-06, 5.453574e-06, 5.437835e-06, 4.086476e-06, 
    4.786887e-06, 4.182504e-06, 2.878138e-06, 3.782181e-06, 1.145049e-06,
  5.347704e-06, 4.085904e-06, 2.885241e-06, 5.298196e-06, 5.838259e-06, 
    5.31224e-06, 2.335769e-06, 3.813735e-06, 6.001011e-06, 8.73268e-06, 
    5.168458e-06, 3.856182e-06, 2.900376e-06, 4.431109e-06, 1.202479e-06,
  7.47599e-06, 3.645993e-06, 4.943034e-06, 4.658318e-06, 4.887381e-06, 
    4.545584e-06, 3.757936e-06, 2.514156e-06, 5.177075e-06, 2.982183e-06, 
    4.049026e-06, 3.184649e-06, 2.858831e-06, 3.626728e-06, 2.899023e-06,
  7.907459e-06, 4.428761e-06, 5.2797e-06, 5.481633e-06, 6.571915e-06, 
    4.847187e-06, 6.798251e-06, 2.871811e-06, 3.415923e-06, 3.263399e-06, 
    2.807997e-06, 3.544267e-06, 3.374749e-06, 3.755189e-06, 3.725542e-06,
  6.291099e-06, 3.809983e-06, 3.323264e-06, 5.804348e-06, 6.257555e-06, 
    5.737399e-06, 4.353304e-06, 3.29307e-06, 3.154738e-06, 3.12521e-06, 
    4.218317e-06, 2.828291e-06, 4.17126e-06, 5.2517e-06, 4.688764e-06,
  6.903504e-06, 2.773308e-06, 1.525082e-06, 2.588517e-06, 4.191827e-06, 
    4.159586e-06, 3.064854e-06, 2.437998e-06, 1.790283e-06, 3.747974e-06, 
    3.302816e-06, 4.15661e-06, 4.038503e-06, 4.674536e-06, 4.926674e-06,
  7.461963e-06, 2.135314e-06, 1.776541e-06, 1.284621e-06, 2.123874e-06, 
    3.564033e-06, 2.001638e-06, 1.918496e-06, 3.302508e-06, 4.961079e-06, 
    5.621055e-06, 5.990834e-06, 5.214074e-06, 4.870652e-06, 5.294643e-06,
  1.014417e-05, 8.778127e-06, 8.785397e-06, 7.070085e-06, 6.62485e-06, 
    4.153685e-06, 3.942721e-06, 3.776042e-06, 4.233229e-06, 2.399773e-06, 
    2.693583e-06, 2.925962e-06, 4.084113e-06, 5.830293e-06, 4.969505e-06,
  7.480179e-06, 5.652128e-06, 5.499788e-06, 5.367442e-06, 6.341426e-06, 
    3.044903e-06, 3.58177e-06, 5.590711e-06, 5.515023e-06, 3.712752e-06, 
    3.67531e-06, 3.162938e-06, 2.824272e-06, 5.116058e-06, 4.782473e-06,
  7.287636e-06, 7.281144e-06, 5.692591e-06, 2.907474e-06, 2.478236e-06, 
    6.553539e-06, 4.467794e-06, 6.647464e-06, 5.301262e-06, 5.146384e-06, 
    3.859848e-06, 2.983185e-06, 3.892801e-06, 2.082365e-06, 4.800101e-06,
  7.501406e-06, 6.831005e-06, 4.864405e-06, 3.727325e-06, 3.618182e-06, 
    3.643241e-06, 4.225169e-06, 5.103178e-06, 6.312202e-06, 4.902613e-06, 
    3.791906e-06, 3.876782e-06, 2.797184e-06, 2.833716e-06, 3.885743e-06,
  5.037133e-06, 6.318439e-06, 3.560597e-06, 4.235235e-06, 3.859547e-06, 
    2.504198e-06, 3.085041e-06, 1.775194e-06, 3.604074e-06, 6.67559e-06, 
    5.296997e-06, 4.201603e-06, 3.425184e-06, 2.566613e-06, 4.21149e-06,
  2.639381e-06, 6.720232e-06, 3.871167e-06, 4.337214e-06, 3.223706e-06, 
    1.933528e-06, 1.14786e-06, 3.107977e-06, 2.823779e-06, 6.36219e-06, 
    4.542e-06, 3.79486e-06, 2.606691e-06, 2.754463e-06, 1.97324e-06,
  3.442063e-06, 5.979537e-06, 5.267946e-06, 1.973683e-06, 3.998222e-06, 
    2.885406e-06, 2.961532e-06, 3.755853e-06, 2.632666e-06, 5.830129e-06, 
    3.117999e-06, 3.454254e-06, 2.001607e-06, 1.999259e-06, 2.251018e-06,
  3.38429e-06, 7.873332e-06, 5.748721e-06, 5.113297e-06, 3.546109e-06, 
    5.365709e-06, 3.588166e-06, 5.68669e-06, 8.530094e-06, 9.523656e-06, 
    2.149981e-06, 4.228451e-06, 3.702188e-06, 3.91431e-06, 1.688002e-06,
  5.968159e-06, 7.484799e-06, 4.735527e-06, 6.031956e-06, 6.588036e-06, 
    6.420938e-06, 5.8163e-06, 6.123234e-06, 9.3293e-06, 8.468528e-06, 
    6.652326e-06, 7.924396e-06, 1.066551e-05, 1.902879e-06, 1.624252e-06,
  9.804911e-06, 7.898719e-06, 6.665849e-06, 7.718987e-06, 6.717847e-06, 
    7.579093e-06, 8.24833e-06, 8.974992e-06, 1.007469e-05, 8.80582e-06, 
    5.572908e-06, 5.178189e-06, 6.685963e-06, 1.568336e-06, 4.166164e-06,
  8.057013e-05, 8.043124e-05, 6.435793e-05, 4.23045e-05, 2.783952e-05, 
    2.128427e-05, 2.026601e-05, 2.797402e-05, 2.480653e-05, 1.087816e-05, 
    3.249142e-06, 2.317189e-06, 1.563734e-06, 4.227821e-06, 4.350494e-06,
  7.525242e-05, 6.715566e-05, 5.489885e-05, 4.072224e-05, 2.972908e-05, 
    2.49236e-05, 2.596741e-05, 2.751792e-05, 2.061021e-05, 6.242021e-06, 
    2.159352e-06, 1.768505e-06, 3.451633e-06, 4.363767e-06, 4.517174e-06,
  7.135727e-05, 5.233272e-05, 4.213615e-05, 3.045202e-05, 2.71781e-05, 
    2.368222e-05, 2.399771e-05, 2.476341e-05, 1.979838e-05, 4.646202e-06, 
    4.07502e-06, 3.2008e-06, 3.79296e-06, 4.784057e-06, 6.971108e-06,
  6.655348e-05, 4.190958e-05, 3.020826e-05, 2.319248e-05, 1.944512e-05, 
    1.873711e-05, 2.07831e-05, 2.40617e-05, 1.361527e-05, 4.410073e-06, 
    5.250165e-06, 3.84475e-06, 4.5521e-06, 6.923255e-06, 6.70371e-06,
  5.70103e-05, 2.848805e-05, 2.356436e-05, 1.791625e-05, 1.779754e-05, 
    1.86074e-05, 1.963744e-05, 1.821923e-05, 1.001631e-05, 4.620228e-06, 
    4.454286e-06, 3.621228e-06, 4.786665e-06, 5.032556e-06, 7.178556e-06,
  5.122774e-05, 2.477016e-05, 2.195505e-05, 1.821312e-05, 1.771434e-05, 
    1.583569e-05, 1.819967e-05, 1.315712e-05, 1.101617e-05, 3.441801e-06, 
    6.243896e-06, 2.810642e-06, 3.617009e-06, 5.75181e-06, 7.469438e-06,
  4.933929e-05, 2.412846e-05, 2.225476e-05, 1.811103e-05, 1.648971e-05, 
    1.620742e-05, 1.712935e-05, 1.268392e-05, 1.042209e-05, 6.170452e-06, 
    6.027989e-06, 5.191776e-06, 3.075385e-06, 4.226567e-06, 7.327032e-06,
  4.694162e-05, 2.204094e-05, 2.261992e-05, 1.775187e-05, 1.688642e-05, 
    1.709596e-05, 1.460669e-05, 1.340182e-05, 6.581311e-06, 3.371713e-06, 
    5.004021e-06, 3.731875e-06, 2.873338e-06, 3.489193e-06, 5.066387e-06,
  3.884262e-05, 2.252158e-05, 1.990492e-05, 1.82792e-05, 1.543125e-05, 
    1.36671e-05, 1.095393e-05, 8.263461e-06, 8.651364e-06, 6.332164e-06, 
    8.00047e-06, 5.992269e-06, 4.921962e-06, 6.709647e-06, 4.114725e-06,
  2.74803e-05, 1.501289e-05, 1.437233e-05, 1.302392e-05, 1.04238e-05, 
    8.396785e-06, 8.673753e-06, 8.094356e-06, 9.146838e-06, 9.391815e-06, 
    6.634523e-06, 1.031227e-05, 4.458935e-06, 4.340401e-06, 3.21083e-06,
  3.44092e-06, 1.10505e-05, 1.305617e-05, 5.62696e-06, 2.872564e-06, 
    1.252435e-05, 4.862563e-05, 5.522049e-05, 2.232735e-05, 1.017383e-05, 
    3.948344e-06, 3.351865e-06, 7.368492e-06, 9.792489e-06, 1.034552e-05,
  1.987134e-06, 5.248731e-06, 9.225615e-06, 9.933443e-06, 6.967533e-07, 
    6.92116e-06, 3.863983e-05, 4.54501e-05, 1.434172e-05, 1.160188e-05, 
    4.384893e-06, 5.767842e-06, 7.86203e-06, 1.021236e-05, 1.051109e-05,
  8.912347e-07, 9.587972e-07, 8.971793e-06, 9.429882e-06, 3.279576e-06, 
    5.127059e-06, 1.701821e-05, 2.494335e-05, 1.580661e-05, 1.172486e-05, 
    6.561641e-06, 7.706405e-06, 8.833563e-06, 6.168204e-06, 1.04017e-05,
  9.732518e-07, 1.605436e-06, 7.873427e-06, 8.619547e-06, 6.478675e-06, 
    5.159362e-06, 4.350506e-06, 1.166345e-05, 1.559145e-05, 2.145223e-05, 
    9.460437e-06, 7.653672e-06, 8.246822e-06, 8.236056e-06, 9.706646e-06,
  5.561624e-07, 1.587148e-06, 2.500133e-06, 9.953601e-06, 3.655017e-06, 
    1.273026e-06, 1.050506e-06, 6.30748e-06, 1.397188e-05, 2.569936e-05, 
    9.986118e-06, 6.929759e-06, 7.847896e-06, 9.753187e-06, 9.646623e-06,
  3.334609e-07, 1.533563e-06, 5.05462e-07, 7.426449e-06, 3.541604e-06, 
    5.445459e-07, 7.16019e-07, 5.18353e-06, 8.325446e-06, 2.134473e-05, 
    1.070693e-05, 8.658709e-06, 5.536709e-06, 8.287265e-06, 8.745938e-06,
  2.055104e-07, 8.7559e-07, 5.82715e-07, 3.186197e-06, 3.452487e-06, 
    8.535959e-07, 2.248474e-06, 4.416891e-06, 1.176969e-05, 2.422349e-05, 
    1.349641e-05, 6.474488e-06, 5.493966e-06, 6.531408e-06, 7.91298e-06,
  2.353054e-07, 2.716484e-07, 5.907406e-07, 1.297812e-06, 2.859479e-06, 
    8.505175e-07, 6.451548e-06, 2.901689e-06, 1.107291e-05, 2.036112e-05, 
    1.663284e-05, 6.529809e-06, 5.471911e-06, 7.451734e-06, 8.493349e-06,
  1.66412e-07, 3.852773e-07, 7.058387e-07, 5.003944e-07, 2.868419e-06, 
    1.182263e-06, 8.310365e-07, 3.824239e-06, 9.555556e-06, 2.015461e-05, 
    1.952805e-05, 9.312437e-06, 7.558302e-06, 6.797934e-06, 8.923565e-06,
  1.030189e-07, 1.424221e-07, 2.221033e-07, 2.267474e-07, 1.725536e-06, 
    1.385352e-06, 5.743886e-07, 2.337887e-06, 1.163625e-05, 1.811691e-05, 
    1.440662e-05, 1.103613e-05, 1.036587e-05, 8.085373e-06, 9.193443e-06,
  3.675483e-06, 1.365781e-06, 5.991023e-07, 3.223416e-06, 1.169931e-05, 
    1.421086e-05, 1.562883e-05, 1.463204e-05, 8.511635e-06, 4.252501e-06, 
    4.847806e-06, 4.414163e-06, 5.607946e-06, 8.070813e-06, 8.076465e-06,
  5.548837e-06, 2.206868e-06, 1.63409e-06, 3.629724e-07, 5.34004e-06, 
    1.647334e-05, 1.777099e-05, 1.273121e-05, 1.055448e-05, 5.924426e-06, 
    5.667644e-06, 5.54695e-06, 5.53881e-06, 7.139867e-06, 8.246513e-06,
  8.449207e-06, 9.444986e-06, 2.866861e-06, 1.017156e-06, 1.252162e-06, 
    1.211179e-05, 1.965507e-05, 6.873442e-06, 6.361949e-06, 1.014982e-05, 
    7.487552e-06, 7.167417e-06, 6.364437e-06, 7.324746e-06, 8.739477e-06,
  8.261723e-06, 9.97623e-06, 1.042592e-05, 4.030941e-06, 1.907961e-06, 
    3.3579e-06, 1.276229e-05, 5.527627e-06, 6.504728e-06, 1.445074e-05, 
    1.07644e-05, 8.980711e-06, 7.90374e-06, 8.270044e-06, 9.339818e-06,
  8.773592e-06, 3.110362e-06, 1.3193e-05, 8.767036e-06, 4.6657e-06, 
    5.72044e-06, 2.987579e-06, 5.284745e-06, 9.393422e-06, 1.219946e-05, 
    1.335521e-05, 1.100771e-05, 9.826785e-06, 9.500103e-06, 1.079929e-05,
  1.51579e-05, 1.117033e-05, 9.589608e-06, 1.630045e-05, 8.148562e-06, 
    5.553723e-06, 4.280528e-06, 2.834538e-06, 6.175459e-06, 8.506096e-06, 
    1.486575e-05, 1.201021e-05, 1.378979e-05, 1.247188e-05, 1.057028e-05,
  1.313784e-05, 8.757022e-06, 6.732667e-06, 2.016041e-05, 1.562333e-05, 
    1.065279e-05, 8.243966e-06, 8.761282e-06, 6.727621e-06, 8.729311e-06, 
    1.394285e-05, 1.475522e-05, 1.521339e-05, 1.369387e-05, 1.391858e-05,
  1.137083e-05, 1.12811e-05, 7.300525e-06, 1.306197e-05, 1.830785e-05, 
    1.281671e-05, 1.113827e-05, 1.30636e-05, 7.057028e-06, 9.909828e-06, 
    1.500508e-05, 1.449721e-05, 1.737591e-05, 1.674532e-05, 1.523124e-05,
  9.768506e-06, 1.358879e-05, 9.201914e-06, 6.871926e-06, 1.428178e-05, 
    1.591532e-05, 8.819029e-06, 1.420821e-05, 8.195321e-06, 5.727714e-06, 
    1.210158e-05, 1.634015e-05, 2.042078e-05, 1.510242e-05, 1.488154e-05,
  3.33321e-06, 1.087114e-05, 6.867444e-06, 3.724593e-06, 4.60843e-06, 
    8.649998e-06, 1.482238e-05, 7.317953e-06, 8.54414e-06, 8.537729e-06, 
    1.041101e-05, 1.434321e-05, 1.821627e-05, 1.705289e-05, 1.421928e-05,
  3.584683e-06, 1.96965e-06, 4.847393e-08, 4.337181e-08, 1.239908e-08, 
    6.383773e-09, 6.970672e-06, 1.068879e-05, 7.467519e-06, 6.73772e-06, 
    8.187678e-06, 7.448667e-06, 5.822746e-06, 7.445522e-06, 7.109463e-06,
  9.899227e-07, 1.664607e-07, 1.850777e-08, 3.347365e-09, 1.536734e-09, 
    4.430395e-10, 7.872255e-07, 5.726756e-06, 8.798656e-06, 1.0561e-05, 
    9.511203e-06, 1.043027e-05, 7.752523e-06, 7.644945e-06, 8.439542e-06,
  2.109287e-06, 6.809377e-07, 1.889944e-08, 1.728056e-09, 1.082259e-10, 
    4.950871e-10, 1.110077e-10, 3.685614e-07, 3.201377e-06, 1.019671e-05, 
    1.298275e-05, 1.181456e-05, 1.142181e-05, 9.543012e-06, 7.534031e-06,
  7.159568e-07, 1.007368e-06, 8.932053e-07, 5.219342e-09, 2.291264e-10, 
    9.576235e-08, 1.02446e-07, 6.862996e-08, 9.217396e-07, 6.616806e-06, 
    1.297364e-05, 1.319394e-05, 1.266892e-05, 1.143973e-05, 8.354951e-06,
  8.602663e-07, 1.034219e-06, 8.364248e-07, 8.647136e-07, 2.894658e-06, 
    9.091528e-07, 5.88126e-08, 1.93299e-07, 2.754162e-07, 2.078394e-06, 
    7.699985e-06, 1.187733e-05, 1.373105e-05, 1.272352e-05, 1.169454e-05,
  3.02149e-06, 1.357444e-06, 1.587313e-06, 4.492907e-06, 5.430285e-06, 
    3.339203e-06, 2.324021e-07, 7.741386e-09, 1.317648e-06, 1.749202e-06, 
    5.003797e-06, 1.054331e-05, 1.221255e-05, 1.192247e-05, 9.645047e-06,
  8.240116e-06, 5.888794e-06, 7.520035e-06, 5.106121e-06, 5.728757e-06, 
    8.604886e-06, 2.557344e-06, 5.341411e-07, 1.573765e-06, 2.965676e-06, 
    4.644678e-06, 7.346096e-06, 8.336081e-06, 9.767273e-06, 1.058e-05,
  9.516158e-06, 1.097582e-05, 1.007594e-05, 1.260507e-05, 1.059563e-05, 
    1.238986e-05, 9.749768e-06, 4.347759e-06, 3.098117e-06, 3.843561e-06, 
    6.74135e-06, 6.418741e-06, 6.722184e-06, 8.839028e-06, 1.135676e-05,
  1.335965e-05, 1.040597e-05, 1.229415e-05, 1.649144e-05, 1.644265e-05, 
    1.435173e-05, 1.634992e-05, 1.02794e-05, 8.382062e-06, 3.727567e-06, 
    6.628669e-06, 6.865881e-06, 6.161572e-06, 9.71093e-06, 1.07482e-05,
  1.302278e-05, 1.295947e-05, 1.764832e-05, 1.295559e-05, 1.714725e-05, 
    1.715009e-05, 1.83953e-05, 1.794039e-05, 4.910507e-06, 4.231114e-06, 
    5.460644e-06, 5.119794e-06, 7.942329e-06, 8.132575e-06, 6.927078e-06,
  6.44622e-05, 2.694563e-05, 2.430681e-06, 1.312625e-06, 4.53967e-07, 
    2.131913e-07, 2.593834e-06, 1.081644e-05, 1.70545e-05, 1.154662e-05, 
    9.662978e-06, 9.988329e-06, 8.273106e-06, 5.919146e-06, 6.463536e-06,
  1.496116e-05, 3.12227e-06, 4.890707e-07, 1.1749e-07, 2.370164e-08, 
    1.442856e-08, 5.850519e-09, 5.5077e-06, 9.957725e-06, 1.007492e-05, 
    9.829984e-06, 9.451041e-06, 9.184319e-06, 5.756962e-06, 6.45539e-06,
  2.01415e-06, 7.416153e-07, 1.387759e-07, 1.510162e-08, 5.36571e-09, 
    1.097127e-08, 9.989746e-08, 4.718087e-06, 6.289373e-06, 6.967698e-06, 
    8.310844e-06, 9.355386e-06, 7.876628e-06, 7.953804e-06, 6.141205e-06,
  2.586219e-07, 8.108669e-08, 2.028072e-08, 8.041886e-09, 4.457341e-09, 
    3.798796e-09, 2.461112e-09, 1.197607e-06, 3.452163e-06, 4.760441e-06, 
    6.35366e-06, 7.602131e-06, 8.599161e-06, 8.747399e-06, 8.520654e-06,
  6.371319e-08, 3.84824e-08, 8.847122e-09, 5.075209e-09, 1.887893e-09, 
    9.625127e-10, 1.430199e-07, 1.446352e-06, 4.064494e-06, 4.845822e-06, 
    6.106157e-06, 6.698847e-06, 8.077502e-06, 5.931182e-06, 7.79794e-06,
  2.42001e-08, 1.851328e-08, 1.256573e-08, 9.445897e-09, 3.973073e-09, 
    5.874013e-07, 1.163124e-07, 1.565596e-06, 3.796834e-06, 4.721986e-06, 
    6.397693e-06, 6.9322e-06, 6.042792e-06, 5.893263e-06, 6.678985e-06,
  4.432839e-08, 3.694314e-08, 1.72237e-08, 6.634977e-09, 1.454316e-08, 
    1.533669e-07, 3.954965e-07, 1.887852e-06, 2.932046e-06, 3.356869e-06, 
    4.32046e-06, 4.431855e-06, 5.538863e-06, 6.512222e-06, 4.703315e-06,
  4.670848e-08, 3.651902e-08, 6.451024e-08, 9.173891e-09, 2.397324e-07, 
    1.269664e-06, 1.002899e-06, 1.475284e-06, 3.043129e-06, 6.024587e-06, 
    7.634197e-06, 6.165293e-06, 9.430062e-06, 4.711583e-06, 4.466173e-06,
  1.034568e-07, 1.769318e-08, 8.232427e-07, 1.726189e-06, 3.913194e-06, 
    7.231666e-06, 5.995795e-06, 3.768191e-06, 4.060199e-06, 4.420341e-06, 
    1.333406e-06, 2.05068e-06, 6.351301e-06, 4.407652e-06, 8.064689e-06,
  8.7671e-08, 1.536639e-06, 3.561435e-06, 3.723196e-06, 7.695823e-06, 
    8.452898e-06, 7.337224e-06, 5.345876e-06, 2.63308e-06, 3.651305e-06, 
    1.253089e-06, 2.220173e-06, 4.907773e-06, 3.406864e-06, 2.98994e-06,
  0.0001795781, 0.000562014, 0.0007118631, 0.0006971788, 0.0004547602, 
    0.0001864753, 2.805083e-05, 4.778638e-06, 9.494791e-06, 5.074725e-06, 
    6.194037e-06, 9.656448e-06, 9.279359e-06, 7.765131e-06, 7.687021e-06,
  0.0005259693, 0.0008189211, 0.0008504486, 0.0005783903, 0.0003094456, 
    3.309758e-05, 6.153928e-08, 5.571079e-07, 7.754027e-06, 7.804596e-06, 
    7.114953e-06, 1.019713e-05, 9.128687e-06, 7.877169e-06, 8.008428e-06,
  0.0008685727, 0.0008395328, 0.000609248, 0.0003530725, 8.799521e-05, 
    1.089026e-07, 6.017719e-07, 5.974496e-08, 7.084506e-06, 9.391305e-06, 
    9.409112e-06, 7.276562e-06, 9.648455e-06, 8.63454e-06, 8.284731e-06,
  0.0008741818, 0.0005052933, 0.0002501765, 5.43341e-05, 3.032363e-07, 
    4.163467e-08, 5.252178e-08, 4.680469e-07, 6.436212e-06, 5.562557e-06, 
    5.590665e-06, 6.62189e-06, 7.319381e-06, 8.235845e-06, 7.838227e-06,
  0.0004103376, 9.724987e-05, 2.885082e-05, 1.972959e-06, 2.440041e-08, 
    8.29542e-09, 1.420187e-08, 9.745875e-07, 2.649591e-06, 1.22608e-06, 
    3.051617e-06, 3.836384e-06, 4.609687e-06, 4.436431e-06, 5.71371e-06,
  3.351901e-05, 1.246571e-05, 4.791273e-07, 1.748402e-08, 3.159638e-09, 
    2.577276e-09, 1.843649e-09, 2.263899e-09, 2.087894e-06, 1.805679e-06, 
    3.320078e-06, 3.340653e-06, 3.180135e-06, 2.763284e-06, 3.772472e-06,
  3.206605e-07, 3.558175e-07, 1.68866e-08, 1.187761e-08, 4.769801e-09, 
    3.021919e-09, 6.296214e-09, 8.457138e-07, 3.949494e-06, 5.656404e-06, 
    6.626854e-06, 3.060959e-06, 3.452962e-06, 3.128245e-06, 2.883751e-06,
  1.280899e-08, 1.416102e-08, 2.841533e-08, 2.603353e-08, 6.677849e-09, 
    1.227355e-08, 5.926842e-07, 2.428267e-06, 4.691664e-06, 8.592136e-06, 
    5.488274e-06, 6.214872e-06, 5.02582e-06, 1.893417e-06, 2.24602e-06,
  2.097141e-09, 3.060549e-09, 1.482269e-09, 1.601261e-09, 3.393113e-09, 
    5.459433e-07, 1.734111e-06, 3.947389e-06, 8.046453e-06, 8.197582e-06, 
    8.547093e-06, 4.54876e-06, 4.350733e-06, 4.874247e-06, 5.200752e-06,
  6.394103e-08, 8.878976e-07, 1.605117e-06, 1.89185e-06, 1.295575e-06, 
    6.068009e-06, 6.988593e-06, 7.569124e-06, 8.684013e-06, 1.199154e-05, 
    9.045911e-06, 6.779064e-06, 8.90621e-06, 1.815368e-05, 1.46344e-05,
  1.794232e-05, 1.489734e-05, 2.094835e-05, 8.042635e-05, 0.0001231728, 
    0.0001410739, 0.0001534053, 0.0001211853, 9.258163e-05, 6.839943e-05, 
    6.986534e-05, 6.745481e-05, 4.57505e-05, 1.534815e-05, 5.900728e-06,
  8.937351e-06, 1.546968e-05, 0.0001018704, 0.0001966922, 0.0002364872, 
    0.0002326562, 0.0001648065, 0.0001310984, 9.982607e-05, 9.004955e-05, 
    9.22441e-05, 9.077069e-05, 5.12205e-05, 1.134712e-05, 3.990111e-06,
  1.738395e-05, 9.406715e-05, 0.0002160492, 0.0002905631, 0.0002924538, 
    0.0002039479, 0.0001402861, 0.0001116092, 9.253571e-05, 9.268003e-05, 
    9.693423e-05, 8.132004e-05, 3.116319e-05, 5.328895e-06, 3.241421e-06,
  0.0001508726, 0.0002595584, 0.0003079911, 0.0003032859, 0.0002182784, 
    0.0001554624, 0.0001166875, 8.388571e-05, 9.09678e-05, 9.626599e-05, 
    9.33171e-05, 4.956379e-05, 1.43592e-05, 5.141517e-06, 3.752378e-06,
  0.0003560195, 0.0003439041, 0.0002841101, 0.0002158223, 0.0001729162, 
    0.0001337549, 8.783014e-05, 6.759986e-05, 8.951826e-05, 8.717627e-05, 
    5.25092e-05, 1.631775e-05, 1.058661e-05, 5.883395e-06, 5.233289e-06,
  0.000404422, 0.0002784658, 0.0002391277, 0.0001936375, 0.0001592049, 
    0.0001156463, 8.811142e-05, 9.217798e-05, 9.545148e-05, 5.597202e-05, 
    1.736914e-05, 7.160155e-06, 6.324091e-06, 5.569906e-06, 4.659546e-06,
  0.0002763857, 0.0002091326, 0.000219087, 0.0001947821, 0.000151524, 
    0.0001295405, 0.000124262, 9.867539e-05, 4.260583e-05, 8.997793e-06, 
    4.523558e-06, 3.972608e-06, 3.487645e-06, 2.957616e-06, 2.411874e-06,
  0.0002042756, 0.0001981229, 0.0001961663, 0.0001559682, 0.0001352323, 
    0.0001154863, 7.419829e-05, 3.252855e-05, 8.271884e-06, 4.203353e-06, 
    3.643633e-06, 4.80276e-06, 3.120058e-06, 3.124183e-06, 3.685941e-06,
  0.0001034346, 9.463191e-05, 8.13962e-05, 6.78568e-05, 5.102408e-05, 
    2.454119e-05, 6.507121e-06, 1.959775e-06, 5.196756e-06, 5.024545e-06, 
    5.72492e-06, 5.865799e-06, 6.365044e-06, 5.972292e-06, 5.454609e-06,
  6.295892e-06, 8.67176e-06, 8.075644e-06, 5.61706e-06, 1.347705e-06, 
    2.587051e-06, 3.965447e-06, 5.1353e-06, 6.24891e-06, 6.196312e-06, 
    8.857137e-06, 1.176599e-05, 9.132639e-06, 7.086728e-06, 7.856789e-06,
  1.659413e-05, 1.787308e-05, 1.580599e-05, 1.302111e-05, 1.238098e-05, 
    1.218748e-05, 1.1839e-05, 1.04265e-05, 6.525876e-06, 4.637755e-06, 
    3.413097e-06, 1.986684e-06, 4.340512e-06, 1.218832e-05, 2.365175e-05,
  2.452485e-05, 2.076625e-05, 1.614635e-05, 1.388771e-05, 1.243622e-05, 
    1.414051e-05, 1.161127e-05, 1.020361e-05, 7.189921e-06, 4.784263e-06, 
    3.180353e-06, 3.479811e-06, 9.966578e-06, 2.650917e-05, 3.352308e-05,
  3.246702e-05, 2.599819e-05, 1.800577e-05, 1.672403e-05, 1.78546e-05, 
    1.463452e-05, 9.896997e-06, 7.797322e-06, 5.463981e-06, 3.948121e-06, 
    3.194908e-06, 6.651429e-06, 2.442935e-05, 4.145946e-05, 4.346832e-05,
  4.232627e-05, 3.507649e-05, 2.041598e-05, 1.735732e-05, 1.47286e-05, 
    1.256538e-05, 8.222451e-06, 7.087058e-06, 5.846892e-06, 3.350639e-06, 
    4.362429e-06, 2.079916e-05, 4.176307e-05, 4.947578e-05, 4.334879e-05,
  3.916982e-05, 3.788871e-05, 2.949713e-05, 1.63548e-05, 1.521589e-05, 
    1.243649e-05, 8.093655e-06, 6.860216e-06, 5.417368e-06, 6.661035e-06, 
    1.875728e-05, 4.369489e-05, 5.702454e-05, 4.994425e-05, 4.620506e-05,
  2.283268e-05, 2.309313e-05, 2.956495e-05, 2.025535e-05, 1.18711e-05, 
    1.08018e-05, 7.088306e-06, 5.800109e-06, 1.197998e-05, 3.10349e-05, 
    5.340897e-05, 6.502118e-05, 6.61868e-05, 5.35845e-05, 5.700557e-05,
  1.04551e-05, 1.609403e-05, 1.662271e-05, 1.339981e-05, 8.337335e-06, 
    7.044335e-06, 9.267797e-06, 3.310258e-05, 6.450248e-05, 8.301133e-05, 
    8.36447e-05, 7.302456e-05, 6.270251e-05, 6.463934e-05, 6.556878e-05,
  7.746746e-06, 7.118014e-06, 9.831337e-06, 1.21859e-05, 2.330102e-05, 
    4.786386e-05, 8.064354e-05, 0.0001090433, 0.0001221807, 0.0001050304, 
    8.416957e-05, 7.40763e-05, 7.139424e-05, 7.11936e-05, 5.89935e-05,
  2.333967e-05, 2.135827e-05, 4.705849e-05, 8.294763e-05, 0.0001205824, 
    0.0001357194, 0.0001260043, 0.0001114581, 9.469821e-05, 8.27025e-05, 
    8.150974e-05, 7.912747e-05, 7.049285e-05, 5.669862e-05, 3.762615e-05,
  0.0001328395, 0.0001104691, 0.000107932, 7.192857e-05, 6.211937e-05, 
    5.368417e-05, 5.252606e-05, 6.702504e-05, 7.211808e-05, 7.467808e-05, 
    8.142131e-05, 6.378282e-05, 5.044304e-05, 3.512993e-05, 2.091843e-05,
  2.171886e-05, 2.034214e-05, 1.367145e-05, 6.674316e-06, 4.199249e-06, 
    4.031547e-06, 3.247168e-06, 2.767546e-06, 2.16429e-06, 2.262583e-06, 
    2.521925e-06, 3.52724e-06, 3.200381e-06, 2.66675e-06, 2.849675e-06,
  1.391189e-05, 1.599543e-05, 1.181643e-05, 8.66916e-06, 9.343056e-06, 
    7.686542e-06, 6.80374e-06, 6.967976e-06, 4.622881e-06, 5.754845e-06, 
    2.337706e-06, 4.958581e-06, 4.554983e-06, 3.436028e-06, 3.184282e-06,
  1.023531e-05, 1.447791e-05, 1.118622e-05, 1.076675e-05, 1.360968e-05, 
    1.69062e-05, 1.150559e-05, 1.183993e-05, 6.22283e-06, 7.779497e-06, 
    6.505799e-06, 5.431592e-06, 4.10273e-06, 3.204595e-06, 3.445107e-06,
  1.284491e-05, 1.309331e-05, 1.175866e-05, 1.456174e-05, 1.687855e-05, 
    1.602044e-05, 1.534779e-05, 1.494839e-05, 1.252328e-05, 1.05502e-05, 
    8.738302e-06, 6.821673e-06, 4.827761e-06, 3.836605e-06, 3.747014e-06,
  1.364802e-05, 1.38905e-05, 1.379213e-05, 1.590793e-05, 1.719014e-05, 
    2.084717e-05, 1.790237e-05, 1.922272e-05, 1.824971e-05, 1.374916e-05, 
    1.110333e-05, 9.483691e-06, 6.66111e-06, 5.14817e-06, 3.395678e-06,
  1.447593e-05, 1.519003e-05, 1.626184e-05, 1.863481e-05, 2.160744e-05, 
    2.821178e-05, 2.667156e-05, 2.610183e-05, 2.240477e-05, 1.871849e-05, 
    1.574525e-05, 1.06645e-05, 7.885081e-06, 5.886041e-06, 3.977718e-06,
  1.513235e-05, 1.252382e-05, 1.531741e-05, 1.892192e-05, 2.329634e-05, 
    3.304116e-05, 3.71503e-05, 4.184855e-05, 3.309483e-05, 2.463313e-05, 
    2.154621e-05, 1.41799e-05, 8.590879e-06, 6.732503e-06, 3.420879e-06,
  8.763716e-06, 9.62226e-06, 8.687703e-06, 1.133609e-05, 1.41631e-05, 
    2.033185e-05, 2.876481e-05, 4.368238e-05, 4.863282e-05, 4.408853e-05, 
    2.937389e-05, 1.791816e-05, 1.038472e-05, 5.247161e-06, 3.069933e-06,
  6.772829e-06, 6.635163e-06, 4.720286e-06, 3.638474e-06, 6.0426e-06, 
    8.432285e-06, 1.121819e-05, 1.949766e-05, 2.524606e-05, 3.852883e-05, 
    3.107862e-05, 1.777652e-05, 1.030805e-05, 5.125754e-06, 4.350879e-06,
  2.845325e-06, 1.825511e-07, 4.138952e-06, 1.668539e-06, 2.341538e-06, 
    5.070018e-06, 9.903384e-06, 1.328572e-05, 1.624568e-05, 2.666557e-05, 
    3.223807e-05, 1.829291e-05, 1.009506e-05, 5.623621e-06, 2.053821e-05,
  1.937711e-06, 3.68536e-06, 5.39453e-06, 8.694966e-06, 1.086692e-05, 
    1.636824e-05, 1.994229e-05, 2.045345e-05, 2.294724e-05, 2.218005e-05, 
    1.57547e-05, 1.548828e-05, 1.78122e-05, 1.52911e-05, 1.601302e-05,
  5.514002e-06, 6.356764e-06, 8.499235e-06, 1.111056e-05, 1.655449e-05, 
    2.237719e-05, 2.306231e-05, 2.459151e-05, 2.398544e-05, 2.115071e-05, 
    1.64457e-05, 1.260407e-05, 1.385358e-05, 1.721771e-05, 1.940046e-05,
  8.150349e-06, 9.401667e-06, 6.989083e-06, 1.449247e-05, 1.733633e-05, 
    1.651148e-05, 2.313059e-05, 2.63457e-05, 2.827967e-05, 2.764108e-05, 
    1.4618e-05, 1.319588e-05, 7.417618e-06, 8.919274e-06, 9.649643e-06,
  6.6059e-06, 9.210594e-06, 1.063038e-05, 1.137236e-05, 1.33902e-05, 
    1.742619e-05, 1.522169e-05, 1.957023e-05, 2.191366e-05, 1.877314e-05, 
    1.811412e-05, 1.194028e-05, 1.3589e-05, 1.099665e-05, 9.227477e-06,
  8.195687e-06, 7.827138e-06, 6.233942e-06, 6.302126e-06, 5.564482e-06, 
    7.212492e-06, 7.723999e-06, 1.167453e-05, 1.142186e-05, 1.217323e-05, 
    1.285259e-05, 1.27111e-05, 9.542571e-06, 8.689532e-06, 8.780009e-06,
  4.724897e-06, 4.446976e-06, 4.92945e-06, 4.251886e-06, 3.161482e-06, 
    4.455585e-06, 3.190023e-06, 8.038146e-06, 9.059137e-06, 8.997936e-06, 
    1.010462e-05, 9.933768e-06, 1.016845e-05, 9.37763e-06, 8.424567e-06,
  2.711527e-06, 2.560013e-06, 1.606078e-06, 1.322623e-06, 3.095366e-06, 
    5.930376e-06, 8.148157e-06, 1.105954e-05, 1.343777e-05, 1.297778e-05, 
    1.443797e-05, 1.197934e-05, 1.10676e-05, 9.685432e-06, 7.575389e-06,
  9.280295e-07, 7.381704e-07, 1.705174e-06, 4.231064e-06, 7.755753e-06, 
    1.033938e-05, 1.193155e-05, 1.572337e-05, 2.305171e-05, 2.43945e-05, 
    2.392354e-05, 1.995521e-05, 1.545468e-05, 1.037773e-05, 6.158398e-06,
  9.655352e-07, 5.723804e-07, 3.977922e-06, 7.229828e-06, 8.512411e-06, 
    1.425915e-05, 1.424058e-05, 2.009681e-05, 3.122839e-05, 4.347668e-05, 
    4.515903e-05, 3.167723e-05, 2.071348e-05, 1.314609e-05, 7.257457e-06,
  3.309897e-07, 1.658304e-06, 6.924083e-06, 1.047379e-05, 1.639736e-05, 
    1.334892e-05, 2.496422e-05, 7.540162e-05, 0.0001374816, 0.0001889047, 
    0.0001465063, 8.447357e-05, 3.842423e-05, 1.831421e-05, 1.078857e-05,
  3.33784e-06, 3.652193e-06, 3.399657e-06, 1.211848e-06, 2.244876e-07, 
    1.152215e-06, 4.655271e-06, 4.305522e-06, 6.326622e-06, 4.609872e-06, 
    7.562252e-06, 1.113908e-05, 1.020522e-05, 1.039466e-05, 1.117748e-05,
  3.773013e-06, 2.649988e-06, 1.221977e-06, 6.450162e-07, 2.709399e-07, 
    2.88067e-06, 3.224794e-06, 4.356909e-06, 4.90866e-06, 6.023155e-06, 
    5.459247e-06, 8.998406e-06, 9.55668e-06, 7.93951e-06, 6.92707e-06,
  6.131786e-07, 3.948036e-07, 2.236178e-07, 2.322617e-06, 1.737454e-06, 
    3.447574e-06, 4.959069e-06, 4.739611e-06, 4.088503e-06, 6.609463e-06, 
    6.440482e-06, 5.722277e-06, 5.255841e-06, 5.288416e-06, 4.037742e-06,
  3.927623e-07, 6.546296e-07, 1.261349e-06, 2.45219e-06, 2.391308e-06, 
    3.09049e-06, 3.229553e-06, 5.473354e-06, 4.572407e-06, 4.264464e-06, 
    3.431397e-06, 4.362129e-06, 4.805398e-06, 3.33771e-06, 2.712367e-06,
  3.488503e-06, 1.66277e-06, 1.591748e-06, 2.159428e-06, 2.396369e-06, 
    4.768894e-06, 5.82813e-06, 6.105033e-06, 6.408197e-06, 3.877885e-06, 
    4.400747e-06, 4.584444e-06, 4.319355e-06, 3.198679e-06, 4.051213e-06,
  6.494857e-08, 2.851815e-06, 3.452361e-06, 4.990385e-06, 5.144843e-06, 
    4.388219e-06, 5.873305e-06, 8.251885e-06, 1.020529e-05, 9.241143e-06, 
    1.004546e-05, 7.426176e-06, 5.63156e-06, 2.155637e-06, 6.630598e-06,
  1.542825e-06, 2.058838e-06, 2.34969e-06, 3.794798e-06, 6.887659e-06, 
    7.694778e-06, 8.324369e-06, 1.373734e-05, 1.849656e-05, 1.505476e-05, 
    1.680379e-05, 1.568679e-05, 1.204222e-05, 8.189866e-06, 6.887492e-06,
  5.921239e-07, 2.209385e-06, 2.375281e-06, 7.266913e-06, 6.826611e-06, 
    8.992023e-06, 9.006911e-06, 1.979466e-05, 2.392075e-05, 1.883096e-05, 
    1.705961e-05, 1.734094e-05, 1.660907e-05, 1.294943e-05, 1.023152e-05,
  3.694364e-06, 4.753937e-06, 4.676238e-06, 6.029503e-06, 5.284467e-06, 
    8.465712e-06, 1.897388e-05, 2.887895e-05, 1.831649e-05, 1.290528e-05, 
    1.690368e-05, 1.594659e-05, 1.639216e-05, 1.305228e-05, 1.243997e-05,
  6.262035e-06, 5.848238e-06, 4.222298e-06, 3.727146e-06, 6.584581e-06, 
    1.282954e-05, 2.767419e-05, 1.676632e-05, 1.118833e-05, 3.959304e-06, 
    5.880432e-06, 1.123728e-05, 1.632455e-05, 1.781543e-05, 1.543036e-05,
  1.012132e-05, 1.110316e-05, 1.267301e-05, 1.212718e-05, 1.418691e-05, 
    1.2729e-05, 1.10392e-05, 8.93117e-06, 7.568871e-06, 4.247222e-06, 
    5.276226e-06, 4.751756e-06, 4.954966e-06, 4.126864e-06, 3.663501e-06,
  1.337887e-05, 1.095009e-05, 1.043583e-05, 1.253181e-05, 1.543176e-05, 
    1.564334e-05, 1.210928e-05, 1.056776e-05, 8.678143e-06, 2.916733e-06, 
    4.828624e-06, 4.775447e-06, 3.838612e-06, 4.987197e-06, 3.25648e-06,
  1.169778e-05, 1.145885e-05, 1.127884e-05, 1.169433e-05, 1.682858e-05, 
    1.686478e-05, 1.421515e-05, 1.003439e-05, 5.034044e-06, 1.991961e-06, 
    3.559555e-06, 2.882495e-06, 3.377815e-06, 4.131669e-06, 3.487835e-06,
  1.517213e-05, 1.846774e-05, 1.210426e-05, 1.713226e-05, 1.514666e-05, 
    1.628016e-05, 1.228493e-05, 8.708488e-06, 3.447937e-06, 1.326412e-06, 
    1.668224e-06, 4.213325e-06, 1.490698e-06, 2.433635e-06, 4.291413e-06,
  2.113083e-05, 2.187281e-05, 1.627e-05, 1.311456e-05, 1.412634e-05, 
    1.332233e-05, 8.722275e-06, 6.622841e-06, 3.402519e-06, 2.977359e-06, 
    5.311025e-06, 2.468611e-06, 3.256539e-06, 2.308077e-06, 1.985252e-06,
  2.523768e-05, 1.807616e-05, 1.524991e-05, 9.916896e-06, 9.055573e-06, 
    1.136653e-05, 4.707291e-06, 2.040532e-06, 2.200279e-06, 2.975132e-06, 
    4.295341e-06, 5.328936e-06, 5.205251e-06, 4.196273e-06, 3.10558e-06,
  2.308133e-05, 1.527885e-05, 1.249382e-05, 8.299294e-06, 4.688492e-06, 
    4.757292e-06, 3.666714e-06, 4.503871e-06, 5.245523e-06, 5.751898e-06, 
    6.380219e-06, 6.216085e-06, 5.536157e-06, 5.113346e-06, 2.883484e-06,
  1.60186e-05, 1.80516e-05, 9.845228e-06, 6.867926e-06, 6.051258e-06, 
    8.787311e-06, 8.177095e-06, 6.41587e-06, 6.68314e-06, 5.086023e-06, 
    3.428879e-06, 3.151416e-06, 1.332148e-06, 5.343338e-07, 1.105361e-06,
  1.587689e-05, 1.051054e-05, 8.442754e-06, 7.484669e-06, 1.029603e-05, 
    8.524119e-06, 7.798923e-06, 4.075392e-06, 2.09151e-06, 8.901545e-07, 
    8.842189e-07, 1.441938e-08, 1.921177e-08, 1.344689e-08, 1.223626e-07,
  9.815163e-06, 7.451926e-06, 6.969982e-06, 6.719266e-06, 1.107305e-05, 
    1.145013e-05, 7.217644e-06, 2.069447e-06, 8.698007e-07, 2.904711e-07, 
    1.663218e-07, 3.594934e-07, 2.075895e-07, 5.347246e-07, 8.684329e-07,
  1.774513e-05, 1.482437e-05, 1.200125e-05, 8.499116e-06, 5.492588e-06, 
    4.17396e-06, 3.881303e-06, 6.253069e-06, 1.036208e-05, 1.29175e-05, 
    1.370683e-05, 9.536491e-06, 1.224949e-05, 4.997839e-06, 3.273446e-06,
  2.461113e-05, 1.673996e-05, 1.22638e-05, 9.564631e-06, 7.427278e-06, 
    5.806825e-06, 3.670571e-06, 1.070975e-05, 1.52411e-05, 1.644956e-05, 
    1.644894e-05, 1.205051e-05, 1.300929e-05, 5.422401e-06, 3.177266e-06,
  3.553283e-05, 2.443551e-05, 1.709484e-05, 1.521292e-05, 1.049132e-05, 
    7.526453e-06, 9.426691e-06, 1.068226e-05, 1.758567e-05, 1.840355e-05, 
    1.48903e-05, 1.356379e-05, 1.001024e-05, 3.672361e-06, 2.664859e-06,
  3.819264e-05, 2.628672e-05, 2.211433e-05, 1.635276e-05, 1.301964e-05, 
    1.001504e-05, 1.014719e-05, 1.46203e-05, 2.041519e-05, 2.273133e-05, 
    1.554909e-05, 1.056339e-05, 1.06765e-05, 5.357904e-06, 2.23494e-06,
  3.761267e-05, 2.931097e-05, 2.155897e-05, 1.546775e-05, 1.28326e-05, 
    1.385573e-05, 1.559795e-05, 1.873786e-05, 2.292397e-05, 2.011399e-05, 
    1.336361e-05, 9.643433e-06, 8.934378e-06, 4.984211e-06, 2.395714e-06,
  3.715276e-05, 2.848951e-05, 2.24307e-05, 1.849529e-05, 1.588276e-05, 
    1.626412e-05, 2.242416e-05, 2.305198e-05, 2.470312e-05, 2.048803e-05, 
    1.564272e-05, 9.489813e-06, 9.078434e-06, 4.314587e-06, 2.874669e-06,
  3.735465e-05, 3.176444e-05, 2.510768e-05, 2.087579e-05, 1.840483e-05, 
    2.18867e-05, 2.73835e-05, 2.942019e-05, 3.032194e-05, 2.224894e-05, 
    1.615301e-05, 1.205689e-05, 8.028904e-06, 4.725905e-06, 3.159643e-06,
  3.743892e-05, 3.336666e-05, 2.442236e-05, 1.942894e-05, 1.794364e-05, 
    2.559946e-05, 3.202752e-05, 3.04543e-05, 3.014133e-05, 1.988794e-05, 
    1.490186e-05, 1.239442e-05, 8.431948e-06, 6.508782e-06, 1.988536e-06,
  4.742584e-05, 3.519708e-05, 2.858745e-05, 2.609994e-05, 2.032307e-05, 
    3.876214e-05, 3.475158e-05, 3.659817e-05, 2.821145e-05, 1.851242e-05, 
    1.439754e-05, 1.220816e-05, 1.193863e-05, 6.242736e-06, 6.986272e-07,
  5.877632e-05, 3.519702e-05, 2.708448e-05, 3.032647e-05, 4.355601e-05, 
    4.920796e-05, 4.014327e-05, 3.760936e-05, 2.404804e-05, 1.890841e-05, 
    1.413337e-05, 1.151555e-05, 7.334496e-06, 3.065728e-06, 6.382124e-07,
  5.747377e-06, 5.322775e-06, 4.688167e-06, 3.599046e-06, 4.299745e-06, 
    4.362692e-06, 4.46541e-06, 5.127848e-06, 2.822695e-06, 7.031869e-07, 
    2.900621e-07, 7.042524e-07, 1.087073e-05, 2.776728e-05, 3.439084e-05,
  8.491867e-06, 6.417733e-06, 4.480005e-06, 4.407987e-06, 3.455826e-06, 
    3.552265e-06, 6.174703e-06, 4.001546e-06, 2.617222e-06, 7.732293e-07, 
    4.787676e-07, 1.718086e-06, 4.76928e-06, 2.659192e-05, 3.715061e-05,
  1.0731e-05, 8.617245e-06, 6.075971e-06, 5.70396e-06, 3.861511e-06, 
    2.463561e-06, 4.159614e-06, 3.774135e-06, 2.247374e-06, 8.066821e-07, 
    4.51103e-08, 1.140423e-08, 6.696546e-06, 2.255075e-05, 3.70769e-05,
  1.329768e-05, 9.24402e-06, 8.891296e-06, 4.608021e-06, 4.337861e-06, 
    2.23263e-06, 3.34385e-06, 3.804173e-06, 2.688822e-06, 1.737659e-06, 
    9.407755e-08, 2.257609e-07, 4.312026e-06, 1.913722e-05, 3.310568e-05,
  1.743397e-05, 1.238423e-05, 9.358057e-06, 5.98072e-06, 4.057249e-06, 
    4.181277e-06, 2.942241e-06, 2.874576e-06, 1.817071e-06, 1.745485e-06, 
    4.850305e-07, 4.174504e-07, 2.026436e-06, 1.636472e-05, 3.153789e-05,
  2.064797e-05, 1.349097e-05, 1.005178e-05, 8.131131e-06, 5.79836e-06, 
    4.428739e-06, 2.538096e-06, 2.862155e-06, 1.532016e-06, 9.183634e-07, 
    1.084326e-06, 3.382683e-07, 1.798033e-06, 1.169987e-05, 2.416716e-05,
  2.196071e-05, 1.456455e-05, 1.243709e-05, 9.099213e-06, 6.695405e-06, 
    4.607872e-06, 2.45212e-06, 2.72635e-06, 3.286239e-06, 1.000134e-06, 
    1.259117e-06, 7.70745e-07, 3.623316e-06, 1.314589e-05, 1.96888e-05,
  2.039942e-05, 1.560834e-05, 1.367607e-05, 8.624335e-06, 6.760335e-06, 
    4.721178e-06, 2.704811e-06, 2.619909e-06, 2.360141e-06, 7.486495e-07, 
    1.047671e-06, 8.061308e-07, 2.594675e-06, 1.22079e-05, 2.549006e-05,
  2.001042e-05, 1.699204e-05, 1.403475e-05, 1.12416e-05, 7.864322e-06, 
    4.601121e-06, 2.843527e-06, 2.688492e-06, 1.735359e-06, 3.872396e-07, 
    7.058875e-07, 7.197661e-07, 5.827238e-06, 1.283456e-05, 2.545831e-05,
  2.226584e-05, 1.710764e-05, 1.358389e-05, 1.030577e-05, 7.206231e-06, 
    5.288496e-06, 2.867701e-06, 2.070656e-06, 1.853797e-06, 4.126572e-07, 
    5.381436e-07, 1.020618e-06, 7.104949e-06, 1.576513e-05, 2.472919e-05,
  4.53938e-06, 3.728837e-06, 4.164236e-06, 3.990238e-06, 9.712199e-06, 
    8.258031e-06, 9.214697e-06, 1.459287e-05, 1.490276e-05, 6.809286e-06, 
    3.367048e-06, 1.369212e-06, 8.996003e-07, 2.201362e-05, 5.561628e-05,
  4.033569e-06, 5.076224e-06, 4.592342e-06, 5.937779e-06, 9.021426e-06, 
    9.231891e-06, 8.664671e-06, 1.472762e-05, 1.472923e-05, 7.587065e-06, 
    4.11595e-06, 1.257615e-06, 9.492114e-07, 2.705839e-05, 7.013037e-05,
  4.871565e-06, 5.319896e-06, 4.651961e-06, 5.113578e-06, 2.969104e-06, 
    7.658419e-06, 8.534307e-06, 1.20299e-05, 1.536828e-05, 1.048209e-05, 
    4.635031e-06, 7.597497e-07, 9.959622e-07, 2.7919e-05, 8.011262e-05,
  6.851656e-06, 5.067935e-06, 7.942341e-06, 3.797469e-06, 4.627538e-06, 
    7.046628e-06, 6.498329e-06, 1.381143e-05, 1.550209e-05, 1.131208e-05, 
    7.38318e-06, 1.562263e-06, 1.37426e-06, 2.759273e-05, 7.740886e-05,
  8.572929e-06, 6.555433e-06, 6.764327e-06, 3.744803e-06, 4.917155e-06, 
    7.258083e-06, 4.702219e-06, 7.92427e-06, 1.016512e-05, 1.288197e-05, 
    1.019226e-05, 1.044574e-06, 9.591229e-07, 1.688654e-05, 6.176667e-05,
  6.338757e-06, 8.289315e-06, 4.563732e-06, 3.587971e-06, 4.685531e-06, 
    7.043182e-06, 3.999774e-06, 4.692641e-06, 8.186418e-06, 1.361714e-05, 
    1.010726e-05, 1.800765e-06, 8.041636e-07, 8.787883e-06, 5.333658e-05,
  7.79625e-06, 7.816731e-06, 6.741127e-06, 4.353119e-06, 3.511153e-06, 
    7.042377e-06, 3.791895e-06, 7.548304e-06, 1.100547e-05, 1.231184e-05, 
    8.15783e-06, 3.443898e-06, 8.247103e-07, 7.493825e-06, 3.662309e-05,
  8.35002e-06, 6.518923e-06, 6.568177e-06, 4.585543e-06, 4.75898e-06, 
    3.645282e-06, 1.549033e-06, 8.17756e-06, 7.489548e-06, 1.021412e-05, 
    9.587882e-06, 1.897079e-06, 1.372041e-07, 3.873089e-06, 2.248697e-05,
  6.688324e-06, 6.59062e-06, 6.254334e-06, 5.002718e-06, 3.604547e-06, 
    4.039368e-06, 2.160892e-06, 8.086586e-06, 8.786293e-06, 8.126637e-06, 
    7.669131e-06, 1.373616e-06, 7.806785e-08, 3.069989e-06, 2.571792e-05,
  7.216112e-06, 7.124889e-06, 5.557104e-06, 4.80218e-06, 4.034076e-06, 
    3.812347e-06, 1.541208e-06, 7.1463e-06, 7.766183e-06, 5.22319e-06, 
    6.31084e-06, 1.808312e-06, 3.612654e-08, 3.537694e-06, 2.518111e-05,
  2.309331e-06, 4.690012e-07, 9.400628e-07, 2.769156e-06, 5.320636e-06, 
    6.87146e-06, 7.950019e-06, 7.86186e-06, 5.336385e-06, 2.444628e-06, 
    1.252119e-07, 8.722361e-07, 2.818989e-05, 8.473574e-05, 7.740861e-05,
  2.378366e-06, 1.492363e-06, 6.878282e-07, 7.781542e-07, 5.873648e-06, 
    8.079047e-06, 9.021132e-06, 1.002304e-05, 5.403849e-06, 2.216066e-06, 
    2.715245e-08, 3.73387e-06, 4.221025e-05, 0.0001676876, 0.0001003827,
  3.02657e-06, 2.468993e-06, 1.073688e-06, 7.032035e-07, 5.225242e-06, 
    8.901425e-06, 8.732212e-06, 8.801548e-06, 5.427391e-06, 2.671383e-06, 
    1.875116e-07, 1.740536e-05, 8.24428e-05, 0.0001743436, 0.0001031548,
  3.862813e-06, 1.914183e-06, 7.076761e-07, 2.103974e-06, 3.066153e-06, 
    6.360206e-06, 6.241158e-06, 7.578947e-06, 6.388071e-06, 3.819822e-06, 
    3.418619e-06, 4.984696e-05, 0.0001293472, 0.0001852875, 0.0001093661,
  3.833238e-06, 2.585502e-06, 1.249977e-06, 1.528026e-06, 1.196042e-06, 
    3.931844e-06, 5.612447e-06, 7.50625e-06, 8.240199e-06, 4.474752e-06, 
    8.312261e-06, 6.877477e-05, 0.0001614978, 0.0001868938, 0.0001297426,
  2.278606e-06, 2.142407e-06, 7.897309e-07, 1.585414e-06, 1.372691e-06, 
    2.02274e-06, 5.846382e-06, 8.081128e-06, 7.818449e-06, 5.589946e-06, 
    1.116693e-05, 5.15018e-05, 0.0001974231, 0.0001935, 0.0001193413,
  6.420581e-06, 3.9878e-06, 3.481574e-06, 2.019744e-06, 3.969883e-06, 
    3.81254e-06, 7.551238e-06, 1.197354e-05, 1.025395e-05, 8.190523e-06, 
    7.527497e-06, 5.550721e-05, 8.890735e-05, 0.0001210992, 0.0001014491,
  6.46123e-06, 5.690291e-06, 3.05457e-06, 2.130636e-06, 3.743684e-06, 
    2.286175e-06, 7.796352e-06, 1.454231e-05, 1.305747e-05, 1.076308e-05, 
    2.881367e-06, 4.095693e-06, 3.35288e-05, 5.419746e-05, 7.147952e-05,
  5.797039e-06, 5.481474e-06, 2.595587e-06, 2.330818e-06, 5.1451e-06, 
    1.187289e-06, 7.42966e-06, 1.310327e-05, 1.060977e-05, 9.70435e-06, 
    2.978719e-06, 4.758901e-06, 1.559118e-05, 3.120039e-05, 5.013608e-05,
  4.759959e-06, 5.46451e-06, 1.745841e-06, 2.861497e-06, 4.278578e-06, 
    5.115032e-06, 3.377306e-06, 6.978615e-06, 9.638187e-06, 1.299675e-05, 
    4.840215e-06, 1.444347e-06, 9.953034e-06, 1.448085e-05, 3.80861e-05,
  8.992105e-07, 1.888613e-06, 3.345629e-06, 6.043463e-06, 6.109482e-06, 
    6.600414e-06, 7.402165e-06, 7.113585e-06, 4.260835e-06, 2.559083e-06, 
    9.641556e-06, 2.57658e-05, 2.862191e-05, 1.880191e-05, 2.146334e-05,
  2.270538e-06, 1.750585e-06, 1.156519e-06, 1.660146e-06, 5.324714e-06, 
    1.01457e-05, 9.370354e-06, 1.394172e-05, 7.483765e-06, 5.212322e-06, 
    2.118549e-05, 3.722261e-05, 3.222008e-05, 4.667113e-05, 3.232842e-05,
  4.218332e-06, 1.948571e-06, 4.304559e-07, 9.153279e-07, 1.006816e-05, 
    1.768378e-05, 1.748703e-05, 1.155887e-05, 1.257516e-05, 1.349646e-05, 
    1.811783e-05, 3.945646e-05, 4.372455e-05, 5.65097e-05, 2.683954e-05,
  6.300473e-06, 2.766815e-06, 6.660882e-07, 2.604422e-06, 1.662316e-05, 
    2.705071e-05, 1.570708e-05, 1.453465e-05, 1.545229e-05, 2.031414e-05, 
    7.028736e-05, 0.0001109807, 6.807872e-05, 4.748888e-05, 2.593065e-05,
  7.252591e-06, 5.801755e-06, 1.960972e-06, 4.440594e-06, 1.80695e-05, 
    2.622419e-05, 1.854249e-05, 1.239575e-05, 4.14584e-05, 0.0001230146, 
    0.0002740485, 0.0002356947, 9.70799e-05, 5.380834e-05, 3.22385e-05,
  6.833737e-06, 5.680955e-06, 4.375441e-06, 4.725197e-06, 1.089732e-05, 
    1.862456e-05, 1.860748e-05, 1.098224e-05, 0.0001451122, 0.000455658, 
    0.0007228269, 0.0004583942, 0.0001495485, 6.737748e-05, 4.642365e-05,
  5.960459e-06, 8.327179e-06, 5.10418e-06, 3.309365e-06, 3.794432e-06, 
    9.89012e-06, 1.464721e-05, 8.480261e-06, 0.0002036754, 0.0006453471, 
    0.0007352644, 0.0003821418, 0.0001604076, 7.110763e-05, 4.091802e-05,
  5.416714e-06, 9.89279e-06, 6.392581e-06, 3.286094e-06, 3.193037e-06, 
    2.466368e-06, 6.209374e-06, 7.435835e-06, 9.966607e-05, 0.0003889757, 
    0.0003974794, 9.687677e-05, 7.896454e-05, 5.212408e-05, 2.884304e-05,
  5.409714e-06, 7.853119e-06, 6.53142e-06, 4.984272e-06, 1.548589e-06, 
    6.090871e-07, 9.480615e-07, 7.209849e-07, 4.18859e-05, 0.0001743139, 
    9.049606e-05, 1.118564e-05, 2.198721e-05, 3.177764e-05, 2.82583e-05,
  2.257261e-06, 5.865574e-06, 6.468405e-06, 7.720962e-06, 3.9921e-06, 
    1.853764e-06, 1.291127e-06, 9.304054e-07, 1.130371e-05, 8.117865e-05, 
    1.993907e-05, 6.782702e-06, 9.122303e-06, 9.327833e-06, 7.523612e-06,
  2.898205e-08, 2.748249e-07, 1.868005e-06, 1.522141e-05, 1.974142e-05, 
    2.315955e-05, 2.555502e-05, 2.071258e-05, 1.111404e-05, 4.748128e-06, 
    2.756186e-06, 5.515373e-06, 1.516097e-05, 6.544772e-05, 7.541451e-05,
  1.390749e-06, 1.346608e-06, 9.015837e-06, 2.5624e-05, 2.873935e-05, 
    2.664348e-05, 2.140908e-05, 2.917215e-05, 1.243827e-05, 6.078959e-06, 
    4.075237e-06, 6.393061e-06, 4.60811e-05, 0.0001020219, 6.564139e-05,
  6.480204e-06, 6.673827e-06, 1.735108e-05, 3.496102e-05, 2.021013e-05, 
    7.22698e-06, 2.023265e-05, 2.247822e-05, 1.683317e-05, 4.329645e-06, 
    2.12247e-06, 1.773672e-05, 8.113283e-05, 8.782426e-05, 4.301074e-05,
  1.290768e-05, 9.580955e-06, 2.193804e-05, 2.612801e-05, 1.281368e-05, 
    7.487443e-06, 1.057944e-05, 2.332302e-05, 2.862177e-05, 4.147912e-06, 
    3.028409e-06, 6.107891e-05, 0.0001088576, 3.612235e-05, 1.273717e-05,
  2.154502e-05, 1.654741e-05, 1.515284e-05, 1.110697e-05, 7.914885e-06, 
    2.815495e-06, 6.569248e-06, 5.695117e-05, 7.275229e-05, 4.963573e-05, 
    5.373199e-05, 9.345332e-05, 7.764723e-05, 1.54314e-05, 1.962378e-06,
  2.486734e-05, 2.658333e-05, 1.4528e-05, 8.692186e-06, 1.545045e-06, 
    5.125584e-07, 1.815365e-06, 5.73304e-05, 0.0002515833, 0.0002273697, 
    0.0002067024, 7.232293e-05, 1.733928e-05, 1.769815e-06, 1.942665e-06,
  2.766495e-05, 2.975979e-05, 1.968887e-05, 7.092665e-06, 9.244474e-07, 
    9.190794e-07, 3.252659e-07, 2.40217e-05, 0.0002877932, 0.0004939358, 
    0.0003078324, 7.551543e-05, 6.683928e-06, 3.525948e-06, 3.566879e-06,
  1.185513e-05, 1.866533e-05, 3.250936e-05, 1.798551e-05, 8.135208e-06, 
    4.263423e-06, 1.484648e-06, 3.480545e-06, 0.0001466731, 0.0004490566, 
    0.0003648237, 6.240146e-05, 8.760428e-06, 1.760921e-06, 1.804947e-06,
  6.690668e-06, 1.756741e-05, 2.311054e-05, 2.89915e-05, 2.015527e-05, 
    1.045774e-05, 6.280484e-06, 3.82263e-06, 5.479641e-05, 0.0002873472, 
    0.0002939951, 4.945927e-05, 9.972183e-06, 2.494245e-06, 1.30789e-06,
  8.613637e-06, 1.217607e-05, 1.729437e-05, 2.372331e-05, 2.291007e-05, 
    1.974678e-05, 1.32253e-05, 6.886619e-06, 2.124158e-05, 0.0001448252, 
    0.0001703557, 4.787126e-05, 1.006409e-05, 3.424798e-06, 3.303645e-06,
  6.084643e-06, 5.946742e-06, 7.803954e-06, 3.681801e-06, 1.272052e-06, 
    1.747094e-06, 2.962138e-06, 8.767632e-06, 2.316083e-05, 2.053863e-05, 
    1.147963e-05, 2.956588e-06, 8.963122e-06, 5.358757e-05, 7.680857e-05,
  4.872226e-06, 5.367326e-06, 6.054344e-06, 3.32395e-06, 2.269442e-06, 
    1.849405e-06, 2.124349e-06, 6.444517e-06, 3.18469e-05, 3.468667e-05, 
    1.441627e-05, 4.816973e-06, 2.79978e-05, 9.033492e-05, 3.45664e-05,
  5.032367e-06, 4.605839e-06, 6.961678e-06, 2.13907e-06, 2.758542e-06, 
    3.402562e-06, 2.976702e-06, 4.199059e-06, 3.057562e-05, 3.881198e-05, 
    1.458251e-05, 7.561844e-06, 3.943252e-05, 7.189193e-05, 1.302025e-05,
  4.079001e-06, 4.806103e-06, 5.033418e-06, 3.40952e-06, 4.143792e-06, 
    1.997222e-06, 3.191781e-06, 5.330907e-06, 1.596447e-05, 2.832295e-05, 
    1.751826e-05, 1.808608e-05, 4.22969e-05, 4.366931e-05, 3.568374e-06,
  2.86549e-06, 5.017884e-06, 4.557263e-06, 6.092391e-06, 4.658222e-06, 
    5.070132e-06, 3.646638e-06, 2.177536e-06, 2.16622e-05, 4.625968e-05, 
    3.043699e-05, 4.66511e-05, 5.736754e-05, 1.316746e-05, 1.316105e-06,
  2.399285e-06, 4.325111e-06, 6.684049e-06, 7.711629e-06, 7.691212e-06, 
    5.645568e-06, 4.400973e-06, 2.063538e-06, 2.730791e-05, 0.0001114858, 
    0.0001452661, 0.0001551257, 9.389252e-05, 2.352459e-05, 1.292361e-06,
  2.851712e-06, 4.089005e-06, 6.008923e-06, 6.920154e-06, 9.552319e-06, 
    7.434355e-06, 6.669455e-06, 3.059431e-06, 1.333781e-05, 0.0001348563, 
    0.0002793682, 0.0003261892, 0.0002173286, 6.122914e-05, 3.076101e-06,
  4.507004e-06, 2.894684e-06, 6.3921e-06, 7.665729e-06, 8.72208e-06, 
    9.927162e-06, 9.386066e-06, 5.771286e-06, 1.77865e-06, 9.939435e-05, 
    0.0003060413, 0.0004185563, 0.0003324123, 0.0001290074, 1.156754e-05,
  5.811088e-06, 5.403645e-06, 6.241721e-06, 6.996765e-06, 7.968927e-06, 
    1.085539e-05, 1.011173e-05, 8.867376e-06, 2.514823e-06, 4.024007e-05, 
    0.0002228521, 0.0003639927, 0.000342594, 0.0001943957, 4.530265e-05,
  6.767975e-06, 5.947278e-06, 7.038793e-06, 9.069856e-06, 7.110694e-06, 
    8.072292e-06, 1.111664e-05, 1.006935e-05, 5.422578e-06, 8.451681e-06, 
    9.354244e-05, 0.0002069199, 0.0002124066, 0.0001506661, 5.97575e-05,
  2.159999e-06, 1.813048e-06, 2.527767e-06, 3.338715e-06, 3.411674e-06, 
    3.724605e-06, 3.884294e-06, 4.343617e-06, 1.012872e-05, 2.155933e-05, 
    3.871537e-05, 3.507524e-05, 9.438267e-06, 3.830504e-06, 1.781368e-05,
  1.827666e-06, 1.522602e-06, 2.459328e-06, 2.948703e-06, 4.000748e-06, 
    4.611164e-06, 4.113384e-06, 3.421442e-06, 4.309901e-06, 1.565754e-05, 
    2.656349e-05, 3.28524e-05, 3.344522e-05, 2.307349e-05, 2.915729e-05,
  4.600143e-06, 2.226317e-06, 2.940573e-06, 3.176625e-06, 3.864853e-06, 
    3.655404e-06, 3.914003e-06, 2.145028e-06, 1.251832e-06, 1.242644e-06, 
    1.886244e-05, 2.865797e-05, 8.541745e-05, 9.176072e-05, 4.075166e-05,
  5.13436e-06, 5.146393e-06, 3.577405e-06, 3.473026e-06, 3.404361e-06, 
    3.724382e-06, 3.106103e-06, 2.497827e-06, 8.185161e-07, 9.584427e-07, 
    3.539222e-06, 2.54567e-05, 9.644798e-05, 0.0001548288, 7.787573e-05,
  4.748411e-06, 6.580472e-06, 2.520339e-06, 4.048629e-06, 4.433926e-06, 
    3.040021e-06, 3.464675e-06, 3.157308e-06, 7.543248e-07, 2.494974e-07, 
    9.185807e-07, 1.151828e-05, 5.653768e-05, 0.0001125165, 6.207197e-05,
  3.339996e-06, 4.673422e-06, 8.195502e-06, 7.279609e-06, 6.912711e-06, 
    4.459574e-06, 3.410935e-06, 3.333845e-06, 1.594522e-06, 7.913411e-07, 
    2.401066e-07, 4.261259e-06, 3.86642e-05, 8.507228e-05, 5.576226e-05,
  8.786625e-06, 3.760691e-06, 4.662211e-06, 2.872046e-06, 5.65704e-06, 
    4.766701e-06, 4.987799e-06, 3.304094e-06, 2.313295e-06, 3.112329e-07, 
    3.545456e-07, 7.526286e-07, 2.85626e-05, 8.5084e-05, 8.839205e-05,
  6.071954e-06, 7.502812e-06, 4.516687e-06, 2.212178e-06, 2.459723e-06, 
    7.712071e-06, 6.412509e-06, 4.407129e-06, 3.313225e-06, 2.549901e-06, 
    4.238912e-07, 4.807531e-08, 1.385815e-05, 7.877914e-05, 0.000121495,
  5.215605e-06, 3.530422e-06, 6.346871e-06, 4.190347e-06, 3.53442e-06, 
    3.883838e-06, 6.269455e-06, 5.583469e-06, 4.173027e-06, 2.724498e-06, 
    2.220142e-06, 2.379612e-07, 1.763615e-06, 4.037311e-05, 0.0001045807,
  4.274226e-06, 3.019079e-06, 4.096457e-06, 7.657036e-06, 4.903463e-06, 
    4.127325e-06, 3.755226e-06, 2.806673e-06, 3.57623e-06, 3.463143e-06, 
    2.694949e-06, 1.431718e-06, 2.45608e-07, 8.560006e-06, 4.614991e-05,
  1.270431e-06, 1.688437e-06, 2.229498e-06, 3.91306e-06, 3.705938e-06, 
    3.404107e-06, 6.333373e-06, 4.485486e-06, 5.425168e-06, 8.955465e-07, 
    1.097787e-05, 4.57387e-05, 9.815287e-05, 0.0001052706, 7.068076e-05,
  3.265849e-06, 2.682428e-06, 2.925907e-06, 4.481922e-06, 5.028119e-06, 
    4.976282e-06, 3.334614e-06, 4.587593e-06, 4.450013e-06, 4.306861e-07, 
    3.1164e-06, 1.232277e-05, 9.506581e-05, 0.000183256, 0.0001545406,
  5.217034e-06, 3.444492e-06, 3.961354e-06, 4.449952e-06, 5.338524e-06, 
    3.584679e-06, 2.333021e-06, 5.563474e-06, 8.476519e-06, 3.685772e-06, 
    2.309823e-06, 1.228528e-06, 3.433464e-05, 0.0001505213, 0.0001875675,
  6.587057e-06, 2.894361e-06, 1.219801e-05, 1.307557e-05, 3.930638e-06, 
    4.600749e-06, 4.733797e-06, 4.741006e-06, 6.410172e-06, 6.195794e-06, 
    2.097286e-06, 2.200914e-06, 3.209744e-06, 4.341469e-05, 8.641211e-05,
  4.55461e-06, 5.98395e-06, 6.532889e-06, 5.175136e-06, 1.195037e-05, 
    1.46437e-05, 7.784468e-06, 3.170662e-06, 3.503976e-06, 1.857787e-06, 
    4.674613e-06, 2.960745e-06, 2.569202e-06, 1.645815e-06, 1.351755e-05,
  3.523903e-06, 4.19915e-06, 3.642049e-06, 2.688507e-06, 3.05219e-06, 
    3.933547e-06, 8.437102e-06, 6.26567e-06, 4.234055e-06, 9.093881e-07, 
    2.54844e-06, 5.17864e-06, 4.778173e-06, 1.909972e-06, 8.636081e-07,
  5.039692e-06, 4.917087e-06, 4.882017e-06, 4.149189e-06, 3.092576e-06, 
    2.708061e-06, 5.57323e-06, 8.591573e-06, 4.110666e-06, 2.378541e-06, 
    1.232691e-06, 1.188666e-06, 5.92615e-06, 5.248696e-06, 2.699257e-06,
  5.88308e-06, 5.34211e-06, 4.742189e-06, 4.15158e-06, 5.423154e-06, 
    3.737333e-06, 6.507506e-06, 5.848175e-06, 8.444915e-06, 5.115594e-06, 
    8.604608e-07, 1.444461e-06, 1.249603e-06, 8.423723e-06, 3.971103e-06,
  7.89269e-06, 6.915833e-06, 4.908091e-06, 4.620495e-06, 6.166014e-06, 
    3.31353e-06, 5.006829e-06, 5.472548e-06, 4.074059e-06, 6.667135e-06, 
    1.849521e-06, 3.665537e-07, 8.044353e-07, 1.07965e-05, 3.445376e-06,
  8.268846e-06, 6.222921e-06, 6.8708e-06, 5.977674e-06, 5.552817e-06, 
    5.791126e-06, 4.045624e-06, 3.585973e-06, 3.448195e-06, 2.582903e-06, 
    3.501649e-06, 2.173983e-06, 1.625039e-06, 9.404589e-06, 1.951062e-06,
  4.4948e-09, 9.747085e-07, 1.254406e-06, 1.617101e-06, 2.395099e-06, 
    3.896404e-06, 6.104313e-06, 6.345455e-06, 2.605739e-06, 6.731689e-07, 
    5.779141e-06, 3.818229e-06, 6.593627e-06, 2.887608e-05, 5.22802e-05,
  1.282602e-06, 1.731404e-06, 1.925268e-06, 2.968146e-06, 3.708443e-06, 
    3.76808e-06, 6.871815e-06, 5.687552e-06, 3.879793e-06, 1.718388e-06, 
    9.104754e-07, 6.547888e-07, 6.627487e-07, 1.977687e-05, 4.294891e-05,
  2.816843e-06, 6.11705e-06, 3.199705e-06, 1.751828e-06, 3.272852e-06, 
    3.211311e-06, 2.68811e-06, 3.349144e-06, 4.138331e-06, 9.568882e-07, 
    1.926607e-06, 2.955722e-06, 3.875875e-06, 6.840059e-06, 1.255978e-05,
  4.211272e-06, 5.219712e-06, 4.844959e-06, 3.275967e-06, 7.157493e-06, 
    6.940452e-06, 3.617827e-06, 7.657946e-06, 3.60377e-06, 2.446004e-06, 
    3.009955e-06, 2.210749e-06, 3.284884e-06, 3.130745e-06, 3.749591e-06,
  5.94018e-06, 4.385009e-06, 2.786216e-06, 2.230146e-06, 3.011581e-06, 
    2.313885e-06, 2.685282e-06, 4.967141e-06, 3.946569e-06, 4.204433e-06, 
    3.011404e-06, 2.893659e-06, 2.721924e-06, 5.484903e-06, 3.917579e-06,
  6.378754e-06, 5.875754e-06, 3.268102e-06, 2.160229e-06, 2.091522e-06, 
    2.173451e-06, 2.484462e-06, 4.851486e-06, 2.525046e-06, 3.813289e-06, 
    3.476731e-06, 3.012466e-06, 2.576832e-06, 4.346258e-06, 5.92446e-06,
  6.944078e-06, 6.603193e-06, 4.772915e-06, 3.911834e-06, 3.889542e-06, 
    5.355289e-06, 3.383536e-06, 4.112471e-06, 2.674495e-06, 1.544908e-06, 
    5.628281e-06, 3.441942e-06, 3.237358e-06, 2.901021e-06, 6.473137e-06,
  8.909604e-06, 8.770099e-06, 9.196832e-06, 8.399481e-06, 6.832064e-06, 
    4.435134e-06, 3.535069e-06, 7.313091e-06, 5.197457e-06, 4.551519e-06, 
    5.925167e-06, 5.887332e-06, 5.547816e-06, 4.4754e-06, 3.481779e-06,
  3.378004e-06, 2.699133e-06, 3.928969e-06, 5.304959e-06, 3.323769e-06, 
    3.891654e-06, 4.511764e-06, 6.693776e-06, 7.005676e-06, 7.155721e-06, 
    8.086642e-06, 8.616567e-06, 7.492999e-06, 7.026595e-06, 5.856909e-06,
  3.146875e-06, 3.463746e-06, 3.840393e-06, 5.375251e-06, 4.714598e-06, 
    4.452754e-06, 5.869136e-06, 5.743551e-06, 5.898436e-06, 6.186492e-06, 
    6.225016e-06, 8.819354e-06, 8.747289e-06, 6.256114e-06, 9.358893e-06,
  5.324378e-06, 2.114914e-08, 1.080395e-07, 2.721925e-07, 8.712416e-07, 
    2.971865e-06, 2.909933e-06, 3.753415e-06, 5.78155e-06, 4.91227e-06, 
    5.204152e-06, 5.51697e-06, 4.029347e-06, 2.118387e-06, 4.392467e-06,
  7.033456e-06, 8.681675e-08, 8.370126e-09, 2.147136e-08, 2.633954e-06, 
    3.379974e-06, 3.601395e-06, 3.864888e-06, 3.564027e-06, 5.382265e-06, 
    6.659644e-06, 5.169407e-06, 4.662141e-06, 3.371852e-06, 1.409912e-06,
  1.046568e-05, 2.286652e-07, 3.964589e-07, 2.426293e-07, 2.90629e-07, 
    2.391084e-06, 4.22077e-06, 2.447937e-06, 3.838702e-06, 6.25809e-06, 
    6.301405e-06, 7.867359e-06, 5.463642e-06, 5.593773e-06, 3.728157e-06,
  1.233142e-05, 1.000921e-06, 8.352799e-08, 3.243006e-06, 1.020271e-06, 
    1.242048e-09, 1.487419e-06, 5.811368e-06, 4.466276e-06, 3.552229e-06, 
    5.385684e-06, 3.123975e-06, 5.469269e-06, 5.342697e-06, 6.225368e-06,
  1.383719e-05, 3.685669e-06, 4.9202e-07, 1.97019e-06, 1.47267e-06, 
    3.865104e-09, 1.727261e-06, 9.813242e-06, 5.502876e-06, 3.659839e-06, 
    3.736135e-06, 3.957589e-06, 6.542042e-06, 7.160479e-06, 6.82459e-06,
  1.945151e-05, 7.001091e-06, 1.32127e-06, 2.612934e-06, 3.540091e-06, 
    2.786567e-06, 3.277153e-06, 5.926823e-06, 5.93843e-06, 4.017174e-06, 
    5.251524e-06, 4.785757e-06, 8.183602e-06, 9.515948e-06, 7.60555e-06,
  3.26799e-05, 1.402441e-05, 2.037141e-06, 4.726738e-06, 7.033833e-06, 
    6.041209e-06, 9.163356e-06, 4.921137e-06, 4.332457e-06, 3.999538e-06, 
    3.497057e-06, 4.905858e-06, 8.904726e-06, 1.02691e-05, 8.613936e-06,
  3.377768e-05, 1.528714e-05, 4.120197e-06, 3.483698e-06, 5.435919e-06, 
    8.673823e-06, 9.867392e-06, 4.938401e-06, 3.288299e-06, 4.787372e-06, 
    2.827672e-06, 5.471482e-06, 8.940085e-06, 9.072269e-06, 8.739399e-06,
  2.62144e-05, 1.691815e-05, 5.821316e-06, 2.260074e-06, 4.117976e-06, 
    3.202906e-06, 2.096375e-06, 2.467365e-06, 1.168222e-06, 1.966643e-06, 
    3.772e-06, 5.347531e-06, 9.653425e-06, 9.519835e-06, 8.080862e-06,
  2.159619e-05, 1.298877e-05, 6.071473e-06, 5.750124e-06, 7.484666e-06, 
    6.165982e-06, 2.068666e-06, 2.380887e-06, 2.621218e-06, 2.520283e-06, 
    3.795268e-06, 5.318302e-06, 9.466298e-06, 1.000928e-05, 8.712565e-06,
  1.405534e-05, 8.200675e-06, 2.121435e-06, 1.034682e-06, 2.552339e-07, 
    4.299167e-07, 2.196468e-06, 4.153057e-06, 3.293773e-06, 4.021251e-06, 
    3.854099e-06, 6.036369e-06, 1.027629e-05, 1.323748e-05, 1.274038e-05,
  1.149176e-05, 9.542145e-06, 4.086251e-06, 2.812358e-06, 7.828862e-07, 
    5.956193e-08, 1.512957e-06, 1.023804e-05, 4.967342e-06, 6.236082e-06, 
    3.408655e-06, 4.980193e-06, 8.196743e-06, 1.365451e-05, 1.287198e-05,
  7.424504e-06, 1.158483e-05, 7.816966e-06, 1.390689e-06, 2.233124e-07, 
    4.90127e-07, 1.321558e-07, 8.847102e-06, 8.817259e-06, 2.687658e-06, 
    3.341271e-06, 5.834548e-06, 7.071149e-06, 1.157689e-05, 1.107465e-05,
  7.544794e-06, 1.090672e-05, 1.22597e-05, 3.833101e-06, 1.891601e-06, 
    2.169803e-07, 1.562669e-07, 3.871674e-06, 8.930569e-06, 1.671432e-06, 
    4.061748e-06, 3.669083e-06, 6.272395e-06, 1.092124e-05, 9.721088e-06,
  6.351281e-06, 1.435417e-05, 1.497652e-05, 5.147667e-06, 2.521636e-06, 
    2.033627e-07, 4.352689e-07, 2.657712e-06, 6.608995e-06, 2.813294e-06, 
    2.827558e-06, 4.55725e-06, 6.525047e-06, 8.125841e-06, 8.619644e-06,
  6.926592e-06, 1.634828e-05, 1.588759e-05, 8.833244e-06, 3.431569e-06, 
    1.08055e-06, 1.191098e-06, 3.3337e-06, 4.091117e-06, 2.747577e-06, 
    3.846743e-06, 5.992895e-06, 5.032237e-06, 7.670556e-06, 8.845344e-06,
  6.935319e-06, 1.320051e-05, 1.347632e-05, 9.787285e-06, 6.705073e-06, 
    2.92112e-06, 1.497433e-06, 3.54649e-06, 4.151641e-06, 1.561381e-06, 
    2.170153e-06, 2.875631e-06, 4.297046e-06, 8.003723e-06, 8.797579e-06,
  1.063246e-05, 1.131233e-05, 1.235095e-05, 1.048062e-05, 6.655611e-06, 
    2.280703e-06, 1.911118e-06, 3.755443e-06, 3.392101e-06, 2.529359e-06, 
    3.136888e-06, 3.840502e-06, 4.061924e-06, 6.938872e-06, 8.981597e-06,
  1.240627e-05, 1.578857e-05, 2.362273e-05, 2.06575e-05, 1.211618e-05, 
    2.13126e-06, 1.656049e-06, 5.40698e-06, 3.168634e-06, 2.568538e-06, 
    3.537581e-06, 7.729375e-06, 5.465306e-06, 6.788431e-06, 9.215812e-06,
  1.860948e-05, 2.927464e-05, 3.611692e-05, 3.030774e-05, 1.732671e-05, 
    6.217111e-06, 3.308325e-06, 4.32266e-06, 3.063674e-06, 3.232733e-06, 
    1.801588e-06, 7.444425e-06, 6.804246e-06, 7.282263e-06, 1.007339e-05,
  9.693578e-06, 9.067573e-06, 2.652682e-06, 2.954883e-06, 3.073856e-06, 
    3.345346e-06, 4.946687e-06, 5.973958e-06, 2.432959e-06, 4.005068e-06, 
    5.867657e-06, 5.941104e-06, 1.006329e-05, 1.519102e-05, 1.470483e-05,
  1.537302e-05, 6.068065e-06, 2.193214e-06, 4.041495e-06, 2.732038e-06, 
    3.858527e-06, 4.443829e-06, 6.044545e-06, 5.048918e-06, 3.800351e-06, 
    3.113309e-06, 4.719081e-06, 7.631604e-06, 1.210117e-05, 1.093203e-05,
  3.128224e-05, 1.666685e-05, 5.847343e-06, 6.030952e-06, 5.043543e-06, 
    2.764905e-06, 3.979653e-06, 4.659826e-06, 3.282859e-06, 2.950136e-06, 
    2.726135e-06, 4.08741e-06, 5.620307e-06, 9.345239e-06, 1.1154e-05,
  4.527762e-05, 3.072808e-05, 1.52196e-05, 9.389494e-06, 8.033879e-06, 
    4.340406e-06, 1.218659e-06, 3.239968e-06, 3.114132e-06, 3.21719e-06, 
    3.867056e-06, 4.753535e-06, 3.521978e-06, 8.026712e-06, 1.116238e-05,
  4.266045e-05, 3.624499e-05, 2.850312e-05, 1.764286e-05, 1.236587e-05, 
    4.619489e-06, 4.55721e-07, 7.812469e-07, 2.150854e-06, 2.969614e-06, 
    2.846305e-06, 7.154955e-06, 3.26599e-06, 7.202256e-06, 9.627945e-06,
  4.628794e-05, 3.586935e-05, 3.278862e-05, 3.575271e-05, 2.25864e-05, 
    7.093525e-06, 1.815545e-06, 8.047411e-07, 2.201858e-06, 6.111248e-06, 
    2.562393e-06, 4.145936e-06, 7.34182e-06, 5.070256e-06, 9.19267e-06,
  5.693081e-05, 4.459491e-05, 4.208118e-05, 4.361092e-05, 3.837957e-05, 
    1.943165e-05, 2.894722e-06, 3.327405e-06, 7.503086e-07, 3.985282e-06, 
    2.131613e-06, 4.542437e-06, 2.53374e-06, 5.009064e-06, 8.251666e-06,
  3.954556e-05, 3.802329e-05, 3.438622e-05, 3.997182e-05, 3.859304e-05, 
    3.355926e-05, 9.669485e-06, 2.747937e-06, 1.238902e-06, 3.369431e-06, 
    2.297706e-06, 3.695731e-06, 4.237586e-06, 5.196886e-06, 6.44296e-06,
  2.249014e-05, 2.212168e-05, 1.76604e-05, 1.913137e-05, 3.818112e-05, 
    3.783546e-05, 1.918568e-05, 4.175402e-06, 9.114542e-07, 1.765637e-06, 
    7.87761e-06, 1.464498e-06, 3.703117e-06, 6.135781e-06, 6.38919e-06,
  1.391604e-05, 1.430796e-05, 7.492795e-06, 5.623627e-06, 1.222843e-05, 
    2.919319e-05, 3.154413e-05, 1.338261e-05, 3.384216e-06, 4.172736e-07, 
    3.457538e-06, 1.400151e-06, 6.082639e-06, 7.589365e-06, 6.031471e-06,
  6.025215e-06, 6.096825e-06, 5.455532e-06, 9.217623e-06, 7.331148e-06, 
    2.209661e-06, 2.103655e-06, 6.972301e-06, 7.191782e-06, 2.475226e-06, 
    2.61698e-06, 2.240576e-06, 7.263514e-06, 1.218052e-05, 1.1578e-05,
  6.258371e-06, 5.789016e-06, 4.401032e-06, 8.000806e-06, 8.442326e-06, 
    3.098679e-06, 2.729564e-06, 5.48972e-06, 5.430966e-06, 7.507796e-06, 
    4.476079e-06, 3.050375e-06, 5.689417e-06, 1.097223e-05, 9.348653e-06,
  7.719769e-06, 5.8187e-06, 5.078185e-06, 3.636607e-06, 7.160866e-06, 
    5.313896e-06, 5.605932e-06, 4.526079e-06, 5.917261e-06, 3.873452e-06, 
    4.217882e-06, 2.925783e-06, 5.515765e-06, 1.055422e-05, 9.823425e-06,
  1.125825e-05, 8.719366e-06, 4.866116e-06, 6.007775e-06, 8.264245e-06, 
    6.688314e-06, 4.650175e-06, 4.362023e-06, 4.258993e-06, 4.545095e-06, 
    3.103605e-06, 3.919271e-06, 5.605072e-06, 9.561942e-06, 9.22972e-06,
  1.345662e-05, 1.308258e-05, 6.427011e-06, 8.716619e-06, 7.3162e-06, 
    6.19066e-06, 4.321083e-06, 5.492171e-06, 3.973925e-06, 3.634786e-06, 
    2.866641e-06, 3.70231e-06, 5.196698e-06, 9.082632e-06, 7.978247e-06,
  1.218697e-05, 1.309631e-05, 1.117063e-05, 8.806774e-06, 6.560143e-06, 
    5.64167e-06, 4.60327e-06, 5.267194e-06, 2.378402e-06, 1.703228e-06, 
    1.761195e-06, 2.999927e-06, 6.298694e-06, 9.631829e-06, 7.254896e-06,
  8.457378e-06, 1.206829e-05, 1.370502e-05, 9.021421e-06, 9.788141e-06, 
    7.147991e-06, 6.701603e-06, 5.417835e-06, 4.812863e-06, 1.701795e-06, 
    1.514775e-06, 3.237597e-06, 5.453846e-06, 9.727969e-06, 8.965731e-06,
  7.774447e-06, 9.9879e-06, 1.529837e-05, 1.646242e-05, 8.227454e-06, 
    8.787251e-06, 5.336112e-06, 6.171863e-06, 5.588466e-06, 1.304263e-06, 
    5.366999e-07, 1.332487e-06, 5.597556e-06, 9.305414e-06, 7.798757e-06,
  1.436921e-05, 1.466266e-05, 1.506507e-05, 1.405108e-05, 2.037923e-05, 
    1.369382e-05, 6.75142e-06, 7.013379e-06, 5.586267e-06, 4.082723e-06, 
    1.023023e-06, 2.448627e-06, 3.928919e-06, 6.428476e-06, 7.228837e-06,
  2.319663e-05, 2.292701e-05, 2.610604e-05, 1.887423e-05, 1.743559e-05, 
    1.918835e-05, 9.479625e-06, 7.69369e-06, 4.982308e-06, 6.013443e-06, 
    1.373578e-07, 1.042308e-06, 3.889742e-06, 5.428249e-06, 6.941064e-06,
  3.748438e-06, 4.346224e-06, 6.054654e-06, 1.268875e-05, 1.256837e-05, 
    4.685105e-06, 3.126376e-08, 6.425446e-09, 5.10349e-07, 3.367204e-06, 
    1.285483e-06, 3.126976e-06, 8.300023e-06, 1.020492e-05, 7.651373e-06,
  2.106178e-06, 2.738529e-06, 4.430745e-06, 4.532447e-06, 9.774211e-06, 
    5.99596e-06, 2.690254e-06, 2.356354e-09, 1.243098e-07, 1.907404e-06, 
    1.873306e-06, 4.210001e-06, 7.287605e-06, 9.18001e-06, 6.540038e-06,
  3.167465e-06, 1.82667e-06, 1.705661e-06, 5.28583e-06, 9.898949e-06, 
    8.420976e-06, 5.231747e-06, 1.982021e-07, 9.679529e-08, 1.551067e-07, 
    1.528422e-06, 3.266205e-06, 6.766672e-06, 8.333218e-06, 5.881814e-06,
  3.17976e-06, 1.432777e-06, 1.37875e-06, 1.905883e-06, 3.914669e-06, 
    6.154013e-06, 4.890836e-06, 3.592756e-06, 1.135453e-06, 1.61628e-06, 
    6.37886e-07, 2.867685e-06, 8.470672e-06, 8.008921e-06, 5.658578e-06,
  5.030086e-06, 3.432232e-06, 2.109852e-06, 2.05239e-06, 3.426559e-06, 
    3.547449e-06, 3.62394e-06, 3.804544e-06, 3.734317e-06, 2.163574e-06, 
    7.801899e-07, 1.733405e-06, 7.885575e-06, 8.331591e-06, 7.20632e-06,
  4.129785e-06, 3.759843e-06, 2.565972e-06, 1.990074e-06, 1.374229e-06, 
    2.635703e-06, 2.634257e-06, 2.478725e-06, 2.986164e-06, 7.140601e-07, 
    3.717733e-07, 1.124311e-06, 5.865206e-06, 6.541437e-06, 5.89103e-06,
  5.74745e-06, 4.822635e-06, 4.374834e-06, 4.383804e-06, 2.135352e-06, 
    1.833919e-06, 2.270879e-06, 3.438504e-06, 2.745341e-06, 2.817441e-06, 
    4.562911e-07, 1.03868e-06, 4.309446e-06, 5.836569e-06, 6.286547e-06,
  4.800925e-06, 5.122646e-06, 6.430691e-06, 6.723313e-06, 4.152473e-06, 
    2.82286e-06, 1.756563e-06, 3.80678e-06, 3.26092e-06, 2.954181e-06, 
    3.50765e-06, 7.721005e-07, 4.111167e-06, 5.540968e-06, 5.733571e-06,
  2.903627e-06, 4.519379e-06, 8.762526e-06, 9.463931e-06, 5.499197e-06, 
    5.528111e-06, 4.332676e-06, 3.00771e-06, 2.630726e-06, 4.188739e-06, 
    4.673137e-06, 1.763332e-06, 3.705971e-06, 4.765132e-06, 5.754413e-06,
  4.426366e-06, 5.111604e-06, 4.687211e-06, 9.297183e-06, 9.412955e-06, 
    7.748502e-06, 6.239567e-06, 3.521282e-06, 3.747399e-06, 5.075563e-06, 
    3.622755e-06, 3.352526e-06, 4.273815e-06, 5.823796e-06, 5.045453e-06,
  6.123182e-05, 2.322352e-05, 2.416947e-06, 1.219893e-06, 1.691924e-06, 
    1.539652e-06, 4.485383e-06, 4.120599e-06, 5.611134e-06, 1.926549e-06, 
    3.764362e-06, 5.920569e-06, 5.901162e-06, 4.910476e-06, 8.187985e-06,
  7.879793e-05, 3.28295e-05, 4.859958e-06, 1.837612e-06, 2.444783e-06, 
    1.7679e-06, 3.752045e-06, 4.399265e-06, 4.011063e-06, 1.672717e-06, 
    5.210195e-06, 7.184851e-06, 6.866037e-06, 6.536343e-06, 5.094147e-06,
  9.499583e-05, 5.392396e-05, 7.094488e-06, 3.351227e-06, 3.401716e-06, 
    2.106023e-06, 3.311589e-06, 4.557957e-06, 2.959565e-06, 3.639849e-06, 
    5.759148e-06, 8.351903e-06, 7.742444e-06, 5.971323e-06, 5.088605e-06,
  0.0001094639, 7.127097e-05, 1.28083e-05, 4.680325e-06, 4.939452e-06, 
    5.673749e-06, 2.817274e-06, 3.097068e-06, 2.311053e-06, 2.610445e-06, 
    4.557149e-06, 5.124869e-06, 8.213848e-06, 6.364302e-06, 6.882506e-06,
  0.0001160153, 8.000957e-05, 1.854545e-05, 5.151575e-06, 3.302889e-06, 
    1.010515e-05, 6.587994e-06, 5.199088e-06, 3.53097e-06, 1.693482e-06, 
    1.993441e-06, 3.793094e-06, 6.631175e-06, 7.420559e-06, 6.55279e-06,
  0.0001217364, 8.946606e-05, 2.581474e-05, 7.555161e-06, 6.725705e-06, 
    9.101014e-06, 7.806175e-06, 5.477154e-06, 7.455358e-06, 2.857072e-06, 
    2.153772e-06, 3.8905e-07, 2.948778e-06, 5.72865e-06, 5.711167e-06,
  0.0001282921, 9.659631e-05, 3.269024e-05, 6.294108e-06, 5.063938e-06, 
    3.767129e-06, 5.728619e-06, 7.168478e-06, 6.256941e-06, 2.826983e-06, 
    1.994418e-06, 6.911577e-07, 2.029738e-06, 3.655636e-06, 5.466381e-06,
  0.0001305203, 0.0001002163, 3.438128e-05, 6.972209e-06, 3.763516e-06, 
    2.643211e-06, 2.810912e-06, 4.335078e-06, 2.974544e-06, 1.566217e-06, 
    1.627296e-06, 6.65136e-07, 4.290443e-07, 2.603982e-06, 4.137627e-06,
  0.0001308188, 9.880464e-05, 3.467075e-05, 8.816474e-06, 3.049596e-06, 
    2.534474e-06, 2.216092e-06, 2.145544e-06, 3.311447e-06, 1.372705e-06, 
    3.547284e-07, 7.448684e-07, 2.537407e-06, 1.825168e-06, 2.656917e-06,
  0.0001295659, 9.043401e-05, 3.755619e-05, 6.060125e-06, 2.49357e-06, 
    3.472648e-06, 1.204224e-06, 1.833059e-06, 1.245511e-06, 5.429438e-07, 
    3.745113e-07, 4.276338e-07, 1.640191e-07, 1.287844e-06, 2.379054e-06,
  1.2302e-05, 3.385477e-05, 3.640355e-05, 1.651366e-05, 2.422846e-06, 
    8.062564e-08, 1.56058e-06, 1.371559e-06, 1.330542e-06, 2.282337e-06, 
    2.985526e-06, 3.829615e-06, 4.308491e-06, 4.721873e-06, 5.691527e-06,
  9.132214e-06, 2.729891e-05, 4.07089e-05, 2.501496e-05, 4.191234e-06, 
    2.936359e-07, 4.015745e-07, 2.319141e-06, 1.797464e-06, 3.202922e-06, 
    3.6764e-06, 4.377293e-06, 4.090134e-06, 5.075575e-06, 5.083829e-06,
  1.224392e-05, 3.675188e-05, 5.718199e-05, 3.722352e-05, 9.054174e-06, 
    2.68337e-07, 2.857571e-07, 4.475867e-06, 1.816717e-06, 2.193195e-06, 
    5.023044e-06, 4.496638e-06, 4.365252e-06, 4.198194e-06, 3.704283e-06,
  2.072635e-05, 4.86855e-05, 7.752865e-05, 6.359886e-05, 1.585434e-05, 
    5.113697e-07, 1.145748e-07, 1.733384e-06, 2.747661e-06, 2.043933e-06, 
    5.912973e-06, 7.393673e-06, 5.223506e-06, 4.540542e-06, 2.342344e-06,
  2.294708e-05, 4.698931e-05, 9.673255e-05, 0.0001015774, 3.862898e-05, 
    1.430236e-06, 2.04074e-07, 1.35282e-06, 3.222607e-06, 2.353125e-06, 
    6.079307e-06, 1.133116e-05, 7.604918e-06, 5.282041e-06, 2.698384e-06,
  2.887999e-05, 5.475446e-05, 0.0001095099, 0.0001378069, 7.7352e-05, 
    4.179678e-06, 4.227088e-08, 2.184603e-06, 2.234191e-06, 2.707289e-06, 
    8.230759e-06, 1.543697e-05, 8.794391e-06, 4.430228e-06, 2.947196e-06,
  3.583396e-05, 5.685541e-05, 0.0001192167, 0.0001600432, 0.0001074216, 
    1.399573e-05, 2.315161e-07, 2.09065e-06, 1.992856e-06, 2.638569e-06, 
    8.665777e-06, 1.182369e-05, 8.792535e-06, 3.72689e-06, 2.919991e-06,
  3.641495e-05, 5.939452e-05, 0.0001189608, 0.0001685728, 0.0001339682, 
    3.419388e-05, 1.157904e-06, 1.176745e-06, 1.371216e-06, 2.756977e-06, 
    8.210417e-06, 8.429194e-06, 6.169195e-06, 9.057977e-07, 2.254089e-06,
  3.905238e-05, 6.283822e-05, 0.0001117617, 0.0001703493, 0.0001494652, 
    5.711802e-05, 2.120578e-06, 2.007637e-06, 8.622065e-07, 1.872242e-06, 
    7.159042e-06, 5.286477e-06, 3.309327e-06, 9.722789e-07, 1.724937e-06,
  3.505058e-05, 6.270751e-05, 0.0001112977, 0.0001697749, 0.0001584288, 
    7.517102e-05, 2.605629e-06, 1.728634e-06, 1.289552e-06, 2.404817e-06, 
    6.824384e-06, 6.131671e-06, 2.971115e-06, 3.76995e-07, 1.561221e-06,
  1.398255e-05, 1.411464e-05, 1.112919e-05, 8.197265e-06, 5.416543e-06, 
    7.0181e-07, 8.360043e-07, 6.991283e-07, 5.336283e-07, 1.214604e-06, 
    3.18165e-06, 1.588642e-06, 1.492174e-06, 2.00646e-06, 4.180289e-06,
  1.252693e-05, 1.24762e-05, 1.061016e-05, 9.645686e-06, 9.664272e-06, 
    6.492754e-06, 5.088335e-07, 4.075758e-07, 8.247309e-07, 1.017568e-06, 
    2.203088e-06, 2.488588e-06, 1.279495e-06, 1.883802e-06, 2.961234e-06,
  8.202063e-06, 1.089092e-05, 1.07857e-05, 9.060094e-06, 1.098306e-05, 
    6.132644e-06, 4.435694e-07, 6.523424e-07, 5.917549e-07, 5.788534e-07, 
    2.31019e-06, 2.389956e-06, 1.109421e-06, 1.429701e-06, 1.945682e-06,
  8.485505e-06, 9.915387e-06, 1.155838e-05, 7.5843e-06, 9.315991e-06, 
    8.609399e-06, 1.905417e-06, 1.039104e-06, 5.642364e-07, 8.391286e-07, 
    1.936752e-06, 2.645055e-06, 1.689412e-06, 1.473809e-06, 2.476678e-06,
  7.816466e-06, 9.243228e-06, 1.059902e-05, 6.881056e-06, 6.830356e-06, 
    1.169649e-05, 4.38712e-06, 8.620549e-07, 1.086874e-06, 7.641195e-07, 
    1.155735e-06, 2.529686e-06, 2.08127e-06, 1.827122e-06, 2.702134e-06,
  6.383538e-06, 9.627529e-06, 7.36232e-06, 8.742527e-06, 5.702214e-06, 
    8.69174e-06, 7.651427e-06, 1.356424e-06, 8.667336e-07, 5.246469e-07, 
    1.6507e-06, 2.807574e-06, 2.632777e-06, 1.53558e-06, 2.742933e-06,
  5.042461e-06, 6.189126e-06, 4.664796e-06, 6.9575e-06, 4.81914e-06, 
    7.832818e-06, 6.673872e-06, 5.347922e-06, 1.74812e-06, 1.071595e-06, 
    1.353722e-06, 1.501342e-06, 3.009961e-06, 2.817259e-06, 2.789365e-06,
  5.202651e-06, 5.374829e-06, 3.532962e-06, 4.02072e-06, 6.24525e-06, 
    5.705242e-06, 4.774315e-06, 3.977761e-06, 2.301015e-06, 1.340395e-06, 
    6.095675e-07, 1.406932e-06, 4.484343e-06, 3.977695e-06, 1.696142e-06,
  3.942326e-06, 3.781649e-06, 2.497299e-06, 1.488556e-06, 1.062494e-05, 
    5.475255e-06, 5.122127e-06, 3.714628e-06, 5.723348e-07, 1.613288e-06, 
    8.953614e-07, 1.816188e-06, 4.470126e-06, 5.289629e-06, 1.545795e-06,
  4.423277e-06, 3.373944e-06, 2.142048e-06, 1.491173e-06, 9.023289e-06, 
    8.5804e-06, 6.069225e-06, 4.207462e-06, 1.807032e-06, 5.734832e-07, 
    1.366527e-06, 1.733607e-06, 4.815189e-06, 5.811378e-06, 2.883157e-06,
  1.241419e-05, 1.048577e-05, 1.100666e-05, 1.048658e-05, 1.014729e-05, 
    5.650103e-06, 1.502592e-06, 1.115745e-06, 7.221474e-07, 1.796544e-06, 
    1.925524e-06, 1.633026e-06, 2.889172e-06, 4.326965e-06, 3.650031e-06,
  9.729289e-06, 8.095459e-06, 1.101892e-05, 1.044034e-05, 1.040897e-05, 
    1.022967e-05, 1.751421e-06, 1.424005e-06, 1.297349e-06, 1.364924e-06, 
    1.093331e-06, 1.511017e-06, 1.786952e-06, 3.082905e-06, 3.581192e-06,
  6.808677e-06, 8.020354e-06, 1.044243e-05, 1.180702e-05, 1.032474e-05, 
    1.074587e-05, 2.561521e-06, 3.138826e-06, 1.074729e-06, 7.702349e-07, 
    9.756372e-07, 9.769066e-07, 2.620263e-06, 3.420831e-06, 4.113109e-06,
  7.891406e-06, 7.677697e-06, 7.996483e-06, 1.038055e-05, 1.031398e-05, 
    1.043011e-05, 4.168259e-06, 2.8998e-06, 1.208911e-06, 1.048947e-06, 
    8.219203e-07, 1.594257e-06, 2.778265e-06, 3.774914e-06, 3.696641e-06,
  7.914563e-06, 6.491431e-06, 6.878758e-06, 9.434465e-06, 1.101488e-05, 
    1.047357e-05, 1.08289e-05, 1.877066e-06, 1.592126e-06, 7.837667e-07, 
    7.622596e-07, 1.920409e-06, 3.287844e-06, 3.663358e-06, 5.396342e-06,
  8.218885e-06, 7.357188e-06, 6.115114e-06, 9.182386e-06, 9.902566e-06, 
    9.49672e-06, 1.01573e-05, 4.838193e-06, 2.042688e-06, 6.940461e-07, 
    1.087472e-06, 1.090461e-06, 3.577305e-06, 3.709625e-06, 4.594695e-06,
  1.214343e-05, 7.987162e-06, 7.592212e-06, 1.056869e-05, 9.868797e-06, 
    1.017973e-05, 9.525384e-06, 6.445595e-06, 2.025718e-06, 1.100307e-06, 
    9.786936e-07, 1.223593e-06, 2.725144e-06, 4.178331e-06, 5.536766e-06,
  1.194606e-05, 8.285623e-06, 8.615953e-06, 1.025109e-05, 1.016073e-05, 
    1.028194e-05, 9.450187e-06, 8.387405e-06, 3.190092e-06, 2.674261e-06, 
    6.798153e-07, 8.729165e-07, 1.912033e-06, 4.77692e-06, 5.42524e-06,
  1.251199e-05, 9.597666e-06, 8.323437e-06, 1.015283e-05, 9.323749e-06, 
    9.493763e-06, 9.894251e-06, 1.020887e-05, 5.269497e-06, 1.899216e-06, 
    1.876966e-06, 1.867277e-06, 2.696447e-06, 3.702633e-06, 6.049786e-06,
  1.140221e-05, 8.335388e-06, 8.048777e-06, 1.074287e-05, 9.489127e-06, 
    9.827269e-06, 8.448327e-06, 9.625039e-06, 7.118504e-06, 1.971234e-06, 
    1.86544e-06, 1.527985e-06, 3.39179e-06, 3.527764e-06, 5.76309e-06,
  4.567215e-06, 1.147767e-06, 5.178413e-06, 1.524237e-05, 1.670319e-05, 
    1.290409e-05, 4.347477e-06, 1.135873e-06, 5.906473e-07, 2.184771e-06, 
    4.167138e-06, 6.136177e-06, 7.742507e-06, 9.840088e-06, 1.030611e-05,
  5.174956e-06, 2.436401e-06, 3.269652e-06, 1.316097e-05, 1.740572e-05, 
    1.734308e-05, 6.407492e-06, 1.3076e-06, 2.018711e-06, 2.52102e-06, 
    3.023735e-06, 5.140121e-06, 6.840191e-06, 8.971502e-06, 1.06149e-05,
  4.525194e-06, 3.040336e-06, 4.336267e-06, 1.241756e-05, 2.026718e-05, 
    2.1003e-05, 6.421264e-06, 2.692433e-06, 1.932175e-06, 1.938258e-06, 
    3.079697e-06, 4.389484e-06, 5.414563e-06, 6.996493e-06, 8.31034e-06,
  5.029156e-06, 4.853154e-06, 5.091517e-06, 9.204877e-06, 1.668711e-05, 
    1.273096e-05, 8.518366e-06, 4.471423e-06, 3.320303e-06, 2.587966e-06, 
    3.516332e-06, 4.901429e-06, 5.477318e-06, 6.690773e-06, 7.150813e-06,
  8.402337e-06, 6.380531e-06, 5.979612e-06, 7.972932e-06, 1.123684e-05, 
    1.361953e-05, 1.364993e-05, 5.636283e-06, 2.560108e-06, 2.676185e-06, 
    4.504257e-06, 4.662661e-06, 5.262455e-06, 6.160641e-06, 7.728511e-06,
  7.98456e-06, 7.584163e-06, 6.610441e-06, 6.02083e-06, 8.442187e-06, 
    1.007874e-05, 1.307612e-05, 6.777657e-06, 7.196633e-06, 4.540725e-06, 
    4.247369e-06, 4.265539e-06, 3.97834e-06, 5.410091e-06, 6.377408e-06,
  7.4733e-06, 9.712095e-06, 8.816303e-06, 8.474725e-06, 5.826013e-06, 
    6.077101e-06, 1.306075e-05, 9.718318e-06, 5.189971e-06, 3.428886e-06, 
    3.462389e-06, 3.675688e-06, 4.789261e-06, 4.825391e-06, 5.346033e-06,
  7.509623e-06, 8.154838e-06, 9.779183e-06, 7.49932e-06, 6.230154e-06, 
    7.424962e-06, 1.131054e-05, 9.016809e-06, 7.71335e-06, 6.85277e-06, 
    6.988128e-06, 5.983629e-06, 5.680068e-06, 4.643435e-06, 4.673951e-06,
  3.734903e-06, 5.335019e-06, 1.133338e-05, 9.210308e-06, 6.912306e-06, 
    9.866256e-06, 9.953621e-06, 8.748711e-06, 1.018648e-05, 7.879904e-06, 
    6.125231e-06, 4.627025e-06, 5.365941e-06, 4.872798e-06, 4.56974e-06,
  4.468121e-06, 2.863039e-06, 1.033289e-05, 9.105282e-06, 7.382948e-06, 
    7.890709e-06, 1.001895e-05, 8.677896e-06, 9.278664e-06, 7.7781e-06, 
    4.533487e-06, 5.908433e-06, 5.647605e-06, 5.278051e-06, 5.489937e-06,
  4.639131e-06, 6.190467e-06, 1.597714e-06, 5.818528e-07, 4.871613e-06, 
    1.060894e-05, 1.11699e-05, 7.241254e-06, 6.14366e-06, 3.976187e-06, 
    3.845498e-06, 4.94216e-06, 7.253983e-06, 1.109049e-05, 1.135247e-05,
  2.110284e-06, 2.961606e-06, 4.953723e-06, 8.53502e-08, 3.432757e-06, 
    1.278853e-05, 1.390871e-05, 9.444767e-06, 9.29038e-06, 6.033445e-06, 
    4.939927e-06, 5.36968e-06, 6.179169e-06, 1.022433e-05, 1.234868e-05,
  1.265676e-06, 7.592783e-07, 3.548477e-06, 1.643632e-07, 5.144065e-07, 
    1.397816e-05, 2.09169e-05, 1.550255e-05, 1.107924e-05, 6.94975e-06, 
    6.535567e-06, 5.419889e-06, 6.777766e-06, 9.89948e-06, 1.091891e-05,
  6.971253e-07, 1.779102e-06, 1.32859e-06, 3.397729e-06, 1.538081e-07, 
    8.878334e-06, 1.968823e-05, 1.828421e-05, 1.072142e-05, 8.638646e-06, 
    7.102143e-06, 6.146493e-06, 7.311698e-06, 1.090226e-05, 1.05104e-05,
  2.451488e-06, 4.53648e-06, 5.039516e-06, 5.227179e-06, 9.885163e-07, 
    3.287807e-06, 8.844746e-06, 1.227621e-05, 1.352912e-05, 8.483483e-06, 
    8.589666e-06, 6.752915e-06, 8.078478e-06, 9.955428e-06, 9.789879e-06,
  2.345757e-06, 2.752242e-06, 4.814091e-06, 4.617257e-06, 5.241575e-06, 
    1.303961e-06, 2.789009e-06, 9.769074e-06, 1.2163e-05, 8.284742e-06, 
    8.552203e-06, 9.052489e-06, 8.211327e-06, 9.464062e-06, 9.687156e-06,
  3.897943e-06, 1.888432e-06, 2.907711e-06, 4.76316e-06, 4.267695e-06, 
    1.887195e-06, 2.378136e-06, 9.243035e-06, 9.716389e-06, 9.770837e-06, 
    7.86124e-06, 9.652717e-06, 9.328384e-06, 7.79776e-06, 9.572343e-06,
  4.470039e-06, 4.033783e-06, 2.84113e-06, 7.51679e-06, 6.260078e-06, 
    1.559261e-06, 1.143147e-06, 6.985581e-06, 1.138859e-05, 9.507968e-06, 
    9.544065e-06, 9.811549e-06, 9.24978e-06, 8.58641e-06, 8.221084e-06,
  2.539e-06, 4.393349e-06, 1.832714e-06, 6.366782e-06, 8.395932e-06, 
    6.494436e-06, 2.170083e-06, 7.278424e-06, 9.136037e-06, 1.089384e-05, 
    1.007729e-05, 9.387557e-06, 9.388668e-06, 8.841009e-06, 8.668066e-06,
  1.318112e-06, 4.007268e-06, 3.16311e-06, 3.482387e-06, 9.273062e-06, 
    8.25237e-06, 6.081169e-06, 5.202121e-06, 7.313098e-06, 8.743695e-06, 
    9.808231e-06, 9.834757e-06, 1.038363e-05, 8.396998e-06, 9.17729e-06,
  7.15841e-06, 7.630306e-06, 2.708215e-06, 2.064196e-06, 3.132282e-06, 
    7.998326e-06, 1.078943e-05, 1.294053e-05, 9.680182e-06, 4.649866e-06, 
    3.553363e-06, 4.969795e-06, 5.406704e-06, 6.987236e-06, 7.610732e-06,
  5.842625e-06, 3.651964e-06, 8.206085e-06, 3.820894e-06, 2.370865e-06, 
    4.921941e-06, 8.229702e-06, 1.017746e-05, 6.715412e-06, 4.328923e-06, 
    3.854871e-06, 5.631137e-06, 7.347205e-06, 7.223248e-06, 7.77396e-06,
  4.997949e-06, 4.086061e-06, 6.890565e-06, 6.388668e-06, 1.620211e-06, 
    2.177373e-06, 4.56294e-06, 3.492473e-06, 5.670804e-06, 4.52314e-06, 
    3.964115e-06, 5.679811e-06, 6.353272e-06, 7.346334e-06, 6.403527e-06,
  3.090285e-06, 2.992617e-06, 7.618349e-06, 7.422293e-06, 3.203368e-06, 
    1.459377e-06, 3.623309e-06, 3.079842e-06, 3.999147e-06, 3.964803e-06, 
    4.165063e-06, 5.390929e-06, 5.693123e-06, 7.635567e-06, 6.882216e-06,
  1.929472e-06, 3.53516e-06, 5.50277e-06, 6.844894e-06, 4.843718e-06, 
    4.231151e-06, 2.90466e-06, 8.894065e-07, 3.68758e-06, 5.034412e-06, 
    4.562866e-06, 5.632296e-06, 8.150398e-06, 7.717313e-06, 9.351103e-06,
  1.639793e-06, 1.303723e-06, 1.403288e-06, 4.286272e-06, 5.731987e-06, 
    4.170886e-06, 3.013006e-06, 3.296846e-06, 3.65144e-06, 6.285404e-06, 
    4.596924e-06, 6.320955e-06, 7.489083e-06, 8.205973e-06, 9.654923e-06,
  9.627183e-07, 2.081168e-06, 2.730162e-06, 1.917718e-06, 3.956143e-06, 
    1.8304e-06, 1.640767e-06, 1.235179e-05, 3.495106e-06, 4.073274e-06, 
    2.14896e-06, 6.518248e-06, 7.453308e-06, 8.238379e-06, 1.026322e-05,
  1.222742e-06, 1.648968e-06, 5.031619e-06, 2.940609e-06, 3.363074e-06, 
    4.049427e-06, 3.747448e-06, 7.373318e-06, 6.437169e-06, 4.020189e-06, 
    3.426321e-06, 6.15798e-06, 7.850704e-06, 7.779995e-06, 8.131156e-06,
  9.456466e-07, 4.057675e-06, 4.660916e-06, 5.957653e-06, 6.027642e-06, 
    6.803507e-06, 6.85043e-06, 7.701286e-06, 6.496509e-06, 7.742834e-06, 
    3.803072e-06, 5.78258e-06, 6.992743e-06, 8.237904e-06, 9.374229e-06,
  8.479823e-07, 1.908869e-06, 4.686695e-06, 6.062984e-06, 8.560211e-06, 
    9.008776e-06, 1.112938e-05, 7.13693e-06, 7.67362e-06, 1.149302e-05, 
    5.888416e-06, 6.118055e-06, 6.766676e-06, 6.560022e-06, 6.270888e-06,
  1.159508e-05, 1.073517e-05, 5.660293e-06, 4.289216e-06, 2.11045e-06, 
    1.271419e-09, 6.685053e-08, 4.712744e-07, 3.671641e-06, 5.31617e-06, 
    4.691109e-06, 7.811223e-06, 8.29424e-06, 7.836008e-06, 7.501173e-06,
  1.076151e-05, 9.839198e-06, 3.701758e-06, 3.098592e-06, 2.924635e-06, 
    1.432567e-07, 3.033381e-07, 2.034816e-06, 4.576745e-06, 4.082533e-06, 
    5.520768e-06, 6.398933e-06, 5.525044e-06, 7.654538e-06, 7.146303e-06,
  9.288873e-06, 7.917698e-06, 1.026839e-06, 5.927894e-06, 1.249571e-06, 
    1.812524e-06, 2.514159e-06, 4.534956e-06, 4.989015e-06, 3.359305e-06, 
    4.282666e-06, 5.13249e-06, 5.547836e-06, 4.940487e-06, 5.694486e-06,
  8.2443e-06, 7.687608e-06, 2.127601e-06, 5.930837e-06, 4.008781e-06, 
    2.123606e-06, 2.382591e-06, 3.557721e-06, 4.530714e-06, 5.187345e-06, 
    2.744151e-06, 4.455741e-06, 5.777285e-06, 3.970906e-06, 4.92156e-06,
  6.276091e-06, 4.902258e-06, 6.650481e-06, 5.107619e-06, 2.242752e-06, 
    3.842102e-06, 5.277126e-06, 4.959236e-06, 6.117104e-06, 3.553872e-06, 
    2.45056e-06, 3.364568e-06, 3.208233e-06, 4.389491e-06, 5.310828e-06,
  3.002988e-06, 5.363944e-06, 6.942924e-06, 5.437768e-06, 7.164906e-06, 
    7.107215e-06, 8.515623e-06, 6.96447e-06, 6.729363e-06, 3.387216e-06, 
    2.444839e-06, 2.89435e-06, 3.3172e-06, 4.469202e-06, 4.102846e-06,
  2.091324e-06, 6.716687e-06, 6.040862e-06, 6.916441e-06, 6.793338e-06, 
    3.865407e-06, 5.811818e-06, 8.100941e-06, 7.995918e-06, 6.402445e-06, 
    3.425411e-06, 3.583154e-06, 3.738446e-06, 4.282774e-06, 5.404214e-06,
  1.715713e-06, 3.568772e-06, 6.664359e-06, 5.723638e-06, 3.734588e-06, 
    4.210313e-06, 7.599356e-06, 5.296945e-06, 1.080425e-05, 1.111646e-05, 
    9.829648e-06, 8.385869e-06, 6.339519e-06, 5.963816e-06, 5.863958e-06,
  1.226892e-06, 1.999111e-06, 2.338949e-06, 1.24581e-06, 1.107992e-06, 
    3.097081e-06, 3.28667e-06, 5.04835e-06, 8.489244e-06, 1.377096e-05, 
    1.326933e-05, 9.362444e-06, 9.690522e-06, 7.997078e-06, 1.075552e-05,
  1.112317e-06, 6.605831e-07, 6.027004e-07, 1.004007e-06, 2.404195e-07, 
    1.020288e-07, 5.609836e-07, 1.337821e-06, 1.546804e-06, 2.686661e-06, 
    2.444517e-06, 5.485449e-06, 8.758083e-06, 1.715265e-05, 1.557617e-05,
  6.146815e-06, 5.791594e-06, 1.127717e-05, 2.035276e-05, 1.618621e-05, 
    1.309542e-06, 6.550993e-07, 2.697439e-06, 2.348942e-06, 3.875132e-06, 
    5.564873e-06, 5.874141e-06, 5.116378e-06, 6.250942e-06, 7.012979e-06,
  6.390956e-06, 5.733918e-06, 1.572314e-05, 2.539761e-05, 1.191105e-05, 
    1.400851e-06, 5.556294e-07, 2.543504e-06, 2.889169e-06, 5.612067e-06, 
    5.81543e-06, 4.803639e-06, 3.979047e-06, 6.776092e-06, 7.666672e-06,
  8.69034e-06, 1.254106e-05, 1.832465e-05, 1.669875e-05, 7.006449e-06, 
    8.720025e-07, 3.267649e-06, 2.401075e-06, 4.012463e-06, 4.108158e-06, 
    6.788265e-06, 6.48251e-06, 5.346065e-06, 5.29474e-06, 5.619203e-06,
  9.671003e-06, 1.312892e-05, 1.892701e-05, 1.333904e-05, 5.016739e-06, 
    1.021253e-07, 2.717148e-06, 2.111793e-06, 4.140204e-06, 4.403144e-06, 
    7.633777e-06, 6.578276e-06, 5.320675e-06, 5.986506e-06, 5.175357e-06,
  1.424311e-05, 1.917045e-05, 1.722439e-05, 1.41195e-05, 1.582533e-06, 
    2.602449e-06, 3.047702e-06, 4.328107e-06, 6.29086e-06, 5.473608e-06, 
    6.840944e-06, 6.861691e-06, 6.232388e-06, 4.467007e-06, 8.540269e-06,
  1.758691e-05, 2.004174e-05, 1.731046e-05, 8.187718e-06, 1.335007e-07, 
    2.360229e-06, 3.153912e-06, 6.065496e-06, 5.604696e-06, 4.337443e-06, 
    3.610959e-06, 8.392512e-06, 6.302681e-06, 5.904306e-06, 5.160522e-06,
  2.264104e-05, 1.642568e-05, 1.199624e-05, 6.57543e-06, 1.852962e-06, 
    2.692904e-06, 6.664577e-06, 5.462153e-06, 5.121685e-06, 5.523235e-06, 
    4.853948e-06, 7.570413e-06, 6.127768e-06, 6.532328e-06, 4.263073e-06,
  2.075665e-05, 1.156169e-05, 6.885265e-06, 2.214308e-06, 4.703402e-06, 
    6.127109e-06, 7.250476e-06, 7.536508e-06, 3.912151e-06, 4.81157e-06, 
    6.257785e-06, 8.451811e-06, 7.82696e-06, 8.866746e-06, 8.304529e-06,
  1.807263e-05, 8.833008e-06, 3.984084e-06, 2.8294e-06, 4.608897e-06, 
    5.886235e-06, 3.982608e-06, 3.699631e-06, 3.00865e-06, 3.214125e-06, 
    2.75984e-06, 4.831033e-06, 7.104636e-06, 8.261304e-06, 7.643343e-06,
  1.115678e-05, 6.454689e-06, 3.422803e-06, 3.407799e-06, 2.954869e-06, 
    3.74374e-06, 7.445746e-06, 6.947017e-06, 7.906006e-06, 3.380636e-06, 
    1.340292e-06, 9.72092e-07, 4.330774e-07, 1.210076e-07, 4.069791e-06,
  1.243238e-05, 1.075587e-05, 4.675619e-06, 3.079912e-06, 1.526676e-05, 
    2.464574e-05, 2.043611e-05, 4.535941e-06, 1.411137e-06, 4.124173e-06, 
    5.526746e-06, 7.309553e-06, 9.663456e-06, 7.261957e-06, 5.744837e-06,
  1.489895e-05, 1.423277e-05, 6.942196e-06, 6.241378e-06, 1.911848e-05, 
    2.994232e-05, 1.556192e-05, 4.279923e-06, 2.089003e-06, 4.120714e-06, 
    6.792937e-06, 7.731417e-06, 7.935091e-06, 6.719984e-06, 6.374219e-06,
  1.437265e-05, 1.715405e-05, 5.347179e-06, 5.324856e-06, 1.784743e-05, 
    2.255269e-05, 1.440865e-05, 3.659929e-06, 5.250253e-06, 4.672198e-06, 
    6.794507e-06, 5.255525e-06, 5.663829e-06, 6.726808e-06, 7.293937e-06,
  1.202492e-05, 1.114355e-05, 5.361151e-06, 9.578079e-06, 1.776321e-05, 
    1.963278e-05, 1.193064e-05, 3.762541e-06, 6.484941e-06, 1.020464e-05, 
    6.496085e-06, 5.346394e-06, 8.363717e-06, 9.733888e-06, 5.685223e-06,
  9.35239e-06, 1.230514e-05, 9.169279e-06, 1.254445e-05, 1.946513e-05, 
    2.041223e-05, 1.208513e-05, 6.280397e-06, 4.846921e-06, 8.479267e-06, 
    7.313836e-06, 6.286497e-06, 7.442385e-06, 6.686736e-06, 7.384779e-06,
  7.247347e-06, 1.189842e-05, 9.024304e-06, 1.142221e-05, 1.954409e-05, 
    1.583424e-05, 1.026863e-05, 1.008401e-05, 8.258079e-06, 9.076792e-06, 
    6.360519e-06, 5.353008e-06, 3.550008e-06, 2.860509e-06, 5.564226e-06,
  5.095195e-06, 9.122179e-06, 7.266527e-06, 1.366994e-05, 2.124546e-05, 
    1.569703e-05, 8.959501e-06, 6.479575e-06, 1.30361e-05, 1.048371e-05, 
    9.630438e-06, 9.032738e-06, 7.151012e-06, 4.780751e-06, 4.620292e-06,
  6.307715e-06, 5.877168e-06, 7.23373e-06, 1.27326e-05, 1.638303e-05, 
    1.488674e-05, 6.768948e-06, 5.700944e-06, 5.476241e-06, 8.305924e-06, 
    1.108298e-05, 1.487369e-05, 1.576978e-05, 1.419699e-05, 9.396478e-06,
  4.967161e-06, 5.124695e-06, 1.078799e-05, 1.291396e-05, 1.539579e-05, 
    7.141309e-06, 3.965514e-06, 5.291778e-06, 1.520055e-05, 6.844331e-06, 
    1.252308e-05, 1.209025e-05, 1.397066e-05, 1.194872e-05, 9.701307e-06,
  3.932572e-06, 5.848082e-06, 1.267335e-05, 1.12892e-05, 1.12874e-05, 
    9.453987e-06, 9.087822e-06, 6.105303e-06, 7.953201e-06, 1.371522e-05, 
    1.181649e-05, 1.088557e-05, 1.046704e-05, 7.538706e-06, 6.854688e-06,
  6.760632e-06, 5.594545e-06, 2.452601e-06, 3.294002e-06, 1.166614e-05, 
    2.165989e-05, 1.940168e-05, 6.843857e-06, 2.083535e-06, 3.528963e-06, 
    6.293434e-06, 7.148558e-06, 4.677843e-06, 3.862378e-06, 5.170473e-06,
  9.936845e-06, 8.224757e-06, 6.018105e-07, 3.807522e-06, 8.976565e-06, 
    2.32528e-05, 1.832863e-05, 5.043561e-06, 2.256005e-06, 4.168892e-06, 
    7.754462e-06, 8.565143e-06, 5.333495e-06, 3.178489e-06, 4.692566e-06,
  1.223636e-05, 4.764388e-06, 1.955927e-06, 6.244996e-06, 1.313299e-05, 
    2.218805e-05, 1.605283e-05, 4.202853e-06, 2.64455e-06, 8.777103e-06, 
    1.09182e-05, 1.071486e-05, 6.230473e-06, 4.803471e-06, 5.202344e-06,
  1.037131e-05, 7.15032e-06, 4.923821e-06, 9.535791e-06, 8.368045e-06, 
    2.561576e-05, 1.541031e-05, 5.538449e-06, 4.101874e-06, 1.132847e-05, 
    1.491383e-05, 1.278316e-05, 8.303249e-06, 5.461792e-06, 7.792616e-06,
  8.630671e-06, 1.060411e-05, 5.830913e-06, 5.883606e-06, 8.38214e-06, 
    1.824668e-05, 1.66638e-05, 6.528883e-06, 7.468029e-06, 1.352689e-05, 
    1.574412e-05, 1.641327e-05, 1.135749e-05, 5.161143e-06, 6.769262e-06,
  7.033607e-06, 1.125298e-05, 7.847459e-06, 5.309939e-06, 6.763262e-06, 
    1.393762e-05, 1.729254e-05, 7.660149e-06, 1.082158e-05, 1.312425e-05, 
    1.798501e-05, 2.08759e-05, 1.533913e-05, 8.760571e-06, 6.295539e-06,
  4.634407e-06, 5.623057e-06, 1.076309e-05, 6.365313e-06, 6.301259e-06, 
    1.190992e-05, 1.562102e-05, 8.754484e-06, 8.105729e-06, 1.218675e-05, 
    1.521838e-05, 1.655775e-05, 1.532745e-05, 1.024896e-05, 9.000008e-06,
  5.198755e-06, 5.411262e-06, 1.251916e-05, 9.390698e-06, 1.084295e-05, 
    9.722581e-06, 1.249536e-05, 8.455811e-06, 5.900512e-06, 9.567227e-06, 
    9.844354e-06, 1.203758e-05, 1.149629e-05, 1.016672e-05, 1.016875e-05,
  5.81525e-06, 5.923853e-06, 8.242268e-06, 9.095555e-06, 1.16033e-05, 
    7.78122e-06, 1.023131e-05, 8.193475e-06, 1.074326e-05, 6.279653e-06, 
    9.452276e-06, 1.157125e-05, 9.639595e-06, 7.116974e-06, 7.433461e-06,
  6.982722e-06, 5.886775e-06, 7.134895e-06, 1.14744e-05, 1.264963e-05, 
    6.957025e-06, 1.087748e-05, 6.733964e-06, 1.01425e-05, 5.546901e-06, 
    1.022532e-05, 8.925971e-06, 7.269179e-06, 5.586751e-06, 7.979002e-06,
  0.0002317766, 9.525319e-05, 0.0001077011, 2.884522e-05, 1.525852e-05, 
    5.499544e-06, 3.645964e-06, 2.915915e-06, 3.652466e-06, 5.180048e-06, 
    5.430097e-06, 3.158677e-06, 2.147008e-06, 1.563065e-06, 2.304681e-06,
  0.00020175, 0.0001357627, 4.746462e-05, 2.483159e-05, 1.013394e-05, 
    6.641088e-06, 3.074567e-06, 4.387652e-06, 7.699635e-06, 9.53662e-06, 
    8.288297e-06, 4.186939e-06, 2.168161e-06, 1.531098e-06, 2.473192e-06,
  0.0001683106, 0.0001345367, 8.099504e-05, 3.800547e-05, 8.106937e-06, 
    4.648944e-06, 9.078151e-06, 1.402045e-05, 1.66148e-05, 1.380707e-05, 
    9.6355e-06, 5.45783e-06, 2.926284e-06, 2.121455e-06, 3.748896e-06,
  0.0001770823, 0.0001493898, 9.280706e-05, 4.923383e-05, 1.472424e-05, 
    1.480701e-05, 1.975551e-05, 2.143673e-05, 2.245765e-05, 1.725417e-05, 
    1.106952e-05, 7.821199e-06, 5.057237e-06, 3.594224e-06, 4.240218e-06,
  0.0001672139, 0.0001364146, 6.971272e-05, 2.053329e-05, 1.212753e-05, 
    2.628129e-05, 2.28912e-05, 1.642937e-05, 1.843867e-05, 1.690714e-05, 
    1.455123e-05, 1.132407e-05, 8.251343e-06, 4.907659e-06, 4.608609e-06,
  0.0001391886, 0.0001009757, 4.282058e-05, 1.415458e-05, 1.780665e-05, 
    2.336392e-05, 2.222415e-05, 1.465527e-05, 1.068153e-05, 1.202862e-05, 
    1.341205e-05, 1.347143e-05, 9.363573e-06, 6.799964e-06, 4.692006e-06,
  9.946797e-05, 7.005563e-05, 3.000417e-05, 2.015894e-05, 2.277508e-05, 
    2.907106e-05, 1.909826e-05, 1.443004e-05, 1.361138e-05, 7.392438e-06, 
    8.901955e-06, 1.126016e-05, 8.053253e-06, 7.79873e-06, 5.841207e-06,
  4.526855e-05, 3.869187e-05, 2.783378e-05, 1.88328e-05, 2.038638e-05, 
    2.333098e-05, 1.934407e-05, 1.724289e-05, 1.248528e-05, 6.294373e-06, 
    7.791492e-06, 5.354531e-06, 6.351296e-06, 6.581653e-06, 7.54037e-06,
  1.171095e-05, 1.267404e-05, 1.26922e-05, 1.140859e-05, 1.035722e-05, 
    1.450226e-05, 1.559955e-05, 1.360025e-05, 9.44851e-06, 7.032445e-06, 
    6.255081e-06, 4.935417e-06, 4.022773e-06, 5.213567e-06, 5.921926e-06,
  1.288782e-05, 1.088426e-05, 8.699097e-06, 9.10776e-06, 9.495253e-06, 
    7.812808e-06, 7.250724e-06, 7.227651e-06, 5.556502e-06, 6.339996e-06, 
    4.444841e-06, 4.60389e-06, 5.145864e-06, 3.47356e-06, 2.193811e-06,
  3.673614e-05, 2.887308e-05, 1.530803e-05, 1.974009e-05, 1.361663e-05, 
    2.718523e-05, 3.428612e-05, 5.812949e-05, 3.505001e-05, 1.955053e-05, 
    1.425313e-05, 3.892118e-06, 1.100575e-06, 9.844273e-07, 4.469396e-07,
  5.037397e-05, 2.544969e-05, 1.942443e-05, 1.569616e-05, 2.185831e-05, 
    2.625998e-05, 3.665582e-05, 5.522947e-05, 4.701333e-05, 3.090331e-05, 
    1.820918e-05, 2.557441e-06, 6.551986e-07, 1.83625e-07, 5.904369e-07,
  4.904955e-05, 3.534009e-05, 2.802723e-05, 1.830058e-05, 1.577021e-05, 
    3.589074e-05, 4.235292e-05, 4.088481e-05, 4.057392e-05, 2.177756e-05, 
    1.136227e-05, 1.989369e-06, 2.208495e-07, 2.400214e-07, 1.451644e-06,
  4.23667e-05, 4.796633e-05, 5.29725e-05, 2.880848e-05, 2.232355e-05, 
    3.493064e-05, 4.606323e-05, 4.61035e-05, 3.766423e-05, 1.497123e-05, 
    8.633962e-06, 1.424015e-06, 7.942507e-07, 1.801289e-06, 2.321667e-06,
  3.666371e-05, 0.0001041855, 0.00012492, 6.876401e-05, 3.096171e-05, 
    3.513175e-05, 4.10882e-05, 4.343621e-05, 3.377494e-05, 1.574186e-05, 
    3.187202e-06, 2.467049e-06, 1.603129e-06, 2.350047e-06, 6.849356e-07,
  0.0001000162, 0.0001818178, 0.0002086455, 8.452144e-05, 3.271748e-05, 
    3.316303e-05, 3.345275e-05, 4.387762e-05, 3.189715e-05, 1.690968e-05, 
    2.920701e-06, 2.537255e-06, 2.116095e-06, 1.712868e-06, 6.481915e-07,
  0.0002606931, 0.0002877959, 0.0002469854, 9.162731e-05, 3.990093e-05, 
    2.72175e-05, 3.624713e-05, 4.658761e-05, 3.633592e-05, 2.046845e-05, 
    3.73769e-06, 1.704042e-06, 1.597476e-06, 1.418636e-06, 7.187709e-07,
  0.0004545233, 0.0003924262, 0.0002563988, 0.0001042809, 3.647989e-05, 
    6.487287e-05, 2.968535e-05, 3.339961e-05, 3.857799e-05, 1.291057e-05, 
    4.695854e-06, 4.247473e-06, 3.522361e-06, 2.248936e-06, 3.787167e-06,
  0.0005387693, 0.0004072531, 0.0002388509, 0.0001019554, 6.744323e-05, 
    4.340553e-05, 3.226699e-05, 3.687059e-05, 2.828535e-05, 8.827841e-06, 
    4.203901e-06, 4.923056e-06, 6.15777e-06, 9.905515e-06, 6.559286e-06,
  0.0004647532, 0.0003185739, 0.0001660251, 8.439686e-05, 7.796365e-05, 
    6.688836e-05, 3.162286e-05, 2.547953e-05, 1.202104e-05, 4.197944e-06, 
    4.909306e-06, 4.249456e-06, 3.780093e-06, 3.251578e-06, 3.850521e-06,
  8.482596e-07, 6.406486e-07, 5.426635e-07, 2.57549e-07, 7.067123e-07, 
    2.56965e-06, 6.467599e-06, 3.909823e-06, 1.395423e-06, 6.40446e-07, 
    2.142153e-06, 1.418439e-05, 2.471744e-05, 1.582867e-05, 2.075734e-06,
  7.174014e-07, 9.416901e-07, 4.868816e-07, 5.049787e-08, 2.720179e-07, 
    4.901419e-07, 2.062446e-06, 1.838866e-06, 4.665951e-07, 1.199905e-06, 
    3.6664e-06, 2.86326e-05, 3.47345e-05, 1.034041e-05, 1.005699e-06,
  2.529544e-06, 1.010945e-06, 4.83656e-07, 8.237354e-08, 5.319577e-08, 
    9.365155e-08, 3.602948e-07, 4.058977e-07, 2.652506e-07, 4.085182e-07, 
    5.131807e-06, 1.721809e-05, 3.046838e-05, 8.003889e-06, 1.573306e-06,
  5.146715e-06, 2.325887e-06, 1.210057e-06, 4.711096e-07, 3.088547e-07, 
    1.592729e-07, 6.303693e-08, 9.473234e-08, 2.268862e-07, 1.26962e-06, 
    4.911627e-06, 1.565444e-05, 2.26506e-05, 1.028868e-05, 1.425126e-06,
  9.617206e-06, 8.364976e-06, 3.799651e-06, 1.272481e-06, 6.95183e-07, 
    4.260349e-07, 1.591548e-07, 7.151171e-08, 1.366887e-06, 1.300289e-06, 
    4.459437e-06, 9.812631e-06, 1.898005e-05, 1.210373e-05, 2.139825e-06,
  1.451917e-05, 1.138599e-05, 7.153332e-06, 2.131348e-06, 3.149216e-07, 
    4.762887e-07, 5.032347e-07, 2.415759e-07, 6.734214e-07, 1.820172e-06, 
    4.735622e-06, 7.134001e-06, 1.599095e-05, 9.050332e-06, 1.904215e-06,
  1.807281e-05, 1.451491e-05, 1.458235e-05, 4.983532e-06, 9.276068e-07, 
    2.381226e-07, 6.765273e-07, 5.631146e-07, 1.766642e-07, 4.527112e-06, 
    5.807015e-06, 5.38247e-06, 1.179863e-05, 1.039901e-05, 2.655653e-06,
  3.228042e-05, 1.671253e-05, 1.734032e-05, 8.471006e-06, 2.443946e-06, 
    1.064452e-06, 1.168628e-06, 6.018428e-07, 3.241572e-07, 7.947307e-06, 
    5.105255e-06, 4.979654e-06, 1.101775e-05, 3.984713e-06, 2.902263e-06,
  2.803928e-05, 2.406964e-05, 1.911268e-05, 7.462379e-06, 4.081662e-06, 
    1.625339e-06, 5.388037e-07, 1.375668e-06, 3.770586e-06, 8.388219e-06, 
    4.632935e-06, 6.064749e-06, 7.336655e-06, 6.34101e-06, 4.353337e-06,
  2.421465e-05, 2.48143e-05, 1.604017e-05, 1.280905e-05, 6.847599e-06, 
    2.507166e-06, 1.624716e-06, 1.403324e-06, 8.16668e-06, 7.715143e-06, 
    5.47003e-06, 6.301229e-06, 7.841079e-06, 4.24926e-06, 1.602439e-06,
  3.195403e-06, 3.376581e-06, 5.472502e-06, 6.419178e-06, 7.880942e-06, 
    8.411521e-06, 9.625954e-06, 1.005772e-05, 6.865966e-06, 4.335782e-06, 
    1.352425e-06, 7.43169e-06, 1.085329e-05, 2.630301e-05, 1.907364e-05,
  4.08971e-06, 4.897429e-06, 5.932928e-06, 6.712717e-06, 7.560148e-06, 
    8.251539e-06, 8.939257e-06, 9.4561e-06, 8.196708e-06, 4.762579e-06, 
    1.638901e-06, 3.392612e-06, 1.012741e-05, 2.396407e-05, 1.651633e-05,
  1.61442e-06, 2.480268e-06, 5.117884e-06, 8.482231e-06, 8.417507e-06, 
    9.633003e-06, 8.246165e-06, 8.977735e-06, 6.94479e-06, 4.064005e-06, 
    2.815803e-06, 2.37118e-06, 8.029768e-06, 1.626814e-05, 1.619444e-05,
  9.143131e-07, 1.295097e-06, 2.687599e-06, 5.877737e-06, 1.024883e-05, 
    1.147406e-05, 9.963509e-06, 9.535123e-06, 5.901068e-06, 4.453992e-06, 
    3.593507e-06, 2.628816e-06, 2.459349e-06, 1.205611e-05, 1.36012e-05,
  1.803088e-06, 2.035793e-06, 2.433141e-06, 3.080316e-06, 6.958821e-06, 
    1.369686e-05, 1.07193e-05, 1.061764e-05, 6.009496e-06, 5.493108e-06, 
    4.048983e-06, 1.793087e-06, 1.015604e-06, 8.126418e-06, 1.533099e-05,
  3.859608e-06, 3.292219e-06, 2.41289e-06, 1.97392e-06, 7.381954e-06, 
    1.323022e-05, 1.326594e-05, 1.321649e-05, 7.987129e-06, 5.471639e-06, 
    5.066478e-06, 2.490822e-06, 5.854203e-07, 6.286627e-06, 1.336326e-05,
  5.013005e-06, 4.276602e-06, 4.257136e-06, 3.796916e-06, 6.537948e-06, 
    1.4058e-05, 1.43523e-05, 1.501084e-05, 7.509981e-06, 3.803455e-06, 
    4.538233e-06, 5.291881e-06, 1.426251e-06, 3.558697e-06, 1.114486e-05,
  7.112067e-06, 5.625322e-06, 6.638038e-06, 6.267707e-06, 7.661287e-06, 
    1.437478e-05, 1.761762e-05, 1.79446e-05, 1.01497e-05, 6.080066e-06, 
    4.666926e-06, 4.775208e-06, 2.148867e-06, 1.097405e-06, 1.059084e-05,
  8.397767e-06, 7.891236e-06, 7.080924e-06, 7.132426e-06, 1.08347e-05, 
    1.500728e-05, 1.673212e-05, 1.69591e-05, 1.244381e-05, 4.351311e-06, 
    5.22912e-06, 4.640244e-06, 3.490222e-06, 2.642913e-06, 9.466979e-06,
  1.120863e-05, 1.030283e-05, 1.007601e-05, 8.377924e-06, 1.097386e-05, 
    1.219808e-05, 1.609678e-05, 1.577888e-05, 1.436411e-05, 8.518117e-06, 
    5.378619e-06, 5.134841e-06, 5.112534e-06, 2.847763e-06, 8.844052e-06,
  3.95771e-06, 5.007581e-06, 6.93226e-06, 6.725794e-06, 3.829888e-06, 
    6.088159e-06, 9.511838e-06, 1.045769e-05, 9.475307e-06, 1.278251e-05, 
    1.485439e-05, 8.035105e-06, 5.807037e-06, 2.890441e-06, 8.993489e-06,
  2.235448e-06, 5.104514e-06, 5.590143e-06, 5.79873e-06, 2.837954e-06, 
    4.783761e-06, 6.953292e-06, 9.930259e-06, 7.673056e-06, 9.2225e-06, 
    1.360353e-05, 1.642718e-05, 7.722576e-06, 5.090397e-06, 3.63508e-06,
  1.921574e-06, 3.997014e-06, 5.534213e-06, 4.894663e-06, 4.941074e-07, 
    3.592138e-06, 7.137305e-06, 7.590429e-06, 9.813456e-06, 1.050089e-05, 
    1.271734e-05, 1.671306e-05, 1.298033e-05, 7.78243e-06, 2.864536e-06,
  2.152522e-06, 4.471746e-06, 4.791964e-06, 4.801132e-06, 1.797602e-07, 
    1.996297e-06, 6.922232e-06, 6.485767e-06, 9.154172e-06, 9.557923e-06, 
    1.103669e-05, 1.532852e-05, 1.843864e-05, 1.037917e-05, 5.03248e-06,
  1.369869e-06, 3.439516e-06, 4.525669e-06, 5.190367e-06, 6.2453e-07, 
    2.158831e-06, 5.225648e-06, 5.954751e-06, 8.253269e-06, 8.212054e-06, 
    1.12149e-05, 1.501857e-05, 1.744132e-05, 1.544833e-05, 8.432138e-06,
  8.252941e-07, 2.884313e-06, 3.733711e-06, 4.114625e-06, 1.455623e-06, 
    2.019038e-06, 4.610366e-06, 6.936684e-06, 7.022844e-06, 7.691287e-06, 
    1.211993e-05, 1.292839e-05, 1.601289e-05, 1.912115e-05, 1.715814e-05,
  4.187292e-07, 1.795415e-06, 1.80437e-06, 3.09509e-06, 1.840233e-06, 
    2.844027e-06, 6.797937e-06, 7.615035e-06, 7.69373e-06, 7.158456e-06, 
    1.264235e-05, 1.58367e-05, 1.677937e-05, 1.667275e-05, 1.792036e-05,
  7.222147e-07, 1.097613e-06, 1.383306e-06, 1.414829e-06, 1.285598e-06, 
    3.155864e-06, 7.077019e-06, 6.775188e-06, 8.546206e-06, 8.821724e-06, 
    1.00764e-05, 1.487157e-05, 1.720763e-05, 1.853141e-05, 1.77885e-05,
  2.628754e-06, 2.227057e-06, 1.486251e-06, 9.604946e-07, 1.081199e-06, 
    2.723093e-06, 7.527005e-06, 7.406138e-06, 9.376537e-06, 8.406574e-06, 
    8.910173e-06, 1.444983e-05, 1.818392e-05, 2.096566e-05, 1.669818e-05,
  2.207892e-06, 2.382517e-06, 1.636324e-06, 1.077026e-06, 1.095057e-06, 
    2.038652e-06, 5.964037e-06, 8.808751e-06, 8.989103e-06, 8.095482e-06, 
    1.101511e-05, 1.257533e-05, 1.613853e-05, 1.662352e-05, 1.867049e-05,
  6.161472e-07, 3.049749e-06, 4.612124e-06, 7.913654e-06, 8.009229e-06, 
    1.965206e-06, 4.864516e-06, 3.678845e-06, 8.84638e-06, 9.569948e-06, 
    7.372738e-06, 6.362452e-06, 6.51813e-06, 6.843874e-06, 7.032389e-06,
  3.597005e-07, 1.378107e-07, 1.918609e-06, 2.278944e-06, 7.689363e-06, 
    2.875206e-06, 6.457393e-06, 4.265214e-06, 6.166605e-06, 8.737968e-06, 
    9.570839e-06, 9.875487e-06, 8.980135e-06, 8.175587e-06, 8.4722e-06,
  1.237621e-06, 1.241264e-07, 4.552403e-08, 9.954215e-07, 2.180853e-06, 
    8.359289e-06, 9.963998e-06, 4.864272e-06, 3.365386e-06, 7.469897e-06, 
    8.357499e-06, 1.074795e-05, 1.224398e-05, 1.009884e-05, 8.535338e-06,
  3.082323e-06, 4.2486e-07, 3.746853e-07, 3.1294e-07, 3.450373e-07, 
    7.872964e-06, 1.222945e-05, 8.692184e-06, 2.513143e-06, 4.597738e-06, 
    1.20146e-05, 1.253061e-05, 1.148345e-05, 1.316457e-05, 1.071966e-05,
  5.11614e-06, 1.640899e-06, 4.453866e-07, 1.431098e-06, 6.468975e-08, 
    2.628162e-06, 5.521747e-06, 8.392017e-06, 1.023133e-05, 4.382447e-06, 
    5.871921e-06, 1.193881e-05, 1.273657e-05, 1.20729e-05, 1.613478e-05,
  6.576232e-06, 1.31502e-06, 9.109933e-07, 8.42551e-07, 7.344498e-07, 
    8.467234e-07, 1.610915e-06, 4.348907e-06, 1.216878e-05, 5.680194e-06, 
    4.306475e-06, 1.262919e-05, 1.378011e-05, 1.527529e-05, 1.619347e-05,
  4.341294e-06, 2.194062e-06, 1.906745e-06, 8.841827e-07, 5.900635e-07, 
    2.542104e-07, 5.572306e-07, 5.381655e-07, 2.434535e-06, 9.766438e-06, 
    4.561711e-06, 9.803432e-06, 1.640485e-05, 1.68569e-05, 1.804154e-05,
  5.002645e-06, 3.203656e-06, 1.394651e-06, 1.497613e-06, 3.971788e-07, 
    2.993065e-07, 4.925621e-07, 3.208146e-08, 1.279275e-06, 5.202147e-07, 
    1.104232e-05, 4.211236e-06, 9.777724e-06, 1.572033e-05, 1.823525e-05,
  4.249508e-06, 3.178263e-06, 1.496539e-06, 4.764073e-07, 2.096509e-07, 
    4.068486e-07, 5.124219e-07, 8.557937e-08, 1.321645e-07, 1.261208e-07, 
    5.088918e-06, 2.826317e-06, 6.116826e-06, 1.171197e-05, 2.066495e-05,
  6.490899e-06, 4.598153e-06, 1.915324e-06, 7.924323e-07, 2.568451e-07, 
    3.96614e-07, 5.12491e-07, 1.205966e-08, 1.782851e-08, 2.980824e-07, 
    4.392928e-07, 5.73463e-07, 2.175643e-06, 7.313429e-06, 1.798155e-05,
  2.11216e-06, 1.241243e-06, 5.381235e-06, 2.672334e-06, 2.301557e-06, 
    5.792947e-06, 7.406191e-06, 3.843576e-06, 4.689709e-06, 5.612918e-06, 
    5.093443e-06, 6.815905e-06, 7.071659e-06, 7.215886e-06, 8.507322e-06,
  6.412448e-06, 1.324611e-06, 9.721003e-06, 2.496062e-06, 7.079427e-07, 
    2.968855e-06, 2.233106e-06, 3.71354e-06, 5.846308e-06, 6.430398e-06, 
    6.07202e-06, 8.176533e-06, 9.674241e-06, 7.486226e-06, 9.773674e-06,
  1.103292e-05, 3.947912e-06, 8.014446e-06, 5.693944e-06, 2.678409e-06, 
    5.298175e-07, 1.251545e-06, 2.843305e-06, 3.241588e-06, 3.7011e-06, 
    7.056434e-06, 7.24788e-06, 6.845105e-06, 8.257313e-06, 7.723395e-06,
  1.000982e-05, 8.427975e-06, 5.727845e-06, 7.508906e-06, 5.306768e-06, 
    1.842941e-06, 1.709501e-06, 3.203488e-07, 1.434774e-07, 2.047685e-06, 
    2.822727e-06, 3.748556e-06, 5.287379e-06, 5.667972e-06, 8.114493e-06,
  1.104479e-05, 7.04649e-06, 4.493905e-06, 3.020518e-06, 6.759248e-06, 
    1.65401e-06, 3.750157e-06, 1.543057e-06, 3.605566e-07, 1.25634e-06, 
    4.864144e-07, 2.742602e-06, 3.871457e-06, 5.039652e-06, 6.311993e-06,
  1.093062e-05, 8.398307e-06, 6.928082e-06, 5.200299e-06, 6.521812e-06, 
    4.692236e-06, 4.64361e-06, 2.211926e-06, 1.23179e-06, 1.781349e-08, 
    1.417791e-06, 3.457817e-06, 3.241681e-06, 5.239598e-06, 7.103973e-06,
  6.751357e-06, 1.069702e-05, 1.090507e-05, 9.113864e-06, 8.498972e-06, 
    7.581169e-06, 5.75727e-06, 3.272109e-06, 1.46695e-06, 3.442332e-08, 
    1.013427e-06, 1.470435e-06, 2.215912e-06, 6.405045e-06, 6.84877e-06,
  1.021751e-05, 1.495323e-05, 1.170858e-05, 1.375076e-05, 1.126294e-05, 
    1.05872e-05, 5.662067e-06, 3.923054e-06, 1.596019e-06, 1.837087e-07, 
    3.602055e-09, 1.512033e-06, 6.16524e-07, 5.867375e-06, 4.954608e-06,
  4.157797e-06, 1.19196e-05, 1.401986e-05, 1.371186e-05, 1.133297e-05, 
    8.199455e-06, 7.927211e-06, 4.343182e-06, 2.120241e-06, 3.746562e-07, 
    4.73097e-09, 1.225883e-06, 1.273033e-06, 2.699533e-06, 4.853145e-06,
  9.564458e-06, 6.308911e-06, 7.351325e-06, 1.070275e-05, 1.03892e-05, 
    6.456663e-06, 6.51353e-06, 1.946541e-06, 1.506561e-06, 6.841715e-08, 
    5.869035e-09, 4.279943e-10, 2.74813e-06, 2.470179e-06, 4.198954e-06,
  5.348496e-06, 5.090033e-06, 4.838294e-06, 2.366758e-06, 4.951038e-06, 
    4.25514e-06, 4.064796e-06, 1.100019e-06, 2.169767e-06, 2.621771e-06, 
    6.007108e-06, 8.481678e-06, 3.746466e-06, 7.24218e-06, 8.604569e-06,
  1.051289e-05, 5.563974e-06, 8.137845e-06, 4.142103e-06, 4.378871e-06, 
    3.577675e-06, 2.539784e-06, 3.513944e-06, 4.000024e-06, 1.183773e-06, 
    2.096536e-06, 8.498739e-06, 6.248256e-06, 5.937118e-06, 7.505515e-06,
  1.233235e-05, 1.004505e-05, 7.300558e-06, 5.205572e-06, 3.081366e-06, 
    5.733698e-06, 5.939772e-06, 8.285532e-06, 7.80854e-06, 3.523283e-06, 
    6.960033e-07, 1.652992e-06, 7.913916e-06, 8.675888e-06, 8.235416e-06,
  1.19391e-05, 1.02986e-05, 3.967647e-06, 1.699632e-06, 1.235257e-06, 
    4.308412e-06, 3.825127e-06, 2.252927e-06, 3.135596e-06, 9.465931e-06, 
    1.424207e-06, 9.553994e-07, 5.675235e-06, 1.30174e-05, 8.152165e-06,
  1.197477e-05, 1.033695e-05, 6.695282e-06, 2.030368e-06, 1.32089e-06, 
    1.30676e-06, 8.655287e-07, 3.569934e-06, 3.216913e-06, 8.037282e-06, 
    4.904181e-06, 6.779338e-07, 5.264672e-06, 8.343055e-06, 9.854803e-06,
  1.178082e-05, 1.0672e-05, 9.554051e-06, 5.682491e-06, 4.016859e-06, 
    2.125428e-06, 2.697093e-06, 4.812376e-06, 6.628204e-06, 1.186481e-05, 
    4.557876e-06, 1.480933e-06, 3.507211e-06, 7.234633e-06, 6.705563e-06,
  1.243364e-05, 1.22318e-05, 1.079663e-05, 9.647479e-06, 1.130584e-05, 
    7.462284e-06, 6.002459e-06, 6.657001e-06, 6.650754e-06, 8.521241e-06, 
    9.226478e-06, 8.180307e-07, 2.392676e-06, 3.319377e-06, 5.97977e-06,
  9.895735e-06, 9.901643e-06, 1.048426e-05, 1.042313e-05, 1.117844e-05, 
    1.185167e-05, 8.05431e-06, 7.389681e-06, 6.258121e-06, 5.347923e-06, 
    5.216849e-06, 1.330523e-06, 1.820651e-06, 3.703074e-06, 7.107342e-06,
  7.420746e-06, 9.877126e-06, 1.035247e-05, 1.074926e-05, 1.127259e-05, 
    1.274057e-05, 9.503884e-06, 6.754289e-06, 6.685814e-06, 6.88094e-06, 
    4.312019e-06, 2.998385e-06, 2.687269e-06, 3.868265e-06, 6.849639e-06,
  1.271665e-05, 1.143807e-05, 1.222632e-05, 1.410446e-05, 1.293194e-05, 
    1.313313e-05, 1.065237e-05, 8.965108e-06, 8.121735e-06, 8.808358e-06, 
    3.390553e-06, 3.075639e-06, 4.098635e-06, 5.899354e-06, 6.189233e-06,
  7.256323e-06, 9.843268e-06, 1.0948e-05, 1.346976e-05, 8.188105e-06, 
    4.611978e-06, 6.069692e-06, 9.441197e-06, 2.846811e-06, 4.423476e-07, 
    3.264105e-06, 5.47426e-06, 8.582416e-06, 6.12849e-06, 5.22259e-06,
  6.544522e-06, 9.892977e-06, 9.411993e-06, 1.578723e-05, 1.054865e-05, 
    5.00431e-06, 5.477588e-06, 6.750018e-06, 1.333395e-05, 2.907222e-06, 
    1.519638e-07, 2.383756e-06, 7.069326e-06, 9.752e-06, 6.895204e-06,
  8.041627e-06, 8.929883e-06, 1.185327e-05, 1.367912e-05, 1.6039e-05, 
    6.709811e-06, 6.346755e-06, 5.730183e-06, 8.7831e-06, 1.393773e-05, 
    2.751629e-07, 1.542595e-06, 5.283678e-06, 7.717347e-06, 1.056912e-05,
  9.124315e-06, 9.947245e-06, 9.684315e-06, 1.514157e-05, 1.623414e-05, 
    1.20134e-05, 9.35075e-06, 8.746857e-06, 9.513803e-06, 1.411294e-05, 
    4.305708e-07, 1.163754e-06, 4.311666e-06, 7.456511e-06, 1.595449e-05,
  1.030333e-05, 6.550821e-06, 1.302632e-05, 1.462446e-05, 1.704329e-05, 
    1.438096e-05, 1.084973e-05, 9.53231e-06, 1.198215e-05, 1.267881e-05, 
    2.708543e-07, 3.239705e-07, 5.152757e-06, 5.369724e-06, 1.017578e-05,
  1.053433e-05, 9.108193e-06, 1.075233e-05, 1.351333e-05, 1.729726e-05, 
    1.504067e-05, 1.168494e-05, 9.751081e-06, 1.241002e-05, 1.412905e-05, 
    3.882729e-07, 4.274996e-07, 6.364033e-06, 5.583492e-06, 9.971378e-06,
  9.634188e-06, 7.76203e-06, 1.086592e-05, 1.680655e-05, 1.925671e-05, 
    1.627998e-05, 1.221322e-05, 1.00605e-05, 1.141805e-05, 1.144421e-05, 
    9.349364e-07, 8.540665e-07, 8.954484e-06, 8.779832e-06, 1.112314e-05,
  7.176453e-06, 7.345071e-06, 1.073439e-05, 1.533118e-05, 1.750251e-05, 
    1.613172e-05, 1.328237e-05, 1.027218e-05, 6.002135e-06, 8.666413e-06, 
    2.755596e-06, 8.644222e-07, 9.188928e-06, 7.590622e-06, 9.743334e-06,
  5.349995e-06, 6.983205e-06, 1.009145e-05, 1.580606e-05, 1.677442e-05, 
    1.531669e-05, 1.237248e-05, 7.205361e-06, 4.79086e-06, 7.087589e-06, 
    2.300338e-06, 2.650608e-06, 5.757395e-06, 8.510332e-06, 8.753172e-06,
  5.544523e-06, 8.207414e-06, 1.131197e-05, 1.508899e-05, 1.678011e-05, 
    1.43483e-05, 1.11356e-05, 6.139011e-06, 6.959924e-06, 4.2206e-06, 
    4.179574e-06, 3.40842e-06, 4.576595e-06, 5.081029e-06, 7.031442e-06,
  9.309342e-06, 9.67875e-06, 6.806845e-06, 7.240924e-06, 7.163027e-06, 
    4.677863e-06, 4.562671e-06, 4.753251e-06, 4.168294e-06, 2.60942e-06, 
    4.293754e-06, 5.978933e-06, 9.29093e-06, 8.066029e-06, 7.661486e-06,
  2.438269e-06, 9.573794e-06, 8.151818e-06, 9.697963e-06, 7.710335e-06, 
    5.810147e-06, 4.241049e-06, 4.624384e-06, 4.726656e-06, 4.828953e-06, 
    4.913794e-06, 4.902277e-06, 8.894563e-06, 1.031086e-05, 9.638802e-06,
  2.039596e-06, 4.6705e-06, 1.100103e-05, 9.833785e-06, 8.546559e-06, 
    5.607465e-06, 5.387279e-06, 5.858937e-06, 4.525083e-06, 6.090397e-06, 
    4.387422e-06, 5.657161e-06, 6.911238e-06, 1.113948e-05, 1.005257e-05,
  1.872686e-06, 1.213378e-06, 5.065837e-06, 9.224548e-06, 8.327784e-06, 
    7.898336e-06, 6.911141e-06, 6.125562e-06, 5.372819e-06, 5.565846e-06, 
    3.803851e-06, 5.521105e-06, 5.070367e-06, 9.495865e-06, 1.013841e-05,
  1.108379e-06, 1.874023e-06, 9.254227e-07, 5.814696e-06, 9.19505e-06, 
    8.68298e-06, 7.726236e-06, 5.661861e-06, 5.508453e-06, 5.030422e-06, 
    4.121105e-06, 5.044791e-06, 5.572086e-06, 6.737864e-06, 9.152095e-06,
  7.803279e-07, 6.710802e-07, 8.558118e-07, 1.905706e-06, 5.041727e-06, 
    5.22418e-06, 5.860508e-06, 4.816968e-06, 5.708097e-06, 5.151932e-06, 
    4.585127e-06, 3.224329e-06, 5.295361e-06, 5.476688e-06, 8.95128e-06,
  1.014736e-06, 7.359753e-07, 9.741179e-07, 1.237969e-06, 2.974986e-06, 
    3.816281e-06, 5.27759e-06, 5.344629e-06, 4.553376e-06, 4.361939e-06, 
    6.550357e-06, 3.548889e-06, 4.657916e-06, 5.554973e-06, 9.339999e-06,
  2.028882e-06, 1.451136e-06, 5.524061e-07, 3.132938e-07, 1.725136e-06, 
    2.808884e-06, 2.734757e-06, 4.736651e-06, 5.12167e-06, 5.768658e-06, 
    7.750384e-06, 5.805904e-06, 5.085098e-06, 5.668016e-06, 6.864594e-06,
  7.325607e-07, 5.575437e-07, 2.321881e-07, 1.150447e-07, 9.499471e-07, 
    2.246724e-06, 2.721572e-06, 2.80599e-06, 3.947617e-06, 5.9878e-06, 
    8.029591e-06, 7.906691e-06, 6.467724e-06, 5.180716e-06, 6.764729e-06,
  3.52761e-07, 3.501741e-07, 3.290875e-08, 2.06316e-08, 7.608504e-07, 
    1.225275e-06, 1.0058e-06, 2.554672e-06, 2.850596e-06, 5.110107e-06, 
    5.188329e-06, 9.45339e-06, 7.275944e-06, 7.658361e-06, 6.894355e-06,
  2.270275e-08, 5.351343e-09, 7.942029e-10, 2.781204e-09, 8.485856e-10, 
    1.136151e-10, 1.713487e-08, 2.311101e-07, 7.895579e-07, 2.078652e-06, 
    3.500062e-06, 4.373226e-06, 1.030004e-05, 6.262002e-06, 7.404901e-06,
  7.218871e-08, 6.089067e-08, 5.081728e-09, 9.857751e-10, 9.222411e-10, 
    1.698739e-11, 4.045871e-10, 1.29319e-08, 9.812511e-08, 1.357311e-06, 
    1.866503e-06, 2.81937e-06, 9.588821e-06, 1.076889e-05, 9.142272e-06,
  2.226284e-08, 5.397733e-08, 1.328035e-07, 3.682436e-08, 1.684745e-09, 
    7.352584e-12, 2.445791e-10, 7.533682e-09, 1.772503e-07, 1.079375e-06, 
    6.7945e-07, 2.558074e-06, 5.967659e-06, 1.118443e-05, 8.781357e-06,
  7.789792e-09, 8.002986e-09, 1.715562e-08, 1.945284e-09, 1.97433e-09, 
    4.991774e-25, 2.08289e-12, 3.322228e-10, 7.169628e-08, 8.201478e-07, 
    2.235504e-06, 2.733246e-06, 4.239638e-06, 1.366404e-05, 9.85996e-06,
  5.439639e-09, 1.459815e-08, 2.957024e-08, 1.215627e-09, 7.79912e-11, 
    3.906192e-25, 1.150371e-12, 1.881818e-10, 9.187501e-09, 1.784346e-08, 
    2.367219e-06, 2.046776e-06, 3.56117e-06, 1.185973e-05, 1.300186e-05,
  1.628819e-10, 9.176611e-10, 6.306285e-08, 2.038839e-08, 1.306416e-11, 
    2.092701e-25, 2.27349e-25, 2.674143e-10, 9.549735e-09, 1.986351e-08, 
    2.807893e-06, 3.762706e-06, 3.586103e-06, 1.022363e-05, 1.163591e-05,
  5.788231e-10, 9.411723e-10, 3.823236e-08, 2.281378e-08, 1.503102e-11, 
    1.994632e-25, 5.933598e-12, 7.719965e-10, 7.087323e-09, 4.879157e-08, 
    5.75529e-06, 3.010534e-06, 1.558597e-06, 9.18333e-06, 1.199942e-05,
  3.158887e-08, 3.134291e-09, 8.702888e-09, 3.081556e-09, 1.070472e-11, 
    1.740754e-25, 7.030766e-12, 1.295905e-09, 1.826693e-08, 5.329022e-08, 
    5.066297e-06, 5.048156e-06, 3.473323e-06, 7.273002e-06, 7.452916e-06,
  1.31719e-07, 1.436736e-08, 2.13198e-10, 2.179938e-11, 1.057842e-17, 
    6.357661e-13, 1.836398e-10, 1.720915e-08, 7.196474e-08, 2.028906e-07, 
    3.678223e-06, 1.157921e-05, 8.77774e-06, 4.228089e-06, 1.092112e-05,
  1.476833e-08, 4.55228e-09, 1.482578e-08, 3.615107e-09, 1.258294e-08, 
    2.832305e-08, 2.178963e-08, 3.2156e-07, 6.478718e-07, 3.261037e-07, 
    3.177411e-06, 1.546409e-05, 1.840166e-05, 1.345088e-05, 1.633484e-05,
  1.292929e-09, 1.205742e-10, 4.416097e-10, 3.553337e-09, 1.970567e-07, 
    4.716876e-06, 6.827708e-06, 1.200064e-05, 9.6431e-06, 6.903082e-06, 
    6.111889e-06, 2.06614e-05, 1.273027e-05, 8.006278e-06, 5.873524e-06,
  3.362127e-08, 5.075365e-09, 1.505008e-08, 3.783215e-10, 3.175795e-09, 
    8.494766e-08, 1.84992e-06, 9.39288e-06, 1.552575e-05, 1.598657e-05, 
    8.374375e-06, 1.892129e-05, 2.395992e-05, 1.11329e-05, 7.360144e-06,
  5.637156e-09, 7.769992e-09, 1.435287e-09, 2.659241e-10, 7.79531e-11, 
    8.273094e-09, 2.954071e-07, 6.19657e-06, 8.736929e-06, 1.039455e-05, 
    1.508279e-05, 2.601968e-06, 1.33356e-05, 2.030318e-05, 1.267951e-05,
  2.965342e-09, 7.601883e-08, 1.40863e-08, 2.201011e-08, 2.900058e-10, 
    1.548935e-09, 5.374657e-08, 3.345835e-06, 7.556598e-06, 1.005041e-05, 
    2.36648e-05, 1.044718e-05, 3.881221e-06, 1.659737e-05, 2.007473e-05,
  4.569635e-08, 1.419199e-07, 2.246406e-07, 1.777604e-07, 1.010993e-08, 
    4.983227e-09, 3.121106e-09, 7.722217e-07, 6.248789e-06, 8.651785e-06, 
    2.532246e-05, 2.622937e-05, 1.000176e-05, 4.043085e-06, 2.195965e-05,
  5.365943e-07, 4.93305e-07, 3.705682e-07, 2.412457e-07, 1.615916e-07, 
    2.071719e-10, 5.684863e-10, 2.000225e-07, 4.18848e-06, 6.255004e-06, 
    1.083947e-05, 3.3721e-05, 1.604108e-05, 6.75769e-06, 1.515332e-05,
  1.732851e-06, 1.167593e-06, 6.42286e-07, 3.388603e-07, 1.244945e-07, 
    1.750465e-09, 6.211478e-11, 4.662683e-07, 3.120672e-06, 4.713886e-06, 
    9.169344e-06, 2.871817e-05, 3.057144e-05, 1.296436e-05, 1.216128e-05,
  2.472877e-06, 2.025841e-06, 1.53181e-06, 1.53118e-06, 5.713546e-07, 
    6.383964e-08, 2.274005e-10, 1.153274e-07, 9.577773e-07, 2.186388e-06, 
    5.387692e-06, 1.398974e-05, 4.075853e-05, 2.51536e-05, 9.114399e-06,
  2.366007e-06, 2.923083e-06, 2.525887e-06, 2.795039e-06, 6.202882e-07, 
    1.586879e-08, 5.014976e-10, 1.42888e-07, 2.710765e-07, 8.096952e-07, 
    1.707647e-06, 5.692483e-06, 2.182823e-05, 3.230836e-05, 1.181116e-05,
  3.816271e-06, 3.375429e-06, 2.366311e-06, 1.692628e-06, 3.622497e-07, 
    1.827759e-07, 9.132127e-08, 4.202627e-08, 6.38815e-07, 2.492875e-07, 
    2.16449e-07, 8.604104e-07, 6.348665e-06, 4.074786e-05, 2.656899e-05,
  4.841928e-06, 6.668352e-06, 6.572871e-06, 3.549768e-06, 4.680621e-06, 
    4.710366e-06, 5.642549e-06, 6.370028e-06, 1.107407e-05, 7.261581e-06, 
    5.580977e-06, 1.006135e-05, 4.563864e-06, 6.449177e-06, 8.689492e-06,
  2.50756e-06, 7.041866e-06, 1.082958e-05, 7.849908e-06, 3.41876e-06, 
    2.480796e-06, 4.584499e-06, 5.082586e-06, 6.492242e-06, 1.577918e-05, 
    9.456618e-06, 4.01575e-06, 6.990805e-06, 5.073124e-06, 8.289709e-06,
  4.114345e-06, 7.004796e-06, 6.405432e-06, 7.483959e-06, 5.874793e-06, 
    3.339677e-06, 2.863939e-06, 4.768206e-06, 5.753433e-06, 9.181033e-06, 
    1.718679e-05, 5.853153e-06, 6.097403e-06, 6.896454e-06, 1.37987e-05,
  6.130735e-06, 7.104377e-06, 7.520917e-06, 7.936194e-06, 8.697895e-06, 
    4.164561e-06, 3.104045e-06, 3.376651e-06, 4.469161e-06, 7.920736e-06, 
    8.463599e-06, 9.872692e-06, 5.881254e-06, 7.037089e-06, 5.395147e-06,
  8.729371e-06, 5.096575e-06, 6.067066e-06, 8.848515e-06, 1.105396e-05, 
    7.946949e-06, 2.366808e-06, 2.367038e-06, 4.64349e-06, 2.984623e-06, 
    1.055686e-05, 1.318513e-05, 7.924628e-06, 6.848735e-06, 5.340735e-06,
  5.19584e-06, 4.651093e-06, 4.533651e-06, 8.959583e-06, 9.750535e-06, 
    1.106136e-05, 3.08841e-06, 3.092922e-06, 4.024789e-06, 3.610798e-06, 
    9.137509e-06, 5.974646e-06, 1.02026e-05, 7.834632e-06, 7.727373e-06,
  3.912231e-06, 4.009127e-06, 3.632829e-06, 3.582527e-06, 9.997353e-06, 
    1.104411e-05, 8.228163e-06, 4.544857e-06, 3.08859e-06, 3.395775e-06, 
    3.893674e-06, 9.568318e-06, 1.294851e-05, 9.744393e-06, 1.07381e-05,
  7.308959e-06, 2.704901e-06, 2.939279e-06, 3.207184e-06, 5.383593e-06, 
    7.085054e-06, 1.251714e-05, 9.300259e-06, 3.608131e-06, 1.958916e-06, 
    3.22098e-06, 5.830236e-06, 1.197789e-05, 1.317587e-05, 1.596037e-05,
  5.175231e-06, 2.373601e-06, 1.859577e-06, 3.935798e-06, 5.115804e-06, 
    5.751077e-06, 9.274096e-06, 8.139579e-06, 4.414688e-06, 2.34633e-06, 
    3.033291e-06, 3.987968e-06, 5.487954e-06, 1.446786e-05, 1.569646e-05,
  4.820299e-06, 3.737544e-06, 2.274084e-06, 3.507864e-06, 4.277388e-06, 
    5.200254e-06, 4.406946e-06, 6.267219e-06, 5.544281e-06, 2.996042e-06, 
    3.821124e-06, 3.67301e-06, 2.115796e-06, 5.932013e-06, 1.287396e-05,
  7.404163e-06, 2.970299e-06, 8.923626e-07, 2.850723e-06, 4.179003e-06, 
    3.023782e-06, 6.172984e-06, 6.126108e-06, 7.667578e-06, 1.305476e-05, 
    7.558854e-06, 6.925705e-06, 1.024788e-05, 1.066541e-05, 1.109149e-05,
  7.930324e-06, 5.39752e-06, 3.671281e-07, 1.55777e-06, 3.720631e-06, 
    4.667167e-06, 8.185429e-06, 7.173069e-06, 6.753547e-06, 1.019629e-05, 
    9.342823e-06, 1.091035e-05, 9.019183e-06, 1.044905e-05, 1.130452e-05,
  8.758814e-06, 5.985304e-06, 4.074917e-07, 3.235988e-07, 7.047704e-07, 
    3.612839e-06, 7.862489e-06, 8.601256e-06, 6.766857e-06, 6.33307e-06, 
    1.044237e-05, 1.131609e-05, 9.919065e-06, 1.010495e-05, 1.013403e-05,
  8.316833e-06, 6.697351e-06, 2.677972e-07, 5.179314e-07, 6.197531e-07, 
    2.365243e-06, 8.119035e-06, 1.082482e-05, 8.379854e-06, 9.128186e-06, 
    7.718789e-06, 1.162713e-05, 1.093796e-05, 1.020636e-05, 1.07786e-05,
  7.610367e-06, 5.070107e-06, 1.538477e-07, 4.45201e-07, 1.294669e-06, 
    3.117111e-06, 8.048287e-06, 7.021876e-06, 6.916664e-06, 9.376823e-06, 
    8.239485e-06, 6.753859e-06, 1.032743e-05, 1.165957e-05, 1.164873e-05,
  5.470039e-06, 2.049259e-06, 2.983431e-07, 7.828967e-07, 2.102637e-06, 
    4.513005e-06, 9.055258e-06, 7.8978e-06, 7.900242e-06, 8.1143e-06, 
    9.431454e-06, 8.628914e-06, 9.420853e-06, 1.226213e-05, 1.275976e-05,
  1.324859e-06, 4.347591e-07, 2.506697e-07, 1.080349e-06, 3.241396e-06, 
    7.746629e-06, 1.157782e-05, 7.230887e-06, 9.236847e-06, 6.580985e-06, 
    9.547457e-06, 9.026614e-06, 9.79427e-06, 1.002069e-05, 1.213393e-05,
  1.700882e-07, 3.083392e-07, 1.132135e-06, 2.0875e-06, 4.443609e-06, 
    1.033707e-05, 6.880015e-06, 8.653759e-06, 8.266706e-06, 7.913212e-06, 
    6.641073e-06, 1.043339e-05, 9.687699e-06, 1.032032e-05, 1.219975e-05,
  1.856443e-07, 5.131496e-07, 1.242071e-06, 2.038086e-06, 4.589858e-06, 
    9.141881e-06, 3.247583e-06, 6.194101e-06, 6.266602e-06, 1.061835e-05, 
    9.504528e-06, 1.165235e-05, 1.069819e-05, 1.030866e-05, 1.292351e-05,
  3.018397e-07, 1.131936e-06, 1.89926e-06, 2.919236e-06, 5.102934e-06, 
    4.580848e-06, 4.066853e-06, 6.215749e-06, 6.461402e-06, 1.588054e-05, 
    1.161139e-05, 1.091685e-05, 1.188863e-05, 1.066038e-05, 1.113149e-05,
  4.154024e-06, 5.380044e-06, 7.427055e-07, 4.747355e-08, 2.337807e-07, 
    1.17788e-06, 1.867478e-06, 7.0093e-06, 9.974597e-06, 7.777361e-06, 
    4.996482e-06, 8.29304e-06, 9.460528e-06, 1.041354e-05, 9.726186e-06,
  3.024325e-06, 3.566943e-06, 7.498078e-07, 8.901608e-08, 4.959928e-08, 
    8.33364e-07, 5.698719e-07, 2.73538e-06, 6.217505e-06, 6.364587e-06, 
    5.532283e-06, 8.611408e-06, 9.512611e-06, 9.893373e-06, 9.981094e-06,
  2.019708e-06, 1.190005e-06, 2.849788e-06, 1.028559e-07, 7.220799e-09, 
    3.532939e-07, 4.534595e-07, 1.336766e-06, 4.352995e-06, 6.699053e-06, 
    6.277602e-06, 7.497256e-06, 7.724959e-06, 1.065336e-05, 1.026396e-05,
  1.995501e-06, 2.986922e-07, 1.342509e-06, 9.586816e-08, 5.237351e-09, 
    1.587784e-07, 4.751886e-07, 7.534469e-07, 3.212413e-06, 5.142583e-06, 
    6.548733e-06, 9.575453e-06, 1.043575e-05, 1.006813e-05, 1.018051e-05,
  2.336601e-06, 3.686033e-07, 1.900029e-07, 8.833753e-08, 7.771248e-09, 
    7.611757e-08, 2.052233e-07, 6.594352e-07, 3.508817e-06, 1.102781e-05, 
    6.578359e-06, 1.159082e-05, 1.665567e-05, 1.007335e-05, 1.049703e-05,
  3.635127e-06, 6.263337e-07, 7.680384e-08, 1.432072e-07, 1.018933e-08, 
    8.12886e-09, 2.217641e-07, 3.887862e-07, 1.326154e-06, 9.878696e-06, 
    7.659644e-06, 7.592137e-06, 1.121852e-05, 1.440892e-05, 9.913028e-06,
  3.723235e-06, 8.114761e-07, 6.236944e-08, 3.66201e-08, 2.090121e-09, 
    2.675876e-09, 1.065432e-07, 6.540487e-09, 2.972976e-07, 6.376751e-06, 
    6.063772e-06, 3.834145e-06, 4.900822e-06, 1.071933e-05, 1.113449e-05,
  2.085608e-06, 8.501848e-07, 1.003214e-07, 4.115441e-08, 3.957346e-09, 
    1.966766e-09, 1.756166e-08, 2.96484e-09, 7.218085e-08, 9.002035e-07, 
    1.210349e-06, 2.813714e-06, 5.199211e-06, 1.069417e-05, 1.084524e-05,
  2.916757e-06, 1.328802e-06, 3.027909e-07, 9.836945e-08, 1.007784e-08, 
    9.821856e-09, 1.70744e-08, 5.173324e-09, 8.34991e-08, 2.543412e-07, 
    8.934883e-07, 2.185183e-06, 1.34041e-05, 9.268193e-06, 1.04792e-05,
  3.183154e-06, 1.404973e-06, 3.271608e-07, 2.972911e-08, 1.340178e-08, 
    2.192315e-09, 5.596695e-08, 3.251008e-08, 4.767294e-08, 4.372149e-08, 
    8.308098e-07, 6.422315e-06, 2.059999e-05, 8.786567e-06, 9.513198e-06,
  5.975605e-06, 5.685813e-06, 4.410144e-06, 4.781058e-06, 3.58961e-06, 
    3.245595e-06, 3.767736e-06, 1.513954e-06, 4.756244e-07, 2.789939e-07, 
    2.276892e-06, 3.732206e-06, 9.923349e-06, 8.37775e-06, 7.94333e-06,
  5.679251e-06, 6.227119e-06, 3.982084e-06, 5.086762e-06, 5.596639e-06, 
    5.184326e-06, 4.421252e-06, 4.057399e-06, 1.80223e-06, 9.718675e-07, 
    1.267781e-06, 3.081883e-06, 1.001801e-05, 8.726641e-06, 7.616678e-06,
  4.547027e-06, 4.714834e-06, 6.867723e-06, 6.643011e-06, 6.336218e-06, 
    4.630109e-06, 5.826449e-06, 3.455793e-06, 2.82034e-06, 6.876476e-07, 
    5.506757e-07, 2.186345e-06, 7.240343e-06, 8.932754e-06, 8.069958e-06,
  5.759717e-06, 4.575634e-06, 7.168643e-06, 8.918852e-06, 6.7744e-06, 
    6.798043e-06, 5.391492e-06, 4.953168e-06, 3.705483e-06, 2.312532e-06, 
    1.666606e-06, 1.441117e-06, 2.309231e-06, 1.092454e-05, 8.734417e-06,
  4.951843e-06, 5.313094e-06, 7.511626e-06, 9.58388e-06, 7.980902e-06, 
    5.908263e-06, 7.690436e-06, 6.188332e-06, 2.916273e-06, 3.464919e-06, 
    1.321801e-06, 2.531793e-07, 1.66513e-06, 9.539436e-06, 1.002587e-05,
  3.04357e-06, 7.714782e-06, 7.989721e-06, 9.959806e-06, 9.512671e-06, 
    6.62218e-06, 8.504132e-06, 7.141321e-06, 3.265058e-06, 4.379373e-06, 
    1.892448e-06, 2.807355e-07, 1.43341e-06, 8.151185e-06, 1.150888e-05,
  3.009274e-06, 7.553048e-06, 5.95335e-06, 7.743986e-06, 9.074377e-06, 
    7.458648e-06, 7.285279e-06, 6.887581e-06, 4.477846e-06, 4.293409e-06, 
    1.433176e-06, 7.157631e-07, 1.662587e-06, 1.005426e-05, 1.062383e-05,
  4.12381e-06, 7.366422e-06, 6.322205e-06, 6.099519e-06, 7.869357e-06, 
    5.040044e-06, 6.913342e-06, 5.794851e-06, 4.384287e-06, 5.155451e-06, 
    1.936701e-06, 7.383822e-07, 2.064494e-06, 1.302694e-05, 8.778634e-06,
  4.549137e-06, 6.253862e-06, 5.991749e-06, 6.466148e-06, 5.839339e-06, 
    6.180027e-06, 6.262458e-06, 5.171913e-06, 4.010214e-06, 4.05734e-06, 
    2.428879e-06, 1.119166e-06, 9.344384e-07, 1.429798e-05, 1.04269e-05,
  2.065244e-06, 3.321684e-06, 4.158811e-06, 4.056842e-06, 4.62248e-06, 
    4.428406e-06, 5.579105e-06, 5.603996e-06, 5.277932e-06, 6.218203e-06, 
    2.366728e-06, 1.995212e-06, 3.363237e-07, 1.062792e-05, 1.201347e-05,
  7.918722e-06, 9.718881e-06, 7.173503e-06, 1.604031e-05, 1.535889e-05, 
    1.258816e-05, 1.129645e-05, 9.177862e-06, 9.147874e-06, 1.343122e-05, 
    1.230679e-05, 8.97024e-06, 8.280225e-06, 9.35682e-06, 1.061422e-05,
  7.361214e-06, 6.268573e-06, 5.250138e-06, 1.106082e-05, 1.644456e-05, 
    1.401214e-05, 1.340641e-05, 1.042011e-05, 1.203845e-05, 1.311258e-05, 
    1.23079e-05, 1.41703e-05, 7.610214e-06, 9.783572e-06, 1.12324e-05,
  5.254994e-06, 6.488733e-06, 3.861428e-06, 8.376552e-06, 1.485531e-05, 
    1.645069e-05, 1.620846e-05, 1.370328e-05, 1.087567e-05, 1.183082e-05, 
    1.28987e-05, 1.471181e-05, 9.49127e-06, 7.689211e-06, 1.047825e-05,
  6.689098e-06, 7.260606e-06, 3.631392e-06, 4.76117e-06, 1.017873e-05, 
    1.543624e-05, 1.503337e-05, 1.145912e-05, 1.00875e-05, 1.273706e-05, 
    1.388432e-05, 1.346935e-05, 1.000609e-05, 8.287716e-06, 9.40146e-06,
  6.247914e-06, 8.226569e-06, 1.891997e-06, 3.2424e-06, 7.938046e-06, 
    1.286446e-05, 1.621258e-05, 1.542717e-05, 1.346581e-05, 1.207524e-05, 
    1.231085e-05, 1.023568e-05, 1.217382e-05, 9.930593e-06, 9.215606e-06,
  6.160411e-06, 7.259386e-06, 9.358912e-07, 4.006293e-06, 7.061687e-06, 
    9.784713e-06, 1.202812e-05, 1.490249e-05, 1.462527e-05, 1.131463e-05, 
    1.012985e-05, 8.968811e-06, 1.352469e-05, 1.097137e-05, 9.575082e-06,
  6.955324e-06, 6.244113e-06, 6.183421e-07, 3.742553e-06, 5.432885e-06, 
    1.015969e-05, 1.311964e-05, 1.377002e-05, 1.753738e-05, 1.414223e-05, 
    1.004175e-05, 1.157701e-05, 1.151427e-05, 1.091573e-05, 9.759865e-06,
  6.899038e-06, 6.99425e-06, 1.24309e-06, 2.548141e-06, 4.607144e-06, 
    6.764785e-06, 9.969393e-06, 1.286726e-05, 1.500507e-05, 1.106257e-05, 
    1.184247e-05, 1.170827e-05, 1.150273e-05, 1.298965e-05, 9.238086e-06,
  4.904259e-06, 2.502993e-06, 2.222563e-06, 2.017399e-06, 3.822708e-06, 
    5.559902e-06, 8.205443e-06, 1.095984e-05, 1.44565e-05, 1.467947e-05, 
    1.165209e-05, 1.017762e-05, 9.813389e-06, 1.279417e-05, 9.587715e-06,
  2.236192e-06, 3.355018e-06, 2.822957e-06, 3.45936e-06, 2.811971e-06, 
    5.003452e-06, 6.243224e-06, 9.055624e-06, 1.188549e-05, 1.453725e-05, 
    1.601148e-05, 1.104698e-05, 1.008614e-05, 1.305618e-05, 1.186639e-05,
  1.145612e-05, 5.546342e-06, 9.774097e-06, 1.349917e-05, 1.516372e-05, 
    1.167967e-05, 9.402916e-06, 6.869493e-06, 7.681638e-06, 8.507155e-06, 
    9.48611e-06, 9.388939e-06, 1.075352e-05, 9.716839e-06, 9.96886e-06,
  1.587098e-05, 1.301327e-05, 8.550625e-06, 1.474709e-05, 1.521551e-05, 
    1.717703e-05, 1.40381e-05, 9.071347e-06, 8.797141e-06, 8.595286e-06, 
    8.159267e-06, 1.07091e-05, 1.00274e-05, 9.905289e-06, 9.589796e-06,
  6.836161e-06, 1.195953e-05, 6.769188e-06, 1.069105e-05, 1.745767e-05, 
    1.991488e-05, 1.723777e-05, 1.334859e-05, 6.573601e-06, 6.686797e-06, 
    7.250479e-06, 8.732454e-06, 8.863725e-06, 9.491671e-06, 9.22809e-06,
  5.732619e-06, 9.074658e-06, 1.192767e-05, 1.088637e-05, 1.142486e-05, 
    1.363358e-05, 1.484517e-05, 1.590842e-05, 1.058868e-05, 8.113563e-06, 
    8.463571e-06, 7.821394e-06, 8.784372e-06, 9.746288e-06, 9.6588e-06,
  6.824222e-06, 6.052531e-06, 7.741188e-06, 9.93978e-06, 1.301305e-05, 
    1.177071e-05, 1.475283e-05, 1.783549e-05, 1.690963e-05, 9.152801e-06, 
    8.828673e-06, 6.527548e-06, 7.047515e-06, 9.679334e-06, 1.004085e-05,
  6.136511e-06, 5.276108e-06, 5.864534e-06, 6.508314e-06, 1.265665e-05, 
    1.322055e-05, 1.524291e-05, 1.496836e-05, 1.612841e-05, 1.547028e-05, 
    1.014872e-05, 7.116766e-06, 8.37885e-06, 5.299215e-06, 8.928788e-06,
  3.598321e-06, 5.713714e-06, 4.180918e-06, 4.809584e-06, 4.780152e-06, 
    8.920712e-06, 1.46899e-05, 1.350028e-05, 1.449095e-05, 1.671464e-05, 
    9.977552e-06, 7.414761e-06, 6.70003e-06, 6.868216e-06, 5.389704e-06,
  3.284609e-06, 4.088204e-06, 6.053203e-06, 4.811776e-06, 5.683446e-06, 
    3.851327e-06, 5.914792e-06, 1.411632e-05, 1.515024e-05, 1.514041e-05, 
    1.475063e-05, 7.50442e-06, 4.480296e-06, 5.649198e-06, 4.807689e-06,
  3.548574e-06, 3.771327e-06, 4.786139e-06, 5.479546e-06, 5.304987e-06, 
    6.40738e-06, 4.997103e-06, 6.653393e-06, 1.456515e-05, 1.716026e-05, 
    1.779099e-05, 8.539317e-06, 8.514085e-06, 5.837524e-06, 5.921667e-06,
  3.598193e-06, 4.750336e-06, 4.367953e-06, 4.649608e-06, 4.967681e-06, 
    5.466275e-06, 7.230012e-06, 3.806161e-06, 6.221778e-06, 1.049899e-05, 
    1.58635e-05, 1.375961e-05, 1.176503e-05, 8.379767e-06, 6.905742e-06,
  5.366362e-06, 4.393495e-06, 5.408499e-06, 6.328398e-06, 7.040715e-06, 
    7.35074e-06, 5.254262e-06, 6.007492e-06, 6.896645e-06, 6.790468e-06, 
    8.298763e-06, 8.602195e-06, 7.761412e-06, 8.512378e-06, 8.216321e-06,
  4.973517e-06, 4.933191e-06, 5.587944e-06, 6.378739e-06, 7.685035e-06, 
    7.403367e-06, 6.144361e-06, 5.782637e-06, 6.461412e-06, 6.844779e-06, 
    7.109245e-06, 7.64767e-06, 8.465066e-06, 8.579304e-06, 8.514329e-06,
  5.966403e-06, 5.411537e-06, 5.010557e-06, 5.634292e-06, 7.380845e-06, 
    6.874086e-06, 5.997945e-06, 7.000639e-06, 6.168405e-06, 6.85639e-06, 
    6.819138e-06, 7.853748e-06, 7.054727e-06, 7.594643e-06, 9.537131e-06,
  5.32137e-06, 5.098776e-06, 6.288697e-06, 6.54593e-06, 8.250986e-06, 
    7.700296e-06, 8.085893e-06, 7.859976e-06, 8.025238e-06, 7.679334e-06, 
    7.830842e-06, 7.519089e-06, 6.125352e-06, 7.445144e-06, 1.222206e-05,
  6.200599e-06, 3.872025e-06, 6.750019e-06, 5.308749e-06, 8.110556e-06, 
    8.208603e-06, 9.368027e-06, 8.69564e-06, 8.019211e-06, 7.756448e-06, 
    6.848671e-06, 8.409673e-06, 6.876424e-06, 7.112688e-06, 1.572459e-05,
  5.058141e-06, 5.201539e-06, 6.222438e-06, 6.417567e-06, 8.506936e-06, 
    5.202828e-06, 7.165427e-06, 8.751379e-06, 1.114033e-05, 1.216153e-05, 
    7.828072e-06, 7.592294e-06, 8.30235e-06, 6.901296e-06, 1.820827e-05,
  6.497665e-06, 5.65621e-06, 7.582943e-06, 5.716536e-06, 7.267946e-06, 
    7.779186e-06, 6.655023e-06, 8.947331e-06, 9.764827e-06, 1.782661e-05, 
    1.263942e-05, 7.710725e-06, 8.227827e-06, 6.476475e-06, 5.681648e-06,
  9.46095e-06, 5.763892e-06, 6.381018e-06, 4.249034e-06, 7.462565e-06, 
    6.954786e-06, 6.489959e-06, 8.88838e-06, 5.980041e-06, 6.128331e-06, 
    1.533787e-05, 1.237124e-05, 1.190058e-05, 8.626113e-06, 9.603065e-06,
  1.071569e-05, 9.548309e-06, 8.84979e-06, 8.071297e-06, 4.690701e-06, 
    6.536266e-06, 5.043422e-06, 5.585e-06, 7.827484e-06, 6.85314e-06, 
    5.690482e-06, 1.020841e-05, 2.01837e-05, 1.761695e-05, 1.066613e-05,
  1.082557e-05, 9.70419e-06, 1.372014e-05, 1.476049e-05, 8.778264e-06, 
    6.905883e-06, 6.45977e-06, 3.741807e-06, 7.560639e-06, 6.209111e-06, 
    5.686206e-06, 7.5838e-06, 6.481911e-06, 2.306245e-05, 2.015016e-05,
  4.179092e-06, 3.58496e-06, 4.358505e-06, 6.644583e-06, 7.325531e-06, 
    5.233069e-06, 7.211323e-06, 6.20563e-06, 8.001343e-06, 8.73709e-06, 
    8.193964e-06, 9.504953e-06, 1.211341e-05, 1.015968e-05, 1.089802e-05,
  3.910277e-06, 3.695437e-06, 5.670163e-06, 5.776561e-06, 6.989811e-06, 
    5.79901e-06, 5.681064e-06, 7.582348e-06, 8.398127e-06, 7.061203e-06, 
    9.862408e-06, 1.103832e-05, 9.253999e-06, 1.337591e-05, 1.188464e-05,
  4.502539e-06, 3.218706e-06, 3.900607e-06, 3.475185e-06, 6.337995e-06, 
    6.453099e-06, 4.582083e-06, 6.00352e-06, 5.817346e-06, 7.649322e-06, 
    8.809485e-06, 8.935e-06, 8.446367e-06, 1.08398e-05, 1.331651e-05,
  7.782525e-06, 3.049082e-06, 2.034116e-06, 3.333535e-06, 5.789119e-06, 
    8.328017e-06, 8.370302e-06, 6.483703e-06, 7.10585e-06, 8.041489e-06, 
    7.991292e-06, 6.445099e-06, 8.957055e-06, 1.20589e-05, 1.322506e-05,
  5.275218e-06, 6.259283e-06, 3.363721e-06, 4.435765e-06, 6.738539e-06, 
    1.016617e-05, 1.032456e-05, 1.012737e-05, 7.14169e-06, 5.326417e-06, 
    7.549894e-06, 8.242869e-06, 8.816302e-06, 1.343556e-05, 1.407807e-05,
  4.062603e-06, 4.081013e-06, 4.35862e-06, 6.492335e-06, 8.414728e-06, 
    9.14757e-06, 8.65554e-06, 1.537282e-05, 5.420465e-06, 5.592557e-06, 
    7.06197e-06, 1.114782e-05, 1.454987e-05, 6.333434e-06, 1.657584e-05,
  3.345506e-06, 2.778172e-06, 1.868507e-06, 4.521987e-06, 7.006668e-06, 
    1.028456e-05, 1.337805e-05, 7.380964e-06, 7.186527e-06, 6.974944e-06, 
    5.888605e-06, 1.069232e-05, 1.724511e-05, 1.862913e-05, 1.782724e-05,
  3.599641e-06, 4.232334e-06, 3.345699e-06, 4.768334e-06, 6.354566e-06, 
    8.176747e-06, 8.936962e-06, 7.997098e-06, 1.420126e-05, 1.425443e-05, 
    7.165108e-06, 1.208454e-05, 1.527658e-05, 1.553748e-05, 2.353277e-05,
  4.438461e-06, 4.783891e-06, 5.948363e-06, 6.193755e-06, 4.293814e-06, 
    5.132338e-06, 4.771921e-06, 9.836793e-06, 1.172709e-05, 1.282992e-05, 
    1.406195e-05, 1.413945e-05, 1.328394e-05, 2.559421e-05, 2.227368e-05,
  7.281048e-06, 7.481668e-06, 6.650036e-06, 1.534237e-05, 5.354164e-06, 
    6.070293e-06, 5.225167e-06, 3.213438e-06, 6.252503e-06, 7.668956e-06, 
    9.941467e-06, 1.580957e-05, 1.262502e-05, 1.140484e-05, 1.692233e-05 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
