netcdf atmos_daily.00010101-00010701.pr.tile3 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pr(time, grid_yt, grid_xt) ;
		pr:_FillValue = 1.e+20f ;
		pr:missing_value = 1.e+20f ;
		pr:units = "kg m-2 s-1" ;
		pr:long_name = "Precipitation" ;
		pr:cell_methods = "time: mean" ;
		pr:cell_measures = "area: area" ;
		pr:time_avg_info = "average_T1,average_T2,average_DT" ;
		pr:standard_name = "precipitation_flux" ;
		pr:interp_method = "conserve_order1" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:00 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile3.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile3.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.0008770345, 0.4596241, 0.9892928, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.01035247, 0.004304647, 0.6546783, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.8534847, 0.8118016, 0.9951549, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9894952, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4452189, 0.3028796, 0.7140614, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9903189, 0.3150955, 0.0007410151, 0, 0.02645395, 
    0.9012984, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.681631, 0, 0, 0, 0.004980796, 0.7708192, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5536854, 0, 0, 0, 0.004666397, 0.9395298, 1,
  1, 1, 1, 1, 1, 1, 1, 0.9995009, 0.3626226, 0, 0, 0, 0, 0.8367797, 1,
  1, 1, 1, 1, 1, 0.8451425, 0.7016711, 0.3953246, 0, 0, 0, 0, 0.006316811, 
    0.8673657, 1 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pr =
  1.66021e-10, 1.42997e-09, 1.327988e-08, 3.989395e-08, 1.575848e-07, 
    4.657797e-07, 4.610174e-07, 1.387621e-07, 9.510071e-08, 3.266056e-07, 
    1.735931e-09, 5.40166e-10, 3.325655e-10, 5.679277e-11, 2.007392e-11,
  2.04674e-10, 3.151667e-09, 3.775034e-09, 1.019665e-08, 8.123922e-08, 
    2.415199e-07, 1.60483e-07, 2.412571e-08, 2.180288e-09, 7.433865e-10, 
    6.144271e-10, 6.763583e-10, 2.37619e-11, 9.076426e-11, 1.217465e-09,
  1.361956e-09, 1.793585e-09, 1.038679e-09, 2.205657e-09, 3.963862e-09, 
    6.982167e-08, 2.638548e-08, 4.059408e-09, 2.189206e-10, 4.332609e-09, 
    6.933538e-09, 4.381168e-09, 7.612032e-10, 5.943356e-09, 5.304796e-09,
  1.046716e-08, 5.72574e-09, 8.641879e-09, 3.868204e-08, 1.231656e-08, 
    7.940228e-09, 6.551531e-09, 3.049356e-08, 4.902777e-10, 1.002119e-08, 
    2.305938e-08, 2.156453e-08, 6.265333e-09, 3.484289e-08, 8.10105e-08,
  2.358808e-07, 4.435491e-08, 6.429575e-09, 4.938261e-08, 3.056677e-08, 
    1.117067e-08, 1.677122e-08, 6.096855e-09, 7.333566e-09, 4.223911e-09, 
    4.337366e-09, 6.675765e-09, 2.329678e-09, 3.057889e-09, 1.542222e-06,
  1.41698e-05, 3.868995e-06, 1.108495e-07, 1.0504e-08, 3.78585e-08, 
    3.63505e-08, 1.960907e-08, 4.641018e-09, 8.209579e-10, 1.093058e-10, 
    1.456677e-09, 5.414612e-09, 1.810268e-08, 1.539902e-07, 1.17162e-05,
  5.48099e-06, 3.429445e-06, 8.251172e-07, 1.450621e-07, 7.895087e-08, 
    4.104816e-08, 8.153823e-09, 3.359003e-09, 1.037313e-09, 7.92648e-11, 
    5.514067e-09, 2.830008e-09, 1.024376e-08, 2.19294e-05, 6.930329e-06,
  3.661083e-06, 3.821117e-06, 1.547147e-06, 4.264546e-07, 9.910512e-08, 
    7.958521e-07, 2.24587e-08, 6.806661e-09, 2.001016e-10, 7.896336e-11, 
    1.34325e-09, 5.788486e-09, 1.907837e-08, 4.224302e-05, 4.159398e-06,
  2.682192e-06, 7.187205e-06, 2.282978e-06, 8.91991e-08, 1.885093e-07, 
    9.871701e-07, 1.058039e-07, 9.782869e-10, 1.316461e-09, 4.857685e-09, 
    8.070518e-09, 6.038048e-08, 6.499948e-08, 1.409407e-05, 1.538428e-06,
  3.255736e-06, 1.490688e-05, 3.062733e-06, 1.874302e-08, 8.604603e-09, 
    8.065189e-09, 8.852583e-09, 2.081551e-09, 1.865696e-08, 4.107099e-08, 
    1.321195e-07, 1.132321e-06, 5.367535e-06, 2.131857e-05, 2.589612e-05,
  1.554111e-10, 4.53467e-10, 5.597391e-10, 5.245566e-10, 2.135177e-10, 
    7.926407e-11, 6.975558e-11, 6.625543e-10, 1.448484e-09, 1.866117e-09, 
    4.58083e-10, 3.110069e-10, 7.798622e-10, 6.09528e-10, 1.294533e-09,
  3.616579e-09, 2.65588e-09, 4.688295e-10, 6.186344e-10, 3.117502e-09, 
    2.216963e-09, 8.805564e-10, 1.178821e-09, 9.056877e-09, 4.206245e-09, 
    8.777338e-10, 4.997133e-10, 1.208569e-09, 6.589546e-10, 2.681154e-10,
  1.695033e-07, 1.852294e-08, 3.064816e-09, 2.859035e-09, 9.913657e-09, 
    1.056163e-08, 4.047562e-09, 4.154701e-09, 1.788841e-08, 6.411108e-09, 
    1.839374e-09, 1.367727e-09, 1.785429e-09, 1.278723e-09, 1.304809e-10,
  1.121495e-07, 1.000984e-07, 7.439459e-08, 1.068986e-07, 7.245065e-08, 
    7.567135e-08, 4.48535e-08, 3.485136e-08, 4.175669e-08, 1.299347e-08, 
    8.526382e-09, 6.952593e-09, 4.301842e-09, 3.472752e-09, 5.857499e-09,
  6.972718e-08, 9.933291e-08, 8.266563e-08, 1.89278e-07, 2.118673e-07, 
    2.093447e-07, 1.330151e-07, 6.442878e-08, 4.058096e-08, 9.770349e-09, 
    2.947096e-09, 1.47973e-09, 1.553252e-09, 1.680778e-09, 1.109373e-07,
  9.814681e-07, 3.575404e-07, 4.657617e-08, 3.342017e-08, 1.145776e-07, 
    2.004561e-07, 1.842923e-07, 6.809712e-08, 3.364655e-08, 1.258858e-08, 
    4.220244e-09, 2.748803e-09, 1.695096e-09, 2.309102e-10, 1.802584e-07,
  3.056912e-06, 4.687928e-07, 3.528928e-08, 1.174668e-08, 3.980411e-08, 
    1.178355e-07, 2.879429e-07, 9.983839e-08, 1.523843e-08, 7.184678e-09, 
    3.959953e-09, 3.098784e-09, 3.535648e-09, 1.71238e-07, 2.322529e-07,
  4.397198e-07, 3.071487e-08, 4.14144e-09, 5.668821e-09, 1.33123e-08, 
    2.95639e-08, 3.681419e-08, 1.708668e-07, 1.612507e-08, 4.227432e-09, 
    2.408714e-09, 3.256465e-09, 4.277649e-09, 2.445575e-06, 3.272151e-08,
  1.062995e-09, 2.360324e-09, 1.065336e-09, 2.946555e-09, 3.569868e-09, 
    9.571531e-08, 5.080347e-09, 2.273744e-09, 1.066382e-09, 3.373569e-09, 
    3.047573e-09, 9.582367e-09, 5.991229e-08, 2.236075e-06, 4.815856e-08,
  5.958752e-08, 4.182712e-09, 6.864647e-10, 9.013066e-10, 2.390542e-09, 
    2.019156e-09, 1.458626e-09, 9.428253e-10, 1.728687e-09, 3.820825e-09, 
    6.618687e-09, 6.328305e-09, 1.020658e-06, 6.948925e-06, 5.093007e-06,
  9.753556e-10, 1.763498e-09, 6.777747e-09, 1.211269e-08, 4.90411e-09, 
    1.57027e-08, 7.257756e-08, 7.021084e-08, 8.23182e-08, 1.834948e-07, 
    9.077469e-08, 3.778096e-08, 7.332183e-09, 5.117926e-09, 5.213824e-09,
  1.497255e-09, 4.920103e-09, 8.125559e-09, 8.084734e-09, 7.238189e-08, 
    7.988614e-08, 1.373147e-07, 1.481631e-07, 3.49941e-07, 2.717976e-07, 
    1.240861e-07, 3.833157e-08, 1.054946e-08, 9.483837e-09, 9.727249e-09,
  2.425643e-08, 4.165705e-08, 2.769907e-08, 5.154407e-08, 1.646968e-07, 
    1.300322e-07, 1.962251e-07, 2.792085e-07, 5.751127e-07, 2.475182e-07, 
    1.103922e-07, 9.039894e-08, 4.041221e-08, 1.659711e-08, 2.026247e-08,
  3.955023e-07, 5.688604e-08, 2.656595e-07, 5.154283e-07, 2.864993e-07, 
    2.044227e-07, 1.903214e-07, 2.935766e-07, 4.126681e-07, 2.622972e-07, 
    1.71449e-07, 8.522924e-08, 7.034315e-08, 3.943856e-08, 3.939727e-08,
  1.935203e-07, 3.72127e-08, 4.129383e-08, 5.170944e-08, 6.509711e-08, 
    9.23586e-08, 9.953955e-08, 1.529013e-07, 1.804799e-07, 1.087622e-07, 
    6.933234e-08, 4.835881e-08, 4.282811e-08, 4.73268e-08, 8.002178e-08,
  4.20822e-06, 7.454668e-07, 3.387304e-08, 9.721839e-08, 1.495425e-07, 
    5.069192e-08, 6.118214e-08, 8.538475e-08, 1.031571e-07, 1.018016e-07, 
    7.165336e-08, 3.763577e-08, 4.449095e-08, 5.930662e-08, 2.076031e-07,
  4.097274e-06, 8.186111e-07, 7.352214e-07, 6.804479e-07, 2.764056e-07, 
    4.316092e-08, 2.345729e-08, 2.909007e-08, 4.738664e-08, 4.090094e-08, 
    3.611959e-08, 2.363737e-08, 4.551316e-08, 1.162496e-07, 1.097686e-07,
  2.492451e-07, 6.958366e-08, 3.232065e-07, 1.050693e-07, 4.713119e-07, 
    8.957944e-07, 1.105319e-07, 7.092102e-09, 6.683091e-09, 7.353838e-09, 
    7.55781e-09, 1.018178e-08, 2.803064e-08, 2.578181e-07, 2.404466e-08,
  1.055461e-07, 6.795169e-08, 1.97179e-08, 2.841211e-08, 5.228756e-07, 
    4.507259e-06, 5.916081e-07, 2.684593e-09, 2.341893e-09, 2.331294e-09, 
    2.30764e-09, 3.22027e-09, 1.512581e-08, 2.142444e-08, 1.602881e-08,
  3.91858e-05, 2.744112e-05, 8.476393e-06, 1.19299e-07, 1.446872e-07, 
    6.239669e-08, 7.464015e-08, 2.285744e-09, 7.116742e-08, 7.334501e-08, 
    5.405429e-09, 4.857669e-09, 5.99942e-09, 1.126917e-08, 1.439433e-08,
  1.527111e-09, 1.542703e-09, 1.778468e-09, 6.506418e-10, 9.986127e-10, 
    4.177417e-09, 3.527331e-08, 1.076766e-07, 2.071859e-06, 1.502517e-06, 
    7.325965e-07, 6.768795e-07, 5.063827e-07, 1.954466e-07, 8.175626e-09,
  1.54576e-08, 4.128559e-09, 3.504613e-09, 4.01883e-08, 2.061827e-08, 
    5.194506e-06, 8.939559e-06, 6.714132e-06, 7.421615e-06, 2.775746e-06, 
    1.078055e-06, 7.092942e-07, 5.757631e-07, 3.821123e-07, 4.933538e-09,
  5.005903e-06, 4.391849e-06, 1.959284e-08, 4.365889e-09, 1.366e-05, 
    1.320352e-05, 1.16026e-05, 1.519898e-05, 1.71692e-05, 8.073293e-06, 
    2.694759e-06, 1.008414e-06, 4.120584e-07, 2.684571e-07, 4.903364e-09,
  2.692939e-05, 1.289693e-05, 2.347477e-06, 1.573995e-05, 2.449797e-05, 
    2.792287e-05, 2.49864e-05, 2.121455e-05, 1.63631e-05, 7.916853e-06, 
    7.094201e-06, 3.7282e-06, 9.023216e-07, 1.17972e-07, 1.179374e-08,
  3.955452e-05, 1.545109e-05, 7.099379e-07, 2.041374e-06, 2.28002e-05, 
    4.371388e-05, 4.16174e-05, 2.493372e-05, 1.130135e-05, 1.157158e-05, 
    2.259463e-08, 1.266484e-08, 9.307147e-09, 1.134316e-08, 2.151501e-07,
  4.739345e-05, 1.687907e-05, 2.778316e-06, 1.973605e-07, 7.729075e-06, 
    2.746863e-05, 4.231461e-05, 9.782497e-06, 6.295476e-08, 1.773695e-07, 
    2.119507e-06, 2.098064e-06, 2.207706e-08, 1.936682e-08, 2.156208e-06,
  5.582917e-05, 4.779119e-05, 2.912123e-05, 2.816551e-05, 4.676861e-05, 
    8.648535e-05, 9.128186e-05, 6.943988e-06, 2.662454e-06, 1.017175e-05, 
    1.921293e-05, 1.004452e-05, 4.067542e-07, 2.939267e-06, 2.857945e-06,
  4.402061e-05, 7.324159e-05, 5.895355e-05, 5.210662e-05, 0.0001014075, 
    0.0001705605, 0.0001240624, 2.940296e-05, 1.307483e-05, 8.047231e-06, 
    1.833703e-05, 2.296943e-05, 1.877018e-06, 3.747318e-05, 1.306059e-06,
  7.909923e-05, 0.000128062, 8.538599e-05, 5.956387e-05, 0.0001186587, 
    0.0001625919, 0.0001027768, 3.338283e-05, 6.274228e-06, 7.040936e-06, 
    1.02032e-05, 3.666545e-05, 2.30639e-05, 2.418904e-05, 4.877753e-07,
  8.090132e-05, 0.0001321072, 0.0001136217, 5.994216e-05, 0.0001168695, 
    0.0001360861, 0.000119799, 4.145408e-05, 3.88417e-05, 2.527538e-05, 
    8.403139e-06, 4.971779e-06, 1.547563e-05, 2.230108e-05, 1.904208e-06,
  6.553607e-07, 3.50951e-06, 2.890472e-07, 1.203989e-06, 1.454522e-07, 
    2.631325e-07, 4.618714e-06, 6.040244e-06, 1.469487e-05, 8.342593e-06, 
    5.352597e-06, 9.734068e-06, 1.509629e-05, 7.852615e-06, 1.881826e-09,
  4.420242e-07, 1.850761e-06, 2.486454e-06, 4.000174e-06, 2.946065e-06, 
    6.170803e-06, 1.234123e-05, 1.758653e-05, 1.428918e-05, 5.237488e-06, 
    2.010192e-06, 5.831859e-06, 1.041105e-05, 5.586558e-06, 2.242629e-09,
  3.913465e-05, 4.661302e-05, 2.514423e-06, 7.992176e-06, 3.311324e-05, 
    2.292439e-05, 1.847607e-05, 2.832953e-05, 2.519328e-05, 7.741911e-06, 
    4.649271e-06, 3.434716e-06, 3.769809e-06, 2.502149e-06, 2.666461e-09,
  0.0001285492, 4.019061e-05, 1.614597e-05, 3.049706e-05, 2.192278e-05, 
    1.891055e-05, 2.941491e-05, 4.613051e-05, 2.483631e-05, 9.568934e-06, 
    1.425326e-05, 1.186638e-05, 4.202367e-06, 1.088153e-06, 2.347456e-07,
  7.510296e-05, 3.233566e-05, 7.533206e-06, 7.962667e-06, 1.303732e-05, 
    1.761876e-05, 3.509572e-05, 4.484262e-05, 2.961801e-05, 2.200332e-05, 
    1.471353e-07, 3.355725e-08, 1.71456e-06, 3.691162e-07, 3.614125e-07,
  2.218928e-05, 2.920038e-05, 1.391702e-05, 1.376161e-05, 1.834085e-05, 
    2.250523e-05, 2.538981e-05, 2.28762e-05, 8.81811e-06, 1.407023e-06, 
    4.549593e-06, 1.117984e-05, 1.197659e-07, 4.752752e-07, 1.804616e-05,
  1.015668e-05, 9.389236e-06, 6.504125e-06, 1.504314e-05, 1.97154e-05, 
    1.98711e-05, 1.942754e-05, 1.608308e-06, 5.962528e-07, 1.152993e-06, 
    6.050604e-06, 1.957277e-05, 4.774256e-06, 4.966614e-05, 2.054971e-05,
  3.265182e-05, 3.598744e-05, 1.080484e-05, 6.618214e-06, 1.868241e-05, 
    2.500646e-05, 1.330047e-05, 5.162227e-06, 3.044139e-06, 2.040318e-06, 
    3.483354e-06, 2.180734e-05, 1.891236e-05, 0.0001180913, 9.234515e-06,
  6.693284e-05, 8.543689e-05, 4.773029e-05, 3.322556e-05, 5.114342e-05, 
    6.87568e-05, 2.88537e-05, 8.470036e-06, 1.672554e-06, 2.464524e-06, 
    2.095589e-06, 3.932179e-06, 1.685465e-05, 2.489738e-05, 4.178379e-07,
  3.231559e-05, 0.0001261095, 8.086667e-05, 4.126427e-05, 6.685801e-05, 
    4.904854e-05, 2.711289e-05, 3.042659e-06, 3.312689e-06, 3.682509e-06, 
    3.223096e-06, 4.102208e-06, 8.905879e-06, 1.254721e-05, 1.305046e-05,
  6.897509e-06, 1.772337e-06, 1.03667e-06, 2.206631e-06, 5.875235e-07, 
    1.993878e-06, 4.732164e-06, 2.062555e-06, 5.561606e-06, 6.016823e-06, 
    4.216693e-06, 1.36633e-06, 4.350476e-07, 1.715277e-07, 2.377851e-10,
  1.148169e-05, 9.385292e-06, 2.69736e-07, 1.751301e-06, 1.268045e-06, 
    3.950036e-06, 5.466058e-06, 4.492173e-06, 1.356495e-05, 1.125937e-05, 
    9.170937e-06, 4.888443e-06, 2.264567e-06, 9.482807e-07, 7.114901e-10,
  4.641466e-05, 3.601625e-05, 2.153485e-06, 5.224482e-06, 7.155015e-06, 
    3.350376e-06, 2.375158e-06, 7.289904e-06, 2.473579e-05, 2.683412e-05, 
    3.325232e-05, 2.896957e-05, 1.392245e-05, 3.76499e-06, 8.635965e-09,
  6.869302e-05, 1.578638e-05, 7.067742e-06, 1.425542e-05, 1.140926e-05, 
    1.486316e-05, 1.278801e-05, 2.455981e-05, 4.985167e-05, 6.411858e-05, 
    9.27919e-05, 7.036098e-05, 4.416823e-05, 1.872136e-05, 1.716889e-06,
  8.675076e-05, 1.48587e-05, 8.255541e-07, 2.459672e-06, 3.454028e-06, 
    1.103292e-05, 2.186856e-05, 4.223071e-05, 8.007768e-05, 0.0001093268, 
    1.038727e-05, 3.999543e-05, 7.755019e-05, 3.267208e-05, 4.934373e-05,
  2.323886e-05, 1.567136e-05, 1.53362e-06, 1.508782e-06, 1.67488e-06, 
    4.910914e-06, 1.295827e-05, 2.614708e-05, 3.759679e-05, 1.153043e-05, 
    8.113124e-05, 0.0001161433, 8.021721e-05, 0.0001147909, 8.787876e-05,
  1.555456e-05, 1.527764e-05, 1.401429e-06, 4.532518e-06, 1.124866e-05, 
    1.497959e-05, 4.167936e-05, 2.821953e-05, 3.404327e-05, 3.037152e-05, 
    4.129051e-05, 7.414876e-05, 8.261814e-05, 0.0002121034, 7.231364e-05,
  2.374816e-05, 5.079743e-05, 2.100398e-05, 2.208728e-05, 2.731557e-05, 
    5.536967e-05, 5.605139e-05, 4.902093e-05, 3.26001e-05, 9.943498e-06, 
    1.0628e-05, 2.084791e-05, 5.126293e-05, 0.0002139064, 3.0712e-05,
  5.975952e-05, 9.653387e-05, 4.610911e-05, 3.511939e-05, 0.000113391, 
    0.0001086323, 8.39582e-05, 5.574153e-05, 3.225038e-06, 4.786274e-06, 
    2.028785e-06, 2.791748e-06, 8.808882e-06, 6.49475e-05, 2.475825e-05,
  0.000100984, 0.0001337004, 7.543057e-05, 4.73783e-05, 0.0001028823, 
    0.000102067, 4.211438e-05, 3.649202e-06, 6.93038e-06, 3.022946e-06, 
    1.213227e-06, 2.162975e-06, 2.166735e-06, 1.389654e-05, 1.25342e-05,
  9.24206e-06, 7.201873e-06, 1.074561e-05, 6.61169e-06, 1.366307e-06, 
    2.155673e-06, 8.646563e-06, 5.149617e-06, 3.86493e-05, 3.089432e-05, 
    1.247763e-05, 9.11259e-06, 5.122244e-06, 3.078366e-06, 4.424017e-08,
  2.808274e-06, 1.432834e-05, 2.210802e-05, 6.702863e-05, 5.215421e-05, 
    3.017459e-05, 2.168457e-05, 2.261802e-05, 6.026352e-05, 3.161885e-05, 
    1.262682e-05, 8.132424e-06, 6.980901e-06, 9.452996e-06, 4.967151e-07,
  6.634535e-05, 2.671801e-05, 1.28022e-05, 6.487322e-05, 0.0001085104, 
    3.572529e-05, 4.467142e-06, 3.753263e-05, 6.858871e-05, 3.848612e-05, 
    4.487809e-05, 3.370074e-05, 2.592545e-05, 2.461913e-05, 4.824518e-08,
  0.0001539851, 1.440979e-05, 1.917796e-05, 4.542146e-05, 2.56425e-05, 
    1.504482e-05, 1.274526e-05, 2.725415e-05, 5.989598e-05, 5.510498e-05, 
    8.623661e-05, 7.652923e-05, 7.143769e-05, 3.932344e-05, 4.211925e-06,
  0.0001936095, 2.84949e-05, 1.344945e-05, 2.515318e-05, 1.83218e-05, 
    2.216188e-05, 2.811754e-05, 3.410782e-05, 4.892137e-05, 4.441895e-05, 
    1.546038e-06, 3.048765e-05, 0.0001407121, 8.149045e-05, 0.0001088904,
  4.018789e-05, 4.251432e-05, 1.360661e-05, 3.385926e-05, 3.991985e-05, 
    2.359429e-05, 1.352344e-05, 8.545391e-06, 8.975919e-06, 9.511749e-07, 
    4.339542e-05, 0.0001120234, 0.0002004122, 0.0002348248, 0.0001251964,
  1.700253e-05, 2.078832e-05, 6.413984e-06, 1.570054e-05, 2.784965e-05, 
    1.819584e-05, 9.257992e-06, 6.65842e-06, 7.076028e-06, 1.740544e-05, 
    2.982269e-05, 6.830304e-05, 0.0002657058, 0.0004431485, 0.0001467942,
  2.523709e-05, 4.574591e-05, 2.135206e-05, 1.624027e-05, 4.446168e-05, 
    4.237367e-05, 1.16988e-05, 4.901335e-06, 1.654105e-05, 2.648363e-05, 
    3.60651e-05, 7.995024e-05, 0.0002896054, 0.0004969227, 6.660887e-05,
  7.435928e-05, 0.0001096922, 5.056563e-05, 2.536416e-05, 6.955076e-05, 
    0.0001133061, 4.675819e-05, 1.818295e-05, 7.367965e-06, 4.36997e-05, 
    6.314174e-05, 0.0001210338, 0.0003012134, 0.0003703446, 0.000127607,
  0.0001212195, 0.0001452349, 5.570001e-05, 9.946774e-06, 4.13279e-05, 
    5.434015e-05, 5.374459e-05, 1.123692e-05, 5.167551e-05, 9.829447e-05, 
    0.000108821, 0.000108074, 0.0001836126, 0.0002237663, 0.0001313537,
  2.876816e-05, 2.075358e-05, 0.0001261586, 0.0001005934, 4.067328e-05, 
    7.264662e-05, 0.0001391716, 0.0001484887, 0.0002245698, 0.0001259965, 
    3.764543e-05, 1.104844e-05, 1.445516e-06, 1.21805e-06, 1.54865e-09,
  1.343402e-05, 1.362828e-05, 5.18605e-05, 0.0001994162, 0.0001218448, 
    9.969686e-05, 0.0001333165, 0.0001733154, 0.0002301611, 0.0001127129, 
    4.028848e-05, 8.65675e-06, 3.087266e-06, 4.92027e-06, 2.731309e-07,
  8.212943e-05, 1.78621e-05, 2.47117e-06, 7.565055e-05, 0.0001250976, 
    9.135441e-05, 5.568561e-05, 0.0001767084, 0.0002086198, 0.0001059983, 
    7.242538e-05, 6.056984e-05, 3.425504e-05, 1.522231e-05, 2.563384e-07,
  9.471705e-05, 1.792316e-05, 2.927577e-05, 9.14435e-05, 9.653753e-05, 
    8.048087e-05, 6.519409e-05, 8.551228e-05, 0.0001042172, 8.431591e-05, 
    0.0001709703, 0.0002867918, 0.0002184122, 9.996746e-05, 1.874434e-05,
  4.608923e-05, 1.317352e-05, 2.168454e-05, 6.016569e-05, 9.82132e-05, 
    0.0001111448, 6.168305e-05, 5.665222e-05, 7.046351e-05, 0.0001044565, 
    7.937143e-05, 0.0003303204, 0.0005211012, 0.0002717226, 0.0001962676,
  6.670336e-06, 8.747285e-06, 6.115909e-06, 3.70558e-05, 8.715522e-05, 
    7.508639e-05, 4.917346e-05, 4.729295e-05, 7.033536e-05, 2.18484e-05, 
    0.0001126148, 0.0003330361, 0.0004812843, 0.000399398, 0.000179458,
  6.763677e-06, 1.032374e-05, 4.410621e-06, 1.046652e-05, 4.313622e-05, 
    4.152721e-05, 5.542215e-05, 1.926856e-05, 2.951265e-05, 1.849952e-05, 
    3.060262e-05, 7.953357e-05, 0.0002651159, 0.0004284357, 0.000154182,
  1.522451e-05, 2.878267e-05, 1.54e-05, 2.313825e-05, 3.714574e-05, 
    5.02436e-05, 3.292325e-05, 1.853045e-05, 3.808509e-05, 1.761617e-05, 
    2.508986e-05, 2.734372e-05, 9.424317e-05, 0.0003551615, 5.78588e-05,
  2.474517e-05, 4.654691e-05, 4.448199e-05, 6.385783e-05, 9.129562e-05, 
    0.0001073045, 8.378731e-05, 8.913992e-05, 1.604627e-05, 3.746538e-05, 
    3.193123e-05, 3.814834e-05, 9.154556e-05, 0.0002126593, 9.558813e-05,
  1.314621e-05, 3.842087e-05, 4.490985e-05, 8.064188e-05, 0.0001488357, 
    0.0001845547, 0.0001524847, 4.266599e-05, 6.745006e-05, 6.494809e-05, 
    8.899409e-05, 0.000113674, 0.000159458, 0.0001827356, 0.0001839106,
  5.472549e-06, 1.68998e-05, 5.392068e-05, 5.52463e-05, 2.859682e-07, 
    7.039099e-06, 9.072644e-06, 3.892999e-06, 9.794588e-06, 2.21906e-05, 
    1.459915e-05, 1.470448e-05, 5.781813e-06, 5.515225e-06, 4.057064e-08,
  2.052516e-06, 7.149487e-07, 5.03396e-06, 8.25842e-06, 8.171359e-06, 
    7.109617e-06, 7.836152e-06, 3.382601e-06, 9.606892e-06, 1.016501e-05, 
    9.06128e-06, 1.324833e-05, 7.591592e-06, 7.914563e-06, 5.61668e-10,
  2.754216e-06, 1.491806e-07, 4.34143e-08, 5.506057e-06, 2.85053e-05, 
    8.708536e-06, 2.04065e-06, 4.872641e-06, 1.574117e-05, 1.951253e-05, 
    2.834358e-05, 3.26038e-05, 1.27533e-05, 5.909495e-06, 4.909789e-09,
  1.300299e-05, 1.436932e-06, 7.258355e-07, 1.740341e-06, 4.08043e-06, 
    3.204967e-06, 3.741665e-06, 8.223074e-06, 1.942265e-05, 4.69918e-05, 
    7.792268e-05, 5.201676e-05, 2.96418e-05, 2.105263e-05, 1.951284e-06,
  1.421852e-05, 1.296273e-06, 3.169094e-07, 9.7954e-07, 2.030609e-06, 
    4.305124e-06, 1.067174e-05, 1.913055e-05, 4.807687e-05, 6.309672e-05, 
    4.766992e-05, 3.785626e-05, 6.738047e-05, 2.903752e-05, 3.264357e-05,
  6.902373e-06, 3.001533e-06, 4.09069e-07, 3.267916e-06, 3.621676e-06, 
    8.418499e-06, 1.478699e-05, 3.179281e-05, 4.289207e-05, 5.742344e-05, 
    7.738305e-05, 5.988562e-05, 4.74355e-05, 9.103264e-05, 6.269256e-05,
  6.52983e-06, 4.719274e-06, 4.156486e-06, 3.891732e-06, 1.107879e-05, 
    8.645929e-06, 1.573178e-05, 2.60519e-05, 4.625114e-05, 2.78368e-05, 
    1.186489e-05, 1.35833e-05, 2.332984e-05, 0.000119796, 5.167301e-05,
  1.086928e-05, 1.032369e-05, 6.795597e-06, 8.610183e-06, 1.393901e-05, 
    7.554168e-06, 7.218037e-06, 1.173685e-05, 2.460404e-05, 5.495746e-06, 
    4.062861e-06, 8.410192e-06, 1.261624e-05, 8.974028e-05, 1.354255e-05,
  2.055824e-05, 2.492158e-05, 1.786605e-05, 2.072157e-05, 1.298109e-05, 
    1.481498e-05, 1.971874e-05, 1.758677e-05, 5.554499e-06, 3.766695e-06, 
    6.377139e-06, 1.265715e-05, 1.270731e-05, 2.03394e-05, 1.316767e-05,
  3.306238e-05, 2.881612e-05, 2.367214e-05, 1.69008e-05, 8.611007e-06, 
    9.863331e-06, 1.549448e-05, 3.25912e-06, 3.243198e-06, 2.705942e-06, 
    9.128285e-06, 1.03266e-05, 1.318078e-05, 7.357812e-06, 8.749864e-06,
  0.0001580086, 0.0001102663, 0.0001635701, 0.0001291647, 7.449561e-05, 
    9.040629e-05, 0.0001230214, 9.317737e-05, 0.0001401984, 6.963499e-05, 
    2.247765e-05, 8.055131e-06, 4.282918e-07, 1.841017e-06, 2.851499e-07,
  9.840159e-05, 0.0001381864, 0.000170209, 0.0002870527, 0.0002292588, 
    0.0001713182, 0.0001211627, 0.0001153079, 0.000144482, 7.704778e-05, 
    1.607605e-05, 5.28832e-06, 1.509097e-06, 5.270546e-06, 9.410916e-09,
  0.0003739761, 0.0002645137, 0.0001956803, 0.0003267736, 0.000327319, 
    0.0001967284, 9.665707e-05, 0.0001465285, 0.000144393, 6.17238e-05, 
    1.07692e-05, 4.867372e-06, 5.307278e-06, 3.515227e-06, 1.305178e-08,
  0.000419867, 0.000153161, 9.561999e-05, 0.0002109006, 0.0002064863, 
    0.0001350518, 0.0001163873, 0.0001491128, 0.000110407, 4.373052e-05, 
    2.317885e-05, 3.265839e-05, 3.248023e-05, 1.203778e-05, 4.903015e-07,
  0.0004152653, 0.0001344319, 1.598031e-05, 1.729343e-05, 1.809646e-05, 
    3.744259e-05, 6.301241e-05, 8.37443e-05, 5.806642e-05, 3.108638e-05, 
    1.250272e-06, 1.413679e-05, 8.890233e-06, 2.042625e-05, 2.776359e-05,
  0.0001989572, 0.0001060082, 1.283119e-05, 2.245527e-05, 4.17827e-05, 
    2.739308e-05, 1.934517e-05, 1.305697e-05, 3.083727e-06, 1.21822e-06, 
    1.997555e-05, 3.46581e-05, 4.8302e-05, 4.335355e-05, 3.347889e-05,
  7.99202e-05, 6.028735e-05, 2.524727e-05, 4.099267e-05, 7.774487e-05, 
    7.001806e-05, 4.100649e-05, 7.111667e-06, 2.190862e-06, 1.359546e-05, 
    3.328191e-05, 6.435151e-05, 4.677842e-05, 9.578836e-05, 2.887622e-05,
  8.273066e-05, 8.133195e-05, 4.673806e-05, 3.215632e-05, 6.991744e-05, 
    7.66951e-05, 4.609473e-05, 4.079046e-06, 7.33728e-06, 1.815732e-05, 
    7.472761e-05, 8.610442e-05, 5.662716e-05, 0.0001260917, 1.027949e-05,
  0.0001922519, 0.0001519558, 7.253603e-05, 3.291372e-05, 5.983323e-05, 
    9.882796e-05, 4.500322e-05, 1.56956e-05, 7.882892e-06, 2.861519e-05, 
    4.291525e-05, 5.484896e-05, 4.538994e-05, 4.294379e-05, 6.767742e-07,
  0.0002502112, 0.000220951, 0.0001093051, 5.753152e-05, 9.850659e-05, 
    9.437223e-05, 6.189617e-05, 3.065046e-05, 4.559872e-05, 3.546035e-05, 
    1.859337e-05, 1.669605e-05, 3.831572e-05, 3.820086e-05, 1.096044e-05,
  0.000158057, 0.0001442917, 0.0001075114, 9.563734e-05, 4.225152e-05, 
    3.699359e-05, 7.815901e-05, 4.489615e-05, 0.0002177682, 0.0001429942, 
    4.281731e-05, 1.18455e-05, 5.385719e-07, 3.967973e-06, 3.2389e-08,
  0.0001056005, 0.0002515569, 0.0002057287, 0.0003691019, 0.0003145234, 
    0.0003131881, 0.0002583966, 0.0002957185, 0.000328017, 0.0001859735, 
    5.282955e-05, 5.672992e-06, 1.747591e-06, 6.412292e-06, 1.136239e-07,
  0.0003338169, 0.0003600384, 0.0003143616, 0.0004488005, 0.0004946812, 
    0.0003544881, 0.0002188086, 0.0002916812, 0.0002774295, 0.0001355384, 
    3.758131e-05, 8.839568e-06, 8.964118e-06, 7.305029e-06, 1.0526e-08,
  0.0005182751, 0.000305167, 0.0002480661, 0.0002909144, 0.0002781574, 
    0.0001936005, 0.0001413954, 0.0001717575, 0.0001358925, 5.622329e-05, 
    1.459571e-05, 3.353156e-05, 5.697662e-05, 3.38861e-05, 3.906851e-06,
  0.000553768, 0.0003019363, 0.0001303104, 0.0001210623, 7.347816e-05, 
    5.357654e-05, 6.000851e-05, 5.456785e-05, 3.455775e-05, 5.186422e-06, 
    7.900582e-08, 4.678719e-06, 2.765321e-05, 5.326239e-05, 9.655266e-05,
  0.0003018336, 0.0002525725, 0.0001876473, 0.0001489129, 0.0001535637, 
    0.0001152097, 7.757099e-05, 3.164808e-05, 1.377631e-05, 3.176523e-06, 
    1.223954e-05, 4.362155e-05, 0.0001793645, 0.0002281809, 0.0001208343,
  0.0001651574, 0.0001932883, 0.0001978907, 0.0001498115, 0.0002345939, 
    0.0002137984, 0.0002357297, 0.0001962585, 0.0001491626, 0.0001055303, 
    9.573706e-05, 0.0001811463, 0.0003694333, 0.0003861462, 9.618371e-05,
  0.0001715305, 0.0001984005, 0.0001517736, 0.0001727034, 0.0002172114, 
    0.000283158, 0.0003385271, 0.0003646406, 0.0003440981, 0.0001736323, 
    0.0001859564, 0.0003087227, 0.0002498594, 0.0003533751, 5.821661e-06,
  0.0001750179, 0.0001793008, 0.0001551808, 0.0001421209, 0.0001867409, 
    0.0002475695, 0.0002720587, 0.0002977886, 0.0001978126, 0.0001510004, 
    0.0001711776, 0.0002773624, 0.0002569185, 0.0001573427, 2.553658e-08,
  0.0001197424, 0.000174236, 0.000178728, 0.0001630549, 0.0001979837, 
    0.0002170628, 0.0002299171, 0.0001960281, 0.0002172927, 0.0001682231, 
    0.0001161864, 0.0001482385, 0.0002304369, 0.0001781846, 8.442115e-05,
  4.079791e-06, 1.360159e-05, 1.480881e-05, 2.028262e-05, 1.288645e-05, 
    2.972664e-05, 7.288832e-05, 0.0001045935, 0.0002482028, 0.0002238851, 
    9.247976e-05, 3.338931e-05, 2.263806e-06, 1.35132e-06, 3.731338e-08,
  7.480899e-07, 1.626857e-06, 3.218385e-06, 1.590667e-05, 5.696241e-05, 
    5.264135e-05, 5.844006e-05, 0.0001094799, 0.0002008999, 0.0001832983, 
    0.0001071486, 2.911807e-05, 9.673627e-06, 6.143704e-06, 3.434597e-07,
  4.133914e-07, 4.62754e-06, 1.741376e-07, 6.696923e-06, 4.279708e-05, 
    3.416836e-05, 3.197253e-05, 8.607343e-05, 0.0001696937, 0.0001675155, 
    0.0001290448, 6.153839e-05, 3.737306e-05, 1.597484e-05, 3.379976e-06,
  1.061792e-06, 6.803254e-06, 1.326509e-05, 1.471266e-05, 2.44433e-05, 
    3.439643e-05, 4.186857e-05, 9.786833e-05, 0.0001613237, 0.000120033, 
    0.0001368191, 0.0001266455, 7.184017e-05, 6.39331e-05, 3.731155e-05,
  5.024499e-07, 1.610721e-06, 7.860017e-06, 1.248517e-05, 1.629574e-05, 
    2.476547e-05, 3.85298e-05, 7.541051e-05, 0.0001084648, 0.0001892151, 
    0.0002000303, 0.0001792086, 0.0002354202, 0.0001064112, 7.23888e-05,
  1.260766e-06, 4.217887e-07, 1.062387e-06, 2.501091e-06, 5.440719e-06, 
    1.659968e-05, 3.715523e-05, 7.747128e-05, 0.0001343465, 0.0001614874, 
    0.0001395093, 0.0001565466, 0.0001632341, 0.0001287991, 9.782355e-05,
  8.621683e-06, 1.931627e-06, 2.501417e-07, 4.969042e-06, 4.467504e-06, 
    7.187702e-06, 2.438996e-05, 4.765323e-05, 6.978431e-05, 5.875175e-05, 
    3.436325e-05, 4.660079e-05, 6.682862e-05, 0.0001461703, 6.520023e-05,
  1.625029e-05, 1.34696e-05, 1.821765e-06, 2.887012e-06, 5.998921e-06, 
    4.75233e-06, 7.71105e-06, 1.37764e-05, 4.155442e-05, 3.833672e-05, 
    4.192687e-05, 6.659772e-05, 8.373936e-05, 0.0001291658, 3.577503e-05,
  3.576323e-05, 2.607e-05, 5.756504e-06, 5.277529e-06, 1.138292e-05, 
    1.939972e-05, 1.531216e-05, 1.680678e-05, 2.137687e-05, 5.362123e-05, 
    5.942996e-05, 7.135645e-05, 9.008508e-05, 0.0001199062, 5.24022e-05,
  5.171453e-05, 3.543488e-05, 9.33538e-06, 3.006812e-06, 1.222625e-05, 
    1.937373e-05, 2.88783e-05, 2.084104e-05, 7.465536e-05, 6.812799e-05, 
    6.613301e-05, 7.140201e-05, 7.864661e-05, 4.700074e-05, 3.739528e-05,
  2.450884e-05, 1.289287e-05, 4.832441e-05, 0.0001033976, 6.149359e-05, 
    0.0001017944, 0.0001417533, 0.0001271474, 0.000142603, 6.963593e-05, 
    2.014299e-05, 7.3116e-06, 5.312215e-06, 5.075859e-06, 7.213916e-07,
  1.002179e-05, 3.518887e-05, 5.144237e-05, 0.0002362296, 0.0001981482, 
    0.0001697089, 0.0001785984, 0.0002226061, 0.0002026471, 9.010013e-05, 
    4.477185e-05, 2.705453e-05, 1.176095e-05, 4.92704e-06, 1.609575e-06,
  0.000207434, 0.0001992631, 3.580774e-05, 0.0002050561, 0.0002886879, 
    0.0002038633, 9.962485e-05, 0.0002548202, 0.0002383898, 0.0001327849, 
    9.981272e-05, 9.686932e-05, 6.032478e-05, 2.415108e-05, 5.723323e-07,
  0.0004107008, 0.0001624517, 4.885874e-05, 0.0001296875, 0.0001574274, 
    0.0001267888, 0.0001259371, 0.000209754, 0.0001888646, 0.0001278747, 
    0.0001238772, 0.0001962224, 0.0002086367, 0.0001088916, 4.011649e-05,
  0.0003507031, 0.0001306881, 2.31953e-05, 3.695034e-05, 6.346325e-05, 
    0.0001137816, 0.0001246567, 0.0001198692, 0.0001084318, 7.512968e-05, 
    5.724055e-06, 5.478803e-05, 0.0002909437, 0.0003249093, 0.0001596211,
  0.0001056882, 7.697483e-05, 2.913348e-05, 3.738509e-05, 6.458307e-05, 
    7.546428e-05, 6.990301e-05, 3.895838e-05, 2.391576e-05, 8.86928e-06, 
    6.218303e-05, 0.000194186, 0.0004938306, 0.0004488481, 0.0002123544,
  5.997031e-05, 6.38533e-05, 3.642455e-05, 3.940057e-05, 6.864976e-05, 
    6.862633e-05, 5.495506e-05, 3.812276e-05, 4.010817e-05, 7.552793e-05, 
    0.0001587848, 0.0002425865, 0.0003242457, 0.0004151406, 0.0001572201,
  8.30773e-05, 0.0001048254, 6.884774e-05, 3.965983e-05, 9.736523e-05, 
    0.000193826, 0.0002054558, 0.0001664686, 0.0001318054, 8.049889e-05, 
    0.0001090981, 0.0001343355, 0.0001038446, 0.0002094887, 4.913705e-05,
  0.0001941762, 0.000276087, 0.0002251355, 0.0001967229, 0.0003718146, 
    0.0004969219, 0.0003388801, 0.0002414293, 5.61415e-05, 6.617372e-05, 
    8.21112e-05, 9.493241e-05, 6.58378e-05, 0.0001122294, 1.254156e-05,
  0.0003590942, 0.0004954281, 0.0004353484, 0.0003816989, 0.0004033354, 
    0.0003977046, 0.0002850263, 9.033093e-05, 5.387146e-05, 6.588564e-05, 
    6.074068e-05, 8.055918e-05, 0.0001152054, 8.086066e-05, 2.193437e-05,
  1.609245e-07, 1.453441e-07, 1.95182e-06, 3.829038e-07, 8.223396e-07, 
    1.070779e-05, 6.635499e-05, 8.381002e-05, 0.0001182278, 6.814038e-05, 
    1.685136e-05, 3.734236e-06, 8.127778e-08, 6.695456e-08, 4.158232e-11,
  8.748167e-09, 1.626363e-06, 2.67554e-06, 1.236568e-05, 3.36968e-05, 
    6.276293e-05, 7.953598e-05, 0.0001007106, 0.0001178887, 6.482163e-05, 
    1.667573e-05, 3.981771e-06, 2.382253e-06, 1.933488e-06, 6.916493e-12,
  8.55756e-06, 2.882192e-05, 1.317991e-05, 3.921681e-05, 0.0001447261, 
    9.514377e-05, 3.063665e-05, 0.0001094338, 0.0001143155, 4.969284e-05, 
    3.23669e-05, 5.774786e-05, 5.611961e-05, 2.869926e-05, 3.306602e-08,
  6.447132e-05, 5.323128e-06, 6.07112e-06, 6.614676e-05, 7.311986e-05, 
    3.873212e-05, 2.052178e-05, 6.073768e-05, 5.327419e-05, 3.139675e-05, 
    8.543312e-05, 0.000249926, 0.0002561036, 0.0001249181, 2.174581e-05,
  9.450359e-05, 7.111058e-06, 5.218732e-07, 4.319052e-07, 3.158573e-07, 
    4.498693e-06, 5.533421e-06, 1.04602e-05, 2.017814e-05, 5.667166e-05, 
    2.112892e-05, 0.0002750112, 0.000426164, 0.0002433949, 0.0001669984,
  5.448974e-05, 1.38583e-05, 3.263666e-07, 1.268255e-07, 4.091674e-07, 
    5.651906e-07, 2.15041e-06, 4.6284e-06, 2.197924e-05, 0.0001518956, 
    0.0004268468, 0.0004344671, 0.000315231, 0.0003269884, 0.0002548369,
  2.024689e-05, 9.436546e-06, 4.009194e-07, 1.295801e-07, 1.148388e-07, 
    3.081832e-07, 8.38152e-06, 5.953184e-05, 0.0002964707, 0.0003663554, 
    0.00017014, 0.0001212738, 0.0001315246, 0.000246391, 0.0001301587,
  3.297437e-05, 1.395647e-05, 2.426195e-06, 8.6618e-08, 2.269745e-05, 
    0.0001166315, 0.0001565014, 0.0001844206, 0.0003029552, 0.0002340255, 
    0.0001752705, 0.000156518, 0.0001098852, 0.0001291188, 3.196833e-05,
  7.163196e-05, 9.392513e-05, 9.216759e-05, 0.000109141, 0.0002169743, 
    0.0002622825, 0.0002256763, 0.0001692868, 0.0001432818, 0.0002408879, 
    0.0001487539, 9.540938e-05, 5.537061e-05, 3.162039e-05, 9.102615e-06,
  0.0001752221, 0.0002641895, 0.0002490001, 0.0002604263, 0.0002565693, 
    0.0002260773, 0.0001892611, 0.0001382807, 0.0001221308, 0.0001028739, 
    4.13038e-05, 1.523962e-05, 5.518782e-06, 4.180125e-06, 2.730655e-06,
  3.839885e-06, 8.825497e-07, 1.197811e-05, 2.86255e-06, 2.085928e-07, 
    3.146979e-08, 8.597969e-08, 1.668507e-06, 1.192589e-05, 1.579526e-05, 
    8.602222e-06, 1.127646e-06, 2.411653e-07, 5.676036e-07, 4.284943e-10,
  2.360255e-07, 7.566305e-06, 6.79414e-06, 7.959163e-06, 4.876556e-06, 
    1.331803e-06, 2.804838e-06, 8.137218e-06, 2.299449e-05, 2.544123e-05, 
    1.333492e-05, 3.941614e-06, 2.611785e-06, 1.431689e-06, 2.271431e-10,
  5.195118e-05, 4.147341e-05, 1.675217e-05, 2.83753e-05, 2.982384e-05, 
    7.586721e-06, 3.221048e-06, 1.064755e-05, 3.902817e-05, 3.431452e-05, 
    2.337349e-05, 2.191197e-05, 1.647238e-05, 6.599607e-06, 3.872733e-09,
  7.815169e-05, 2.634042e-05, 1.144484e-05, 2.785253e-05, 1.188476e-05, 
    9.269664e-06, 7.64889e-06, 2.03694e-05, 3.294514e-05, 2.853377e-05, 
    5.237688e-05, 9.094532e-05, 0.000104446, 6.236836e-05, 1.203256e-06,
  7.457594e-05, 4.246169e-05, 5.826519e-06, 1.0426e-05, 7.882991e-06, 
    8.546854e-06, 1.132286e-05, 2.097263e-05, 2.57135e-05, 3.158999e-05, 
    1.868176e-05, 6.827569e-05, 0.0001086581, 0.0001177749, 0.0001465387,
  3.179319e-05, 2.877257e-05, 3.905341e-06, 6.812507e-06, 1.040195e-05, 
    1.144098e-05, 8.566106e-06, 1.142434e-05, 1.176956e-05, 4.172489e-06, 
    1.972018e-05, 2.9968e-05, 7.360072e-05, 0.0002104036, 0.0002669218,
  1.752547e-05, 1.7929e-05, 1.819085e-05, 4.719653e-06, 1.675077e-05, 
    1.533236e-05, 1.266225e-05, 1.640846e-05, 5.823957e-06, 3.938962e-06, 
    2.527206e-06, 4.174954e-06, 2.894677e-05, 0.0003617424, 0.0002520242,
  2.175851e-05, 2.850515e-05, 2.028134e-05, 2.655415e-05, 2.279427e-05, 
    3.14651e-05, 1.880666e-05, 9.307042e-06, 1.17129e-05, 1.164223e-05, 
    2.010616e-05, 2.437466e-05, 6.402891e-05, 0.0002833868, 0.0001285304,
  3.255195e-05, 2.931027e-05, 3.049478e-05, 3.14683e-05, 3.392826e-05, 
    5.988738e-05, 4.809658e-05, 2.594411e-05, 2.814411e-05, 0.0001358141, 
    0.0001112301, 6.655317e-05, 8.572728e-05, 9.697179e-05, 9.74879e-05,
  1.42839e-05, 2.571834e-05, 2.316281e-05, 1.597568e-05, 3.486517e-05, 
    6.559702e-05, 9.927731e-05, 0.0001250942, 0.0001281301, 6.153581e-05, 
    4.465059e-05, 3.766347e-05, 3.115555e-05, 2.415249e-05, 1.742131e-05,
  4.465293e-06, 1.747901e-06, 1.944997e-05, 9.103755e-06, 4.430055e-06, 
    9.295966e-07, 1.266187e-07, 1.879023e-09, 2.101687e-10, 3.810239e-10, 
    1.595687e-09, 1.479286e-10, 6.959028e-14, 7.356536e-11, 4.729254e-11,
  7.647097e-06, 1.248376e-05, 5.837989e-06, 8.280715e-06, 8.388414e-06, 
    1.000675e-05, 4.265426e-06, 4.976203e-07, 1.535704e-07, 1.342957e-06, 
    6.037947e-07, 6.784565e-08, 2.698766e-10, 2.068338e-10, 6.88494e-10,
  2.335021e-05, 7.637836e-05, 3.316834e-05, 3.024554e-05, 5.067577e-05, 
    2.581343e-05, 4.37565e-06, 5.060496e-06, 5.489127e-06, 3.073122e-06, 
    1.297488e-06, 5.171214e-08, 6.983748e-09, 7.041356e-09, 6.57266e-09,
  7.054467e-06, 1.015049e-05, 1.554367e-05, 6.054189e-05, 4.0465e-05, 
    2.075099e-05, 1.124723e-05, 9.99683e-06, 5.751641e-06, 1.303542e-06, 
    7.435773e-08, 9.917486e-09, 3.365849e-08, 4.819853e-08, 7.06159e-08,
  1.589194e-05, 6.884749e-06, 2.169559e-06, 7.068639e-06, 5.092888e-06, 
    2.733755e-06, 2.199482e-06, 2.64505e-06, 1.731273e-06, 5.677594e-07, 
    4.812731e-08, 1.006722e-09, 6.518816e-10, 4.72772e-08, 2.548679e-06,
  3.094543e-05, 9.377054e-06, 6.932718e-07, 3.721864e-08, 3.407229e-08, 
    1.98295e-08, 1.210833e-08, 2.440734e-07, 4.555039e-07, 1.888565e-07, 
    4.010424e-09, 2.9098e-09, 7.047248e-10, 2.201778e-07, 5.985817e-06,
  7.953761e-06, 3.892312e-06, 5.789585e-07, 1.386942e-08, 4.429044e-10, 
    1.50192e-10, 1.58313e-11, 2.529546e-09, 6.153711e-09, 3.113766e-09, 
    7.826496e-10, 3.825905e-09, 1.201873e-08, 3.726127e-06, 1.505072e-06,
  3.977199e-06, 8.733201e-07, 1.645098e-07, 1.183528e-08, 9.673111e-10, 
    6.615304e-11, 4.416179e-12, 3.57885e-11, 2.73113e-09, 1.177591e-09, 
    5.187963e-11, 1.175798e-09, 6.788786e-09, 8.796274e-06, 5.687929e-07,
  5.228463e-06, 1.924922e-06, 5.35308e-07, 1.132784e-07, 1.321235e-09, 
    1.822255e-09, 8.208377e-10, 6.404966e-12, 1.013476e-10, 1.764359e-10, 
    1.927157e-10, 2.917701e-09, 1.968598e-08, 1.25058e-06, 3.718311e-07,
  1.123925e-05, 2.213834e-05, 3.786226e-06, 2.86273e-07, 7.036121e-10, 
    5.808402e-14, 1.08755e-12, 2.995897e-10, 2.550369e-09, 1.67089e-09, 
    7.704958e-09, 1.348909e-07, 5.199348e-07, 3.476077e-07, 4.026375e-08,
  5.269914e-11, 1.39716e-11, 6.144068e-14, 5.337334e-12, 2.228573e-10, 
    9.233862e-08, 1.090285e-07, 4.995434e-09, 5.193357e-10, 1.413555e-10, 
    4.320439e-08, 4.162246e-10, 2.296476e-14, 1.143516e-29, 5.951166e-29,
  8.406249e-09, 2.111654e-09, 1.156226e-10, 7.994322e-10, 8.843412e-08, 
    1.33303e-06, 4.427887e-06, 1.903135e-06, 1.79511e-06, 3.654802e-06, 
    9.236509e-07, 1.891547e-08, 2.310855e-10, 6.414341e-13, 8.726184e-27,
  1.262204e-06, 4.0766e-06, 3.599033e-07, 3.866516e-08, 1.153123e-06, 
    5.257779e-06, 6.871209e-06, 9.802335e-06, 7.235956e-06, 3.342178e-06, 
    1.195392e-06, 8.349761e-08, 2.609954e-09, 1.684298e-10, 1.122397e-13,
  1.233232e-05, 8.91869e-06, 1.766125e-06, 5.29682e-06, 4.698717e-06, 
    3.525768e-06, 3.843541e-06, 5.787172e-06, 6.187965e-06, 1.665406e-06, 
    1.322383e-07, 6.560667e-09, 8.283629e-10, 2.918553e-10, 5.329127e-10,
  9.824739e-05, 2.514061e-05, 1.306219e-06, 1.426338e-06, 1.200169e-06, 
    3.721245e-07, 6.97427e-07, 1.146019e-06, 1.148482e-06, 6.032231e-07, 
    9.142421e-08, 5.035107e-09, 5.770018e-10, 1.387233e-11, 4.625223e-09,
  7.553183e-05, 2.531538e-05, 1.372166e-06, 4.641881e-08, 2.606665e-08, 
    1.451643e-08, 5.900712e-09, 7.159704e-09, 4.258433e-09, 3.009358e-09, 
    3.326754e-09, 3.422109e-09, 2.111479e-10, 3.151822e-11, 2.436668e-06,
  1.849896e-05, 1.643674e-05, 4.774003e-06, 1.83525e-06, 2.296036e-06, 
    2.167258e-08, 1.624655e-08, 1.649517e-09, 4.283556e-10, 6.163497e-08, 
    2.235665e-08, 6.138952e-08, 4.357979e-08, 3.327185e-08, 2.100237e-06,
  3.099862e-05, 2.374602e-05, 1.672519e-05, 9.321357e-06, 7.903183e-06, 
    6.470729e-06, 2.73128e-06, 1.088692e-06, 3.621815e-06, 9.893447e-06, 
    1.004716e-05, 1.402097e-05, 4.855786e-07, 4.014839e-05, 4.967567e-06,
  5.400822e-05, 0.0001102224, 6.473633e-05, 4.177442e-05, 5.196422e-05, 
    7.334016e-05, 2.974857e-05, 4.156634e-05, 8.545221e-05, 9.538844e-05, 
    6.132563e-05, 7.500414e-05, 7.127682e-05, 7.017826e-05, 2.397608e-06,
  6.413011e-05, 0.0001640202, 9.671125e-05, 5.405245e-05, 9.756692e-05, 
    7.859839e-05, 7.705883e-05, 8.229847e-05, 7.218657e-05, 1.852337e-05, 
    8.335851e-06, 6.018791e-06, 1.583555e-05, 3.171902e-05, 1.255234e-05,
  1.009121e-06, 1.22238e-08, 5.233819e-09, 4.294048e-09, 1.403808e-10, 
    1.320198e-15, 3.82557e-26, 2.846746e-26, 1.746669e-26, 5.895475e-20, 
    2.780478e-08, 5.893945e-10, 1.314054e-12, 2.471897e-18, 2.810838e-27,
  3.395536e-06, 2.331485e-06, 5.202641e-06, 6.731164e-08, 1.649382e-07, 
    2.128621e-08, 1.306741e-09, 1.659608e-08, 5.454175e-07, 3.089996e-06, 
    2.186598e-06, 1.959953e-07, 3.858035e-10, 1.1685e-16, 4.305434e-26,
  0.0001193121, 0.0001201045, 8.759153e-06, 5.708469e-06, 9.161477e-06, 
    2.066834e-06, 1.19831e-06, 8.578385e-07, 1.694499e-06, 2.12881e-06, 
    1.99606e-06, 2.130721e-07, 1.34983e-08, 2.735659e-10, 1.071821e-13,
  0.0001736483, 8.797431e-05, 5.699358e-05, 4.335996e-05, 2.075831e-05, 
    7.992554e-06, 1.734758e-06, 4.70059e-07, 2.810702e-07, 1.817006e-06, 
    2.511301e-07, 1.282182e-08, 2.588723e-09, 3.990289e-11, 1.242693e-09,
  0.0002726308, 0.0001004707, 3.522646e-05, 3.38814e-05, 1.486319e-05, 
    6.598008e-06, 1.205264e-06, 1.153007e-07, 3.713591e-08, 9.361373e-08, 
    5.978257e-08, 3.039915e-10, 3.152527e-10, 1.599299e-09, 5.996394e-09,
  0.0001918279, 0.0001382638, 4.428246e-05, 3.11693e-05, 3.073509e-05, 
    7.540071e-06, 2.539094e-06, 1.766854e-07, 5.273261e-11, 5.699149e-12, 
    1.520974e-08, 3.277534e-10, 5.494371e-12, 2.631416e-09, 1.369765e-06,
  0.000149089, 0.0001431157, 7.737172e-05, 6.053306e-05, 5.071381e-05, 
    3.511949e-05, 2.693025e-06, 7.785721e-09, 5.124515e-10, 2.661915e-09, 
    5.493299e-09, 1.576554e-09, 2.979925e-10, 2.459416e-07, 9.225296e-07,
  0.0001913935, 0.0002013989, 0.0001177543, 8.273547e-05, 0.0001032845, 
    0.0001070876, 3.966414e-05, 1.845035e-06, 2.522404e-08, 3.214958e-09, 
    4.225791e-08, 7.658119e-09, 3.163689e-09, 4.629069e-06, 8.312629e-07,
  0.0001987142, 0.0002291574, 0.0001683888, 8.976769e-05, 0.0001121064, 
    0.0001561625, 9.529097e-05, 3.667633e-05, 2.692088e-07, 9.323826e-06, 
    9.620902e-06, 1.582187e-05, 9.572776e-06, 1.048057e-05, 1.538508e-06,
  0.0002037823, 0.0003298139, 0.0001574926, 6.813709e-05, 9.651508e-05, 
    0.0001098126, 0.0001147992, 8.258533e-05, 0.0001072774, 8.276122e-05, 
    2.76076e-05, 2.792852e-05, 4.618506e-05, 4.082353e-05, 3.074719e-05,
  9.115339e-06, 1.179354e-05, 8.361095e-06, 8.401003e-06, 2.360953e-06, 
    1.411217e-06, 3.265379e-06, 6.841067e-06, 3.574234e-05, 4.009659e-05, 
    1.566935e-05, 5.294813e-06, 3.854593e-07, 9.178081e-08, 4.807552e-14,
  7.091675e-06, 1.248239e-05, 1.164876e-05, 1.784771e-05, 2.911461e-05, 
    2.288164e-05, 1.798555e-05, 1.944662e-05, 5.323397e-05, 4.599852e-05, 
    1.994968e-05, 6.639397e-06, 6.067824e-07, 1.837083e-07, 1.491414e-10,
  2.548331e-05, 2.282742e-05, 7.60242e-06, 2.680172e-05, 7.742729e-05, 
    5.040584e-05, 2.262089e-05, 2.728404e-05, 5.315197e-05, 3.427049e-05, 
    1.919289e-05, 9.776731e-06, 4.94139e-06, 1.956307e-06, 7.248942e-08,
  4.870271e-05, 1.026895e-05, 1.583016e-05, 3.0975e-05, 4.505084e-05, 
    4.984222e-05, 5.326263e-05, 4.213759e-05, 3.86707e-05, 2.470627e-05, 
    1.732445e-05, 1.795822e-05, 2.5252e-05, 1.694769e-05, 1.69691e-06,
  4.434734e-05, 1.537401e-05, 1.168117e-05, 1.808652e-05, 2.337463e-05, 
    4.231868e-05, 4.209841e-05, 3.525339e-05, 2.994448e-05, 1.662321e-05, 
    6.515418e-06, 7.923379e-05, 0.0001403635, 9.324597e-05, 0.0001035919,
  5.599111e-05, 3.150473e-05, 7.026819e-06, 1.90897e-05, 2.526966e-05, 
    4.362418e-05, 4.363407e-05, 2.71866e-05, 7.901363e-06, 4.483534e-06, 
    4.935825e-05, 6.172823e-05, 9.14124e-05, 0.0001225626, 0.0001301356,
  5.820421e-05, 2.84771e-05, 8.641861e-06, 1.162004e-05, 2.366098e-05, 
    2.159001e-05, 2.903674e-05, 1.649405e-05, 2.080915e-05, 4.519748e-05, 
    5.169706e-05, 3.116019e-05, 4.065095e-05, 0.000150686, 0.0001246862,
  5.545517e-05, 3.226701e-05, 8.948537e-06, 9.394435e-06, 1.531912e-05, 
    3.303067e-05, 3.856679e-05, 5.158348e-05, 6.213033e-05, 8.027035e-05, 
    4.482524e-05, 4.014823e-05, 5.862189e-05, 0.0001410778, 5.621038e-05,
  9.813534e-05, 0.0001099685, 4.231968e-05, 3.698701e-05, 6.90302e-05, 
    7.867889e-05, 6.060232e-05, 5.667383e-05, 6.504932e-05, 7.176639e-05, 
    5.127742e-05, 4.723103e-05, 5.260947e-05, 8.181821e-05, 1.901513e-05,
  0.0002183258, 0.0002038241, 0.0001194181, 6.84302e-05, 7.68083e-05, 
    8.465158e-05, 7.313613e-05, 3.332493e-05, 5.541181e-05, 4.518369e-05, 
    5.377369e-05, 5.837396e-05, 4.502778e-05, 3.222652e-05, 7.450632e-06,
  4.623606e-08, 9.769377e-09, 1.165598e-09, 4.965829e-10, 9.367686e-09, 
    4.950684e-08, 1.404113e-07, 2.646135e-07, 2.010725e-06, 1.768433e-06, 
    5.171339e-07, 1.422083e-07, 1.309115e-07, 2.204814e-07, 8.0178e-08,
  2.203657e-06, 5.331441e-08, 2.798326e-08, 2.966767e-08, 8.738295e-08, 
    5.121377e-07, 2.177803e-06, 3.285874e-06, 1.534707e-05, 9.565431e-06, 
    1.76295e-06, 2.489441e-07, 1.160311e-07, 1.157546e-07, 2.433046e-08,
  3.511144e-05, 5.164053e-05, 1.645007e-06, 3.565818e-07, 5.080357e-06, 
    7.943182e-06, 6.319525e-06, 1.841532e-05, 2.089399e-05, 1.010284e-05, 
    2.015053e-06, 6.947594e-07, 3.403165e-07, 8.639775e-08, 3.773674e-09,
  0.0001171462, 5.286609e-05, 2.300732e-05, 2.828228e-05, 1.368872e-05, 
    9.408961e-06, 1.127471e-05, 1.526474e-05, 1.19192e-05, 4.014198e-06, 
    2.258404e-06, 3.972037e-06, 3.365057e-06, 4.981266e-07, 7.520171e-09,
  0.0001291713, 4.802267e-05, 6.163054e-06, 3.446124e-06, 1.424077e-06, 
    1.209284e-06, 1.787786e-06, 3.189437e-06, 2.64586e-06, 1.346973e-06, 
    3.974537e-09, 2.153119e-09, 4.077475e-07, 8.617933e-08, 2.003632e-07,
  0.0001349072, 5.794441e-05, 2.112528e-05, 1.592088e-05, 1.229712e-05, 
    2.718928e-06, 2.007503e-06, 1.462939e-06, 4.788934e-07, 4.585453e-06, 
    6.094739e-07, 2.999931e-06, 1.320564e-06, 2.689814e-06, 7.275793e-06,
  0.0001553623, 0.000121692, 0.0001090302, 0.0001150386, 0.0001200208, 
    0.0001053687, 4.741846e-05, 3.430622e-05, 0.0001114925, 9.265292e-05, 
    3.603347e-05, 5.154996e-06, 7.431789e-06, 8.817778e-05, 2.317621e-05,
  0.0001923828, 0.0002177961, 0.0001736016, 0.0001336821, 0.0001350604, 
    0.0001562049, 0.000151169, 0.0001373413, 0.000191966, 8.14732e-05, 
    3.151123e-05, 6.858022e-05, 0.0001047959, 0.0003058676, 6.889924e-05,
  0.0001976846, 0.0002524544, 0.0001639477, 9.263084e-05, 7.958036e-05, 
    9.227259e-05, 7.786822e-05, 8.852343e-05, 7.272793e-05, 3.664085e-05, 
    1.989655e-05, 3.098047e-05, 0.0001196305, 0.0002474329, 4.737262e-05,
  0.0001042263, 0.000139701, 0.0001228943, 6.447506e-05, 6.608305e-05, 
    5.556731e-05, 4.826039e-05, 3.830456e-05, 2.579241e-05, 3.08429e-05, 
    1.932416e-05, 2.688731e-05, 7.43563e-05, 0.0001062449, 6.729285e-05,
  3.516567e-06, 4.072329e-06, 1.421373e-05, 7.181186e-07, 5.117047e-07, 
    1.323626e-08, 9.121083e-11, 4.602612e-11, 5.66848e-08, 2.30787e-08, 
    1.678365e-09, 2.919041e-11, 1.82409e-09, 1.286802e-08, 8.220637e-12,
  5.066027e-06, 2.630215e-05, 3.530164e-05, 3.572256e-05, 1.829031e-05, 
    7.285495e-06, 1.529784e-06, 4.008239e-07, 3.183551e-07, 1.747343e-07, 
    7.985726e-09, 2.952343e-09, 9.637155e-09, 1.698521e-08, 9.953172e-11,
  7.82045e-05, 0.0001530602, 3.627936e-05, 0.0001142501, 0.0001415902, 
    5.880378e-05, 7.302688e-06, 2.23085e-06, 1.383796e-06, 4.570902e-07, 
    1.039331e-08, 1.14966e-08, 2.545708e-08, 2.617979e-08, 5.399699e-10,
  0.000212916, 0.0001264013, 8.642775e-05, 0.000157756, 0.0001590766, 
    6.121182e-05, 3.431621e-05, 9.339957e-06, 1.929332e-06, 2.955765e-07, 
    1.932866e-08, 3.01151e-08, 1.258532e-07, 1.275571e-07, 2.406809e-10,
  0.0003092164, 0.0001764843, 4.01945e-05, 2.715696e-05, 2.11654e-05, 
    1.879608e-05, 1.9136e-05, 9.478795e-06, 1.213082e-06, 6.06647e-08, 
    7.4052e-11, 5.160059e-09, 2.683834e-09, 6.772971e-10, 1.566634e-06,
  0.000343985, 0.0002074742, 8.745347e-05, 4.414167e-05, 3.30798e-05, 
    3.710118e-05, 1.762282e-05, 6.73773e-06, 2.792044e-07, 7.503357e-07, 
    2.070019e-07, 2.622723e-06, 8.500397e-07, 3.661838e-07, 9.523346e-06,
  0.0001870881, 0.0001681386, 0.0001783205, 0.0001362745, 0.0001290824, 
    9.088015e-05, 4.615506e-05, 1.358006e-05, 9.424493e-06, 1.982353e-05, 
    4.61408e-07, 4.680832e-07, 3.088305e-08, 1.582939e-05, 1.308098e-05,
  0.0001431919, 0.0001419522, 0.0001031479, 0.0001028189, 0.0001305641, 
    0.0001528863, 0.0001224679, 6.774021e-05, 5.525113e-05, 1.120668e-05, 
    6.752592e-07, 7.906724e-07, 2.608767e-06, 3.947113e-05, 9.570871e-06,
  0.0001477749, 0.000187751, 0.0001539829, 9.237527e-05, 8.527843e-05, 
    0.0001059391, 0.0001041608, 0.0001260702, 0.0001171272, 7.995378e-05, 
    4.237295e-05, 3.642928e-05, 3.302738e-05, 4.025301e-05, 1.652432e-05,
  0.0001362711, 0.0002068193, 0.0002238072, 0.0001933437, 0.0001495905, 
    0.0001206073, 0.0001310415, 9.868954e-05, 0.0001365091, 0.0001022806, 
    5.019604e-05, 4.313552e-05, 5.536186e-05, 4.897563e-05, 3.21304e-05,
  0.0001551377, 0.0001544041, 8.208332e-05, 7.890834e-05, 4.22871e-05, 
    5.328726e-05, 8.407861e-05, 0.0001331831, 0.0002056042, 0.0001642866, 
    6.27563e-05, 2.188318e-05, 1.184268e-05, 1.564266e-05, 4.862347e-07,
  7.375095e-05, 0.0001570341, 0.000105501, 0.000124044, 0.0001099959, 
    7.837061e-05, 8.484904e-05, 0.000105577, 0.0001620936, 0.0001439641, 
    6.710638e-05, 2.507846e-05, 1.281167e-05, 8.099534e-06, 3.788238e-08,
  0.000168247, 0.0001636729, 8.993348e-05, 0.0001805826, 0.0002089002, 
    0.0001149935, 5.091508e-05, 6.900724e-05, 0.0001203233, 0.0001011796, 
    6.801847e-05, 4.921955e-05, 3.337682e-05, 1.557572e-05, 3.843332e-08,
  0.0002152361, 0.0001590491, 0.0001370861, 0.000158821, 0.0001374719, 
    9.395013e-05, 6.494993e-05, 8.028778e-05, 8.509481e-05, 6.376486e-05, 
    6.938598e-05, 9.341972e-05, 7.999197e-05, 5.660991e-05, 1.505884e-05,
  0.0001570444, 0.0001186919, 0.0001062278, 0.0001074312, 7.861533e-05, 
    7.415598e-05, 6.539511e-05, 7.897006e-05, 6.281513e-05, 9.102694e-05, 
    0.0001112769, 0.0001180286, 0.0001780249, 0.000102724, 9.104906e-05,
  6.89688e-05, 9.361809e-05, 0.000114147, 0.0001083052, 8.69143e-05, 
    6.524842e-05, 7.372771e-05, 7.280969e-05, 9.273705e-05, 8.687329e-05, 
    5.827257e-05, 8.011311e-05, 0.0001160847, 0.000215265, 0.0001147615,
  3.100037e-05, 4.796337e-05, 5.288081e-05, 5.394651e-05, 5.582394e-05, 
    8.58354e-05, 0.0001283003, 0.000151444, 0.0001437503, 7.195829e-05, 
    2.716918e-05, 2.143405e-05, 4.364959e-05, 0.0001979374, 0.0001078824,
  1.245325e-05, 1.435935e-05, 1.075767e-05, 1.8467e-05, 2.018294e-05, 
    4.511074e-05, 0.0001093067, 0.0001232529, 0.0001437445, 6.00393e-05, 
    4.306405e-05, 4.092973e-05, 3.839954e-05, 0.0001358447, 4.179183e-05,
  6.952003e-06, 1.242926e-05, 1.357731e-05, 3.421845e-05, 3.118078e-05, 
    4.628831e-05, 7.432827e-05, 0.0001162274, 8.493598e-05, 6.122905e-05, 
    5.362167e-05, 6.051797e-05, 6.21846e-05, 5.841599e-05, 3.933667e-05,
  6.136381e-06, 1.669674e-05, 3.996798e-05, 6.664837e-05, 7.832245e-05, 
    7.990028e-05, 9.190402e-05, 5.759573e-05, 3.02082e-05, 3.197645e-05, 
    3.875601e-05, 5.574034e-05, 7.100042e-05, 9.519718e-05, 7.339482e-05,
  0.0002217244, 0.0003193864, 0.0003214022, 0.0003234255, 0.0002225847, 
    0.0001858995, 0.000181694, 0.0001948802, 0.0002798506, 0.0002188814, 
    7.905575e-05, 1.845727e-05, 2.209985e-06, 3.808394e-07, 6.818784e-09,
  9.212983e-05, 0.0001782294, 0.0002189656, 0.0002070162, 0.0002417874, 
    0.0002330722, 0.0002128627, 0.0002224383, 0.0002469499, 0.0002117323, 
    9.641015e-05, 3.535138e-05, 1.057817e-05, 3.07314e-06, 1.187055e-07,
  3.829694e-05, 4.889677e-05, 8.401535e-05, 0.0001179296, 0.0001582955, 
    0.0001654982, 0.0001462018, 0.0001810218, 0.0001964027, 0.0001466444, 
    8.222192e-05, 4.885227e-05, 2.032911e-05, 5.721639e-06, 1.396413e-07,
  4.000171e-05, 2.504437e-05, 3.149005e-05, 6.252847e-05, 9.421654e-05, 
    0.0001109867, 0.0001179399, 0.0001349724, 0.0001327254, 7.941123e-05, 
    6.034587e-05, 4.540037e-05, 2.751802e-05, 1.689003e-05, 9.249603e-06,
  3.651408e-05, 2.868268e-05, 3.098471e-05, 4.9517e-05, 7.466356e-05, 
    9.51075e-05, 0.0001015592, 0.0001061365, 0.0001103438, 0.0001408007, 
    8.818042e-05, 4.566089e-05, 0.000127996, 4.661304e-05, 5.574639e-05,
  1.803112e-05, 2.287245e-05, 3.954118e-05, 4.843263e-05, 6.588941e-05, 
    8.367182e-05, 0.000101919, 0.0001354609, 0.0002272427, 0.0002294291, 
    9.235233e-05, 2.232132e-05, 8.636253e-06, 3.209278e-05, 7.147387e-05,
  2.572195e-05, 1.850584e-05, 3.028621e-05, 2.559623e-05, 2.93308e-05, 
    4.178465e-05, 7.227518e-05, 0.00012774, 0.0001489419, 7.026763e-05, 
    1.534901e-05, 3.743094e-06, 7.218543e-07, 1.328749e-05, 1.952637e-05,
  1.646052e-05, 1.102964e-05, 1.471801e-05, 1.448005e-05, 7.966088e-06, 
    1.404089e-05, 2.305637e-05, 3.962214e-05, 8.643753e-05, 2.532904e-05, 
    8.888668e-06, 7.190899e-06, 2.295947e-06, 6.442429e-06, 3.233564e-06,
  1.016778e-05, 1.147286e-05, 1.901433e-05, 2.722963e-05, 1.56613e-05, 
    2.338265e-05, 3.907531e-05, 6.960484e-05, 4.506695e-05, 8.696526e-06, 
    4.929352e-06, 5.350613e-06, 2.245859e-06, 1.352221e-06, 6.026817e-07,
  2.097026e-06, 9.029261e-06, 5.270015e-05, 7.616472e-05, 7.118186e-05, 
    6.471949e-05, 9.119385e-05, 5.305849e-05, 2.340982e-05, 7.908535e-06, 
    3.749321e-06, 6.384172e-06, 7.258841e-06, 1.264664e-06, 2.762036e-07,
  0.0002153508, 0.0001383759, 9.251449e-05, 7.346829e-05, 5.736247e-05, 
    6.345269e-05, 8.356944e-05, 9.618538e-05, 0.0001442793, 0.0001086005, 
    3.673414e-05, 1.522667e-05, 8.068029e-06, 1.012402e-05, 2.924853e-07,
  7.125444e-05, 3.21384e-05, 1.334855e-05, 2.729545e-05, 2.991749e-05, 
    3.844802e-05, 4.738748e-05, 6.107953e-05, 0.0001313754, 0.0001291502, 
    6.067872e-05, 3.092993e-05, 1.523931e-05, 1.998892e-05, 3.56432e-06,
  7.428331e-05, 6.623387e-05, 2.997178e-05, 2.022302e-05, 2.354391e-05, 
    2.597904e-05, 2.827069e-05, 6.10822e-05, 0.00012234, 0.0001263111, 
    9.667718e-05, 6.905726e-05, 4.989177e-05, 4.365655e-05, 2.845145e-05,
  4.749096e-05, 2.644484e-05, 1.661065e-05, 1.965536e-05, 2.086443e-05, 
    2.876524e-05, 3.364573e-05, 4.664094e-05, 7.29809e-05, 9.898824e-05, 
    0.0001369653, 0.000133665, 9.516216e-05, 7.885281e-05, 6.05136e-05,
  1.354018e-05, 9.818781e-06, 8.528146e-06, 1.012049e-05, 1.77152e-05, 
    2.139054e-05, 2.79531e-05, 3.411676e-05, 8.430772e-05, 0.0002107321, 
    0.0002068924, 9.068293e-05, 9.567518e-05, 3.995037e-05, 2.68443e-05,
  3.848568e-06, 3.405764e-06, 4.431956e-06, 8.373355e-06, 1.620384e-05, 
    1.748245e-05, 2.216138e-05, 4.925862e-05, 0.0001404868, 0.0001082182, 
    5.728452e-05, 2.898125e-05, 1.051661e-05, 3.319194e-06, 7.769567e-06,
  1.005544e-06, 1.054159e-06, 6.170922e-06, 1.027314e-05, 1.710251e-05, 
    1.903085e-05, 3.29487e-05, 6.058684e-05, 6.838046e-05, 3.73261e-05, 
    1.842033e-05, 1.152213e-05, 1.879907e-06, 8.197119e-06, 2.533364e-06,
  5.642711e-07, 1.155961e-06, 6.268822e-06, 1.870667e-05, 2.13197e-05, 
    2.599302e-05, 2.337697e-05, 3.150217e-05, 5.852534e-05, 2.810894e-05, 
    1.328601e-05, 8.609511e-06, 2.559487e-06, 1.149675e-05, 1.887843e-06,
  1.398971e-07, 2.737655e-06, 1.784766e-05, 3.924768e-05, 4.19604e-05, 
    4.353588e-05, 4.456966e-05, 6.209299e-05, 3.012451e-05, 2.145898e-05, 
    1.171698e-05, 1.376266e-05, 1.236703e-05, 8.641024e-06, 5.70647e-07,
  3.635599e-07, 3.678987e-06, 4.400963e-05, 7.176676e-05, 7.857778e-05, 
    6.913247e-05, 7.784484e-05, 3.341611e-05, 2.461553e-05, 1.711276e-05, 
    1.529134e-05, 2.251627e-05, 2.181489e-05, 9.121333e-06, 2.928848e-06,
  2.592888e-05, 5.170674e-06, 3.097254e-06, 1.250859e-05, 2.385737e-05, 
    4.578516e-05, 8.647886e-05, 0.0001464855, 0.0001920931, 0.0001507673, 
    0.0001137762, 0.0001122272, 0.0001141227, 6.811089e-05, 3.961937e-05,
  1.376589e-06, 1.182304e-06, 3.086941e-06, 1.784029e-05, 3.989241e-05, 
    6.23114e-05, 0.0001055001, 0.0001498157, 0.0001430946, 0.0001157036, 
    9.208078e-05, 7.92766e-05, 5.821647e-05, 2.468907e-05, 1.51725e-05,
  3.308233e-06, 4.766016e-06, 3.445563e-06, 5.921425e-06, 1.641524e-05, 
    3.31686e-05, 5.218908e-05, 6.098103e-05, 5.395766e-05, 4.425445e-05, 
    3.573419e-05, 2.614447e-05, 1.074316e-05, 8.53987e-06, 1.87366e-06,
  1.088194e-06, 5.255982e-06, 3.877733e-06, 7.459204e-06, 7.701196e-06, 
    9.98507e-06, 1.202985e-05, 1.136724e-05, 1.517334e-05, 4.188694e-05, 
    6.667218e-05, 4.826512e-05, 1.412662e-05, 1.610326e-05, 1.108455e-06,
  7.670092e-07, 4.39706e-06, 4.789654e-06, 4.63072e-06, 3.39356e-06, 
    5.891389e-06, 1.141235e-05, 1.49885e-05, 4.621107e-05, 0.0001203139, 
    4.269693e-05, 1.614391e-05, 6.536861e-05, 1.348228e-05, 1.662808e-05,
  9.018762e-07, 9.626122e-06, 8.016044e-06, 8.014727e-06, 5.185378e-06, 
    7.801831e-06, 1.220982e-05, 2.061862e-05, 6.801441e-05, 4.59244e-05, 
    5.816142e-05, 4.675086e-05, 2.368674e-05, 1.989542e-05, 2.103169e-05,
  1.381256e-06, 6.973218e-06, 8.597121e-06, 5.262612e-06, 3.624194e-06, 
    1.809918e-06, 4.541983e-06, 8.19208e-06, 1.633266e-05, 5.036778e-05, 
    5.501097e-05, 3.730676e-05, 1.821138e-05, 5.675346e-05, 9.301641e-06,
  3.183228e-08, 1.154555e-06, 4.730814e-06, 4.271095e-06, 1.759067e-06, 
    2.18495e-06, 3.071667e-06, 3.795441e-06, 3.303228e-05, 3.604926e-05, 
    4.099757e-05, 2.986464e-05, 1.964492e-05, 4.560501e-05, 4.24365e-06,
  7.353864e-08, 8.466399e-07, 5.848751e-06, 1.512301e-05, 1.223996e-05, 
    1.622158e-05, 1.513945e-05, 1.647979e-05, 1.596524e-05, 4.42225e-05, 
    3.729189e-05, 3.165982e-05, 2.45517e-05, 1.435699e-05, 1.743483e-06,
  4.011137e-06, 3.719128e-06, 1.337688e-05, 1.935589e-05, 2.582566e-05, 
    4.027689e-05, 3.598749e-05, 2.129648e-05, 4.607705e-05, 5.205893e-05, 
    4.335992e-05, 2.887834e-05, 2.367031e-05, 6.372584e-06, 3.973315e-06,
  1.691281e-05, 1.030608e-05, 4.924622e-06, 1.841761e-05, 1.404574e-05, 
    1.887786e-05, 5.08964e-05, 5.744758e-05, 5.685226e-05, 2.468964e-05, 
    5.8733e-06, 3.860658e-06, 3.076299e-06, 2.957696e-06, 1.634446e-06,
  9.485715e-06, 2.669855e-06, 1.087158e-06, 2.42878e-05, 2.40121e-05, 
    1.721575e-05, 2.810491e-05, 6.513268e-05, 6.160257e-05, 3.042676e-05, 
    8.950104e-06, 2.508814e-06, 9.572311e-07, 2.162481e-06, 8.709492e-07,
  1.997097e-05, 6.764886e-06, 5.062987e-06, 1.309608e-05, 2.233366e-05, 
    1.807521e-05, 1.740991e-05, 4.615376e-05, 6.35505e-05, 4.011057e-05, 
    2.15158e-05, 1.015286e-05, 3.3856e-06, 1.468824e-06, 4.049925e-07,
  4.021105e-05, 1.819607e-05, 2.715391e-05, 4.758364e-05, 3.972293e-05, 
    3.536673e-05, 3.315746e-05, 5.466854e-05, 7.004155e-05, 6.734161e-05, 
    5.647017e-05, 3.951705e-05, 1.680168e-05, 9.81057e-06, 1.918925e-06,
  9.367679e-06, 1.404411e-05, 2.419271e-05, 4.420257e-05, 5.669619e-05, 
    5.971284e-05, 5.892156e-05, 7.71211e-05, 9.4241e-05, 8.94532e-05, 
    1.281245e-06, 2.243268e-05, 8.395921e-05, 1.759256e-05, 2.128964e-05,
  1.39575e-06, 5.010829e-06, 1.220876e-05, 4.215247e-05, 6.495963e-05, 
    7.062762e-05, 7.097986e-05, 7.440625e-05, 8.519363e-05, 6.55815e-06, 
    6.67947e-05, 0.0001701509, 8.769608e-05, 4.982261e-05, 2.072452e-05,
  1.38692e-05, 9.750283e-06, 8.919011e-06, 2.741507e-05, 5.299352e-05, 
    5.509397e-05, 5.087847e-05, 4.724761e-05, 4.459809e-05, 3.154822e-05, 
    0.0001293798, 0.0002034165, 0.0001594053, 0.0001357519, 1.442112e-05,
  2.989263e-05, 4.751707e-05, 3.484196e-05, 5.43182e-05, 8.317483e-05, 
    7.91948e-05, 5.523012e-05, 5.824463e-05, 7.038286e-05, 7.47241e-05, 
    0.000139093, 0.0001767173, 0.0002010833, 0.0001556774, 1.559649e-05,
  7.444039e-05, 0.0001104088, 9.326774e-05, 0.0001312997, 0.0001967345, 
    0.0002053567, 0.0001533723, 0.0001506077, 8.92363e-05, 0.0002023397, 
    0.0001757668, 0.0001691883, 0.0002007915, 0.0001729016, 2.357579e-05,
  5.783554e-05, 0.0001494123, 0.0001683532, 0.0002008803, 0.0002656716, 
    0.0002945373, 0.0002779199, 0.0001156036, 0.0002458128, 0.0002346454, 
    0.0001816043, 0.0001851485, 0.0001960605, 0.0001949487, 7.747376e-05,
  5.929816e-05, 2.615877e-05, 5.107453e-05, 0.0001082708, 6.047959e-05, 
    4.443612e-05, 8.759251e-05, 0.0001317327, 0.0001770348, 0.0001168937, 
    5.371205e-05, 3.682601e-05, 1.627701e-05, 1.423768e-05, 3.065205e-07,
  1.486978e-05, 6.846251e-06, 5.588099e-06, 4.643562e-05, 2.679961e-05, 
    1.714912e-05, 3.033423e-05, 8.972397e-05, 0.0001396513, 9.21136e-05, 
    5.954175e-05, 4.248583e-05, 3.041713e-05, 2.846117e-05, 6.627378e-07,
  2.673588e-05, 5.854291e-06, 6.028083e-07, 2.920934e-06, 8.551619e-06, 
    9.937003e-06, 9.060169e-06, 4.91716e-05, 0.0001060537, 8.345137e-05, 
    9.187645e-05, 7.968832e-05, 4.051474e-05, 3.057957e-05, 4.075773e-07,
  1.679808e-05, 1.813833e-05, 3.002566e-05, 5.301116e-05, 6.712622e-05, 
    6.674642e-05, 4.70103e-05, 5.542046e-05, 8.526017e-05, 0.0001014529, 
    0.0001829874, 0.0002309349, 0.0001407026, 8.025989e-05, 1.079528e-05,
  8.435896e-06, 1.094922e-05, 1.729028e-05, 5.714846e-05, 5.625702e-05, 
    7.157275e-05, 7.424523e-05, 8.090522e-05, 8.79623e-05, 0.0001168808, 
    1.902601e-05, 0.0001441129, 0.0005701132, 0.0002025733, 0.0001246352,
  9.448437e-06, 1.824968e-05, 2.705657e-05, 4.506332e-05, 5.750159e-05, 
    5.157719e-05, 5.308369e-05, 6.70786e-05, 5.112993e-05, 1.910023e-05, 
    0.0001092698, 0.0002256505, 0.0003006969, 0.0002973314, 0.0001736946,
  2.888185e-05, 3.766877e-05, 4.795891e-05, 4.21931e-05, 3.41243e-05, 
    2.226491e-05, 2.240922e-05, 2.235633e-05, 1.141583e-05, 3.25434e-05, 
    8.342027e-05, 0.0001029666, 0.0001290653, 0.0002963621, 0.0001092783,
  4.886575e-05, 4.912415e-05, 4.337898e-05, 4.102499e-05, 2.180363e-05, 
    2.08739e-05, 2.113795e-05, 2.321505e-05, 5.713433e-05, 5.786816e-05, 
    9.1339e-05, 7.171251e-05, 7.152835e-05, 0.0001915131, 8.11927e-05,
  5.935885e-05, 5.568046e-05, 4.921049e-05, 5.442026e-05, 5.868874e-05, 
    7.235509e-05, 8.024308e-05, 9.569435e-05, 4.499478e-05, 9.579023e-05, 
    6.639479e-05, 7.005093e-05, 6.79588e-05, 0.000149862, 3.571887e-05,
  3.488124e-05, 4.263624e-05, 4.885485e-05, 2.976086e-05, 3.089438e-05, 
    0.000106615, 0.0001479278, 5.589595e-05, 5.98359e-05, 5.489206e-05, 
    4.541608e-05, 4.722469e-05, 4.600874e-05, 3.643159e-05, 2.791632e-05,
  1.836883e-13, 1.577014e-24, 5.35946e-27, 1.185294e-16, 3.662383e-30, 
    1.264928e-29, 1.912002e-28, 1.274472e-12, 9.532251e-11, 5.775648e-09, 
    3.956255e-07, 6.837568e-06, 7.320386e-06, 8.452509e-06, 1.180994e-06,
  4.56571e-12, 6.865595e-12, 1.070401e-15, 2.560999e-12, 3.166211e-11, 
    2.769968e-10, 2.096943e-10, 6.066901e-10, 5.507368e-09, 4.701282e-08, 
    6.177161e-07, 3.843128e-06, 4.817455e-06, 9.049746e-06, 3.407821e-07,
  2.130928e-07, 5.643583e-10, 6.549067e-09, 1.455032e-08, 1.376777e-08, 
    3.800503e-08, 2.596489e-08, 6.220687e-08, 2.584215e-07, 1.720646e-06, 
    8.536554e-06, 1.646482e-05, 1.110306e-05, 1.131745e-05, 3.879843e-07,
  1.725511e-06, 1.584941e-08, 2.363141e-08, 1.708438e-06, 1.995221e-06, 
    1.820376e-06, 1.536907e-06, 2.410059e-06, 2.910731e-06, 8.992176e-06, 
    4.394581e-05, 6.195411e-05, 6.214291e-05, 3.876991e-05, 7.682294e-06,
  2.589784e-07, 7.519374e-09, 3.922198e-08, 2.907469e-06, 3.351781e-06, 
    2.410058e-06, 6.138544e-06, 7.9121e-06, 7.203255e-06, 1.09811e-05, 
    1.462262e-06, 6.072249e-05, 0.0002437148, 5.578802e-05, 6.9457e-05,
  1.578295e-08, 4.109757e-09, 4.752769e-10, 1.159261e-06, 5.130296e-06, 
    1.852837e-06, 4.701027e-06, 5.60964e-06, 5.936904e-06, 3.005756e-06, 
    4.953209e-05, 0.000109355, 0.0001023946, 0.0001199135, 6.309718e-05,
  3.666577e-08, 1.670466e-08, 1.366929e-09, 8.555533e-07, 3.371138e-06, 
    3.690996e-06, 4.305349e-06, 5.24282e-06, 3.084642e-06, 1.34047e-05, 
    3.609377e-05, 4.830025e-05, 4.382502e-05, 0.0001128636, 3.274865e-05,
  7.127495e-08, 3.177479e-08, 4.825876e-09, 3.180348e-07, 2.487487e-06, 
    3.676885e-06, 2.717141e-06, 4.012452e-06, 1.276009e-05, 2.212341e-05, 
    4.255284e-05, 2.106264e-05, 2.361129e-05, 5.470788e-05, 1.406614e-05,
  1.463212e-06, 4.136234e-07, 2.388273e-08, 5.765013e-07, 1.836292e-06, 
    7.518056e-06, 8.227689e-06, 9.952573e-06, 3.116056e-06, 5.19399e-05, 
    2.827888e-05, 4.898897e-06, 1.009618e-05, 1.884976e-05, 6.336571e-06,
  4.232531e-06, 2.477321e-06, 3.558658e-07, 1.511142e-09, 1.252306e-07, 
    3.451339e-07, 3.668272e-06, 6.326687e-06, 2.778226e-05, 2.232e-05, 
    5.706371e-06, 2.825122e-06, 6.873405e-06, 5.934039e-06, 6.539958e-06,
  1.425498e-08, 1.34959e-08, 1.866636e-08, 4.323002e-07, 4.186016e-07, 
    2.500032e-07, 1.707323e-07, 3.199127e-08, 3.95202e-08, 5.274092e-08, 
    4.629297e-08, 2.225502e-08, 2.618705e-08, 1.114077e-07, 2.8956e-07,
  6.088103e-07, 1.936239e-08, 1.701093e-08, 2.350539e-07, 3.609543e-07, 
    2.25962e-07, 1.793283e-07, 1.409307e-07, 1.400103e-07, 8.507769e-08, 
    7.72871e-08, 6.513154e-08, 4.104651e-08, 5.880232e-07, 4.26917e-07,
  1.03576e-05, 1.712806e-05, 3.296076e-07, 5.284907e-07, 6.844129e-07, 
    3.60418e-07, 2.947152e-07, 2.87618e-07, 2.265963e-07, 1.589058e-07, 
    1.006226e-07, 2.681377e-07, 9.643907e-07, 1.093533e-06, 7.877034e-07,
  8.517128e-05, 8.909873e-06, 3.275947e-06, 3.176101e-06, 1.585286e-06, 
    8.259266e-07, 5.948851e-07, 4.86039e-07, 2.752867e-07, 1.542001e-07, 
    9.156898e-08, 2.967241e-07, 6.059641e-06, 7.376963e-06, 9.59407e-06,
  0.0001880015, 2.973455e-05, 8.060527e-06, 7.926626e-06, 4.617845e-06, 
    1.31202e-06, 5.088785e-07, 3.219623e-07, 1.850465e-07, 9.914277e-08, 
    1.191413e-08, 4.057857e-09, 7.615479e-06, 1.861719e-05, 5.057884e-05,
  0.0001578917, 6.135876e-05, 2.049147e-05, 1.690308e-05, 1.625222e-05, 
    7.288794e-06, 1.97963e-06, 3.797098e-07, 1.637888e-07, 2.375921e-09, 
    1.611839e-08, 1.449e-06, 1.566916e-05, 7.971236e-05, 3.786039e-05,
  5.420192e-05, 5.99145e-05, 3.4721e-05, 4.640832e-05, 5.098127e-05, 
    3.282021e-05, 1.073561e-05, 1.486801e-06, 1.064072e-09, 6.760343e-10, 
    1.385112e-09, 4.170619e-06, 9.062081e-06, 7.611916e-05, 2.22785e-05,
  2.957735e-05, 6.251612e-05, 3.618485e-05, 3.764211e-05, 6.382075e-05, 
    4.910696e-05, 1.389894e-05, 2.204013e-06, 2.355426e-08, 2.77153e-09, 
    6.675199e-07, 2.928704e-06, 4.4414e-06, 3.783562e-05, 1.397861e-06,
  6.898421e-05, 7.498056e-05, 3.45432e-05, 1.509501e-05, 3.349773e-05, 
    4.629174e-05, 8.887007e-06, 5.006531e-06, 1.589487e-08, 1.751906e-08, 
    2.140009e-06, 2.049027e-07, 5.029739e-06, 5.743879e-06, 1.063426e-07,
  8.60009e-05, 7.890246e-05, 3.645064e-05, 6.864826e-06, 9.147554e-06, 
    3.435976e-06, 3.941329e-06, 8.816316e-07, 1.558479e-06, 2.281746e-07, 
    1.142514e-06, 2.994127e-07, 4.06345e-06, 4.413636e-07, 3.90576e-07,
  0.0001304962, 2.086506e-05, 6.161428e-06, 8.881066e-06, 9.388763e-06, 
    1.262113e-05, 1.638087e-05, 9.844777e-06, 8.966138e-06, 5.049676e-06, 
    1.811559e-06, 6.592362e-07, 6.110923e-07, 4.346051e-07, 2.645709e-07,
  0.0001019884, 3.207056e-05, 7.452002e-06, 1.331778e-05, 1.414939e-05, 
    2.230094e-05, 3.735175e-05, 2.398628e-05, 2.147785e-05, 9.708317e-06, 
    2.467338e-06, 8.726017e-07, 8.322265e-07, 4.766347e-07, 3.416061e-07,
  0.0002130586, 0.0001818983, 5.67496e-05, 2.823395e-05, 3.445389e-05, 
    3.536691e-05, 2.311726e-05, 2.283902e-05, 2.012749e-05, 8.078365e-06, 
    2.019994e-06, 6.360122e-07, 8.513794e-07, 6.819852e-07, 5.294469e-07,
  0.0003148175, 0.0001036789, 6.661934e-05, 7.603862e-05, 3.995921e-05, 
    3.235408e-05, 4.389776e-05, 3.975916e-05, 1.256296e-05, 1.863887e-06, 
    8.931115e-07, 8.021181e-07, 1.047746e-06, 9.241462e-07, 1.233452e-06,
  0.0002216951, 9.792631e-05, 2.791123e-05, 3.731879e-05, 5.416143e-05, 
    8.791065e-05, 0.0001138563, 8.865081e-05, 2.246863e-05, 5.827544e-06, 
    2.473877e-09, 6.372097e-09, 4.984344e-07, 2.313678e-07, 4.766848e-07,
  0.0001059189, 0.0001009797, 3.316531e-05, 4.782073e-05, 9.991491e-05, 
    0.0001795355, 0.0002085274, 0.0001333358, 3.953027e-05, 4.335049e-08, 
    1.123014e-08, 9.942591e-09, 1.041665e-08, 2.563353e-07, 5.418224e-08,
  6.817433e-05, 7.60276e-05, 5.842775e-05, 5.825281e-05, 0.0001101894, 
    0.0001703704, 0.0001763245, 0.0001062461, 6.072867e-06, 8.858797e-07, 
    5.758119e-07, 4.737145e-09, 1.018153e-08, 6.272329e-07, 2.81797e-08,
  6.615036e-05, 8.617514e-05, 7.573488e-05, 5.704162e-05, 5.662848e-05, 
    6.11926e-05, 5.347175e-05, 4.623859e-05, 1.709647e-05, 1.034327e-06, 
    1.566075e-06, 1.186956e-06, 1.088231e-08, 5.68486e-06, 4.896236e-07,
  8.107052e-05, 8.332441e-05, 7.75777e-05, 6.444119e-05, 3.54326e-05, 
    2.313203e-05, 9.025623e-06, 1.100337e-05, 7.592381e-06, 7.902645e-06, 
    3.608754e-06, 4.539539e-06, 1.657496e-06, 4.561534e-06, 3.435527e-08,
  9.182638e-05, 7.565676e-05, 7.036055e-05, 5.842188e-05, 5.321739e-05, 
    3.044006e-05, 1.610997e-05, 1.113241e-06, 5.093159e-06, 7.142219e-06, 
    5.639716e-06, 6.928014e-06, 9.689632e-06, 3.835627e-06, 2.2075e-06,
  5.051999e-05, 4.297006e-05, 1.645312e-05, 6.335322e-06, 2.973846e-06, 
    6.15836e-06, 3.673894e-05, 5.31691e-05, 7.543249e-05, 4.091031e-05, 
    1.750223e-05, 1.519032e-05, 1.073008e-05, 6.925755e-06, 1.914056e-05,
  1.906217e-05, 6.990247e-06, 1.610086e-06, 6.590089e-06, 7.033788e-06, 
    2.403553e-05, 5.157479e-05, 7.492854e-05, 8.769668e-05, 4.589152e-05, 
    2.203133e-05, 1.583881e-05, 1.091436e-05, 7.179235e-06, 1.509773e-05,
  5.132332e-05, 1.445626e-05, 2.396239e-06, 6.960095e-06, 2.943661e-05, 
    4.386618e-05, 5.622449e-05, 7.810217e-05, 6.282978e-05, 2.820945e-05, 
    1.798137e-05, 1.264912e-05, 1.144957e-05, 7.680994e-06, 1.110283e-05,
  0.0001046344, 1.823203e-05, 5.372509e-06, 1.567989e-05, 2.367684e-05, 
    5.060427e-05, 9.00954e-05, 9.787269e-05, 4.541285e-05, 1.26497e-05, 
    1.077817e-05, 8.615566e-06, 9.229264e-06, 7.31555e-06, 1.216698e-05,
  6.338969e-05, 4.131385e-05, 1.972656e-05, 1.241216e-05, 1.677165e-05, 
    3.973663e-05, 7.56189e-05, 8.782977e-05, 6.117198e-05, 8.848547e-05, 
    3.829833e-05, 1.682305e-05, 2.843756e-05, 4.498573e-06, 1.222456e-05,
  1.400182e-05, 3.539741e-05, 4.091633e-05, 3.105996e-05, 3.115518e-05, 
    3.229659e-05, 4.543014e-05, 8.313909e-05, 0.0001519957, 0.0001428316, 
    9.832057e-05, 4.184054e-05, 4.54875e-06, 1.557092e-06, 9.861586e-06,
  4.205773e-06, 1.969408e-05, 5.456719e-05, 7.77104e-05, 9.061758e-05, 
    8.773938e-05, 6.690899e-05, 5.0964e-05, 5.431576e-05, 2.996858e-05, 
    1.958329e-05, 9.955847e-06, 1.916613e-06, 1.75671e-06, 5.878916e-06,
  3.708472e-07, 5.470124e-06, 2.853878e-05, 6.717623e-05, 9.244417e-05, 
    9.658756e-05, 6.295725e-05, 2.791412e-05, 5.089085e-05, 1.011356e-05, 
    1.301303e-05, 6.38601e-06, 1.204676e-06, 8.217553e-06, 7.9738e-06,
  2.117585e-07, 2.1661e-06, 9.354621e-06, 2.900877e-05, 3.743328e-05, 
    5.699251e-05, 5.068079e-05, 6.386524e-05, 1.05659e-05, 1.138154e-05, 
    8.357981e-06, 8.974682e-06, 1.385739e-06, 4.902076e-06, 3.409504e-06,
  1.040717e-07, 1.276683e-06, 1.104142e-05, 1.433039e-05, 3.210274e-05, 
    3.827686e-05, 4.867089e-05, 1.832386e-05, 1.431886e-05, 6.183021e-06, 
    9.432495e-06, 1.277355e-05, 4.66735e-06, 4.157841e-06, 2.441087e-06,
  2.220918e-05, 1.520668e-06, 2.645501e-06, 1.140668e-06, 2.372666e-06, 
    8.022921e-06, 1.183928e-05, 6.442121e-06, 2.918083e-05, 2.215424e-05, 
    1.184608e-05, 2.889447e-05, 3.668348e-05, 4.021507e-05, 1.784047e-05,
  1.336777e-05, 4.104378e-06, 1.437825e-07, 2.377076e-07, 2.693183e-07, 
    3.059074e-06, 1.21348e-05, 1.165065e-05, 2.107563e-05, 2.084674e-05, 
    1.332022e-05, 3.218553e-05, 4.423091e-05, 3.993657e-05, 1.866221e-05,
  5.741056e-06, 1.953451e-06, 7.450943e-08, 7.965441e-08, 1.880602e-06, 
    3.509214e-06, 9.470913e-06, 1.977126e-05, 2.388938e-05, 1.883946e-05, 
    2.177673e-05, 3.159723e-05, 4.342284e-05, 4.946281e-05, 2.261029e-05,
  2.256752e-05, 8.956138e-07, 1.020725e-06, 5.184454e-06, 7.313524e-06, 
    1.225102e-05, 1.630389e-05, 3.657683e-05, 3.018228e-05, 1.614462e-05, 
    3.000074e-05, 2.855393e-05, 2.436759e-05, 2.256376e-05, 2.422966e-05,
  1.750344e-05, 1.580633e-06, 5.369949e-07, 3.687704e-06, 6.934578e-06, 
    9.968695e-06, 2.084051e-05, 3.197672e-05, 3.169333e-05, 9.3718e-05, 
    0.0001060492, 0.0001030173, 0.0001031302, 1.711756e-05, 2.460083e-05,
  6.754651e-06, 4.864422e-06, 1.201334e-06, 3.145052e-06, 8.211171e-06, 
    9.331311e-06, 1.611995e-05, 3.50784e-05, 7.88016e-05, 0.0001020528, 
    9.518819e-05, 9.285401e-05, 4.944271e-05, 1.899927e-05, 1.98693e-05,
  1.266286e-06, 1.745366e-06, 3.54335e-08, 1.834225e-06, 5.897365e-06, 
    5.610845e-06, 7.906856e-06, 1.615373e-05, 3.631768e-05, 2.335158e-05, 
    1.45153e-05, 3.251758e-05, 2.43991e-05, 2.07118e-05, 8.066001e-06,
  3.550073e-07, 3.18807e-07, 2.31793e-08, 3.567698e-07, 9.658984e-07, 
    4.759862e-06, 3.894977e-06, 4.511669e-06, 1.914361e-05, 1.532035e-06, 
    7.1606e-06, 3.689068e-05, 3.974454e-05, 4.432706e-05, 2.684313e-06,
  1.714524e-09, 1.560919e-07, 5.740022e-07, 1.429298e-06, 1.260363e-06, 
    5.092169e-06, 8.81937e-06, 1.316125e-05, 3.076399e-06, 4.069361e-07, 
    3.528511e-06, 3.834284e-05, 5.604108e-05, 1.79338e-05, 8.888011e-06,
  1.581676e-10, 3.936086e-09, 2.359926e-08, 2.986376e-07, 6.12587e-07, 
    3.854084e-06, 9.189055e-06, 6.171733e-06, 5.703565e-06, 2.529361e-06, 
    3.281685e-06, 4.589262e-05, 5.794414e-05, 2.162211e-05, 5.347022e-06,
  0.0003086874, 7.320422e-05, 5.547611e-05, 4.748419e-05, 3.159424e-05, 
    2.104085e-05, 1.735195e-05, 1.014196e-05, 1.762965e-05, 1.662235e-05, 
    5.93452e-06, 4.521251e-06, 6.759346e-06, 1.154044e-05, 3.316624e-06,
  0.0002300328, 0.0002836277, 6.974226e-05, 3.570002e-05, 3.267046e-05, 
    3.056483e-05, 2.308123e-05, 1.208473e-05, 1.83103e-05, 8.098342e-06, 
    7.130437e-06, 3.607612e-06, 7.250634e-06, 1.135753e-05, 6.650589e-06,
  0.0001339216, 0.000383076, 0.0002731071, 6.518983e-05, 4.515164e-05, 
    2.484197e-05, 6.113482e-06, 6.757419e-06, 7.992731e-06, 4.035032e-06, 
    4.597397e-06, 2.597061e-06, 5.488347e-06, 1.458772e-05, 6.375737e-06,
  0.0001120912, 0.0001023398, 0.000160054, 0.0001520476, 5.311401e-05, 
    2.727873e-05, 1.402661e-05, 5.732481e-06, 4.053939e-06, 1.636392e-06, 
    1.508665e-06, 4.49728e-07, 2.034155e-06, 4.759459e-06, 1.629506e-05,
  9.301849e-05, 5.146666e-05, 5.271309e-05, 5.976798e-05, 4.556043e-05, 
    2.674061e-05, 1.30361e-05, 7.318396e-06, 2.198113e-06, 3.013653e-06, 
    1.232249e-07, 1.254214e-06, 7.449723e-06, 4.566425e-06, 2.994456e-05,
  4.620136e-05, 4.33907e-05, 3.408416e-05, 3.812066e-05, 4.167173e-05, 
    2.936191e-05, 1.577304e-05, 6.127233e-06, 4.87423e-06, 2.151741e-06, 
    1.796427e-05, 9.061282e-06, 6.217733e-06, 6.473444e-07, 2.512305e-05,
  2.051369e-05, 1.56637e-05, 1.163066e-05, 8.456507e-06, 1.037147e-05, 
    1.075411e-05, 8.439675e-06, 3.653123e-06, 3.576012e-06, 3.359081e-06, 
    5.583526e-08, 8.596481e-07, 1.586667e-06, 4.165716e-06, 9.683033e-06,
  4.003497e-06, 6.805319e-06, 4.953454e-06, 2.583456e-06, 1.799028e-06, 
    7.523789e-07, 9.158705e-07, 3.883533e-06, 2.660109e-05, 7.754329e-06, 
    1.600881e-07, 6.224615e-07, 2.182001e-06, 1.769871e-05, 3.279023e-06,
  3.003644e-06, 5.111992e-06, 2.19012e-06, 6.042968e-07, 1.397789e-06, 
    2.083314e-07, 3.456673e-07, 1.222116e-06, 4.863906e-07, 2.170346e-05, 
    4.017177e-07, 5.954586e-07, 4.134242e-06, 2.172574e-05, 2.874805e-05,
  6.428207e-08, 1.094789e-06, 1.76823e-07, 6.286152e-08, 8.021898e-08, 
    5.614799e-09, 1.62216e-09, 5.76762e-08, 1.113424e-05, 1.476752e-05, 
    3.25356e-06, 4.879571e-06, 1.806116e-05, 3.560845e-05, 3.391814e-05,
  0.0001747497, 0.0001278447, 5.187443e-05, 3.136238e-05, 1.81381e-05, 
    2.024524e-05, 1.130513e-05, 7.354906e-06, 2.155264e-06, 5.787305e-06, 
    9.040304e-06, 1.5801e-05, 2.117969e-05, 2.559514e-05, 5.44294e-05,
  0.0001280255, 0.0001668981, 1.96495e-05, 1.43762e-05, 2.9936e-05, 
    3.060585e-05, 1.831079e-05, 5.021829e-06, 1.50153e-06, 3.290133e-06, 
    4.025724e-06, 1.053058e-05, 1.070893e-05, 2.027606e-05, 2.887255e-05,
  8.844649e-05, 0.0001522541, 9.299093e-05, 3.280537e-05, 4.535408e-05, 
    3.843265e-05, 1.358825e-05, 1.022812e-05, 1.045863e-05, 3.003588e-06, 
    1.935897e-06, 1.399944e-06, 4.686111e-06, 2.387883e-05, 1.087786e-05,
  4.499961e-05, 2.218594e-05, 3.796998e-05, 9.435668e-05, 5.395992e-05, 
    6.220597e-05, 5.296033e-05, 2.809805e-05, 9.015187e-06, 3.780394e-06, 
    9.860742e-07, 1.28966e-07, 3.44397e-07, 6.429197e-06, 9.190157e-06,
  5.2503e-05, 1.276602e-05, 3.166805e-06, 1.012599e-05, 1.644767e-05, 
    3.306766e-05, 4.967645e-05, 2.826085e-05, 9.000093e-06, 4.33486e-06, 
    3.323352e-08, 1.606206e-08, 2.805479e-07, 3.232595e-07, 1.381019e-05,
  2.710471e-05, 1.058162e-05, 4.087226e-06, 7.423329e-06, 1.576186e-05, 
    2.42149e-05, 3.001757e-05, 1.640243e-05, 1.121852e-05, 6.249889e-08, 
    2.074801e-07, 1.367355e-08, 2.19327e-08, 1.350898e-07, 1.445473e-05,
  4.713408e-06, 4.306496e-06, 1.109623e-05, 9.925437e-06, 7.271258e-06, 
    9.747831e-06, 1.077196e-05, 6.855179e-06, 1.038925e-05, 2.5463e-06, 
    5.398434e-09, 1.08846e-08, 1.885423e-08, 9.638116e-08, 2.175585e-06,
  9.298049e-07, 3.221639e-06, 8.07156e-06, 6.026794e-06, 3.079834e-06, 
    1.964155e-06, 2.276733e-06, 4.454894e-06, 1.648488e-05, 3.991954e-06, 
    1.328419e-07, 1.489502e-08, 3.347581e-08, 4.270756e-08, 6.607024e-09,
  2.065398e-08, 1.707789e-06, 5.421595e-06, 2.508237e-06, 3.039312e-06, 
    4.498959e-06, 1.308647e-06, 8.692156e-07, 4.790051e-06, 2.451773e-05, 
    4.094475e-07, 4.394917e-08, 2.69047e-08, 2.094444e-08, 4.092584e-09,
  3.751766e-09, 1.457449e-06, 1.780398e-06, 1.556582e-06, 1.142694e-07, 
    1.265666e-08, 1.536269e-08, 1.87731e-06, 1.379929e-05, 2.840519e-05, 
    6.778666e-06, 2.220539e-08, 1.005249e-07, 7.316244e-07, 4.49833e-07,
  9.845011e-05, 0.0001343929, 0.0001959247, 0.0001535568, 7.152313e-05, 
    2.314054e-05, 1.633667e-06, 7.369891e-08, 4.205831e-06, 1.859587e-06, 
    7.278669e-07, 1.004637e-05, 2.407416e-05, 2.976959e-05, 4.143066e-05,
  0.0001194579, 0.0001610593, 0.0002365901, 0.0002143976, 0.0002099297, 
    0.0001273525, 4.924772e-05, 1.259228e-05, 1.251066e-05, 5.21983e-06, 
    6.369737e-07, 2.91825e-06, 1.531895e-05, 1.65466e-05, 1.618144e-05,
  0.000142846, 0.0001760936, 0.000193471, 0.0001830983, 0.000232025, 
    0.0001619855, 7.379134e-05, 3.914459e-05, 3.210635e-05, 1.20958e-05, 
    1.75807e-06, 1.539197e-06, 1.266731e-05, 2.526464e-05, 1.144037e-05,
  0.0001000762, 5.248006e-05, 6.614233e-05, 0.0001193, 0.0001151446, 
    0.0001049304, 8.375585e-05, 6.114657e-05, 4.416926e-05, 1.866667e-05, 
    2.94903e-06, 3.955597e-07, 1.574653e-06, 6.954573e-06, 2.261129e-05,
  0.0001028767, 3.215926e-05, 1.234775e-05, 2.439408e-05, 3.217333e-05, 
    3.137729e-05, 3.253543e-05, 2.928397e-05, 2.344327e-05, 7.312162e-06, 
    4.492288e-09, 1.247732e-08, 1.318062e-07, 2.662957e-07, 2.511048e-05,
  6.151897e-05, 4.863744e-05, 3.588527e-05, 2.902456e-05, 2.38642e-05, 
    6.703513e-06, 3.127306e-06, 2.674617e-06, 2.394019e-06, 1.453146e-08, 
    1.008946e-07, 8.018608e-08, 2.908977e-08, 1.202924e-07, 3.018892e-05,
  2.526806e-05, 3.663396e-05, 4.66403e-05, 3.385621e-05, 1.917104e-05, 
    3.447231e-06, 2.984513e-06, 6.62386e-07, 1.260585e-07, 2.260584e-08, 
    5.465102e-08, 6.437574e-08, 6.169088e-08, 1.084134e-07, 4.754609e-06,
  5.136744e-06, 9.590854e-06, 1.216762e-05, 8.864202e-06, 4.940671e-06, 
    3.969742e-06, 4.186081e-06, 3.682517e-06, 3.967475e-06, 1.670109e-08, 
    2.480238e-08, 5.743359e-08, 8.324589e-08, 8.336549e-08, 4.290847e-08,
  1.172425e-06, 1.372752e-06, 4.790247e-06, 5.293353e-06, 4.264097e-06, 
    7.004187e-06, 3.287812e-06, 1.458792e-06, 2.423199e-08, 7.810885e-09, 
    9.981283e-09, 5.42747e-08, 1.383349e-07, 9.136512e-08, 2.622409e-08,
  2.766484e-07, 1.12501e-07, 1.400562e-07, 5.609401e-07, 5.253148e-07, 
    3.175254e-08, 4.680981e-07, 2.703927e-09, 1.193868e-07, 4.844005e-09, 
    7.898993e-08, 4.863083e-08, 5.534336e-08, 5.403278e-08, 3.612809e-08,
  0.0002758583, 0.0001817796, 0.0001990645, 0.0001274806, 6.853975e-05, 
    2.848475e-05, 1.428953e-05, 1.37262e-06, 4.022677e-06, 4.546538e-06, 
    4.767962e-06, 4.667934e-06, 4.640938e-06, 1.548484e-05, 6.072283e-06,
  0.0002488232, 0.0002540901, 0.0002062035, 0.0001585769, 0.0001249307, 
    7.2349e-05, 3.208993e-05, 9.36075e-06, 1.152162e-05, 1.332476e-05, 
    1.293455e-05, 1.113119e-05, 7.513579e-06, 6.639226e-06, 4.386662e-06,
  0.0002630636, 0.000292786, 0.000197235, 0.0001462278, 0.0001198546, 
    7.315796e-05, 2.559881e-05, 1.453925e-05, 2.764082e-05, 2.403151e-05, 
    2.609682e-05, 2.193078e-05, 2.3245e-05, 1.960801e-05, 1.063084e-05,
  0.0002770225, 0.0001139954, 0.0001319655, 0.0001335654, 8.071381e-05, 
    5.028533e-05, 3.131322e-05, 2.344046e-05, 3.068912e-05, 3.875018e-05, 
    4.356181e-05, 3.464006e-05, 3.236379e-05, 2.677026e-05, 2.997974e-05,
  0.0002411535, 0.0001065128, 5.794725e-05, 5.562594e-05, 3.403533e-05, 
    2.024456e-05, 2.407358e-05, 1.886882e-05, 2.854043e-05, 2.669048e-05, 
    9.58031e-07, 5.136283e-07, 1.14508e-05, 2.541822e-06, 1.874527e-05,
  0.0002211133, 0.0001682652, 9.537629e-05, 7.327845e-05, 5.135403e-05, 
    2.403079e-05, 1.641268e-05, 9.009796e-06, 1.289667e-05, 3.050622e-06, 
    2.271891e-05, 1.460883e-06, 6.807898e-08, 9.00187e-07, 1.16845e-05,
  0.0002135311, 0.0002321911, 0.0001976972, 0.0001346672, 6.480281e-05, 
    2.365527e-05, 1.683234e-05, 1.570011e-05, 3.871941e-05, 1.205335e-05, 
    3.11037e-08, 1.83324e-08, 2.037655e-08, 1.613599e-06, 1.487954e-06,
  0.0002673778, 0.0002877809, 0.0002629417, 0.0001591151, 5.536868e-05, 
    2.235424e-05, 2.320798e-05, 2.976754e-05, 4.091288e-05, 3.779298e-06, 
    1.420955e-06, 2.431643e-06, 6.919318e-07, 7.951052e-06, 1.453864e-06,
  0.0001883088, 0.0001887736, 0.0001703734, 9.378969e-05, 2.876849e-05, 
    2.279646e-05, 2.597663e-05, 5.325496e-05, 2.742392e-05, 4.204663e-06, 
    1.681639e-06, 3.706138e-06, 1.958024e-06, 3.666029e-06, 8.166812e-06,
  1.595894e-05, 2.969732e-05, 4.2736e-05, 2.657764e-05, 2.452551e-05, 
    1.450485e-05, 4.074426e-05, 2.76495e-05, 1.264152e-05, 3.733201e-06, 
    1.484701e-06, 1.150229e-06, 1.366445e-06, 3.144899e-06, 4.283124e-06,
  0.0001580896, 0.0001446341, 0.000139832, 0.0001263386, 6.572568e-05, 
    6.727335e-05, 6.789653e-05, 3.233585e-05, 4.158889e-05, 2.294564e-05, 
    1.11672e-05, 5.302816e-06, 1.404253e-06, 1.948339e-06, 1.349198e-06,
  9.168194e-05, 0.0001304627, 0.0001719458, 0.0001487569, 0.000133088, 
    0.0001270992, 0.0001123083, 8.600006e-05, 6.921968e-05, 2.858274e-05, 
    1.480875e-05, 1.251393e-05, 8.641584e-06, 3.106403e-06, 5.502862e-06,
  0.0001601626, 5.73594e-05, 7.110197e-05, 0.0001049262, 0.0001488138, 
    0.0001098386, 9.237964e-05, 0.000121287, 9.139054e-05, 3.452644e-05, 
    2.317538e-05, 2.418393e-05, 2.426392e-05, 1.517429e-05, 1.888602e-05,
  8.774066e-05, 4.846196e-05, 3.720532e-05, 7.243848e-05, 9.224112e-05, 
    9.989122e-05, 0.0001379268, 0.0001587314, 0.0001210225, 5.425913e-05, 
    4.534389e-05, 3.83271e-05, 4.153145e-05, 3.678527e-05, 3.599451e-05,
  4.99113e-05, 2.382611e-05, 2.972519e-05, 4.91038e-05, 6.882983e-05, 
    9.876501e-05, 0.0001335228, 0.0001566352, 0.0001270822, 0.0001109947, 
    6.568082e-05, 6.615937e-05, 8.486742e-05, 1.565716e-05, 4.357942e-05,
  5.059686e-06, 1.50067e-05, 2.191074e-05, 4.691071e-05, 8.436893e-05, 
    7.548741e-05, 8.161206e-05, 9.079879e-05, 0.0001485673, 0.0001749011, 
    0.0001623515, 0.0001094026, 5.410825e-05, 4.610282e-05, 4.872768e-05,
  6.853057e-06, 1.578742e-05, 2.936335e-05, 6.997911e-05, 7.40979e-05, 
    4.157317e-05, 4.507187e-05, 6.671258e-05, 9.999184e-05, 5.305207e-05, 
    3.125069e-05, 4.670041e-05, 4.469539e-05, 7.226413e-05, 4.684541e-05,
  1.229517e-05, 2.276057e-05, 5.883106e-05, 6.514577e-05, 3.755568e-05, 
    2.112698e-05, 2.345212e-05, 2.712931e-05, 4.336293e-05, 2.21225e-05, 
    1.500478e-05, 1.744588e-05, 1.770496e-05, 5.541712e-05, 2.304144e-05,
  2.278544e-06, 3.974596e-06, 2.038378e-05, 2.390267e-05, 1.455386e-05, 
    1.602538e-05, 2.427756e-05, 4.369243e-05, 2.553162e-05, 1.044188e-05, 
    4.06031e-06, 1.214063e-06, 1.246127e-07, 9.475531e-06, 1.21683e-05,
  3.497351e-07, 7.186016e-06, 2.327704e-05, 3.407285e-05, 3.971303e-05, 
    3.2119e-05, 3.702318e-05, 2.274879e-05, 1.378539e-05, 9.335949e-06, 
    4.175241e-06, 2.707553e-06, 1.305508e-06, 1.295352e-06, 1.603156e-06,
  4.629272e-05, 4.491301e-05, 3.412442e-05, 3.465754e-05, 3.077784e-05, 
    4.281172e-05, 5.994214e-05, 5.885899e-05, 0.0001249154, 9.847814e-05, 
    4.095869e-05, 2.930808e-05, 1.501115e-05, 1.156442e-05, 4.092244e-07,
  6.507178e-06, 1.611859e-05, 1.359407e-05, 2.010836e-05, 1.425113e-05, 
    2.320473e-05, 4.815156e-05, 6.556635e-05, 0.0001561698, 0.0001096803, 
    6.651683e-05, 5.530278e-05, 4.956318e-05, 2.898936e-05, 1.317962e-06,
  1.149381e-07, 1.370855e-07, 3.413503e-07, 1.614374e-07, 6.830975e-06, 
    1.408799e-05, 1.605835e-05, 6.059029e-05, 0.0001423227, 0.0001209891, 
    0.0001095441, 0.0001065662, 0.000107137, 8.310902e-05, 4.590191e-05,
  8.660975e-08, 6.068684e-07, 6.168744e-07, 1.015154e-05, 1.221601e-05, 
    1.307108e-05, 1.507498e-05, 3.740116e-05, 8.396432e-05, 9.612403e-05, 
    0.000144454, 0.0001511787, 0.0001097399, 8.503306e-05, 3.973123e-05,
  2.443565e-08, 1.145124e-06, 4.964905e-06, 1.155163e-05, 1.188234e-05, 
    1.382129e-05, 1.986219e-05, 3.359457e-05, 5.928832e-05, 0.00015086, 
    0.0001951245, 0.0001373053, 0.0001148497, 3.395243e-05, 2.616842e-05,
  7.085421e-08, 2.234494e-06, 3.572018e-06, 8.523787e-06, 9.067891e-06, 
    1.476151e-05, 1.870181e-05, 2.872872e-05, 7.44893e-05, 8.290871e-05, 
    6.246552e-05, 5.228211e-05, 4.271593e-05, 3.789205e-05, 3.965406e-05,
  1.005534e-06, 1.353315e-06, 4.60721e-06, 5.574841e-06, 9.38512e-06, 
    1.117551e-05, 2.375487e-05, 3.153232e-05, 3.049663e-05, 1.832963e-05, 
    1.526194e-05, 3.173284e-05, 2.363322e-05, 6.444289e-05, 5.303323e-05,
  1.298604e-07, 1.105812e-06, 4.508699e-06, 7.660784e-06, 9.323132e-06, 
    6.823606e-06, 1.63672e-05, 1.985541e-05, 3.247555e-05, 1.601519e-05, 
    3.283396e-05, 5.189485e-05, 3.042218e-05, 6.030205e-05, 1.356521e-05,
  3.442032e-07, 3.109112e-06, 1.122401e-05, 1.970969e-05, 2.977067e-05, 
    3.648398e-05, 3.240971e-05, 2.633829e-05, 1.471884e-05, 2.814515e-05, 
    3.595766e-05, 4.091675e-05, 3.517957e-05, 3.88628e-05, 1.146065e-05,
  2.718207e-07, 8.818338e-06, 2.34583e-05, 3.086874e-05, 5.200321e-05, 
    6.755025e-05, 5.752038e-05, 1.434399e-05, 3.467898e-05, 4.92003e-05, 
    4.113486e-05, 3.385366e-05, 3.040264e-05, 1.093599e-05, 3.638013e-06,
  2.178123e-05, 1.923545e-05, 1.051345e-07, 5.282883e-07, 1.680174e-07, 
    4.583726e-07, 5.157058e-06, 7.238161e-06, 2.039194e-05, 2.768508e-05, 
    2.153056e-05, 1.773199e-05, 1.844742e-05, 2.416035e-05, 1.210914e-05,
  2.02798e-06, 3.623363e-06, 2.728153e-07, 1.491994e-06, 2.014003e-06, 
    2.096726e-06, 6.238989e-06, 8.018328e-06, 9.710511e-06, 1.099942e-05, 
    1.2728e-05, 1.242487e-05, 1.640607e-05, 1.530942e-05, 1.371463e-05,
  1.045262e-06, 6.255897e-06, 5.454272e-06, 1.765128e-06, 4.982161e-06, 
    5.178749e-06, 6.950395e-06, 1.161724e-05, 1.886235e-05, 1.959565e-05, 
    1.989829e-05, 1.569463e-05, 1.104105e-05, 1.182224e-05, 7.288724e-06,
  4.238957e-07, 7.008824e-06, 1.389009e-05, 2.235459e-05, 2.726044e-05, 
    3.332368e-05, 2.604901e-05, 2.545157e-05, 2.704389e-05, 3.028473e-05, 
    6.74213e-05, 6.113144e-05, 3.341115e-05, 2.014339e-05, 4.916251e-06,
  6.65991e-06, 6.965331e-06, 1.276566e-05, 3.012942e-05, 2.313828e-05, 
    3.67592e-05, 3.774603e-05, 4.131603e-05, 4.897447e-05, 3.560058e-05, 
    6.678148e-06, 3.875639e-05, 0.0001070662, 1.451409e-05, 7.183911e-06,
  7.602173e-06, 1.210986e-05, 1.947277e-05, 2.300059e-05, 2.734425e-05, 
    3.954172e-05, 5.049752e-05, 4.628019e-05, 4.256527e-05, 4.320387e-06, 
    3.156109e-05, 0.0001029453, 6.84575e-05, 5.015199e-05, 2.282474e-05,
  1.446307e-05, 1.345712e-05, 1.834514e-05, 2.257683e-05, 3.49265e-05, 
    1.674852e-05, 3.130616e-05, 2.893058e-05, 2.445965e-05, 1.379553e-05, 
    5.912774e-05, 9.871962e-05, 0.000104667, 0.0001586119, 1.931847e-05,
  2.223675e-05, 2.019811e-05, 2.119715e-05, 2.47835e-05, 1.787844e-05, 
    2.623745e-05, 2.956982e-05, 3.820384e-05, 5.780162e-05, 3.218716e-05, 
    7.485577e-05, 7.183715e-05, 0.0001147066, 0.0001945667, 1.0775e-05,
  2.254119e-05, 2.789151e-05, 3.731362e-05, 5.535766e-05, 8.895529e-05, 
    0.0001200203, 0.0001147564, 0.0001565212, 2.026243e-05, 9.989646e-05, 
    5.929561e-05, 4.421484e-05, 0.0001036089, 0.0001357763, 1.574342e-05,
  7.972569e-06, 2.568427e-05, 4.745992e-05, 5.448575e-05, 7.33889e-05, 
    0.0001177372, 0.0001363015, 3.316597e-05, 9.85588e-05, 0.0001118593, 
    5.442203e-05, 3.553559e-05, 6.075768e-05, 6.743721e-05, 3.08465e-05,
  6.685286e-09, 4.618533e-09, 3.770551e-10, 2.220433e-08, 1.276885e-08, 
    1.112704e-08, 3.36904e-08, 2.382906e-06, 1.56412e-05, 3.273458e-05, 
    2.943049e-05, 2.951464e-05, 2.084198e-05, 1.067432e-05, 2.803604e-06,
  1.902637e-28, 4.673429e-27, 5.526592e-12, 3.630657e-11, 2.671182e-10, 
    1.03983e-09, 2.710545e-09, 9.976004e-08, 4.054677e-06, 1.277099e-05, 
    1.637099e-05, 1.651163e-05, 1.345013e-05, 1.16381e-05, 1.004123e-06,
  5.048367e-28, 7.251031e-13, 4.058095e-10, 2.527671e-09, 1.800226e-08, 
    1.056353e-07, 1.452547e-07, 1.422738e-07, 4.624087e-07, 8.002895e-06, 
    2.722112e-05, 3.058117e-05, 1.452021e-05, 2.185785e-05, 4.613406e-07,
  4.32988e-27, 2.510752e-11, 6.144067e-09, 2.441943e-07, 2.314111e-07, 
    1.014151e-06, 4.597503e-06, 4.921821e-06, 8.579228e-06, 2.505746e-05, 
    7.6512e-05, 0.0001157459, 6.918984e-05, 3.838281e-05, 4.972468e-06,
  1.383143e-11, 2.60969e-10, 1.959215e-08, 1.566239e-06, 2.723519e-06, 
    6.704474e-06, 7.602197e-06, 1.6536e-05, 2.365411e-05, 4.226416e-05, 
    6.068732e-06, 8.215938e-05, 0.0002508896, 6.715877e-05, 9.711176e-05,
  1.004561e-10, 2.024004e-09, 8.807815e-08, 3.343949e-06, 4.597384e-06, 
    6.282419e-06, 9.271906e-06, 1.969825e-05, 1.917679e-05, 1.183211e-06, 
    3.115037e-05, 7.463287e-05, 0.0001133639, 0.0001817198, 9.812137e-05,
  2.509705e-11, 3.549646e-09, 1.91311e-07, 2.460306e-06, 2.61695e-06, 
    2.204561e-06, 6.920413e-06, 1.523669e-05, 1.442996e-05, 2.718216e-05, 
    3.615879e-05, 3.494109e-05, 6.70228e-05, 0.0002016771, 0.0001058438,
  7.579558e-11, 1.584116e-09, 7.701277e-07, 2.579068e-07, 9.255038e-07, 
    1.367153e-06, 3.526853e-06, 1.498608e-05, 4.515753e-05, 3.148693e-05, 
    3.816573e-05, 2.224193e-05, 3.425068e-05, 0.0001398648, 6.253946e-05,
  1.781865e-10, 4.240562e-11, 1.945049e-09, 2.090847e-08, 4.274179e-07, 
    3.965977e-06, 1.698795e-05, 2.888036e-05, 1.668226e-05, 5.756526e-05, 
    5.168676e-05, 4.030059e-05, 4.2595e-05, 7.303791e-05, 2.487998e-05,
  5.228074e-09, 1.787861e-10, 4.815173e-10, 2.243896e-08, 2.08248e-07, 
    1.156929e-06, 6.115202e-06, 7.99702e-06, 3.798732e-05, 4.733707e-05, 
    3.543021e-05, 2.865421e-05, 3.094257e-05, 2.04425e-05, 6.551704e-06,
  1.288347e-11, 1.10175e-10, 3.506018e-10, 1.479285e-09, 2.646249e-09, 
    4.355063e-09, 4.80327e-08, 1.51111e-08, 4.505758e-09, 9.296978e-08, 
    9.791642e-07, 1.459332e-06, 1.548898e-07, 3.907583e-07, 5.469862e-08,
  3.384467e-09, 4.765439e-10, 9.471889e-10, 4.39203e-09, 6.697479e-09, 
    2.229978e-08, 2.169299e-07, 1.838749e-07, 1.401171e-07, 4.464583e-07, 
    1.554785e-06, 1.554208e-06, 3.463582e-07, 7.054841e-07, 3.281536e-07,
  1.11062e-07, 2.97839e-06, 1.466223e-07, 1.530834e-08, 8.681027e-08, 
    7.961932e-08, 2.541275e-07, 6.766362e-07, 1.493781e-06, 1.749585e-06, 
    3.228345e-06, 4.873021e-06, 2.202976e-06, 2.340475e-06, 2.784599e-07,
  6.315888e-06, 1.629201e-06, 9.616419e-07, 2.830237e-06, 1.700626e-06, 
    8.472001e-07, 1.326408e-06, 4.00424e-06, 1.317027e-05, 2.095259e-05, 
    5.2958e-06, 4.092068e-06, 1.725334e-06, 5.411107e-06, 2.232058e-06,
  2.045646e-05, 5.037679e-06, 1.561565e-07, 1.429739e-07, 1.251337e-07, 
    4.889781e-08, 3.955476e-07, 5.661785e-06, 1.632171e-05, 3.001976e-05, 
    5.162725e-09, 1.853233e-07, 1.639957e-06, 1.788324e-06, 5.237175e-06,
  9.977944e-06, 1.521351e-06, 5.716174e-08, 3.748347e-09, 1.690953e-08, 
    4.379116e-08, 1.210827e-07, 6.648063e-07, 5.412301e-06, 2.333163e-06, 
    6.963339e-06, 2.606474e-06, 9.538275e-08, 7.670223e-06, 7.952794e-06,
  1.02574e-06, 2.089848e-07, 1.551256e-08, 3.739125e-09, 1.534614e-08, 
    4.203347e-08, 3.124947e-08, 4.150042e-08, 1.594273e-08, 3.112666e-06, 
    1.837763e-05, 1.585188e-05, 3.509168e-06, 4.96156e-05, 8.53967e-06,
  6.090817e-07, 5.57828e-06, 4.655844e-07, 1.392247e-08, 1.70469e-08, 
    2.311927e-08, 7.686155e-09, 3.488439e-09, 1.262805e-09, 1.126015e-08, 
    8.122608e-06, 2.226614e-05, 5.259354e-05, 7.129126e-05, 1.25434e-06,
  2.116882e-05, 2.094446e-05, 6.328177e-06, 1.723066e-07, 4.939077e-07, 
    1.698305e-06, 2.06809e-07, 1.306749e-07, 2.019389e-09, 9.795323e-09, 
    2.094716e-07, 5.555644e-06, 3.78705e-05, 4.640371e-05, 2.201847e-07,
  5.389837e-05, 5.783401e-05, 1.941482e-05, 9.224904e-07, 3.96527e-07, 
    1.373385e-06, 5.023022e-07, 2.925304e-07, 1.878294e-07, 1.234078e-07, 
    5.473846e-07, 1.043172e-06, 5.936484e-06, 1.434397e-05, 5.573302e-06,
  3.933339e-08, 4.312063e-07, 2.187938e-09, 4.261702e-09, 7.226225e-08, 
    2.632904e-07, 9.924779e-07, 1.850409e-08, 1.085038e-07, 1.673265e-06, 
    2.304054e-06, 2.199615e-07, 1.163671e-07, 2.093019e-06, 1.706885e-08,
  2.801362e-06, 2.599673e-06, 9.206085e-07, 5.472162e-07, 6.755403e-07, 
    1.575125e-06, 6.367941e-06, 3.319881e-06, 4.87863e-06, 6.165136e-06, 
    4.017568e-06, 1.051657e-06, 1.779408e-07, 7.887209e-07, 6.296861e-08,
  5.930449e-05, 5.664193e-05, 1.309933e-05, 1.112244e-05, 1.896438e-05, 
    9.581292e-06, 2.879019e-06, 6.213915e-06, 1.453768e-05, 5.456655e-06, 
    2.603691e-06, 9.471401e-07, 2.512788e-07, 2.087094e-07, 3.229971e-07,
  0.0002844668, 4.461674e-05, 1.633074e-05, 3.424065e-05, 1.928978e-05, 
    1.19419e-05, 7.949732e-06, 9.203975e-06, 5.899225e-06, 9.075264e-07, 
    3.090751e-07, 4.631296e-07, 3.390284e-07, 2.499644e-07, 7.044137e-07,
  0.0003182657, 8.224725e-05, 1.041406e-05, 9.507931e-06, 8.978209e-06, 
    1.156082e-05, 1.288255e-05, 9.196475e-06, 2.428762e-06, 1.013151e-06, 
    4.307334e-10, 9.575924e-10, 3.447657e-08, 7.395157e-09, 9.940769e-07,
  0.0001668372, 0.0001080278, 1.647294e-05, 2.950906e-05, 4.643018e-05, 
    4.19235e-05, 2.84347e-05, 1.308252e-05, 6.677801e-06, 2.583333e-07, 
    9.90247e-08, 6.433703e-09, 1.004833e-08, 2.190841e-08, 3.246517e-06,
  6.945173e-05, 7.60406e-05, 4.430371e-05, 5.810881e-05, 9.354451e-05, 
    7.640903e-05, 4.0047e-05, 1.535105e-06, 1.415656e-07, 9.246797e-07, 
    1.116784e-06, 5.875279e-07, 2.300154e-08, 1.140685e-06, 1.260578e-06,
  4.42057e-05, 8.830641e-05, 4.838318e-05, 3.83096e-05, 5.033912e-05, 
    6.232626e-05, 2.601995e-05, 1.666648e-05, 3.67415e-06, 7.604141e-06, 
    1.75718e-05, 1.189299e-05, 4.738528e-07, 3.425578e-05, 1.303453e-06,
  7.822722e-05, 9.789765e-05, 5.594021e-05, 4.732706e-05, 6.579357e-05, 
    8.028543e-05, 3.320738e-05, 1.481179e-05, 6.598407e-06, 3.465015e-05, 
    2.323215e-05, 2.860123e-05, 1.533498e-05, 2.802013e-05, 3.448888e-08,
  8.364362e-05, 8.093204e-05, 7.26749e-05, 5.756156e-05, 6.63651e-05, 
    5.989185e-05, 5.17148e-05, 1.583386e-05, 3.166042e-05, 2.557545e-05, 
    1.021032e-05, 5.253117e-06, 1.398526e-05, 2.191044e-05, 5.335624e-06,
  0.0001205748, 1.350194e-05, 4.891613e-06, 1.531728e-07, 6.921351e-08, 
    3.560993e-08, 4.517674e-07, 2.586708e-07, 2.382226e-06, 3.898546e-06, 
    2.369809e-06, 1.745536e-06, 5.265492e-08, 1.844201e-08, 2.573967e-08,
  3.827058e-05, 3.711123e-05, 7.342384e-06, 5.147479e-06, 3.420361e-07, 
    4.761538e-07, 8.041697e-06, 4.530839e-06, 6.768622e-06, 3.215023e-06, 
    1.234876e-06, 1.73091e-06, 6.096091e-08, 3.232422e-08, 4.490061e-08,
  0.0001505776, 0.0001682935, 4.140808e-05, 1.839803e-05, 9.78179e-06, 
    2.611358e-06, 3.218838e-06, 8.01437e-06, 1.197108e-05, 3.908234e-06, 
    1.627717e-06, 1.036537e-06, 1.981064e-07, 9.810584e-08, 4.12169e-08,
  0.0001983542, 6.244642e-05, 5.730761e-05, 7.289877e-05, 2.007855e-05, 
    6.310625e-06, 4.571984e-06, 1.0134e-05, 5.883959e-06, 2.517771e-06, 
    2.250198e-07, 3.347463e-07, 4.778805e-07, 3.333548e-07, 2.02178e-07,
  0.0001718949, 3.47596e-05, 8.786707e-06, 7.939249e-06, 3.535421e-06, 
    1.645434e-06, 2.194164e-06, 5.882634e-06, 9.258245e-06, 3.773638e-06, 
    3.763699e-08, 2.196366e-09, 1.370346e-07, 4.09174e-08, 1.436456e-07,
  9.500521e-05, 4.113086e-05, 1.258774e-05, 6.38669e-06, 5.635234e-06, 
    2.765853e-06, 2.309392e-06, 1.763589e-06, 4.029104e-06, 3.418985e-06, 
    5.026245e-06, 6.14865e-08, 5.559553e-09, 6.087504e-09, 2.728633e-07,
  3.36451e-05, 2.384951e-05, 1.301708e-05, 1.09846e-05, 2.137345e-05, 
    9.309722e-06, 2.789002e-06, 1.350942e-06, 3.400483e-08, 3.132267e-06, 
    1.289823e-05, 2.619107e-06, 4.066748e-08, 2.509123e-06, 1.90623e-06,
  1.629575e-05, 3.134158e-05, 1.715292e-05, 7.932092e-06, 1.43126e-05, 
    1.590541e-05, 1.207662e-05, 8.157284e-06, 1.880285e-07, 2.590027e-08, 
    4.405836e-08, 1.294439e-06, 1.09045e-07, 5.472947e-05, 1.822828e-06,
  0.0001000427, 4.920203e-05, 2.594962e-05, 5.754776e-06, 8.876043e-06, 
    1.195305e-05, 6.54575e-06, 1.715547e-06, 8.96144e-08, 1.259484e-07, 
    8.648863e-08, 9.279731e-07, 2.483222e-06, 1.565213e-05, 5.153617e-08,
  0.0001767922, 0.0001109501, 9.495865e-06, 9.788355e-07, 3.277484e-06, 
    1.972666e-06, 1.380415e-06, 1.876705e-07, 5.204653e-07, 3.448636e-07, 
    3.590855e-08, 2.635351e-09, 1.258369e-07, 2.958606e-06, 9.20955e-08,
  0.0003097159, 5.099682e-05, 2.055932e-05, 1.530083e-07, 6.894366e-08, 
    1.150714e-07, 4.112932e-07, 2.665244e-07, 6.972415e-07, 7.556295e-07, 
    7.650851e-07, 2.092342e-07, 2.567352e-08, 1.931177e-09, 2.746136e-07,
  0.0003442422, 0.0002679533, 2.772067e-05, 2.425012e-05, 4.728648e-06, 
    2.354629e-06, 1.49672e-06, 7.010992e-07, 1.113982e-06, 2.480753e-06, 
    2.653096e-06, 8.268936e-07, 2.878007e-08, 2.344111e-09, 4.47189e-08,
  0.0004840132, 0.0004142165, 0.0001631987, 4.950365e-05, 4.261558e-05, 
    6.417092e-06, 1.702414e-06, 1.458732e-06, 1.724014e-06, 2.041738e-06, 
    2.811363e-06, 3.588212e-07, 4.556609e-08, 4.562378e-09, 1.305632e-07,
  0.0005313223, 0.0001829379, 0.0001431915, 9.359157e-05, 3.759086e-05, 
    1.538632e-05, 6.76131e-06, 3.062012e-06, 8.106128e-07, 6.111492e-07, 
    3.358533e-07, 8.725584e-08, 1.353715e-08, 3.855599e-09, 1.677272e-07,
  0.0005673215, 0.0001208359, 1.481655e-05, 1.144709e-05, 9.109138e-06, 
    1.004106e-05, 9.042197e-06, 2.419334e-06, 2.317259e-07, 7.418256e-07, 
    4.395313e-10, 2.396323e-10, 6.789347e-10, 1.073555e-09, 2.978221e-07,
  0.0004536888, 0.0001554778, 6.68107e-06, 6.146019e-06, 1.852462e-05, 
    1.121186e-05, 5.837422e-06, 9.706944e-07, 4.492079e-08, 3.031407e-10, 
    7.083265e-09, 1.869467e-09, 4.764294e-10, 3.727123e-09, 5.398495e-07,
  0.0002012939, 0.0001295399, 2.985995e-05, 3.644941e-05, 6.356387e-05, 
    3.733892e-05, 2.139467e-05, 9.12829e-07, 7.706997e-09, 3.490067e-09, 
    2.803482e-08, 1.277128e-08, 1.625823e-09, 7.63507e-09, 9.072188e-09,
  0.0001055165, 0.0001207333, 0.0001026104, 0.0001236166, 0.0001838418, 
    0.0001422401, 5.091392e-05, 8.188263e-06, 5.681219e-07, 8.576126e-09, 
    2.663695e-08, 1.579616e-08, 6.520781e-09, 3.709371e-08, 1.438896e-10,
  0.0002075069, 0.0001142097, 9.727795e-05, 0.0001290675, 0.0001755376, 
    0.0001924455, 6.092864e-05, 6.855399e-06, 7.361375e-09, 5.147664e-09, 
    1.711897e-09, 1.868385e-09, 3.10618e-09, 1.254742e-09, 1.216055e-10,
  0.0001256262, 0.000155229, 0.0001076034, 9.40017e-05, 0.0001276459, 
    6.147575e-05, 2.261105e-05, 7.754516e-06, 6.5476e-06, 1.950983e-07, 
    6.649986e-09, 4.31648e-09, 3.893766e-09, 1.764582e-09, 3.842589e-10,
  0.0001664286, 4.455891e-05, 5.290714e-05, 3.522032e-05, 8.957369e-06, 
    1.351236e-05, 2.101366e-05, 4.894564e-06, 7.594683e-06, 2.187437e-06, 
    1.207725e-06, 1.255795e-06, 1.700606e-06, 9.831999e-06, 4.019405e-05,
  0.0001027105, 4.333933e-05, 7.56271e-06, 4.39026e-06, 1.220904e-05, 
    1.924146e-05, 2.073207e-05, 1.070168e-05, 5.863199e-06, 2.049145e-06, 
    1.492506e-06, 1.145501e-06, 1.028046e-06, 2.181663e-06, 2.03669e-06,
  0.0001424596, 0.0001421035, 3.126105e-05, 4.050779e-06, 1.286433e-05, 
    1.567416e-05, 8.104491e-06, 7.354415e-06, 9.14737e-06, 3.978478e-06, 
    1.701851e-06, 4.374747e-07, 1.059786e-06, 2.926031e-06, 1.60942e-06,
  0.000138335, 2.811924e-05, 1.725884e-05, 1.636458e-05, 8.640626e-06, 
    1.005903e-05, 1.222856e-05, 1.019349e-05, 7.382152e-06, 1.179628e-06, 
    3.353854e-06, 2.300599e-06, 1.299609e-06, 2.005599e-06, 1.073027e-05,
  9.726761e-05, 2.420028e-05, 3.588149e-06, 2.280203e-06, 6.226187e-06, 
    1.502747e-05, 1.282063e-05, 6.659472e-06, 3.061933e-06, 6.076169e-06, 
    1.441298e-08, 9.370742e-09, 2.227602e-07, 1.668898e-07, 8.332528e-06,
  5.045941e-05, 4.542169e-05, 1.69248e-05, 1.230122e-05, 4.323048e-05, 
    6.375711e-05, 3.152419e-05, 8.900637e-06, 8.318166e-06, 2.915173e-08, 
    2.566152e-09, 1.883336e-09, 3.273996e-08, 1.220436e-07, 7.692418e-06,
  2.828381e-05, 3.875556e-05, 3.317734e-05, 3.831951e-05, 7.440306e-05, 
    0.0001097898, 8.381496e-05, 1.007306e-05, 1.65948e-06, 3.4316e-07, 
    2.510692e-09, 6.040502e-09, 2.182463e-08, 1.795313e-07, 3.436266e-07,
  9.985318e-06, 1.831724e-05, 2.158274e-05, 3.52829e-05, 8.264217e-05, 
    0.0001024604, 7.217875e-05, 2.710444e-05, 2.896508e-06, 4.570386e-07, 
    2.433569e-08, 3.53699e-09, 1.29733e-08, 1.486285e-07, 3.528297e-08,
  6.235083e-06, 1.031555e-05, 7.536656e-06, 1.623216e-05, 4.628095e-05, 
    4.897964e-05, 3.412542e-05, 1.609631e-05, 1.539946e-06, 1.836768e-06, 
    2.092639e-08, 3.703671e-09, 4.851741e-09, 6.320837e-09, 1.068511e-09,
  9.576762e-06, 1.014333e-05, 7.945074e-06, 1.039293e-05, 2.545505e-05, 
    3.15636e-05, 2.694863e-05, 1.051183e-05, 2.084856e-05, 7.41819e-06, 
    6.204714e-07, 1.404657e-08, 1.533946e-09, 1.651667e-09, 3.520137e-10,
  1.35956e-05, 6.858083e-06, 2.630314e-05, 2.422333e-05, 2.467919e-06, 
    3.97366e-07, 1.563126e-06, 1.384212e-07, 6.946217e-06, 5.711277e-06, 
    2.81266e-06, 3.467376e-06, 7.872217e-06, 1.778008e-05, 1.981838e-05,
  1.099632e-05, 4.392154e-05, 2.048262e-05, 1.485654e-05, 5.202454e-06, 
    4.807618e-07, 4.195739e-06, 6.713042e-07, 5.183147e-06, 8.584728e-06, 
    5.097912e-06, 1.984363e-06, 1.686316e-06, 2.870586e-06, 2.493246e-06,
  5.869681e-05, 3.098296e-05, 2.50358e-05, 1.269802e-05, 6.835036e-06, 
    2.812603e-06, 4.662858e-06, 3.039405e-06, 2.716146e-06, 7.302544e-06, 
    8.606322e-06, 4.242541e-06, 2.065826e-06, 1.430012e-05, 3.703353e-06,
  4.680518e-05, 1.488666e-05, 1.293946e-05, 1.833846e-05, 1.461939e-05, 
    9.362014e-06, 1.395611e-05, 1.199984e-05, 9.664121e-06, 1.190465e-05, 
    3.5202e-05, 1.12907e-05, 2.278486e-06, 6.535507e-06, 2.623567e-05,
  3.773295e-05, 1.851952e-05, 9.830822e-06, 1.166838e-05, 6.416362e-06, 
    2.616166e-05, 2.912259e-05, 3.759782e-05, 2.867073e-05, 3.245619e-05, 
    9.791815e-06, 1.660281e-05, 1.262606e-05, 2.166899e-06, 1.763686e-05,
  6.823052e-06, 1.095473e-05, 5.080797e-06, 1.358144e-05, 1.509092e-05, 
    1.365847e-05, 1.893455e-05, 2.357848e-05, 4.420558e-05, 4.052381e-06, 
    4.014208e-05, 4.316143e-05, 2.30219e-06, 1.875201e-07, 1.247003e-05,
  5.057891e-06, 7.893705e-06, 1.191013e-05, 1.826442e-05, 3.233059e-05, 
    1.802312e-05, 2.049927e-05, 2.641338e-05, 2.152536e-05, 1.774716e-05, 
    6.974747e-06, 1.286707e-05, 1.136039e-06, 8.957047e-07, 2.419946e-06,
  4.98688e-06, 1.496395e-05, 1.901242e-05, 2.194442e-05, 1.91259e-05, 
    1.393587e-05, 1.345077e-05, 3.24773e-05, 2.271907e-05, 1.699611e-05, 
    8.568074e-06, 7.112576e-06, 7.096086e-07, 1.317754e-06, 5.820319e-07,
  1.155969e-05, 2.424773e-05, 2.430484e-05, 2.080337e-05, 1.786042e-05, 
    1.70744e-05, 2.793918e-05, 2.053147e-05, 2.990015e-05, 3.033518e-05, 
    1.367652e-05, 8.494681e-06, 3.80678e-06, 3.052342e-06, 2.496962e-06,
  7.748961e-06, 2.639515e-05, 2.20618e-05, 9.77689e-06, 9.568835e-06, 
    5.81369e-06, 1.450993e-05, 2.870425e-05, 3.416296e-05, 1.789457e-05, 
    1.171306e-05, 1.257291e-05, 1.075454e-05, 9.876404e-06, 2.644397e-06,
  4.646753e-06, 4.553382e-06, 1.108467e-08, 9.326024e-09, 1.42518e-10, 
    1.951435e-11, 9.24241e-10, 8.817719e-09, 5.608911e-08, 6.172783e-07, 
    2.831781e-06, 6.321073e-06, 1.83369e-05, 2.582463e-05, 1.121961e-05,
  9.791976e-06, 4.890324e-06, 2.364379e-07, 2.161365e-07, 1.51198e-09, 
    2.309058e-10, 1.915444e-10, 3.93688e-10, 7.43863e-08, 2.677839e-07, 
    3.333208e-06, 1.199731e-05, 2.608412e-05, 2.365363e-05, 1.544954e-05,
  2.468794e-05, 4.576324e-07, 4.003365e-07, 9.162547e-08, 4.165767e-08, 
    1.16405e-08, 2.182163e-08, 5.416854e-09, 1.730656e-07, 1.978263e-06, 
    1.898703e-05, 2.894261e-05, 5.224794e-05, 5.718003e-05, 3.761239e-05,
  4.593674e-05, 2.309952e-06, 6.002567e-07, 2.570075e-06, 4.708252e-06, 
    1.336999e-06, 6.053638e-07, 2.181007e-07, 6.480636e-08, 6.108508e-06, 
    6.253587e-05, 6.377857e-05, 5.560937e-05, 4.852907e-05, 6.689892e-05,
  6.837356e-05, 1.044518e-05, 7.762941e-07, 1.061643e-06, 1.322908e-06, 
    1.260202e-06, 9.775881e-06, 4.097588e-06, 2.618954e-06, 2.348457e-06, 
    2.319625e-06, 3.094501e-05, 9.98043e-05, 2.7091e-05, 4.18489e-05,
  4.05893e-05, 1.05812e-05, 7.245175e-07, 1.453822e-07, 1.874138e-06, 
    1.448296e-06, 2.363156e-06, 1.117184e-06, 1.627228e-06, 2.48651e-07, 
    2.578334e-06, 2.389278e-05, 3.069241e-05, 5.181831e-06, 2.208881e-05,
  7.542728e-06, 4.672383e-06, 9.509826e-07, 1.401718e-06, 1.069335e-06, 
    8.357753e-07, 2.233601e-06, 1.47999e-06, 3.005622e-07, 5.313756e-07, 
    3.256993e-06, 4.536843e-06, 9.103463e-06, 1.465131e-05, 1.198458e-05,
  9.14329e-07, 4.926628e-06, 2.391369e-06, 1.001137e-06, 1.048043e-06, 
    7.281715e-07, 2.800488e-07, 6.535964e-07, 1.906899e-07, 1.139805e-06, 
    2.949639e-06, 1.12161e-06, 4.1015e-06, 2.679952e-05, 1.307009e-05,
  2.194084e-06, 8.645529e-06, 5.32964e-06, 8.924676e-07, 1.518854e-06, 
    2.355585e-06, 1.8191e-07, 5.803381e-09, 3.820963e-08, 2.194719e-07, 
    2.459833e-06, 1.949605e-06, 6.818801e-06, 1.127039e-05, 1.516237e-05,
  6.588244e-07, 9.76233e-06, 4.836181e-06, 7.640628e-07, 2.238307e-06, 
    4.698653e-08, 4.449958e-10, 1.161861e-10, 5.831109e-08, 3.758462e-07, 
    1.163843e-06, 5.051973e-06, 2.796493e-06, 1.017937e-05, 1.153584e-05,
  1.710601e-09, 2.191091e-10, 2.376781e-10, 1.343694e-09, 1.969075e-09, 
    6.370809e-10, 6.401859e-11, 1.093873e-10, 5.238921e-09, 3.578966e-08, 
    1.585083e-06, 1.241283e-05, 2.96135e-05, 2.984161e-05, 1.823551e-05,
  6.619334e-09, 9.905436e-09, 1.272635e-09, 1.607961e-09, 6.078869e-10, 
    6.343058e-10, 2.160899e-09, 7.76172e-10, 1.664153e-07, 4.994996e-08, 
    1.593451e-07, 6.083368e-06, 2.615373e-05, 2.337306e-05, 1.62205e-05,
  3.242887e-06, 1.872422e-06, 1.205355e-07, 2.184223e-07, 2.746111e-07, 
    3.114433e-07, 3.390678e-08, 4.290474e-07, 2.390925e-06, 1.155475e-06, 
    2.364458e-06, 1.99501e-06, 2.295159e-05, 3.247252e-05, 1.643273e-05,
  5.298226e-06, 1.588567e-06, 1.853708e-06, 4.755253e-06, 2.473482e-06, 
    3.831383e-06, 1.785765e-06, 3.434793e-06, 7.424217e-06, 8.963416e-06, 
    3.772388e-06, 7.738059e-07, 3.00016e-06, 1.25147e-05, 3.576863e-05,
  2.30755e-05, 4.155416e-07, 1.037676e-07, 3.68381e-07, 2.595688e-07, 
    1.105619e-06, 4.874337e-06, 3.031316e-06, 7.304086e-06, 2.081016e-06, 
    8.057378e-09, 6.663555e-10, 3.047159e-08, 3.664595e-06, 1.602682e-05,
  1.364032e-05, 4.742973e-06, 1.057593e-07, 2.079903e-06, 2.890611e-06, 
    2.346669e-06, 2.308858e-06, 2.090453e-06, 3.171587e-06, 1.108522e-09, 
    1.361435e-08, 2.092087e-09, 2.787058e-09, 2.713049e-06, 1.471238e-05,
  1.348731e-06, 6.896786e-07, 6.156399e-08, 8.001732e-08, 1.21642e-06, 
    3.15619e-06, 4.818214e-06, 1.424064e-06, 1.526269e-08, 1.14348e-07, 
    6.58412e-09, 9.129017e-09, 9.204121e-09, 8.231186e-07, 1.591242e-06,
  5.534585e-06, 3.693527e-06, 4.621967e-06, 7.840308e-07, 6.984359e-07, 
    2.054371e-06, 3.738674e-06, 4.261983e-06, 5.619156e-08, 3.277903e-07, 
    1.176312e-08, 4.585641e-11, 1.766291e-08, 8.966936e-07, 2.581485e-08,
  3.133409e-05, 4.105417e-05, 1.226119e-05, 8.1436e-06, 1.362636e-05, 
    9.623847e-06, 5.646777e-06, 7.788016e-06, 1.975834e-07, 2.972731e-07, 
    5.579398e-08, 1.37774e-11, 5.536352e-09, 1.068891e-06, 2.005412e-07,
  3.233728e-05, 6.311759e-05, 3.438073e-05, 9.517442e-06, 1.011404e-05, 
    6.189853e-06, 5.878052e-06, 1.421928e-07, 7.56037e-07, 7.513957e-07, 
    1.242772e-07, 4.05445e-10, 1.265062e-09, 6.289664e-08, 3.350536e-07,
  5.452736e-08, 5.785405e-08, 6.913466e-08, 8.097836e-08, 8.251374e-08, 
    1.913788e-07, 4.526656e-07, 1.400716e-07, 1.177189e-06, 6.259764e-06, 
    1.105838e-05, 4.944144e-06, 1.316966e-05, 2.199175e-05, 7.904947e-06,
  7.494101e-08, 5.649401e-08, 6.171438e-08, 7.925503e-08, 1.90985e-07, 
    1.415041e-06, 4.730206e-06, 4.490628e-06, 3.302095e-06, 7.676668e-06, 
    1.302226e-05, 9.444267e-06, 1.260096e-05, 1.515018e-05, 2.08611e-06,
  1.137991e-07, 1.13715e-06, 1.517306e-07, 3.757923e-08, 3.539491e-06, 
    4.170813e-06, 3.283193e-06, 5.283888e-06, 9.611829e-06, 1.588251e-05, 
    3.571099e-05, 2.092874e-05, 1.618688e-05, 1.625729e-05, 1.204333e-06,
  5.662495e-07, 7.489758e-08, 3.940925e-06, 1.432663e-05, 1.271046e-05, 
    1.038184e-05, 1.195538e-05, 6.356668e-06, 1.038522e-05, 2.594815e-05, 
    4.665384e-05, 2.156225e-05, 1.006657e-05, 8.912737e-06, 1.576251e-05,
  1.278627e-06, 3.05956e-08, 7.307256e-08, 3.539344e-07, 8.174224e-07, 
    2.042978e-06, 9.293317e-06, 9.636994e-06, 1.188386e-05, 1.280531e-05, 
    1.522969e-06, 6.117357e-08, 1.684094e-08, 4.894771e-07, 1.810029e-05,
  4.308554e-06, 4.686187e-07, 1.072448e-06, 2.20539e-06, 6.167936e-06, 
    5.750327e-06, 9.327163e-06, 6.036813e-06, 5.753783e-06, 4.378359e-07, 
    5.632442e-08, 1.145135e-08, 1.517595e-09, 1.678115e-07, 1.933456e-05,
  4.630103e-06, 4.862992e-06, 1.232254e-06, 8.732104e-07, 5.266741e-06, 
    6.964883e-06, 1.805053e-05, 5.899068e-06, 3.183664e-06, 8.987009e-07, 
    1.079046e-08, 5.267689e-09, 7.450629e-10, 4.274735e-08, 1.177744e-06,
  1.364164e-05, 1.284797e-05, 9.157527e-06, 4.801325e-06, 6.762457e-06, 
    1.295969e-05, 1.531322e-05, 1.922716e-05, 1.250773e-05, 1.54741e-07, 
    8.195327e-09, 6.663929e-09, 4.043073e-09, 1.933557e-08, 7.051055e-09,
  1.643048e-05, 2.410735e-05, 1.540943e-05, 1.093602e-05, 2.537472e-05, 
    2.000398e-05, 1.907068e-05, 2.237164e-05, 1.150396e-06, 9.483736e-07, 
    5.525754e-07, 6.445275e-09, 4.533273e-09, 4.916984e-09, 3.89551e-09,
  3.825669e-06, 1.16701e-05, 9.574177e-06, 6.084135e-06, 8.029171e-06, 
    7.953339e-06, 2.30807e-06, 1.714752e-07, 2.096099e-06, 1.506368e-06, 
    9.398599e-08, 6.573589e-09, 5.015516e-09, 6.691725e-09, 7.315959e-10,
  1.047135e-07, 1.920302e-07, 2.364774e-07, 5.828596e-07, 1.61433e-06, 
    1.358471e-06, 3.484988e-06, 6.911849e-07, 1.707878e-06, 1.976401e-06, 
    6.088462e-06, 2.520193e-05, 2.092441e-05, 2.81824e-05, 1.670592e-05,
  7.564363e-08, 9.54192e-08, 1.337283e-07, 9.039684e-08, 1.718921e-06, 
    2.534446e-06, 7.070705e-06, 4.970691e-06, 1.841335e-06, 1.32481e-06, 
    3.913046e-06, 1.796934e-05, 2.68165e-05, 1.872952e-05, 3.507804e-06,
  1.368493e-07, 3.567234e-06, 6.472417e-07, 1.805724e-07, 3.860039e-06, 
    2.466813e-06, 1.433705e-06, 1.679954e-06, 3.195301e-06, 6.337007e-06, 
    1.495137e-05, 1.988887e-05, 2.603208e-05, 1.699809e-05, 2.850523e-06,
  1.238026e-06, 3.116239e-08, 1.922843e-06, 9.58706e-06, 4.031654e-06, 
    2.793825e-06, 3.255872e-06, 3.39752e-06, 9.547387e-06, 3.162842e-05, 
    6.160138e-05, 4.070354e-05, 3.053743e-05, 6.78529e-06, 1.514235e-05,
  3.291798e-06, 5.096217e-07, 3.317644e-07, 2.222707e-06, 3.035631e-06, 
    1.163897e-06, 5.600522e-06, 1.041164e-05, 3.362808e-05, 7.953867e-05, 
    2.23362e-06, 8.177472e-08, 7.692383e-06, 5.034289e-07, 2.325977e-05,
  1.155786e-06, 1.130316e-06, 3.638524e-06, 4.660571e-06, 6.193761e-06, 
    2.969705e-06, 7.383912e-06, 1.288089e-05, 5.242541e-05, 1.476996e-05, 
    5.722909e-07, 1.30668e-07, 3.252026e-07, 6.155603e-07, 1.303868e-05,
  1.302305e-06, 1.633401e-06, 4.171641e-06, 4.591718e-06, 9.05012e-06, 
    6.797311e-06, 1.122236e-05, 1.590703e-05, 1.812746e-05, 6.494126e-06, 
    5.949731e-08, 1.862283e-07, 1.132115e-07, 7.01174e-06, 2.690955e-06,
  2.372418e-08, 3.683776e-09, 1.674946e-06, 1.355614e-06, 4.827954e-06, 
    1.202795e-05, 1.827198e-05, 2.128572e-05, 1.335651e-05, 6.943003e-06, 
    6.608366e-08, 1.01446e-07, 2.531198e-07, 1.154743e-05, 7.572535e-07,
  1.476434e-08, 2.997067e-09, 3.689891e-08, 1.004381e-07, 1.006233e-06, 
    1.03066e-05, 1.862529e-05, 1.354859e-05, 8.734719e-06, 4.067329e-06, 
    1.328355e-06, 3.757827e-07, 1.097942e-07, 2.078964e-06, 2.247251e-07,
  1.118828e-08, 3.5835e-09, 2.348433e-09, 3.755014e-07, 1.390489e-06, 
    9.819656e-07, 1.425621e-06, 1.325638e-06, 3.544053e-06, 1.64609e-06, 
    4.564592e-07, 1.208385e-07, 1.414179e-07, 4.394676e-07, 2.224864e-07,
  3.290158e-07, 3.344648e-07, 1.56361e-07, 4.387172e-07, 1.695004e-06, 
    2.928562e-06, 7.047106e-06, 2.099034e-06, 1.975222e-06, 3.014714e-06, 
    2.914574e-06, 1.322122e-05, 1.833738e-05, 2.672052e-05, 2.265365e-05,
  2.636585e-07, 1.333124e-07, 6.684864e-08, 1.227124e-07, 3.137236e-06, 
    3.802763e-06, 3.825656e-06, 3.643784e-06, 1.372161e-06, 1.374114e-06, 
    2.410669e-06, 5.498513e-06, 1.449249e-05, 2.71682e-05, 1.8413e-05,
  2.251411e-07, 2.012504e-06, 1.149999e-06, 2.069416e-08, 3.64841e-06, 
    1.394429e-06, 4.272434e-07, 5.820379e-07, 1.051935e-06, 3.475979e-06, 
    9.601584e-06, 1.457372e-05, 1.55354e-05, 2.678055e-05, 2.271936e-05,
  9.70619e-09, 4.683437e-08, 3.014113e-07, 7.556016e-07, 1.102341e-07, 
    2.902841e-07, 6.489811e-07, 1.241802e-06, 2.749601e-06, 1.004996e-05, 
    4.649767e-05, 4.425504e-05, 3.806968e-05, 3.222676e-05, 3.939947e-05,
  1.241426e-07, 1.45896e-06, 3.179575e-08, 1.089073e-08, 2.147386e-08, 
    9.06368e-09, 2.872745e-07, 2.18334e-06, 7.175106e-06, 1.430676e-05, 
    6.984168e-07, 4.660321e-06, 5.527824e-05, 3.039351e-05, 8.775193e-05,
  2.115474e-08, 9.918462e-08, 1.4285e-06, 2.046485e-09, 3.206743e-08, 
    1.129455e-09, 2.976938e-08, 1.862689e-06, 2.695921e-05, 8.304937e-06, 
    8.324887e-06, 1.927699e-06, 2.265709e-06, 6.964276e-05, 9.912916e-05,
  9.756193e-08, 2.052942e-08, 5.952144e-07, 3.098575e-07, 2.094329e-07, 
    4.051094e-07, 5.618708e-06, 1.815012e-05, 3.091936e-05, 1.729853e-06, 
    5.398161e-07, 7.488414e-08, 1.295223e-07, 9.716192e-05, 8.454222e-05,
  1.570855e-08, 5.692494e-09, 2.687865e-08, 2.779561e-07, 1.404111e-06, 
    3.520457e-06, 9.007705e-06, 1.663839e-05, 1.545943e-05, 6.595029e-07, 
    4.735591e-07, 1.788829e-07, 1.043846e-07, 1.953662e-05, 5.71587e-06,
  5.446653e-09, 7.755238e-09, 2.077794e-08, 3.802399e-08, 5.729741e-07, 
    6.8316e-06, 9.944986e-06, 1.084177e-05, 7.844009e-07, 4.888468e-07, 
    4.38269e-07, 3.321543e-07, 2.579281e-09, 2.811587e-07, 5.080188e-07,
  9.324863e-09, 1.467197e-08, 2.785455e-08, 8.02644e-07, 2.337939e-06, 
    2.243479e-06, 5.13168e-06, 5.189136e-07, 5.50017e-07, 1.255627e-06, 
    1.199967e-06, 1.062622e-07, 8.027764e-09, 8.83448e-08, 7.452297e-08,
  1.925321e-08, 8.811276e-08, 1.524385e-07, 8.758951e-08, 1.184528e-07, 
    2.233326e-06, 9.488371e-06, 1.090574e-05, 2.0411e-05, 3.676184e-05, 
    1.722921e-05, 1.03947e-05, 9.56744e-06, 1.581588e-05, 2.654123e-05,
  4.036576e-08, 8.470386e-08, 8.689654e-08, 1.19106e-07, 2.670251e-06, 
    8.335684e-06, 1.399975e-05, 1.621227e-05, 4.144749e-05, 3.393904e-05, 
    1.938263e-05, 2.241998e-05, 3.169456e-05, 4.010199e-05, 6.881683e-05,
  2.521333e-07, 7.120353e-07, 4.640803e-07, 1.065562e-06, 5.036863e-06, 
    3.502732e-06, 3.538397e-06, 8.880711e-06, 3.828339e-05, 4.114484e-05, 
    4.477391e-05, 5.405596e-05, 7.175042e-05, 9.1822e-05, 0.0001927204,
  5.362662e-07, 3.047938e-07, 1.892618e-06, 5.619062e-06, 3.736257e-06, 
    4.34247e-06, 3.893923e-06, 5.176433e-06, 1.75016e-05, 3.574759e-05, 
    6.868437e-05, 8.419404e-05, 8.460476e-05, 8.738181e-05, 6.546047e-05,
  3.502989e-07, 2.918696e-07, 4.774524e-07, 1.164128e-07, 3.902917e-07, 
    7.186261e-07, 2.66313e-06, 7.46694e-06, 1.748402e-05, 4.353136e-05, 
    3.82504e-05, 9.398696e-05, 0.0001206677, 5.059445e-05, 5.693891e-05,
  2.088984e-07, 2.488173e-07, 3.204763e-07, 2.308435e-07, 4.034988e-08, 
    7.913559e-07, 3.72232e-06, 7.650779e-06, 4.700477e-05, 3.136452e-05, 
    2.686148e-05, 2.638328e-05, 3.037337e-05, 7.926256e-05, 7.369227e-05,
  5.280874e-07, 5.892961e-07, 9.068328e-07, 2.835719e-06, 1.838367e-06, 
    5.328099e-06, 1.582608e-05, 2.298204e-05, 3.049949e-05, 4.65181e-06, 
    9.119197e-07, 1.172029e-06, 3.308528e-06, 8.493973e-05, 3.682732e-05,
  8.457549e-07, 1.013483e-05, 1.387626e-05, 2.350999e-06, 2.80133e-07, 
    1.197872e-06, 1.440432e-05, 1.729037e-05, 2.078448e-05, 5.367277e-06, 
    4.540137e-06, 4.726007e-06, 3.732785e-06, 3.633424e-05, 3.753982e-06,
  6.535733e-06, 1.454871e-05, 1.163852e-05, 6.505375e-07, 7.006261e-07, 
    4.765981e-06, 4.79124e-06, 1.415386e-05, 8.68776e-06, 7.744102e-06, 
    9.93382e-06, 1.057511e-05, 6.012991e-07, 2.455686e-06, 5.279446e-06,
  1.210267e-05, 1.784627e-05, 7.683834e-06, 1.209218e-06, 1.43584e-06, 
    8.513469e-07, 1.286627e-06, 2.675061e-06, 9.948496e-06, 1.193207e-05, 
    9.630553e-06, 5.617259e-06, 1.421748e-06, 1.40388e-06, 1.044976e-05,
  9.758762e-06, 3.233523e-05, 6.439223e-05, 0.0001417674, 0.0002306244, 
    0.0002641972, 0.0002723632, 0.0002260307, 0.0002029348, 9.46042e-05, 
    3.538026e-05, 1.992006e-05, 1.903259e-05, 2.023634e-05, 4.790768e-05,
  2.023197e-05, 1.312549e-05, 3.004846e-05, 0.0001251757, 0.0002513142, 
    0.0003301568, 0.0003492021, 0.0003363727, 0.0002874197, 0.0001616455, 
    7.988176e-05, 4.918708e-05, 2.956555e-05, 1.761216e-05, 1.424813e-05,
  1.319557e-05, 2.913933e-05, 2.374724e-05, 3.315549e-05, 0.0001393009, 
    0.0001950449, 0.0002428487, 0.0003244262, 0.0003258935, 0.0002218643, 
    0.0001556877, 0.0001246922, 0.0001045397, 8.89755e-05, 0.0001167433,
  3.158828e-05, 1.623622e-05, 2.372678e-05, 4.42427e-05, 4.532054e-05, 
    6.147907e-05, 9.445012e-05, 0.0001422246, 0.0001887157, 0.0001646342, 
    0.0001902289, 0.0001683636, 0.0001349726, 0.0001602153, 0.0001928409,
  2.461356e-05, 2.226428e-05, 1.895952e-05, 1.618433e-05, 1.459453e-05, 
    1.782355e-05, 2.289586e-05, 2.305339e-05, 3.537365e-05, 8.729561e-05, 
    0.0001085019, 8.482515e-05, 8.836772e-05, 6.487968e-05, 8.479684e-05,
  6.450818e-06, 1.089219e-05, 1.013179e-05, 1.440402e-05, 1.860942e-05, 
    1.22418e-05, 1.327163e-05, 1.860731e-05, 3.413938e-05, 1.790307e-05, 
    1.319284e-05, 6.582011e-06, 3.68259e-06, 2.835907e-05, 4.164547e-05,
  7.492462e-06, 8.680518e-06, 2.042911e-05, 2.147876e-05, 1.098566e-05, 
    5.924784e-06, 8.650377e-06, 1.905109e-05, 2.537044e-05, 1.794658e-05, 
    8.512312e-06, 5.277955e-06, 8.958908e-06, 1.952137e-05, 1.107124e-05,
  1.711816e-06, 8.752637e-06, 2.229097e-05, 1.147116e-05, 1.79295e-06, 
    2.489511e-07, 3.632678e-06, 1.448119e-05, 5.344677e-05, 2.656418e-05, 
    1.982238e-05, 1.252504e-05, 1.625047e-05, 2.62775e-05, 3.313502e-06,
  5.167807e-06, 1.186556e-05, 1.727032e-05, 5.516331e-06, 2.715477e-07, 
    1.597199e-06, 2.256158e-06, 2.566399e-05, 2.379636e-05, 3.190144e-05, 
    2.614061e-05, 1.493652e-05, 3.096197e-06, 3.528606e-06, 5.613367e-06,
  3.65856e-06, 1.038136e-05, 1.200504e-05, 6.877967e-07, 4.180736e-08, 
    2.983367e-07, 6.381134e-06, 8.227175e-06, 3.089615e-05, 3.644748e-05, 
    2.429537e-05, 9.382897e-06, 3.791766e-07, 4.354398e-07, 2.636735e-06,
  3.060213e-11, 1.976639e-10, 2.697969e-09, 1.830232e-08, 3.259117e-08, 
    6.461951e-07, 1.236273e-05, 3.765991e-05, 0.0001212979, 0.0001564811, 
    0.000121613, 0.0001174244, 9.129829e-05, 9.302215e-05, 0.0002562538,
  1.021653e-11, 4.088507e-12, 3.725776e-10, 1.181618e-08, 1.446589e-08, 
    1.723512e-07, 5.00586e-06, 2.708993e-05, 0.0001083721, 0.0001838388, 
    0.0002354119, 0.000232646, 0.0001556083, 9.002505e-05, 0.0001986598,
  2.193787e-27, 7.201902e-14, 2.09609e-10, 1.910159e-09, 3.40166e-08, 
    8.962422e-08, 8.619228e-07, 1.185449e-05, 5.886425e-05, 0.0001183486, 
    0.0001973516, 0.0002247444, 0.0001835256, 0.000190244, 0.0002348169,
  9.221669e-27, 3.963062e-14, 9.487524e-10, 3.658317e-07, 2.681343e-07, 
    4.320243e-06, 3.929385e-06, 5.007262e-06, 2.027591e-05, 8.086213e-05, 
    0.0001688784, 0.0001689214, 0.0001284083, 0.0001956384, 0.0002087446,
  1.776346e-14, 1.636147e-29, 6.859562e-13, 1.180902e-09, 2.657086e-07, 
    5.899508e-06, 1.610674e-05, 2.970522e-05, 6.872815e-05, 0.0001033384, 
    3.816411e-05, 5.800516e-05, 0.0001761771, 0.0001487441, 0.000106974,
  8.608968e-11, 4.084779e-14, 2.539894e-12, 6.460391e-10, 1.177983e-07, 
    4.532639e-06, 2.306845e-05, 6.552111e-05, 9.603798e-05, 2.796528e-05, 
    1.388735e-05, 3.280112e-06, 1.514034e-05, 3.665559e-05, 6.483516e-05,
  7.954724e-10, 7.011174e-13, 1.460171e-11, 1.23297e-10, 4.676589e-09, 
    4.943146e-07, 1.471854e-05, 3.247698e-05, 4.554989e-05, 2.982631e-05, 
    6.838959e-06, 1.213384e-06, 7.55085e-07, 1.418486e-05, 1.440614e-05,
  2.31672e-09, 4.863775e-11, 4.957558e-16, 5.676931e-12, 4.860855e-09, 
    4.215571e-07, 5.297324e-06, 2.286789e-05, 7.914663e-05, 2.908854e-05, 
    4.391579e-06, 1.162533e-09, 9.310064e-08, 5.962118e-07, 6.377296e-06,
  3.602887e-10, 1.002234e-09, 1.213416e-10, 6.342583e-11, 7.50427e-09, 
    4.455255e-07, 5.934243e-06, 1.917802e-05, 1.140079e-05, 1.28757e-05, 
    5.858388e-06, 6.009525e-08, 1.653348e-09, 5.751471e-08, 1.305227e-06,
  1.046207e-09, 4.922243e-09, 2.325054e-09, 1.136124e-09, 1.885796e-08, 
    3.271503e-07, 5.474702e-06, 2.855855e-06, 4.6717e-06, 2.801146e-06, 
    1.489241e-06, 1.383663e-11, 9.805647e-14, 6.785785e-10, 2.141562e-08,
  7.160004e-10, 2.329971e-10, 8.031705e-10, 1.052191e-09, 6.258822e-09, 
    3.030851e-07, 3.657576e-06, 6.568312e-06, 1.67927e-05, 4.083611e-05, 
    6.092236e-05, 8.295508e-05, 7.065212e-05, 4.40445e-05, 5.262519e-05,
  1.176276e-09, 1.746439e-09, 1.94341e-09, 1.651799e-09, 7.679639e-09, 
    2.149058e-07, 2.035082e-06, 3.153925e-06, 8.364964e-06, 1.946113e-05, 
    5.640258e-05, 7.160465e-05, 5.011701e-05, 3.053834e-05, 6.979436e-05,
  2.817669e-09, 2.151694e-08, 2.099946e-08, 1.723307e-08, 1.480845e-08, 
    2.41312e-08, 9.39171e-07, 4.345317e-06, 5.062613e-06, 1.062493e-05, 
    3.427035e-05, 4.797924e-05, 2.867394e-05, 5.162029e-05, 5.432931e-05,
  3.360591e-08, 5.76059e-08, 2.150502e-07, 1.746544e-07, 7.235956e-08, 
    1.068037e-07, 3.079281e-07, 4.330389e-07, 1.047975e-06, 1.723851e-05, 
    5.925335e-05, 8.417362e-05, 3.899441e-05, 7.757067e-05, 2.46749e-05,
  3.153599e-08, 1.354142e-07, 5.278951e-07, 4.674254e-07, 2.560691e-07, 
    1.000967e-07, 7.862971e-07, 3.999857e-06, 1.213266e-05, 3.383352e-05, 
    7.05316e-06, 3.124518e-05, 7.988661e-05, 7.740786e-05, 2.408415e-05,
  7.788714e-09, 1.371431e-07, 3.515712e-07, 1.234931e-06, 7.854919e-07, 
    3.878485e-07, 2.696131e-07, 3.812572e-06, 1.631372e-05, 5.688564e-06, 
    1.911249e-05, 8.21091e-06, 1.222115e-05, 5.481151e-05, 2.186558e-05,
  1.689828e-08, 1.182062e-07, 5.320449e-07, 1.567681e-06, 2.023802e-06, 
    1.068018e-06, 5.633827e-07, 1.104094e-06, 4.382304e-06, 7.836371e-06, 
    1.05705e-05, 4.462473e-06, 4.985934e-06, 3.531445e-05, 1.440031e-05,
  1.354977e-08, 1.34585e-07, 8.361451e-07, 1.306498e-06, 2.498387e-06, 
    2.016414e-06, 1.126138e-06, 6.512669e-07, 3.510113e-06, 3.662803e-06, 
    1.911281e-06, 5.085799e-07, 3.424046e-06, 3.69788e-05, 3.503407e-06,
  1.401116e-08, 6.01417e-07, 9.278024e-07, 1.512046e-06, 2.684172e-06, 
    2.47155e-06, 1.385641e-06, 7.611904e-07, 7.639512e-08, 8.571195e-07, 
    1.753266e-07, 9.692248e-10, 9.51544e-07, 8.374936e-07, 3.766609e-07,
  4.946189e-08, 7.04828e-07, 1.441052e-06, 2.058827e-06, 3.701213e-06, 
    2.937714e-06, 1.726232e-06, 3.887157e-07, 2.824713e-07, 9.425081e-08, 
    3.664195e-08, 4.754269e-09, 7.033513e-10, 2.209194e-08, 1.567921e-08,
  3.345146e-05, 1.010318e-05, 6.754484e-06, 6.409954e-06, 1.202143e-06, 
    4.959282e-07, 3.820772e-07, 2.142756e-07, 1.758035e-06, 4.074846e-06, 
    3.590122e-06, 5.06039e-06, 2.98549e-06, 8.563609e-06, 2.143739e-06,
  3.499057e-05, 2.041553e-05, 4.31078e-06, 1.520731e-06, 1.092223e-06, 
    9.341255e-07, 1.642273e-06, 1.50826e-06, 2.358869e-06, 1.599065e-06, 
    6.51974e-07, 1.046917e-06, 6.904367e-07, 1.233682e-06, 6.973967e-06,
  0.0001423574, 6.799892e-05, 2.085889e-05, 6.095313e-06, 7.073276e-06, 
    1.968319e-06, 1.119132e-06, 1.328182e-06, 2.271363e-06, 1.058609e-06, 
    5.055259e-07, 4.152116e-07, 1.666118e-07, 1.210367e-06, 5.624317e-06,
  0.0001770653, 4.795995e-05, 3.154171e-05, 2.893307e-05, 1.144744e-05, 
    5.600738e-06, 3.30548e-06, 2.140262e-06, 1.082829e-06, 4.617754e-07, 
    1.648866e-06, 7.627575e-07, 5.036129e-07, 6.215117e-06, 2.521506e-06,
  0.0001430663, 5.430447e-05, 3.542749e-05, 3.547192e-05, 1.873391e-05, 
    8.066082e-06, 4.624202e-06, 3.550002e-06, 3.295359e-06, 3.871754e-06, 
    8.751783e-08, 3.015677e-07, 1.386037e-06, 5.593573e-06, 4.006472e-06,
  7.865151e-05, 8.300888e-05, 9.984026e-05, 0.000103824, 7.51267e-05, 
    4.080053e-05, 2.614201e-05, 1.395592e-05, 1.214147e-05, 1.096346e-05, 
    1.381136e-05, 3.929488e-06, 7.384705e-07, 1.209287e-05, 1.302186e-05,
  5.848077e-05, 0.0001013902, 0.0001254637, 0.0001205683, 8.783094e-05, 
    8.152505e-05, 7.896321e-05, 6.989353e-05, 8.308562e-05, 3.751303e-05, 
    1.112009e-05, 9.370889e-06, 5.723309e-06, 2.815608e-05, 8.674902e-06,
  5.762267e-05, 7.641989e-05, 7.131236e-05, 5.526837e-05, 4.695495e-05, 
    4.551706e-05, 6.318187e-05, 7.000756e-05, 8.455538e-05, 3.245485e-05, 
    1.561783e-05, 1.524149e-05, 1.61776e-05, 4.705186e-05, 3.998556e-06,
  4.944398e-05, 3.074585e-05, 2.074354e-05, 3.006705e-05, 3.060387e-05, 
    4.373259e-05, 5.184635e-05, 7.712205e-05, 3.880892e-05, 1.756499e-05, 
    8.142938e-06, 7.97153e-06, 1.911598e-05, 3.005543e-05, 9.927079e-06,
  3.088199e-05, 1.272328e-05, 2.791003e-05, 4.76866e-05, 5.899384e-05, 
    4.979875e-05, 5.369058e-05, 3.507597e-05, 1.646253e-05, 7.044333e-06, 
    8.971724e-06, 6.758921e-06, 6.14887e-06, 8.706671e-06, 1.041063e-05,
  0.0003406292, 0.0002723966, 0.0002788801, 0.000277918, 0.0002544141, 
    0.0003120953, 0.000268797, 0.0002077965, 0.000175328, 0.000101197, 
    4.324322e-05, 2.574507e-05, 2.137382e-05, 1.091394e-05, 3.227443e-06,
  0.0001571622, 0.0001774125, 0.0002684952, 0.0003003441, 0.0003462723, 
    0.0003139543, 0.0002631899, 0.0002149754, 0.0001864742, 0.0001182868, 
    7.961818e-05, 6.464445e-05, 5.375478e-05, 3.39473e-05, 4.230207e-05,
  0.0001175521, 0.0001258288, 0.0001603575, 0.000218412, 0.0002097111, 
    0.0001919523, 0.000179618, 0.0001961273, 0.0001584018, 9.888157e-05, 
    7.762331e-05, 8.009723e-05, 7.238454e-05, 5.250446e-05, 4.817263e-05,
  4.691436e-05, 4.17449e-05, 7.974586e-05, 0.0001128062, 0.0001017608, 
    0.0001055281, 0.0001243068, 0.0001587376, 0.0001256824, 7.97904e-05, 
    9.864494e-05, 0.0001150637, 8.038962e-05, 5.347506e-05, 2.265684e-05,
  9.260615e-06, 1.925756e-05, 4.136726e-05, 6.17174e-05, 6.196538e-05, 
    7.097864e-05, 8.46886e-05, 9.516998e-05, 9.448879e-05, 0.0001324847, 
    0.0001145156, 0.0001224598, 0.0001039504, 2.223056e-05, 2.146108e-05,
  1.510432e-06, 7.789231e-06, 2.004368e-05, 3.176695e-05, 4.578163e-05, 
    6.459317e-05, 8.66375e-05, 9.756776e-05, 0.0001450612, 0.0001564619, 
    0.0001258359, 4.905926e-05, 2.141216e-05, 3.099335e-05, 4.082107e-05,
  4.170038e-07, 2.348387e-06, 8.565055e-06, 6.463663e-06, 1.27728e-05, 
    2.742636e-05, 5.928171e-05, 7.748891e-05, 0.0001040159, 5.487512e-05, 
    2.442032e-05, 2.429864e-05, 2.636181e-05, 5.048757e-05, 4.411352e-05,
  2.872236e-08, 1.265369e-06, 5.275399e-06, 4.218942e-06, 1.718328e-06, 
    3.674453e-06, 1.399693e-05, 2.343797e-05, 3.2904e-05, 8.932227e-06, 
    8.906771e-06, 9.909107e-06, 6.643026e-06, 1.669285e-05, 1.1373e-05,
  1.611761e-08, 5.979792e-07, 4.788734e-06, 2.998759e-06, 3.248648e-06, 
    1.094881e-05, 2.013363e-05, 3.935104e-05, 1.053928e-05, 5.06986e-06, 
    6.965735e-06, 1.248178e-05, 6.26584e-06, 1.204483e-05, 2.344192e-05,
  4.149191e-08, 4.906743e-07, 4.419831e-06, 6.827588e-06, 8.164633e-06, 
    1.450087e-05, 2.476361e-05, 1.187487e-05, 5.18202e-06, 5.189596e-06, 
    1.086803e-05, 1.160207e-05, 3.398191e-06, 1.173104e-06, 3.399311e-06,
  9.307938e-07, 1.766756e-07, 4.478876e-06, 6.129428e-06, 3.956054e-06, 
    1.753642e-05, 1.869059e-05, 1.539014e-05, 3.492722e-05, 2.265994e-05, 
    1.041308e-05, 6.567621e-06, 7.265511e-06, 1.490584e-05, 1.790132e-05,
  2.278227e-07, 1.633453e-06, 2.024428e-06, 9.432577e-06, 1.003012e-05, 
    2.140085e-05, 2.123341e-05, 1.602013e-05, 1.767628e-05, 1.172381e-05, 
    6.164972e-06, 3.541124e-06, 4.026379e-06, 8.32363e-06, 8.277233e-06,
  1.961712e-05, 1.012766e-05, 9.121445e-07, 8.287002e-06, 3.264241e-05, 
    2.069576e-05, 8.172175e-06, 2.387178e-05, 1.860041e-05, 7.246185e-06, 
    1.974346e-06, 1.386295e-06, 1.812859e-06, 4.845602e-06, 1.19634e-06,
  1.85969e-05, 1.479204e-06, 1.000611e-06, 3.044203e-06, 5.859733e-06, 
    6.744957e-06, 6.811963e-06, 1.782213e-05, 1.486058e-05, 8.381215e-06, 
    6.738217e-06, 3.840128e-06, 4.026611e-06, 3.962549e-06, 9.554807e-07,
  2.731265e-06, 9.31795e-07, 8.836193e-07, 1.659482e-06, 1.722731e-06, 
    2.633159e-06, 4.379009e-06, 6.321033e-06, 8.897807e-06, 1.003528e-05, 
    1.370951e-07, 1.853041e-06, 6.67999e-06, 1.331229e-06, 3.043174e-06,
  1.587086e-07, 1.314799e-07, 1.72489e-07, 4.1053e-07, 5.840635e-07, 
    8.157267e-07, 1.190159e-06, 1.651266e-06, 1.576644e-06, 1.096294e-07, 
    4.52805e-06, 1.199769e-06, 3.671224e-08, 3.903647e-06, 5.458213e-06,
  9.32902e-07, 1.357091e-07, 7.939258e-08, 2.438917e-07, 1.930903e-07, 
    3.062412e-07, 2.670187e-06, 3.092848e-07, 1.555053e-06, 3.281025e-06, 
    3.895612e-06, 6.814637e-07, 9.841635e-09, 1.911666e-05, 9.541025e-06,
  5.039446e-06, 2.999027e-06, 1.038457e-06, 2.066739e-07, 9.180563e-07, 
    3.099405e-06, 5.96591e-06, 4.627913e-06, 9.8628e-06, 8.523127e-06, 
    4.011193e-06, 4.892324e-06, 9.857865e-07, 3.089766e-05, 7.741615e-06,
  1.902083e-05, 1.895961e-05, 4.596075e-06, 2.952865e-06, 4.267432e-05, 
    9.907871e-05, 6.659912e-05, 3.479916e-05, 1.506802e-05, 1.987218e-05, 
    9.459745e-06, 1.053047e-05, 1.196692e-05, 2.907507e-05, 1.076965e-05,
  4.134961e-05, 4.532149e-05, 2.670375e-05, 4.40384e-05, 0.0001617637, 
    0.0002103102, 0.0001778586, 7.885004e-05, 8.354693e-05, 5.637025e-05, 
    3.56403e-05, 3.8824e-05, 4.502991e-05, 3.94238e-05, 1.639155e-05,
  1.256814e-05, 1.29597e-05, 7.076176e-05, 8.277393e-05, 5.273695e-05, 
    7.976909e-05, 0.0001581051, 0.0002577491, 0.0004023897, 0.0002686234, 
    0.0001372646, 7.090611e-05, 4.895731e-05, 2.829074e-05, 3.077442e-06,
  2.689558e-06, 1.646528e-05, 5.814504e-05, 0.0001608299, 0.0001351788, 
    0.0001275107, 0.0001726584, 0.0002754581, 0.000380158, 0.0002797942, 
    0.0001833084, 0.0001156793, 7.831043e-05, 4.927051e-05, 7.001655e-06,
  0.0001011724, 2.643868e-05, 8.336968e-06, 5.662755e-05, 0.0001719858, 
    0.0001198554, 8.699027e-05, 0.0002219993, 0.0002861602, 0.0002023244, 
    0.0001397478, 0.0001138557, 7.401291e-05, 3.762296e-05, 3.495298e-07,
  0.000143657, 3.61805e-05, 5.812946e-05, 0.0001184418, 0.000144753, 
    0.0001185952, 9.523351e-05, 0.000144954, 0.0001835336, 0.0001718104, 
    0.0002657539, 0.0002739352, 0.0001665725, 5.810595e-05, 1.072269e-05,
  9.379491e-05, 7.236401e-05, 0.0001017695, 0.0001602952, 0.0001490769, 
    0.0001511537, 0.0001272785, 0.0001364202, 0.0001574986, 0.0002246838, 
    0.0001356743, 0.0002802481, 0.0004884622, 0.000163644, 8.150027e-05,
  2.893319e-05, 6.452372e-05, 9.810666e-05, 9.766371e-05, 0.0001007932, 
    0.0001088868, 0.0001106026, 0.000117433, 0.0001197432, 5.787572e-05, 
    0.0001457893, 0.000244556, 0.0002580159, 0.0003156649, 0.0001823156,
  2.103354e-05, 6.126773e-05, 6.285313e-05, 5.567571e-05, 4.377547e-05, 
    3.032171e-05, 5.891874e-05, 4.868678e-05, 5.659195e-05, 6.327965e-05, 
    9.14053e-05, 0.0001138752, 0.0001588266, 0.0003582451, 0.0001881866,
  5.081278e-05, 6.840438e-05, 5.849989e-05, 3.956045e-05, 4.509771e-05, 
    4.044705e-05, 5.852156e-05, 3.977898e-05, 6.775176e-05, 7.655664e-05, 
    6.682361e-05, 8.443795e-05, 0.0001364342, 0.0002669594, 0.0001334651,
  6.725252e-05, 0.000107136, 8.648051e-05, 9.362397e-05, 0.0001079667, 
    0.0001093637, 8.546974e-05, 0.0001176702, 5.793155e-05, 9.624028e-05, 
    5.250244e-05, 4.622394e-05, 0.0001074525, 0.0001744308, 0.0001519315,
  5.383847e-05, 0.0001078287, 0.00013166, 0.0001379707, 0.0001505771, 
    0.000168135, 0.0001619898, 9.221554e-05, 8.865113e-05, 6.513453e-05, 
    3.699058e-05, 3.48675e-05, 5.084653e-05, 8.730715e-05, 8.719345e-05,
  2.36462e-05, 3.462068e-05, 6.482423e-05, 3.820787e-05, 1.108453e-05, 
    1.203599e-06, 1.193922e-06, 3.578428e-06, 2.210288e-05, 4.639193e-05, 
    6.058268e-05, 7.168115e-05, 6.03771e-05, 2.920725e-05, 1.280079e-05,
  9.68998e-06, 7.461254e-06, 9.380332e-06, 5.979493e-06, 2.10697e-06, 
    8.10879e-07, 5.246418e-07, 2.757552e-07, 8.034746e-07, 3.834968e-06, 
    9.45252e-06, 1.401891e-05, 8.708008e-06, 6.534844e-06, 2.406939e-06,
  2.30572e-07, 6.264945e-08, 2.675916e-08, 4.774007e-08, 5.088798e-08, 
    4.787377e-08, 5.747188e-08, 7.208214e-08, 4.896353e-07, 4.637596e-06, 
    1.606444e-05, 1.133778e-05, 3.519656e-06, 6.102396e-06, 1.039001e-07,
  1.461138e-08, 1.324515e-07, 1.380283e-07, 3.230886e-07, 3.861801e-07, 
    1.867303e-06, 4.290832e-06, 2.940777e-06, 1.124449e-05, 3.797836e-05, 
    6.751453e-05, 8.406273e-05, 3.316375e-05, 3.161816e-05, 3.45779e-06,
  5.861283e-08, 1.369288e-06, 1.166683e-06, 8.900383e-07, 1.078345e-06, 
    2.517904e-06, 4.471183e-06, 9.55841e-06, 2.468973e-05, 7.134024e-05, 
    2.843596e-05, 3.245441e-05, 0.0001038979, 3.22844e-05, 4.025691e-05,
  2.570007e-08, 1.160879e-06, 1.052441e-06, 6.066799e-07, 1.150174e-06, 
    1.820085e-06, 1.247182e-06, 5.899655e-06, 1.466061e-05, 2.071416e-05, 
    3.61243e-05, 1.400606e-05, 1.196007e-05, 4.550549e-05, 4.479616e-05,
  2.412757e-08, 7.100019e-07, 7.268558e-07, 6.699362e-07, 1.280095e-07, 
    8.284468e-07, 5.151842e-07, 2.696552e-06, 1.321584e-05, 2.98812e-05, 
    1.406679e-05, 6.459588e-07, 9.074336e-08, 1.627605e-05, 1.728181e-05,
  1.434029e-08, 7.607266e-08, 7.67002e-07, 8.193909e-07, 1.915952e-07, 
    3.806535e-07, 7.645859e-07, 1.40545e-06, 2.183007e-05, 2.986071e-05, 
    5.697504e-06, 1.084232e-06, 5.808307e-07, 1.863233e-05, 4.870218e-06,
  9.524443e-09, 4.59799e-08, 5.845164e-07, 6.122571e-07, 1.167239e-06, 
    2.335113e-06, 3.158676e-06, 3.39575e-06, 5.002085e-06, 1.830722e-05, 
    2.040624e-06, 3.781522e-06, 7.208041e-06, 8.868464e-06, 7.019152e-07,
  8.314234e-09, 3.497334e-08, 4.541169e-08, 7.454464e-08, 5.299041e-07, 
    1.164266e-06, 2.087733e-06, 2.087698e-06, 1.121396e-05, 8.718221e-06, 
    1.089171e-06, 1.082706e-06, 5.388465e-06, 3.766122e-06, 1.434149e-06,
  9.289299e-09, 1.032123e-08, 3.837769e-09, 1.798623e-09, 1.016024e-09, 
    6.071971e-10, 8.095331e-10, 2.317353e-08, 6.068709e-07, 8.719576e-08, 
    3.239881e-09, 1.427113e-09, 1.459083e-07, 1.304136e-07, 1.597671e-08,
  1.801822e-08, 1.106281e-08, 1.249259e-08, 1.725448e-08, 4.313802e-07, 
    8.695101e-07, 1.206122e-06, 1.142117e-06, 9.987054e-07, 1.95789e-07, 
    3.526095e-08, 3.841189e-08, 1.353925e-07, 2.27619e-07, 2.082873e-08,
  2.999797e-08, 7.522753e-08, 4.318218e-08, 3.697376e-08, 1.25772e-06, 
    1.217506e-06, 1.462356e-06, 2.537806e-06, 2.860784e-06, 1.718784e-06, 
    6.139209e-07, 3.663397e-07, 1.00044e-07, 1.306116e-07, 8.948494e-09,
  9.247297e-08, 3.260894e-08, 4.971985e-07, 1.371965e-06, 1.179236e-06, 
    1.870376e-06, 3.005787e-06, 4.053342e-06, 5.069665e-06, 4.058974e-06, 
    2.342894e-06, 1.526059e-06, 8.782283e-07, 3.02791e-07, 2.147317e-07,
  5.603975e-08, 7.327142e-08, 1.714267e-07, 4.828193e-07, 5.91046e-07, 
    9.176e-07, 1.726549e-06, 2.640565e-06, 4.639913e-06, 3.557461e-06, 
    3.209501e-08, 4.699107e-09, 1.228547e-06, 1.750346e-07, 4.140979e-07,
  6.696287e-08, 1.945168e-07, 3.467144e-08, 7.310406e-07, 1.143381e-06, 
    1.547961e-06, 1.055309e-06, 6.674532e-07, 2.563722e-07, 7.473979e-08, 
    3.488436e-08, 2.812491e-09, 1.042863e-08, 7.612723e-08, 2.400737e-06,
  1.496335e-07, 1.124076e-06, 6.465613e-08, 7.18989e-07, 1.308058e-06, 
    2.252149e-06, 1.449147e-06, 6.624782e-07, 3.078232e-07, 6.135131e-08, 
    1.592593e-08, 1.519428e-08, 2.71451e-08, 2.367835e-06, 6.383517e-07,
  2.443183e-08, 2.852222e-07, 6.436887e-07, 7.512976e-07, 1.767919e-06, 
    4.53585e-06, 4.934352e-06, 2.598274e-06, 3.377154e-07, 6.104729e-08, 
    2.874267e-08, 2.004395e-07, 6.189438e-07, 8.519417e-06, 1.698593e-06,
  2.919566e-08, 2.056745e-06, 7.135953e-07, 5.225708e-07, 8.247655e-06, 
    2.746725e-05, 2.341207e-05, 9.793122e-06, 1.627368e-07, 5.68498e-08, 
    2.689813e-08, 5.005784e-07, 6.633144e-06, 9.899597e-06, 4.630255e-07,
  2.492086e-06, 1.445285e-06, 1.32255e-06, 1.30933e-06, 1.361009e-05, 
    1.641345e-05, 1.344745e-05, 4.233977e-07, 8.303366e-08, 3.112811e-08, 
    8.834125e-08, 1.700954e-07, 4.930764e-06, 1.09925e-05, 4.715052e-06,
  8.024724e-09, 1.664663e-08, 2.549251e-08, 4.783089e-08, 1.042589e-07, 
    1.88443e-07, 1.044645e-05, 6.395768e-06, 3.875058e-05, 3.900464e-05, 
    3.110576e-05, 2.109109e-05, 1.022313e-05, 4.812726e-06, 8.612724e-08,
  1.647198e-08, 2.713834e-08, 5.117349e-08, 1.492238e-07, 1.571293e-06, 
    9.709856e-06, 2.067599e-05, 2.233486e-05, 2.457573e-05, 1.862695e-05, 
    2.419596e-05, 2.570249e-05, 1.620392e-05, 6.191886e-06, 1.108497e-07,
  4.50949e-08, 1.630847e-06, 6.129666e-07, 8.74402e-07, 1.448684e-05, 
    1.502677e-05, 1.719876e-05, 1.969812e-05, 1.968946e-05, 1.302026e-05, 
    1.888648e-05, 1.803457e-05, 1.041349e-05, 2.908969e-06, 2.396234e-07,
  6.962318e-06, 2.548022e-07, 4.658486e-06, 1.370207e-05, 1.33637e-05, 
    1.327984e-05, 2.002885e-05, 2.386064e-05, 1.901089e-05, 9.151719e-06, 
    1.405861e-05, 9.947058e-06, 5.439617e-06, 2.283337e-06, 2.201564e-06,
  3.197679e-06, 3.69873e-06, 6.211005e-06, 9.082672e-06, 7.982776e-06, 
    8.594267e-06, 1.731759e-05, 2.218508e-05, 2.004211e-05, 1.210019e-05, 
    2.814039e-07, 4.315397e-07, 5.176766e-06, 8.788136e-07, 1.740312e-06,
  1.091412e-06, 5.58637e-06, 8.112264e-06, 1.009222e-05, 8.391856e-06, 
    4.469842e-06, 3.414602e-06, 5.42119e-06, 8.792021e-06, 5.183609e-07, 
    6.250347e-06, 5.588121e-06, 1.984198e-06, 8.277773e-07, 1.745814e-05,
  8.565572e-06, 7.053827e-06, 3.036382e-06, 6.371296e-06, 4.24461e-06, 
    1.124803e-05, 1.259118e-05, 1.728381e-05, 2.394604e-05, 6.54575e-06, 
    2.482341e-06, 2.73288e-06, 2.13557e-06, 3.992199e-06, 5.60633e-06,
  1.231138e-05, 1.730036e-05, 1.318332e-05, 1.266615e-05, 2.132921e-05, 
    3.277458e-05, 3.093353e-05, 4.006039e-05, 4.468695e-05, 6.582085e-06, 
    6.232642e-07, 4.586954e-07, 6.88443e-07, 3.579555e-06, 2.041577e-07,
  1.854946e-05, 2.137614e-05, 1.818635e-05, 3.061451e-05, 4.765981e-05, 
    5.455373e-05, 4.599491e-05, 4.713455e-05, 9.144117e-07, 1.480538e-07, 
    1.532459e-07, 2.382136e-07, 3.355596e-07, 1.519082e-07, 5.286848e-08,
  2.371533e-05, 2.714983e-05, 2.809086e-05, 5.347823e-05, 7.578077e-05, 
    3.467813e-05, 2.225751e-05, 7.805627e-07, 1.278487e-07, 1.052911e-07, 
    9.548739e-08, 8.146545e-08, 4.698305e-08, 8.756309e-08, 4.152672e-08,
  1.062756e-08, 7.685374e-09, 9.91358e-09, 9.964855e-09, 3.138123e-07, 
    1.600822e-08, 8.810925e-06, 1.798736e-05, 4.491136e-05, 6.743355e-05, 
    8.277218e-05, 9.369031e-05, 7.632418e-05, 2.269323e-05, 1.177871e-05,
  1.782365e-06, 1.916572e-08, 4.339557e-09, 4.717818e-09, 1.525062e-08, 
    1.227407e-06, 8.412984e-06, 1.583268e-05, 2.558707e-05, 4.512391e-05, 
    6.102159e-05, 6.435908e-05, 4.497181e-05, 1.524733e-05, 1.573171e-05,
  6.905658e-06, 1.079606e-06, 1.18607e-07, 1.713346e-07, 9.00806e-07, 
    4.065484e-07, 3.071803e-06, 4.644281e-06, 3.187043e-06, 3.664978e-06, 
    7.781945e-06, 1.086075e-05, 4.728482e-06, 6.905195e-06, 6.11451e-07,
  1.335685e-05, 6.342016e-06, 5.926336e-06, 1.036441e-05, 3.621785e-06, 
    6.606228e-06, 5.144906e-06, 4.263123e-06, 6.299106e-06, 1.692998e-05, 
    3.344562e-05, 3.078667e-05, 1.20305e-05, 1.579007e-05, 4.066991e-06,
  2.270283e-05, 6.503737e-06, 4.321575e-06, 3.963677e-06, 5.496887e-06, 
    3.218093e-06, 6.271216e-06, 7.53922e-06, 2.009567e-05, 3.954205e-05, 
    6.639194e-06, 1.191576e-05, 2.692879e-05, 1.869818e-05, 1.019811e-05,
  1.894126e-05, 1.087789e-05, 5.871328e-06, 9.116332e-06, 8.029367e-06, 
    7.187503e-06, 3.634215e-06, 6.939795e-06, 2.195792e-05, 6.929247e-06, 
    2.41658e-05, 1.714033e-05, 1.06152e-05, 4.120731e-05, 1.566024e-05,
  1.236255e-05, 8.211911e-06, 8.957791e-06, 9.587316e-06, 9.815702e-06, 
    9.126424e-06, 8.662222e-06, 1.480963e-05, 1.581211e-05, 4.001875e-06, 
    4.916043e-07, 3.969195e-07, 9.225155e-07, 2.880762e-05, 1.039478e-05,
  9.035194e-06, 1.058123e-05, 1.4556e-05, 1.800262e-05, 2.340608e-05, 
    2.990703e-05, 1.078089e-05, 6.021319e-06, 7.089535e-06, 5.822816e-08, 
    8.702953e-09, 8.420018e-09, 8.00051e-09, 1.07585e-05, 8.120496e-07,
  1.300841e-05, 1.121956e-05, 2.400535e-05, 3.942029e-05, 4.16062e-05, 
    4.03695e-05, 1.595343e-05, 5.297289e-06, 4.694559e-08, 1.453178e-08, 
    3.009836e-07, 5.824628e-08, 1.469546e-08, 8.920964e-08, 5.857508e-08,
  4.443195e-06, 2.201498e-06, 2.648326e-05, 3.167982e-05, 2.582402e-05, 
    8.89166e-06, 7.9109e-06, 7.773062e-07, 5.763252e-07, 1.236839e-06, 
    1.686973e-06, 4.207007e-07, 3.343901e-07, 9.429625e-07, 1.51007e-06,
  4.151506e-05, 3.900773e-05, 2.785448e-05, 1.098798e-05, 3.287819e-06, 
    6.00198e-07, 3.878838e-07, 1.277332e-07, 1.051315e-05, 2.045419e-05, 
    1.726119e-05, 3.117832e-05, 4.825435e-05, 3.185719e-05, 5.22787e-05,
  4.171267e-05, 3.973948e-05, 8.906075e-06, 8.586201e-06, 1.444396e-06, 
    2.27383e-06, 9.646018e-07, 3.747462e-07, 7.4331e-06, 1.319465e-05, 
    8.688945e-06, 1.629338e-05, 2.011385e-05, 6.407238e-06, 2.008598e-05,
  0.0001755057, 9.150445e-05, 2.528726e-05, 7.836674e-06, 2.141464e-05, 
    7.226364e-06, 1.194944e-07, 7.098149e-08, 3.044608e-06, 7.716877e-06, 
    8.059604e-06, 8.290292e-06, 8.528488e-06, 4.026873e-06, 8.444549e-06,
  0.0001249262, 5.02565e-05, 4.27233e-05, 2.971943e-05, 1.330669e-05, 
    8.978674e-06, 6.595086e-06, 2.929303e-06, 1.690622e-06, 2.263318e-06, 
    2.079268e-06, 2.498159e-06, 4.77645e-06, 4.740249e-06, 4.307782e-06,
  0.0001586897, 0.0001030051, 6.473774e-05, 2.54277e-05, 4.366476e-06, 
    3.200008e-06, 2.258971e-06, 1.633609e-06, 2.422447e-06, 8.922051e-06, 
    1.966195e-06, 3.347771e-06, 4.675646e-07, 2.796799e-06, 1.194523e-06,
  0.000180053, 0.00017479, 0.0001260264, 2.557075e-05, 3.133608e-06, 
    1.451527e-06, 1.926822e-06, 5.116572e-07, 1.908724e-06, 4.916696e-07, 
    2.077379e-06, 1.296492e-07, 1.379947e-06, 7.183238e-06, 2.724074e-06,
  0.0001311093, 0.0001333237, 7.729889e-05, 4.269588e-06, 2.625649e-06, 
    3.584129e-06, 2.010061e-06, 2.056129e-06, 1.124894e-06, 3.071503e-06, 
    3.172856e-07, 2.904709e-08, 1.472789e-06, 6.527775e-06, 2.2305e-06,
  4.336616e-05, 6.191141e-05, 2.201605e-05, 1.033314e-05, 1.103775e-05, 
    9.034177e-06, 1.768968e-06, 2.957712e-06, 5.402702e-06, 1.590185e-06, 
    2.310151e-06, 7.80912e-07, 2.458651e-08, 7.215759e-06, 1.089303e-07,
  1.173783e-05, 3.043178e-05, 1.468016e-05, 1.392963e-05, 2.372289e-05, 
    2.219184e-05, 7.677025e-06, 2.327217e-06, 8.921311e-07, 3.841846e-06, 
    4.561188e-06, 1.089784e-06, 1.413792e-08, 1.302233e-07, 3.969734e-08,
  6.504631e-08, 8.178319e-07, 1.11487e-05, 7.407331e-06, 7.49922e-06, 
    2.821424e-06, 2.675864e-06, 2.038055e-06, 9.091856e-06, 6.826584e-06, 
    5.327287e-06, 4.281594e-06, 1.335666e-06, 2.104895e-06, 3.696541e-06,
  2.02178e-05, 6.264736e-05, 0.000100548, 0.000130078, 0.0001262796, 
    0.000107738, 0.0001060714, 9.277536e-05, 0.0001286643, 9.468232e-05, 
    5.68151e-05, 4.222095e-05, 4.4547e-05, 4.487109e-05, 3.443983e-05,
  7.961381e-06, 5.972431e-05, 0.000142794, 0.0001582717, 0.000153942, 
    0.0001122248, 9.138395e-05, 9.088411e-05, 8.179209e-05, 6.163876e-05, 
    3.771281e-05, 1.850967e-05, 2.104463e-05, 2.897096e-05, 2.191294e-05,
  3.636086e-05, 9.572813e-05, 0.0001594076, 0.000163575, 0.000142266, 
    0.0001022869, 7.801679e-05, 6.783084e-05, 4.29485e-05, 2.536384e-05, 
    1.203107e-05, 5.659304e-06, 9.100914e-06, 1.52793e-05, 2.360869e-05,
  4.069067e-05, 3.962106e-05, 6.134825e-05, 0.000122283, 0.0001018294, 
    9.119067e-05, 8.292227e-05, 5.209511e-05, 1.833364e-05, 7.649702e-06, 
    4.519649e-06, 9.774603e-07, 3.305875e-06, 5.785479e-06, 3.154972e-05,
  3.624071e-05, 4.754637e-05, 5.013295e-05, 0.000100933, 0.0001231798, 
    0.0001144379, 8.767067e-05, 5.345262e-05, 2.009748e-05, 7.00604e-06, 
    9.015123e-07, 4.828055e-08, 1.229498e-06, 3.688382e-08, 9.032181e-06,
  1.763963e-05, 2.702938e-05, 8.689473e-05, 0.0001438356, 0.0001434195, 
    0.0001092362, 8.033769e-05, 4.735284e-05, 4.201329e-05, 8.489936e-06, 
    3.539755e-06, 3.825033e-07, 1.190406e-08, 2.79937e-08, 1.484546e-05,
  5.28414e-06, 1.139015e-05, 2.9406e-05, 2.144355e-05, 5.422909e-06, 
    2.865431e-06, 8.454947e-07, 8.18847e-06, 3.34216e-06, 2.430104e-06, 
    3.47905e-08, 2.843573e-08, 1.04404e-09, 1.721991e-07, 3.362542e-06,
  5.245502e-06, 5.411551e-06, 4.124337e-06, 1.045409e-06, 1.441906e-06, 
    2.690267e-07, 1.265256e-07, 1.53853e-06, 3.736307e-06, 5.050648e-07, 
    7.891047e-07, 2.711124e-06, 2.431261e-09, 2.651183e-06, 1.031201e-07,
  4.995968e-07, 5.974278e-06, 4.600163e-06, 5.587077e-06, 4.647522e-06, 
    4.878106e-06, 2.975972e-06, 1.154792e-05, 1.782926e-06, 3.097367e-06, 
    3.407891e-06, 8.626458e-07, 1.37233e-06, 2.947815e-07, 7.462065e-08,
  2.855884e-07, 1.30745e-06, 5.838227e-06, 6.595403e-06, 1.056128e-05, 
    6.40409e-06, 6.177976e-06, 3.526689e-06, 5.614972e-06, 5.735093e-06, 
    2.625939e-06, 2.259938e-06, 1.023065e-06, 5.73082e-07, 5.270155e-07,
  1.623527e-05, 1.541543e-05, 4.149217e-05, 1.786924e-05, 5.599935e-06, 
    7.730819e-06, 1.633941e-05, 2.399978e-05, 6.382016e-05, 7.099532e-05, 
    6.006606e-05, 0.0001206993, 0.0001002671, 7.139931e-05, 4.837237e-05,
  2.774963e-06, 1.239123e-05, 1.922233e-05, 5.026556e-06, 1.180429e-06, 
    1.669621e-06, 6.391746e-06, 1.309836e-05, 2.933116e-05, 4.899423e-05, 
    8.188812e-05, 9.359067e-05, 9.190568e-05, 3.341631e-05, 2.778678e-05,
  2.568853e-05, 1.174703e-05, 7.510631e-08, 1.729189e-07, 4.326093e-07, 
    3.274001e-07, 2.609098e-06, 6.885087e-06, 1.561216e-05, 2.981625e-05, 
    5.467963e-05, 5.952713e-05, 3.050919e-05, 1.36769e-05, 6.809287e-07,
  5.929977e-05, 6.220819e-06, 3.601432e-06, 3.48387e-06, 3.308752e-06, 
    7.530967e-06, 8.203566e-06, 7.165179e-06, 1.25648e-05, 9.259073e-06, 
    2.388227e-05, 2.058451e-05, 1.412307e-05, 1.869693e-05, 1.2248e-06,
  4.703539e-05, 6.657258e-06, 1.195811e-06, 1.168122e-06, 1.505928e-06, 
    3.28835e-06, 5.589583e-06, 9.36551e-06, 1.198964e-05, 2.115585e-05, 
    2.67184e-05, 1.15216e-05, 1.155558e-05, 3.848398e-06, 3.307589e-06,
  3.736091e-06, 5.737005e-06, 2.198947e-06, 3.259835e-06, 1.092393e-07, 
    1.637451e-06, 2.231585e-06, 4.455028e-06, 2.102246e-05, 1.859897e-05, 
    2.011865e-05, 8.673332e-06, 3.478169e-06, 6.98225e-06, 3.674997e-06,
  5.402035e-06, 6.477193e-06, 1.77481e-06, 1.777941e-06, 2.204818e-07, 
    3.073521e-07, 1.656531e-06, 3.752652e-06, 5.524835e-06, 4.230713e-06, 
    4.056013e-06, 6.399008e-06, 3.442284e-07, 1.374927e-05, 8.352034e-07,
  4.516837e-07, 2.745685e-06, 1.85823e-06, 7.773532e-07, 8.146193e-07, 
    9.270074e-09, 4.652594e-07, 3.851032e-06, 9.019495e-06, 7.151426e-06, 
    8.759806e-06, 1.143842e-05, 3.370929e-06, 1.605604e-05, 2.032284e-07,
  8.014272e-08, 2.289352e-07, 8.757334e-07, 2.99615e-06, 3.281223e-06, 
    6.987336e-08, 9.955435e-07, 2.510183e-06, 1.843221e-06, 7.070876e-06, 
    7.423666e-06, 1.012351e-05, 8.817119e-06, 9.113153e-07, 5.38134e-07,
  1.688546e-08, 2.194116e-07, 8.892808e-07, 5.672146e-07, 2.078749e-06, 
    7.548896e-07, 1.514035e-07, 1.907331e-06, 7.634221e-06, 5.887253e-06, 
    6.683181e-06, 6.496696e-06, 6.922266e-06, 4.236378e-06, 6.492953e-06,
  8.39209e-05, 2.050798e-05, 4.854831e-05, 4.562697e-05, 3.025657e-06, 
    1.618029e-06, 1.263632e-06, 3.937149e-07, 6.735446e-06, 1.11513e-05, 
    8.89885e-06, 1.093675e-05, 2.114102e-05, 4.838064e-05, 1.269292e-05,
  5.46025e-05, 5.876552e-05, 7.519196e-05, 4.506195e-05, 1.754917e-05, 
    1.420487e-05, 5.977344e-06, 4.381101e-06, 1.436721e-05, 8.691688e-06, 
    2.567484e-06, 2.731168e-06, 8.836687e-06, 2.199664e-05, 4.6461e-06,
  0.0001390468, 9.878242e-05, 5.867593e-05, 6.073802e-05, 9.151758e-05, 
    3.471935e-05, 1.000307e-05, 1.795515e-05, 2.003807e-05, 5.98097e-06, 
    6.941187e-07, 3.525911e-07, 3.505637e-07, 1.177705e-06, 4.336565e-07,
  0.0001762828, 7.280908e-05, 6.35032e-05, 0.0001035529, 6.189929e-05, 
    5.210402e-05, 3.408895e-05, 3.075464e-05, 1.707163e-05, 4.256686e-06, 
    3.062503e-06, 1.605388e-06, 8.636538e-07, 8.608024e-07, 2.922615e-07,
  0.0001501912, 8.310904e-05, 3.971604e-05, 4.243998e-05, 3.317626e-05, 
    3.35846e-05, 2.178675e-05, 1.621275e-05, 8.501273e-06, 3.511412e-06, 
    1.6151e-08, 3.660585e-07, 1.315435e-06, 1.025572e-06, 2.006537e-06,
  7.457526e-05, 6.847102e-05, 2.868457e-05, 4.424984e-05, 3.681918e-05, 
    2.264225e-05, 4.826052e-06, 5.800908e-07, 1.316045e-06, 8.801662e-08, 
    5.088095e-06, 2.066476e-06, 4.184878e-07, 3.685251e-07, 2.413884e-06,
  7.310819e-05, 8.481326e-05, 9.001883e-05, 0.000105372, 6.187025e-05, 
    1.198406e-05, 1.023561e-06, 5.146848e-06, 1.467965e-05, 4.400235e-06, 
    1.860152e-06, 1.524302e-06, 2.570252e-06, 4.933416e-06, 1.332461e-06,
  0.0001084995, 0.0001431179, 0.0001404397, 9.237989e-05, 3.181442e-05, 
    5.263145e-06, 6.815996e-07, 7.984729e-06, 1.972515e-05, 5.582815e-06, 
    3.059545e-06, 1.671822e-06, 1.918867e-06, 9.138021e-06, 2.044386e-07,
  0.0001575547, 0.0001376372, 8.478687e-05, 3.047049e-05, 4.593825e-06, 
    1.251684e-06, 3.202941e-06, 9.368867e-06, 4.339603e-06, 5.382379e-06, 
    2.838902e-06, 3.323337e-06, 2.559498e-06, 5.32506e-07, 6.957308e-07,
  7.22222e-05, 2.979012e-05, 7.758955e-06, 2.820563e-06, 6.040646e-06, 
    4.823199e-06, 1.19935e-05, 4.66031e-06, 2.588494e-06, 2.109487e-06, 
    4.722524e-06, 4.68323e-06, 2.993267e-06, 2.451478e-06, 4.45333e-06,
  6.038678e-05, 0.0001701065, 0.0002210978, 0.0001580403, 0.0001191709, 
    0.0001388503, 0.0002068905, 0.0001737595, 0.0002428576, 0.0001640851, 
    6.076548e-05, 2.750051e-05, 2.078236e-05, 4.420171e-05, 7.035225e-06,
  1.521397e-05, 4.632449e-05, 0.0001210991, 0.000165465, 0.0001266813, 
    0.0001327803, 0.0001534719, 0.0001736323, 0.0002273875, 0.0001488521, 
    8.069906e-05, 4.750052e-05, 4.582692e-05, 8.758617e-05, 1.440263e-05,
  5.03022e-05, 5.323525e-05, 5.141791e-05, 0.0001280753, 0.0001409448, 
    0.000123892, 0.0001112, 0.0002005074, 0.0002456585, 0.0001876759, 
    0.0001490135, 0.0001390194, 0.0001300003, 0.0001197714, 0.0001150278,
  3.396368e-05, 4.287974e-05, 5.789904e-05, 0.0001002681, 8.373676e-05, 
    9.984239e-05, 0.0001188755, 0.0002010279, 0.0002097569, 0.0001912936, 
    0.0002003952, 0.0001711043, 0.0001364649, 0.000122884, 5.165951e-05,
  8.675814e-06, 1.938734e-05, 3.238086e-05, 5.227787e-05, 6.68055e-05, 
    9.370747e-05, 0.0001278179, 0.0001605362, 0.0001871329, 0.0002348654, 
    0.000140568, 9.501456e-05, 0.0001160396, 4.522208e-05, 2.324692e-05,
  3.70483e-06, 1.555277e-05, 2.200859e-05, 4.809002e-05, 0.0001333856, 
    0.0001883044, 0.000209697, 0.0001847674, 0.0002156395, 0.0001202722, 
    4.246434e-05, 2.338186e-05, 2.054916e-05, 3.14383e-05, 4.085573e-05,
  1.367331e-05, 1.309107e-05, 2.420151e-05, 8.062857e-05, 0.0001655332, 
    0.0001780978, 0.0001167667, 9.157485e-05, 9.361425e-05, 1.256099e-05, 
    1.337293e-06, 5.541574e-07, 1.277646e-07, 1.527503e-05, 1.607567e-05,
  8.124927e-06, 1.065828e-05, 3.294724e-05, 5.130224e-05, 4.48031e-05, 
    2.388804e-05, 1.089453e-05, 2.059651e-05, 5.010664e-05, 1.085697e-05, 
    4.896983e-06, 3.52618e-06, 1.217681e-08, 6.550564e-06, 7.27441e-06,
  1.261113e-06, 3.54435e-06, 1.105081e-05, 1.61997e-05, 1.660747e-05, 
    2.515691e-05, 3.151584e-05, 5.55866e-05, 2.304595e-05, 1.194863e-05, 
    9.39824e-06, 8.254791e-06, 3.916709e-07, 6.535638e-06, 9.509241e-06,
  8.186872e-08, 2.988332e-06, 1.604636e-05, 2.091034e-05, 2.770078e-05, 
    3.250978e-05, 3.585791e-05, 2.045228e-05, 1.635224e-05, 1.654805e-05, 
    1.557186e-05, 1.535604e-05, 3.997587e-06, 5.743023e-06, 5.308931e-06,
  3.710335e-07, 3.867021e-07, 5.81308e-07, 5.504371e-08, 4.464521e-09, 
    3.258739e-08, 1.555664e-06, 1.932932e-05, 6.119815e-05, 0.0001181312, 
    9.446044e-05, 9.08349e-05, 0.0001034522, 6.336082e-05, 4.753167e-05,
  1.297315e-07, 3.852511e-10, 4.439957e-11, 2.060815e-09, 2.981274e-09, 
    1.509449e-08, 1.074324e-06, 2.333925e-06, 2.492188e-05, 6.494841e-05, 
    5.212841e-05, 5.112555e-05, 4.115103e-05, 1.981163e-05, 1.162196e-05,
  8.312813e-08, 5.641318e-09, 8.528016e-09, 7.843115e-09, 1.776765e-08, 
    6.635639e-08, 1.124952e-07, 1.394317e-06, 7.796389e-06, 2.205029e-05, 
    3.65757e-05, 4.053628e-05, 2.30002e-05, 1.898221e-05, 7.87927e-06,
  1.273032e-09, 4.287421e-08, 4.535578e-07, 1.679946e-06, 9.551638e-07, 
    3.95716e-06, 5.606677e-06, 2.860262e-06, 2.563977e-06, 1.149265e-05, 
    2.80034e-05, 3.389277e-05, 1.210556e-05, 2.074605e-05, 4.659605e-06,
  3.25563e-08, 2.517326e-06, 1.533116e-06, 2.997974e-06, 1.200228e-06, 
    1.8629e-06, 7.961209e-06, 1.366458e-05, 1.456613e-05, 3.721357e-05, 
    2.588094e-06, 8.041526e-06, 2.845988e-05, 2.123817e-05, 3.211193e-06,
  1.511897e-07, 4.950859e-06, 4.754465e-06, 2.592659e-06, 4.888015e-06, 
    4.749675e-06, 4.405404e-06, 1.087475e-05, 1.735712e-05, 5.187011e-06, 
    4.428431e-06, 3.229556e-06, 5.485883e-06, 2.654314e-05, 9.739681e-06,
  2.021937e-08, 2.257555e-06, 3.255929e-06, 3.178583e-06, 3.821259e-06, 
    6.228172e-06, 6.820967e-06, 1.550129e-05, 8.999396e-06, 3.010396e-06, 
    1.892349e-06, 1.367167e-06, 3.198882e-06, 4.059932e-05, 9.404773e-06,
  1.6721e-08, 1.610993e-06, 3.197689e-06, 1.89801e-06, 5.149531e-06, 
    3.571688e-06, 5.896562e-06, 9.778875e-06, 1.698341e-05, 2.020996e-06, 
    2.45811e-06, 1.533933e-07, 3.936785e-08, 1.852106e-05, 2.006077e-06,
  1.414147e-09, 7.745909e-08, 8.930083e-07, 2.187149e-06, 3.576979e-06, 
    8.90636e-06, 1.190468e-05, 7.61175e-06, 8.221264e-07, 4.817058e-06, 
    4.241957e-06, 2.250507e-06, 4.298892e-09, 1.302803e-07, 5.549327e-08,
  4.319212e-10, 7.555202e-08, 2.748671e-06, 2.621169e-06, 6.887353e-06, 
    7.438639e-06, 5.395151e-06, 2.033672e-06, 1.581632e-06, 4.033554e-06, 
    4.995921e-06, 4.831899e-06, 9.61091e-08, 3.870851e-09, 1.550992e-08,
  5.26597e-08, 1.055651e-06, 3.203654e-06, 9.870729e-09, 1.324875e-08, 
    6.187421e-07, 1.725872e-06, 6.627712e-07, 5.124038e-06, 1.637601e-05, 
    2.169713e-05, 5.04479e-05, 3.453666e-05, 1.776536e-05, 3.043519e-05,
  6.341061e-09, 9.829664e-10, 1.97462e-07, 8.231222e-11, 2.684655e-09, 
    5.210926e-07, 1.514406e-06, 1.349601e-06, 1.071594e-05, 1.262899e-05, 
    1.205039e-05, 2.778849e-05, 1.830179e-05, 8.516422e-06, 1.797542e-05,
  1.165325e-08, 2.945853e-10, 2.048447e-10, 1.160256e-10, 5.584871e-08, 
    2.040104e-08, 5.540266e-09, 2.162537e-08, 4.005392e-06, 1.042764e-05, 
    1.479969e-05, 2.096111e-05, 2.696901e-05, 1.843438e-05, 8.682468e-06,
  1.721402e-07, 6.870731e-09, 1.551054e-09, 3.389506e-09, 3.091281e-09, 
    4.485234e-09, 6.917129e-08, 2.140834e-07, 1.303697e-06, 3.483408e-06, 
    4.537208e-06, 3.200518e-06, 8.868221e-06, 1.555814e-05, 1.668026e-05,
  2.730044e-10, 4.792664e-10, 1.316193e-09, 6.050445e-09, 1.004892e-08, 
    5.421324e-09, 1.943839e-09, 5.896167e-07, 1.827861e-06, 6.971444e-06, 
    1.331967e-08, 5.498818e-09, 1.342657e-06, 5.621437e-07, 8.864329e-06,
  2.674713e-10, 5.591967e-10, 1.018134e-09, 5.761828e-09, 1.712472e-08, 
    2.423548e-08, 1.127317e-08, 8.126634e-08, 3.130898e-08, 3.506717e-08, 
    4.166008e-07, 1.174727e-07, 1.619842e-09, 4.767102e-08, 1.209822e-05,
  4.800833e-10, 8.189658e-10, 4.265565e-10, 1.254445e-09, 2.710543e-09, 
    8.480554e-08, 4.437828e-08, 4.998545e-11, 9.91318e-08, 1.36954e-07, 
    1.045267e-07, 7.616978e-08, 7.904537e-09, 2.250604e-07, 3.765401e-06,
  5.678994e-10, 1.452983e-09, 1.727916e-09, 1.489321e-08, 1.833524e-09, 
    1.324035e-07, 3.603242e-08, 5.253333e-10, 3.009764e-09, 2.571824e-08, 
    2.920253e-08, 6.262513e-08, 9.625284e-07, 1.943789e-06, 8.367157e-08,
  3.820742e-10, 2.019403e-09, 3.465809e-09, 2.064259e-09, 4.257837e-09, 
    3.723385e-08, 5.710721e-08, 7.775327e-08, 1.169988e-09, 2.397062e-08, 
    1.06405e-08, 3.514117e-08, 2.780485e-08, 1.18152e-07, 2.714768e-09,
  1.352336e-10, 1.932324e-09, 4.220873e-09, 3.086632e-09, 3.178256e-09, 
    1.273913e-09, 2.319557e-08, 2.083464e-09, 2.057841e-09, 9.365722e-08, 
    2.618903e-08, 3.246132e-07, 6.261147e-08, 4.395581e-09, 4.7205e-11,
  4.128496e-08, 5.93208e-07, 1.703667e-06, 9.606175e-07, 2.42772e-07, 
    6.956056e-08, 6.680648e-07, 5.287677e-08, 3.087425e-08, 3.880461e-06, 
    1.173472e-05, 5.060106e-05, 3.009349e-05, 1.867619e-05, 5.234067e-05,
  1.464444e-10, 1.558006e-10, 8.018123e-07, 1.674238e-08, 2.024446e-09, 
    7.911987e-09, 9.269171e-08, 1.914857e-07, 6.934837e-09, 3.045257e-07, 
    4.416857e-06, 2.170991e-05, 2.01892e-05, 1.874181e-05, 3.572496e-05,
  1.326001e-09, 4.048313e-10, 8.249057e-09, 1.519691e-09, 4.628103e-08, 
    5.972119e-08, 3.285794e-08, 8.675759e-09, 1.18856e-09, 2.100948e-08, 
    6.050736e-07, 4.095835e-06, 1.821068e-05, 1.480833e-05, 1.058999e-05,
  1.047988e-06, 4.330925e-07, 6.27875e-07, 2.752689e-08, 2.418103e-08, 
    1.583183e-07, 4.761686e-07, 1.122469e-07, 6.631492e-09, 2.031966e-09, 
    6.534149e-07, 8.912447e-08, 2.031668e-06, 5.911435e-06, 5.534359e-06,
  2.490585e-06, 2.40782e-06, 8.968048e-07, 3.682525e-07, 3.812792e-08, 
    9.30433e-08, 6.515619e-07, 1.722898e-06, 1.372463e-07, 1.760911e-09, 
    6.332264e-09, 7.434748e-10, 3.998156e-06, 1.143548e-06, 7.174256e-06,
  7.098469e-07, 5.151244e-06, 1.069926e-07, 2.465631e-07, 5.203871e-08, 
    1.104048e-07, 1.477135e-07, 1.021475e-07, 3.222432e-08, 7.646655e-10, 
    4.935111e-10, 1.357632e-10, 4.450433e-09, 4.61617e-07, 2.63256e-05,
  4.117328e-08, 3.243116e-07, 4.400554e-07, 7.987823e-07, 2.523211e-07, 
    4.927907e-08, 1.255321e-07, 7.252462e-08, 6.709731e-09, 8.060173e-09, 
    6.887892e-09, 2.338609e-09, 1.636639e-09, 3.668186e-06, 1.450048e-05,
  3.609287e-08, 1.445348e-07, 1.293051e-06, 3.679633e-06, 1.613794e-06, 
    2.623188e-06, 1.269759e-07, 4.031455e-08, 6.249355e-09, 2.793241e-08, 
    1.648847e-08, 4.461134e-09, 2.475492e-09, 3.572397e-06, 2.325676e-07,
  5.457994e-08, 1.052849e-07, 1.030311e-06, 7.785983e-06, 1.564753e-05, 
    1.190918e-05, 7.342569e-06, 7.501561e-08, 8.338398e-09, 3.348358e-08, 
    2.9209e-08, 8.692723e-09, 1.42601e-09, 9.31989e-08, 8.466776e-09,
  5.886989e-08, 1.038336e-07, 1.570988e-06, 4.207982e-06, 1.260172e-05, 
    9.441068e-06, 1.360338e-06, 4.485345e-09, 8.720297e-09, 3.53501e-08, 
    1.094188e-08, 1.773993e-08, 6.482115e-09, 6.468139e-10, 2.573961e-10,
  2.468513e-06, 2.412841e-05, 6.203893e-05, 4.376704e-05, 1.862258e-05, 
    3.247801e-06, 1.199427e-07, 3.162497e-10, 3.686316e-08, 2.358527e-07, 
    3.078432e-06, 1.700707e-05, 1.243736e-05, 1.052541e-05, 2.686688e-05,
  5.705392e-06, 1.580406e-05, 6.515664e-05, 8.798573e-05, 3.857989e-05, 
    1.440609e-05, 2.258847e-06, 5.095472e-09, 2.204853e-08, 8.234763e-08, 
    1.047914e-06, 4.174189e-06, 1.073423e-06, 2.539736e-06, 9.408281e-06,
  5.305431e-05, 6.183526e-05, 5.407034e-05, 8.961622e-05, 7.518724e-05, 
    1.630522e-05, 5.194542e-06, 2.570225e-06, 4.692546e-07, 2.298893e-07, 
    1.338896e-06, 1.089039e-07, 8.795826e-08, 4.834408e-07, 1.204839e-07,
  4.848632e-05, 2.114167e-05, 0.0001070806, 0.0001650056, 8.93948e-05, 
    4.305585e-05, 1.391945e-05, 1.060534e-05, 3.702211e-06, 6.248647e-07, 
    2.87969e-07, 9.118595e-08, 1.007961e-06, 8.6762e-07, 1.801323e-08,
  5.325228e-05, 2.611817e-05, 8.356119e-05, 0.0001748727, 0.0001176005, 
    6.587372e-05, 1.972711e-05, 1.17391e-05, 9.741006e-06, 2.931528e-06, 
    5.286796e-09, 6.790665e-10, 9.017431e-09, 4.4071e-09, 5.726189e-08,
  3.564476e-05, 4.540611e-05, 0.0001064595, 0.0001923757, 0.000172411, 
    9.27931e-05, 3.138561e-05, 7.385641e-06, 4.934261e-06, 1.837532e-08, 
    7.701154e-10, 1.804676e-10, 1.270479e-11, 4.056527e-09, 3.737833e-07,
  3.086341e-05, 6.405979e-05, 0.0001276553, 0.0001923376, 0.000142669, 
    8.985523e-05, 4.248559e-05, 7.115627e-06, 1.087832e-05, 1.799865e-06, 
    5.916397e-08, 1.274939e-10, 5.420428e-09, 1.235113e-06, 2.832585e-07,
  3.719132e-05, 8.115047e-05, 9.832062e-05, 0.0001106318, 9.370111e-05, 
    8.426238e-05, 4.923114e-05, 1.36843e-05, 1.282905e-05, 4.263693e-06, 
    2.545911e-06, 6.972529e-10, 1.123579e-09, 6.666879e-07, 5.579183e-08,
  3.905951e-05, 5.693613e-05, 6.802153e-05, 7.910829e-05, 9.533506e-05, 
    9.851078e-05, 6.685383e-05, 3.427635e-05, 7.931876e-06, 1.701647e-05, 
    1.074061e-05, 9.995497e-08, 7.028688e-10, 2.597864e-08, 1.653157e-08,
  3.582093e-05, 4.552564e-05, 5.759688e-05, 6.274284e-05, 6.269716e-05, 
    9.607339e-05, 9.760705e-05, 3.713029e-05, 3.555405e-05, 3.470193e-05, 
    3.154178e-05, 8.256113e-06, 2.161457e-09, 2.301918e-09, 4.232578e-09,
  3.151994e-10, 3.504111e-09, 3.920169e-06, 1.197025e-05, 2.278508e-05, 
    2.433157e-05, 2.203939e-05, 1.499104e-05, 2.516805e-05, 1.896065e-05, 
    1.328758e-05, 1.350016e-05, 6.207264e-06, 4.139386e-06, 4.911665e-07,
  4.970999e-10, 5.058894e-09, 6.747783e-07, 1.249989e-05, 1.924962e-05, 
    2.619341e-05, 3.087873e-05, 2.848449e-05, 3.380206e-05, 3.406017e-05, 
    2.654161e-05, 2.609643e-05, 1.621339e-05, 1.000677e-05, 2.379252e-06,
  3.793434e-07, 4.547879e-07, 2.133418e-07, 1.25531e-07, 1.12155e-05, 
    2.042084e-05, 2.989905e-05, 3.121021e-05, 4.046574e-05, 4.087875e-05, 
    4.717808e-05, 3.994018e-05, 2.398178e-05, 1.222162e-05, 6.182928e-07,
  2.119493e-07, 2.925704e-06, 9.697078e-06, 1.305629e-05, 1.523701e-05, 
    3.626484e-05, 4.547207e-05, 4.610359e-05, 4.292328e-05, 5.035846e-05, 
    0.0001250576, 0.0001076941, 5.760934e-05, 3.56106e-05, 7.739609e-06,
  1.652967e-07, 3.888448e-06, 5.386164e-06, 1.286011e-05, 1.357941e-05, 
    3.137159e-05, 4.632436e-05, 5.915818e-05, 5.89588e-05, 0.0001044239, 
    2.095678e-05, 5.209007e-05, 0.0001160556, 4.149747e-05, 3.216714e-05,
  1.118873e-06, 4.175537e-06, 7.183363e-06, 9.335598e-06, 8.479974e-06, 
    1.751326e-05, 3.604322e-05, 3.546717e-05, 6.780573e-05, 3.149624e-05, 
    4.121733e-05, 6.468111e-05, 4.283187e-05, 7.544197e-05, 2.792077e-05,
  3.671557e-06, 2.522891e-06, 5.856979e-06, 9.758634e-06, 1.235217e-05, 
    3.101675e-05, 2.516839e-05, 1.477981e-05, 1.562463e-05, 1.836955e-05, 
    2.225981e-05, 2.505609e-05, 2.311283e-05, 7.377223e-05, 1.783935e-05,
  1.027843e-06, 4.89069e-06, 6.017398e-06, 9.465973e-06, 1.464619e-05, 
    2.589629e-05, 2.021073e-05, 1.047179e-05, 4.866818e-06, 3.411594e-06, 
    1.150832e-05, 1.905542e-05, 3.145072e-05, 8.220832e-05, 2.618051e-06,
  7.072902e-07, 4.639186e-06, 7.524307e-06, 1.246832e-05, 3.711816e-05, 
    3.326575e-05, 3.594834e-05, 1.512836e-05, 5.381856e-08, 8.191483e-07, 
    4.093306e-06, 1.767863e-05, 3.489749e-05, 4.74501e-05, 3.554567e-06,
  1.430637e-07, 1.341502e-06, 6.303212e-06, 4.034672e-06, 1.579065e-05, 
    4.263377e-05, 2.231527e-05, 4.149729e-07, 5.722234e-09, 2.66255e-08, 
    2.353318e-06, 1.544914e-05, 3.026819e-05, 3.975365e-05, 2.506571e-05,
  1.944516e-09, 4.364702e-11, 7.756013e-07, 2.183816e-09, 9.951369e-09, 
    3.569624e-08, 2.051743e-07, 5.847096e-08, 8.38483e-07, 2.732571e-07, 
    9.510671e-07, 5.142781e-06, 4.209583e-06, 1.437477e-06, 1.477246e-06,
  7.685597e-09, 2.14447e-10, 1.987851e-10, 3.513922e-09, 1.81493e-08, 
    3.167867e-08, 2.528603e-07, 5.202212e-07, 3.460941e-06, 1.12611e-06, 
    2.590535e-07, 1.019241e-06, 1.696544e-06, 2.145374e-06, 3.117711e-06,
  7.760835e-07, 2.138951e-06, 5.780079e-07, 7.635534e-08, 5.189201e-07, 
    4.224167e-07, 2.633738e-07, 8.136297e-07, 1.175765e-05, 5.909527e-06, 
    1.864159e-06, 3.008166e-07, 1.896243e-07, 5.545157e-07, 1.96338e-07,
  9.212237e-07, 3.584053e-07, 5.226016e-07, 2.886013e-06, 3.046331e-06, 
    3.361164e-06, 2.59307e-06, 4.485387e-06, 1.112338e-05, 1.110873e-05, 
    6.727202e-06, 2.39074e-06, 5.205463e-07, 3.22998e-07, 3.356815e-07,
  1.760212e-07, 5.263137e-08, 3.740375e-08, 7.922812e-08, 8.469434e-08, 
    2.840129e-07, 7.233284e-07, 9.685888e-07, 4.679917e-06, 4.759401e-07, 
    3.596449e-08, 2.972017e-08, 2.930867e-06, 5.067277e-06, 1.160043e-05,
  4.344716e-06, 9.688731e-07, 4.002831e-08, 1.522813e-08, 9.220951e-08, 
    6.925476e-07, 7.947767e-08, 1.268206e-07, 1.368778e-07, 3.824859e-08, 
    7.625523e-08, 1.912638e-07, 1.296231e-06, 2.248377e-05, 1.197186e-05,
  3.675993e-06, 1.116344e-06, 1.052612e-07, 4.549028e-08, 5.092992e-08, 
    2.673649e-07, 1.004251e-07, 1.429628e-07, 9.487506e-08, 6.861897e-08, 
    3.676879e-08, 1.590912e-06, 2.351444e-06, 1.664465e-05, 2.89597e-06,
  2.197897e-07, 1.947716e-07, 1.411157e-07, 1.213779e-07, 6.623856e-08, 
    1.046017e-06, 2.36952e-07, 7.860343e-08, 7.815686e-08, 6.009078e-08, 
    1.788748e-07, 1.968657e-06, 2.516347e-06, 8.66768e-06, 2.800854e-07,
  9.09626e-07, 2.806474e-07, 2.103185e-07, 2.667558e-07, 3.630206e-07, 
    1.95676e-06, 1.639881e-06, 7.987905e-07, 4.350274e-08, 2.75331e-07, 
    5.608052e-07, 9.227938e-07, 4.020622e-06, 1.535459e-06, 2.421261e-07,
  5.130292e-07, 1.929317e-06, 6.20375e-07, 1.681794e-07, 1.198184e-07, 
    9.427329e-08, 4.943059e-08, 1.487428e-07, 1.740775e-07, 3.003861e-06, 
    1.814399e-06, 1.378703e-06, 4.181414e-06, 4.62062e-06, 6.415209e-06,
  3.284567e-07, 3.475274e-07, 3.670827e-07, 3.902992e-07, 4.914595e-07, 
    3.308873e-07, 2.758042e-07, 6.316976e-07, 1.587464e-05, 2.284541e-05, 
    1.096437e-05, 2.860112e-06, 4.264842e-07, 2.782483e-07, 7.545909e-09,
  1.181716e-07, 1.462695e-07, 1.88588e-07, 2.203506e-07, 2.532618e-07, 
    4.218415e-07, 6.81005e-07, 4.315545e-06, 4.228574e-05, 3.094455e-05, 
    1.119275e-05, 5.421115e-06, 1.18362e-06, 1.086855e-06, 1.334547e-08,
  1.422048e-07, 2.145538e-06, 5.026627e-07, 1.018945e-07, 4.832727e-06, 
    4.238641e-06, 2.53015e-06, 9.251941e-06, 5.913677e-05, 4.161646e-05, 
    2.075976e-05, 1.469147e-05, 9.814476e-06, 2.402182e-06, 1.967341e-08,
  5.621823e-06, 1.446791e-06, 3.530299e-06, 4.496879e-07, 3.398797e-06, 
    5.006332e-06, 1.093885e-05, 2.365577e-05, 3.679222e-05, 3.486892e-05, 
    2.848047e-05, 2.229935e-05, 3.332731e-05, 2.381432e-05, 7.453758e-08,
  1.594083e-06, 1.032364e-06, 1.686738e-06, 6.114107e-07, 5.18831e-07, 
    7.24596e-06, 1.308291e-05, 2.269698e-05, 1.392155e-05, 2.725958e-06, 
    2.867771e-07, 2.237449e-06, 2.05751e-05, 8.210049e-05, 0.000127352,
  1.482937e-06, 1.161838e-06, 1.845919e-07, 1.293416e-07, 3.354643e-06, 
    8.757292e-06, 1.93599e-05, 4.771251e-05, 5.317937e-05, 8.427787e-07, 
    8.716852e-06, 2.999389e-05, 0.0001423201, 0.0002291697, 0.0001266305,
  5.565877e-06, 2.451657e-06, 1.797483e-07, 1.223986e-07, 2.287656e-07, 
    2.444755e-06, 9.254611e-06, 1.021628e-05, 1.534546e-05, 3.870785e-06, 
    2.615977e-06, 3.311435e-06, 8.085208e-06, 7.568445e-05, 7.280424e-05,
  9.39015e-06, 1.230847e-05, 3.733281e-06, 4.538135e-07, 2.944462e-07, 
    3.786429e-06, 2.598215e-09, 1.564916e-06, 3.492794e-06, 5.292979e-07, 
    2.340608e-07, 1.91409e-07, 2.718096e-07, 3.990602e-05, 4.293485e-06,
  4.437805e-05, 5.297147e-05, 1.760521e-05, 5.376095e-06, 8.813953e-06, 
    1.039611e-05, 5.174973e-06, 7.872679e-06, 9.664701e-08, 2.87467e-07, 
    8.213602e-07, 1.094858e-06, 3.584338e-07, 2.868274e-06, 1.565701e-07,
  9.477579e-05, 0.0001009301, 3.451154e-05, 4.345187e-06, 7.677642e-06, 
    9.85657e-06, 9.498133e-06, 4.572382e-09, 4.105824e-08, 3.563227e-07, 
    1.536198e-06, 1.496062e-06, 6.369743e-07, 1.769242e-06, 4.524833e-07,
  6.338341e-05, 5.269919e-05, 6.23949e-05, 2.929154e-05, 2.262707e-05, 
    3.822823e-06, 8.295105e-06, 1.220565e-05, 6.118878e-05, 0.0001074715, 
    5.962455e-05, 2.738971e-05, 1.342589e-05, 1.644219e-05, 1.058646e-08,
  6.041891e-05, 7.628786e-05, 0.0001203429, 0.0001023631, 1.612182e-05, 
    3.211369e-05, 6.870333e-05, 8.589422e-05, 0.0001442471, 0.000113114, 
    7.002958e-05, 4.190797e-05, 2.98087e-05, 2.542028e-05, 2.522067e-07,
  0.0001601124, 0.0001014582, 7.358135e-05, 8.634007e-05, 5.320799e-05, 
    3.617564e-05, 5.001444e-05, 0.0001208225, 0.0001389136, 0.0001017058, 
    5.516031e-05, 4.347783e-05, 3.777698e-05, 1.732015e-05, 9.82976e-09,
  0.0001777677, 6.919174e-05, 6.936706e-05, 8.33339e-05, 4.967482e-05, 
    2.673861e-05, 3.276346e-05, 4.64767e-05, 5.508953e-05, 3.59799e-05, 
    2.06623e-05, 2.237682e-05, 2.938001e-05, 1.768034e-05, 9.501166e-08,
  0.0001737865, 6.8229e-05, 5.374978e-05, 7.035766e-05, 3.531185e-05, 
    1.962024e-05, 1.793815e-05, 1.550332e-05, 2.029775e-05, 5.356096e-07, 
    2.970641e-08, 5.041411e-06, 1.996489e-05, 5.998564e-05, 0.0001068089,
  7.228812e-05, 9.89725e-05, 5.861883e-05, 9.290261e-05, 7.021449e-05, 
    3.064282e-05, 2.258693e-05, 1.650374e-05, 1.778387e-05, 6.682348e-09, 
    6.178396e-07, 7.987152e-06, 2.357151e-05, 8.632102e-05, 7.06128e-05,
  7.164535e-05, 0.0001007535, 5.525086e-05, 7.989744e-05, 7.033396e-05, 
    3.37992e-05, 2.417676e-05, 1.947471e-05, 3.978666e-06, 1.774322e-09, 
    1.575856e-08, 8.97216e-08, 1.539581e-08, 2.454239e-05, 5.584256e-05,
  0.0001055817, 0.0001289611, 7.009505e-05, 7.327413e-05, 6.789926e-05, 
    4.785241e-05, 2.806679e-05, 2.00552e-05, 3.515077e-06, 1.107786e-09, 
    5.863025e-10, 6.181166e-09, 5.511161e-08, 3.411925e-05, 2.323886e-05,
  0.000129472, 0.0001255698, 0.0001091998, 0.0001262597, 0.0001236007, 
    9.4887e-05, 5.079094e-05, 3.908398e-05, 8.593787e-06, 9.129505e-07, 
    2.843184e-07, 4.602032e-07, 5.253488e-07, 1.709715e-05, 1.196252e-05,
  0.0001445123, 0.0001370501, 0.0001271102, 0.0001831181, 0.0002267677, 
    8.638265e-05, 3.216191e-05, 1.412622e-05, 9.267915e-06, 3.810761e-06, 
    4.295509e-06, 2.818707e-06, 1.632834e-06, 3.617028e-05, 2.360495e-05,
  5.549027e-06, 1.290335e-05, 3.437055e-05, 3.268023e-05, 2.646104e-05, 
    4.620919e-05, 4.973555e-05, 0.0001066084, 0.0001678206, 0.0001571966, 
    0.000102853, 6.983618e-05, 5.993332e-05, 8.038786e-05, 6.508062e-05,
  1.926275e-07, 8.34542e-10, 1.555137e-05, 4.981536e-05, 7.515433e-05, 
    8.299707e-05, 0.0001000817, 0.0001198663, 0.0001873672, 0.0001836542, 
    0.0001366758, 9.355035e-05, 5.824276e-05, 7.746524e-05, 7.099978e-05,
  1.24139e-06, 1.00201e-05, 4.269889e-06, 3.820972e-05, 6.871427e-05, 
    7.97751e-05, 6.224688e-05, 8.027336e-05, 0.0001559094, 0.0001781108, 
    0.0001901304, 0.0001414503, 8.078665e-05, 0.0001151962, 3.937546e-05,
  1.575728e-06, 6.59946e-06, 3.740807e-05, 8.821167e-05, 8.243745e-05, 
    9.815457e-05, 7.112972e-05, 4.301492e-05, 0.0001053268, 0.0002497507, 
    0.0003617999, 0.0003011727, 0.0002226391, 0.0001578747, 0.0001146903,
  2.767246e-06, 6.348847e-06, 2.775547e-05, 8.870081e-05, 8.396348e-05, 
    5.833713e-05, 4.62963e-05, 6.255943e-05, 0.0001237403, 0.0002884739, 
    3.062433e-05, 0.0001466813, 0.0004462072, 0.0003397716, 0.0002072854,
  1.457218e-06, 1.531033e-05, 2.984804e-05, 7.166207e-05, 8.497405e-05, 
    2.32234e-05, 1.98259e-05, 5.964192e-05, 9.66805e-05, 4.327206e-06, 
    1.165365e-05, 1.601288e-05, 0.0001446364, 0.0002892476, 0.0001762292,
  1.272844e-05, 1.068631e-05, 2.367477e-05, 4.4556e-05, 8.12109e-05, 
    3.470587e-05, 1.910142e-05, 3.708737e-05, 1.71782e-05, 3.796621e-06, 
    4.592263e-06, 4.777772e-06, 3.760334e-06, 7.261508e-05, 0.0001050416,
  2.122077e-05, 1.975637e-05, 2.05471e-05, 3.855877e-05, 4.443593e-05, 
    2.161073e-05, 2.685352e-05, 3.301254e-05, 2.188014e-05, 9.37817e-07, 
    2.789152e-06, 4.876208e-06, 1.262309e-08, 3.823456e-05, 8.030063e-05,
  2.396157e-05, 3.198402e-05, 3.881278e-05, 8.748343e-05, 6.658104e-05, 
    4.893793e-05, 4.0372e-05, 5.427508e-05, 5.899257e-07, 5.790338e-07, 
    2.143256e-07, 3.318308e-06, 3.346962e-07, 2.620396e-05, 3.703415e-05,
  3.017588e-05, 3.490736e-05, 5.818993e-05, 0.000116463, 0.0001652328, 
    7.518119e-05, 2.757304e-05, 1.83486e-06, 1.011364e-07, 1.895076e-08, 
    6.873441e-08, 6.371952e-07, 1.803195e-06, 1.115238e-05, 1.643716e-05,
  1.023579e-09, 2.816639e-09, 8.502172e-09, 1.596713e-09, 4.413544e-11, 
    1.851931e-10, 7.219786e-12, 3.057318e-12, 3.044694e-09, 2.848402e-07, 
    6.302031e-06, 2.665968e-05, 1.510308e-05, 3.210371e-05, 8.813353e-05,
  3.19023e-10, 9.528817e-09, 6.519933e-09, 3.751885e-09, 2.843918e-07, 
    6.635942e-10, 6.026806e-11, 2.526938e-11, 3.808128e-09, 1.293231e-07, 
    2.404759e-06, 1.04491e-05, 8.088746e-06, 3.238548e-05, 0.0001169532,
  4.060377e-07, 4.946171e-06, 1.174476e-06, 9.704574e-08, 9.274378e-07, 
    6.664438e-07, 7.159865e-09, 7.865483e-09, 1.733353e-07, 2.412605e-06, 
    1.223843e-05, 1.853657e-05, 1.005709e-05, 5.052037e-05, 4.925069e-05,
  1.530002e-06, 5.825058e-06, 2.238815e-05, 2.331615e-05, 1.231062e-05, 
    6.55093e-06, 4.29024e-06, 1.272842e-06, 3.01783e-06, 1.737168e-05, 
    7.844811e-05, 0.0001115453, 7.588604e-05, 0.0001323687, 9.295918e-05,
  2.06857e-07, 4.653462e-06, 1.111508e-05, 2.844203e-05, 5.387594e-06, 
    3.516936e-06, 8.511412e-06, 6.99831e-06, 1.510669e-05, 4.133139e-05, 
    4.431761e-06, 3.093589e-05, 0.0002749749, 0.0002990172, 0.0001416766,
  1.28164e-07, 3.894767e-06, 8.69883e-06, 1.527374e-05, 2.816262e-05, 
    5.608688e-06, 1.970405e-06, 4.235422e-06, 9.062519e-06, 8.020425e-06, 
    3.912322e-05, 5.399999e-05, 0.00019837, 0.0003932343, 7.707243e-05,
  1.088135e-07, 5.866664e-07, 1.28377e-06, 4.552556e-06, 1.186709e-05, 
    4.371715e-06, 2.362053e-06, 2.014544e-06, 4.770695e-06, 1.025798e-05, 
    6.90431e-06, 2.723295e-05, 9.648957e-05, 8.585974e-05, 4.997869e-05,
  5.132038e-08, 4.738611e-08, 1.06422e-06, 3.289382e-07, 2.33552e-06, 
    2.415285e-06, 1.019088e-06, 1.443926e-06, 1.382129e-05, 3.49832e-07, 
    2.622036e-06, 1.828459e-05, 6.071401e-06, 9.883974e-05, 6.742446e-05,
  5.161381e-08, 1.341785e-06, 1.775687e-06, 9.697778e-07, 8.079525e-07, 
    1.274176e-06, 2.211218e-06, 2.611801e-06, 1.135193e-06, 4.069556e-07, 
    5.59851e-07, 1.037102e-05, 2.749965e-06, 6.670672e-05, 6.052685e-05,
  1.833885e-07, 2.258014e-06, 9.296594e-07, 7.674445e-07, 1.447816e-07, 
    4.425194e-08, 1.006835e-07, 2.153613e-07, 8.17024e-08, 1.069044e-07, 
    1.467653e-07, 5.056775e-06, 3.000114e-06, 3.032962e-05, 6.78729e-05,
  2.485693e-27, 4.888188e-28, 2.914765e-15, 3.541348e-12, 2.646537e-10, 
    1.682629e-09, 3.9057e-09, 1.5042e-08, 1.88148e-06, 3.749297e-06, 
    1.193534e-05, 4.165012e-05, 3.893551e-05, 2.271454e-05, 1.104417e-05,
  1.291514e-32, 6.623578e-31, 1.587927e-27, 4.265284e-15, 3.325752e-12, 
    1.509975e-11, 2.142129e-10, 2.630199e-09, 4.469327e-07, 1.54394e-06, 
    8.553885e-06, 3.155187e-05, 2.873202e-05, 2.185006e-05, 8.25619e-06,
  0, 2.65525e-35, 9.929473e-28, 2.828945e-15, 7.885152e-11, 4.513085e-10, 
    7.254432e-10, 4.684087e-09, 2.485197e-07, 1.655117e-06, 4.163934e-06, 
    9.981537e-06, 1.110889e-05, 2.8763e-05, 9.873496e-06,
  3.378205e-27, 6.179834e-14, 2.941395e-13, 8.29231e-13, 3.630019e-10, 
    1.459049e-07, 1.125944e-07, 8.373593e-08, 1.671826e-06, 1.244805e-05, 
    2.457241e-05, 3.30568e-05, 1.841562e-05, 6.618943e-05, 2.49128e-05,
  6.581677e-14, 4.457285e-13, 7.372049e-13, 2.935611e-13, 1.692995e-11, 
    1.145095e-09, 4.980236e-08, 4.646073e-07, 1.568154e-06, 6.277189e-06, 
    3.265264e-07, 2.150608e-05, 7.784451e-05, 9.105018e-05, 1.388409e-05,
  1.130676e-15, 7.995837e-13, 1.266593e-12, 1.494176e-13, 3.60893e-13, 
    1.010598e-10, 7.329475e-09, 2.926724e-07, 9.741861e-08, 5.952356e-07, 
    1.319111e-05, 1.320697e-05, 5.317672e-05, 0.0001267278, 5.563843e-06,
  2.740364e-11, 8.481619e-25, 8.526333e-26, 2.048335e-26, 1.297855e-14, 
    1.365083e-11, 3.693358e-10, 8.258735e-09, 8.399045e-08, 4.220772e-06, 
    5.416135e-06, 1.942489e-06, 8.532941e-06, 2.614448e-05, 4.576785e-07,
  3.623709e-10, 1.405319e-10, 6.099924e-12, 2.78793e-26, 6.883088e-20, 
    4.570134e-15, 5.10952e-11, 3.310375e-08, 6.689917e-07, 2.062137e-06, 
    9.307993e-07, 1.103151e-07, 7.557703e-07, 7.180811e-06, 2.410264e-07,
  6.97507e-10, 6.502503e-10, 4.699247e-10, 4.139546e-25, 5.617517e-26, 
    2.763912e-25, 3.483671e-14, 1.072268e-09, 4.718526e-08, 2.83301e-07, 
    3.374365e-07, 1.346962e-07, 2.055551e-08, 7.774741e-08, 1.598413e-07,
  2.357861e-09, 3.517387e-10, 1.313064e-09, 2.2518e-10, 1.313113e-17, 
    1.697355e-25, 7.794783e-16, 1.461371e-10, 1.64083e-08, 1.375377e-07, 
    1.944713e-07, 2.252716e-08, 8.606411e-10, 1.550246e-08, 6.440634e-08,
  3.029591e-22, 4.113811e-14, 6.103638e-13, 3.189766e-12, 5.079944e-11, 
    1.431293e-10, 2.054583e-09, 4.070619e-08, 3.605702e-06, 8.962403e-06, 
    1.380282e-05, 3.884042e-05, 3.884952e-05, 1.776135e-05, 1.443854e-05,
  1.459036e-12, 8.421741e-23, 7.526141e-24, 3.056679e-14, 2.206621e-12, 
    6.903001e-14, 2.088513e-11, 3.828004e-09, 7.79802e-07, 1.311719e-06, 
    2.738491e-06, 2.35353e-05, 3.702051e-05, 2.21942e-05, 8.299567e-06,
  1.413065e-09, 4.327211e-17, 2.171091e-23, 7.572887e-13, 1.336713e-11, 
    7.849679e-14, 3.537006e-11, 2.596451e-09, 4.517197e-08, 1.235669e-07, 
    1.317534e-06, 6.452546e-06, 2.354755e-05, 3.116312e-05, 1.238799e-05,
  3.700793e-08, 4.229312e-13, 1.247828e-15, 7.934359e-11, 2.835848e-15, 
    2.133586e-12, 1.406867e-09, 2.404753e-07, 2.529374e-07, 6.44729e-07, 
    2.118726e-07, 1.217617e-07, 3.561576e-06, 1.38978e-05, 3.628505e-05,
  1.171496e-07, 2.779261e-10, 5.055923e-12, 1.728612e-13, 2.787088e-12, 
    3.104992e-12, 4.718241e-12, 1.227904e-11, 2.468867e-10, 1.262609e-08, 
    5.448407e-11, 5.993198e-10, 9.735333e-08, 1.05701e-05, 2.527371e-05,
  1.078549e-07, 1.676755e-08, 2.921434e-10, 3.129218e-11, 1.563319e-11, 
    3.082816e-11, 1.865638e-11, 4.578662e-11, 4.368809e-12, 4.137041e-12, 
    5.868773e-07, 2.612301e-07, 1.646961e-07, 1.166982e-05, 1.314769e-05,
  1.794399e-07, 8.165484e-09, 3.388199e-09, 3.842272e-10, 1.176361e-10, 
    8.876769e-11, 3.964281e-11, 1.58409e-10, 2.463226e-11, 3.294734e-11, 
    1.126528e-07, 7.160241e-09, 1.771895e-08, 1.719803e-06, 5.668635e-06,
  1.586605e-07, 1.726716e-09, 1.523532e-09, 1.104504e-09, 7.057412e-10, 
    2.361518e-10, 6.0424e-10, 6.657274e-10, 2.001499e-12, 1.377057e-10, 
    1.906866e-09, 3.726607e-10, 6.511211e-08, 1.592088e-06, 1.794035e-08,
  4.259488e-06, 7.570883e-08, 2.395703e-09, 1.545336e-09, 4.944567e-09, 
    5.515473e-10, 1.800643e-09, 5.963282e-10, 3.070994e-11, 2.200435e-11, 
    1.016654e-10, 4.114934e-09, 2.165365e-08, 2.461869e-08, 4.786912e-10,
  1.336486e-07, 6.862328e-08, 2.656502e-08, 3.7001e-09, 2.764182e-09, 
    2.1702e-09, 5.380238e-09, 1.287742e-09, 6.122282e-10, 1.29747e-11, 
    2.895347e-11, 4.061876e-10, 1.592226e-09, 1.46895e-11, 3.249056e-10,
  9.81668e-12, 8.744427e-11, 9.723466e-12, 3.23397e-12, 2.678152e-11, 
    6.531739e-08, 7.879286e-07, 1.322145e-07, 1.668483e-06, 6.97339e-06, 
    1.144711e-05, 2.886987e-05, 3.153842e-05, 2.839241e-05, 4.931999e-06,
  1.076514e-09, 4.101746e-09, 2.218643e-09, 1.341542e-09, 6.938903e-10, 
    1.910542e-06, 9.316196e-07, 1.908252e-06, 4.402818e-06, 4.24497e-06, 
    5.442013e-06, 1.249346e-05, 2.900751e-05, 4.746764e-05, 6.653577e-06,
  1.187925e-07, 7.766994e-08, 2.406358e-08, 1.146602e-09, 1.842684e-07, 
    2.661631e-09, 1.279231e-09, 9.120741e-09, 1.771237e-06, 1.076982e-06, 
    1.941581e-06, 1.034904e-06, 8.082301e-06, 3.002033e-05, 1.707325e-05,
  9.455e-07, 4.727767e-08, 2.672865e-07, 3.355648e-08, 5.134695e-07, 
    9.17339e-09, 1.784005e-09, 2.390275e-09, 2.017566e-07, 3.979639e-08, 
    2.855272e-08, 7.633039e-09, 3.030121e-07, 2.259397e-06, 3.03877e-05,
  3.275659e-07, 2.207765e-07, 1.035932e-08, 1.077713e-09, 3.217367e-09, 
    1.322268e-09, 5.987816e-09, 3.035276e-09, 1.110691e-07, 1.676861e-09, 
    1.449956e-09, 4.237108e-10, 2.283271e-09, 8.615736e-09, 2.43393e-05,
  6.225657e-07, 1.656497e-07, 3.360489e-08, 4.252895e-09, 2.868579e-09, 
    2.369417e-09, 2.302472e-09, 2.337965e-09, 2.339498e-09, 8.726569e-10, 
    3.601951e-10, 7.78424e-10, 7.539519e-11, 1.101644e-07, 2.788802e-05,
  2.748642e-06, 2.393718e-07, 1.137181e-07, 3.945725e-08, 1.274879e-08, 
    6.437503e-09, 5.526256e-09, 3.799741e-09, 1.17565e-09, 1.602622e-09, 
    6.781695e-10, 4.811948e-10, 7.753886e-10, 1.359898e-07, 1.208249e-05,
  5.123688e-06, 1.457281e-07, 1.356552e-07, 7.111462e-08, 3.475749e-08, 
    1.250951e-08, 1.155111e-08, 7.913154e-09, 1.317429e-08, 5.124828e-09, 
    9.085546e-10, 4.091588e-10, 2.447215e-09, 1.745422e-06, 1.307137e-07,
  2.073045e-05, 3.847134e-07, 8.567064e-08, 8.11132e-08, 1.457852e-07, 
    2.860556e-08, 2.723106e-08, 2.751502e-08, 1.714145e-08, 4.659048e-09, 
    9.6111e-09, 3.044891e-09, 3.745664e-10, 2.164475e-08, 9.769393e-10,
  1.234638e-05, 7.169475e-07, 9.738964e-08, 6.3613e-08, 6.198181e-08, 
    4.438829e-08, 7.870638e-08, 6.926404e-08, 5.890572e-08, 2.724922e-08, 
    3.397984e-08, 2.596993e-08, 7.983107e-09, 3.097325e-09, 7.050217e-10,
  6.778833e-09, 9.803681e-08, 6.920672e-06, 1.757286e-06, 1.604339e-06, 
    1.180748e-05, 2.296485e-05, 1.238837e-05, 8.337838e-06, 1.751384e-06, 
    2.385927e-07, 1.746981e-08, 4.646387e-06, 9.283773e-06, 1.84342e-05,
  2.788001e-08, 7.344848e-08, 3.872609e-07, 1.140628e-06, 1.520604e-06, 
    1.364373e-05, 2.23847e-05, 1.361784e-05, 6.528471e-06, 8.583702e-07, 
    1.179906e-07, 1.194212e-06, 3.13711e-06, 1.421755e-05, 4.94248e-06,
  5.68606e-06, 1.796857e-05, 2.648268e-06, 2.654077e-08, 2.756404e-06, 
    1.049495e-05, 9.754807e-06, 5.346258e-06, 3.034113e-06, 1.689389e-06, 
    2.209699e-06, 2.41552e-06, 4.865637e-06, 8.209574e-06, 3.609302e-06,
  1.283607e-05, 2.994872e-05, 1.333314e-05, 1.598305e-05, 1.548349e-05, 
    1.617353e-05, 9.718034e-06, 6.031929e-06, 1.563506e-06, 2.053855e-06, 
    1.925365e-06, 1.161002e-06, 1.744723e-06, 1.114491e-06, 9.257333e-06,
  2.566413e-05, 2.498207e-05, 1.211878e-05, 8.981374e-06, 8.764643e-06, 
    4.58571e-06, 7.208283e-06, 8.000722e-06, 8.930732e-07, 3.076636e-08, 
    9.083535e-09, 2.577024e-09, 8.450144e-09, 1.740544e-08, 6.594597e-06,
  9.146287e-06, 1.0428e-05, 8.859321e-06, 4.309456e-06, 4.402574e-06, 
    2.855784e-06, 1.063059e-06, 1.594487e-07, 5.265889e-09, 4.30316e-09, 
    3.84621e-09, 1.940005e-09, 2.979983e-10, 3.456436e-09, 1.060333e-05,
  2.234342e-05, 7.712376e-06, 6.893634e-07, 7.42269e-08, 2.164858e-07, 
    6.325576e-07, 9.585244e-08, 6.35556e-09, 7.177368e-09, 2.555731e-09, 
    6.513609e-10, 2.755526e-09, 1.252947e-09, 5.505216e-09, 6.714486e-07,
  4.3594e-06, 1.087065e-05, 2.881267e-06, 1.005134e-07, 6.325813e-07, 
    1.655556e-06, 6.115287e-08, 1.906688e-08, 8.489133e-08, 4.701279e-11, 
    1.205198e-09, 4.57966e-09, 1.371258e-09, 2.212213e-08, 3.745365e-09,
  3.416676e-05, 1.175273e-05, 2.993361e-06, 4.301712e-07, 2.332588e-06, 
    7.080385e-06, 6.222214e-06, 2.692414e-08, 1.200171e-07, 2.501245e-08, 
    1.690952e-10, 1.770726e-09, 5.323234e-09, 1.112923e-08, 1.930123e-09,
  9.623822e-06, 2.75228e-06, 7.762362e-07, 6.169197e-08, 9.858225e-07, 
    3.433354e-08, 1.117668e-08, 1.457006e-07, 1.368019e-06, 2.607578e-08, 
    1.702228e-09, 1.70241e-08, 4.123768e-09, 8.983845e-09, 3.685492e-09,
  6.298006e-09, 3.123231e-06, 4.154351e-05, 6.395423e-05, 7.3879e-05, 
    5.27599e-05, 4.577906e-05, 3.507449e-05, 6.279266e-05, 6.871635e-05, 
    6.871892e-05, 5.253879e-05, 3.000739e-05, 1.261547e-05, 9.642528e-06,
  6.360052e-08, 1.964434e-06, 4.928507e-05, 9.393045e-05, 9.488128e-05, 
    5.700212e-05, 2.559335e-05, 1.241914e-05, 1.766556e-05, 1.532046e-05, 
    1.167135e-05, 5.745597e-06, 3.148558e-06, 4.591276e-06, 9.232962e-07,
  5.545428e-05, 5.047427e-05, 3.764463e-05, 2.756217e-05, 4.58297e-05, 
    4.899081e-05, 2.860907e-05, 6.25431e-06, 3.620169e-06, 6.814108e-07, 
    2.580318e-07, 3.267676e-07, 2.040667e-06, 4.589949e-06, 8.605434e-07,
  7.035908e-05, 6.373158e-05, 4.55502e-05, 3.650305e-05, 2.277504e-05, 
    3.478595e-05, 3.513598e-05, 9.134211e-06, 1.072257e-06, 3.068968e-08, 
    1.055271e-07, 1.704696e-08, 2.337027e-07, 3.443325e-06, 1.756078e-05,
  5.700814e-05, 4.678469e-05, 3.533521e-05, 3.080424e-05, 2.978627e-05, 
    1.8972e-05, 2.784385e-05, 7.678557e-06, 2.512995e-06, 2.017049e-06, 
    2.003717e-09, 6.749293e-10, 1.042987e-09, 6.976221e-07, 9.61031e-06,
  3.140443e-05, 4.261745e-05, 2.945497e-05, 2.592045e-05, 1.884337e-05, 
    2.370202e-05, 2.556739e-05, 2.66273e-05, 3.608152e-06, 1.688449e-09, 
    1.902677e-09, 1.138488e-09, 6.316724e-10, 3.680683e-08, 6.814498e-06,
  1.997163e-05, 2.449942e-05, 2.951804e-05, 2.6902e-05, 1.427006e-05, 
    2.5508e-05, 3.564189e-05, 1.130494e-05, 6.37949e-09, 4.00472e-09, 
    9.557465e-10, 1.125077e-09, 4.33884e-10, 3.413514e-09, 6.08893e-07,
  1.041597e-05, 2.694422e-05, 2.205455e-05, 1.616222e-05, 1.13146e-05, 
    2.342987e-05, 1.603819e-05, 2.224564e-06, 3.100692e-09, 4.189011e-09, 
    5.281397e-10, 1.23149e-09, 2.395927e-09, 1.538025e-09, 4.509099e-09,
  5.188771e-06, 1.883171e-05, 2.499828e-05, 1.671482e-05, 2.115449e-05, 
    1.383806e-05, 1.483569e-05, 4.835774e-06, 1.410152e-09, 9.624672e-10, 
    1.836728e-10, 3.762628e-10, 2.574614e-09, 1.688622e-09, 3.586141e-10,
  8.971565e-06, 8.724609e-06, 1.401767e-05, 1.022136e-05, 3.837657e-06, 
    1.230368e-07, 4.223477e-07, 3.69845e-08, 6.441056e-08, 2.434352e-10, 
    3.835451e-10, 4.711007e-10, 2.193996e-09, 1.245944e-09, 2.20642e-10,
  1.065024e-06, 2.02976e-06, 4.185603e-06, 6.996602e-07, 2.553817e-08, 
    5.006714e-09, 6.748747e-09, 1.526378e-08, 1.660734e-06, 1.652238e-05, 
    6.823827e-05, 0.0001013293, 7.608809e-05, 3.998158e-05, 5.083975e-05,
  2.492897e-09, 1.202583e-09, 1.484713e-08, 1.345276e-06, 1.224885e-07, 
    9.017055e-08, 4.862614e-09, 1.05511e-08, 3.375626e-07, 1.147091e-07, 
    1.744635e-06, 1.57507e-05, 2.197892e-05, 2.289453e-05, 4.283721e-05,
  7.557526e-06, 1.136487e-09, 6.971835e-08, 1.676877e-07, 9.437343e-07, 
    8.225578e-08, 2.965604e-08, 2.668565e-08, 8.651334e-07, 3.283635e-07, 
    1.035773e-07, 1.029888e-06, 8.134858e-06, 1.610514e-05, 7.917388e-06,
  3.475448e-05, 4.553386e-07, 2.992251e-06, 5.258111e-06, 3.622665e-06, 
    5.30835e-06, 6.722536e-06, 2.41785e-06, 9.1865e-08, 1.608689e-09, 
    2.455131e-07, 3.432017e-07, 3.276662e-07, 4.020448e-06, 1.968056e-05,
  8.291016e-05, 5.31228e-06, 6.535839e-06, 1.286921e-05, 7.661156e-06, 
    3.493482e-06, 4.571701e-06, 8.848423e-06, 3.658535e-06, 2.771808e-08, 
    1.048022e-09, 1.259793e-08, 2.600459e-09, 6.485374e-07, 2.067909e-05,
  5.53083e-05, 3.753429e-05, 1.573901e-05, 2.931322e-05, 2.504036e-05, 
    1.376988e-05, 4.65928e-06, 1.203528e-06, 1.616169e-07, 2.267222e-09, 
    2.434213e-10, 1.023529e-10, 1.441367e-10, 4.955292e-08, 1.415912e-05,
  5.719945e-05, 6.38468e-05, 2.099616e-05, 4.207086e-05, 3.900275e-05, 
    2.839241e-05, 1.175481e-05, 2.19256e-06, 4.731438e-07, 1.206649e-09, 
    8.766733e-11, 1.5767e-10, 1.361323e-09, 1.875502e-08, 1.338316e-06,
  0.0001104458, 0.0001392401, 7.447237e-05, 4.06354e-05, 6.446228e-05, 
    4.360666e-05, 1.345505e-05, 4.615146e-06, 3.134838e-06, 1.502408e-08, 
    2.035847e-09, 1.353451e-11, 5.812635e-11, 4.827032e-10, 1.362837e-08,
  0.0002197659, 0.0002079044, 0.0001171338, 4.9689e-05, 7.865117e-05, 
    7.076794e-05, 1.900793e-05, 1.195437e-05, 1.701521e-06, 6.586067e-07, 
    1.355269e-08, 4.59122e-11, 1.477174e-13, 8.955564e-14, 2.081524e-10,
  0.0001923144, 0.0002314635, 0.0001169117, 3.561631e-05, 3.815896e-05, 
    2.026715e-05, 1.156815e-05, 1.191444e-05, 1.426403e-05, 2.712696e-06, 
    1.002773e-07, 2.81729e-08, 1.756153e-12, 1.442833e-10, 9.39429e-10,
  3.042915e-10, 3.958276e-07, 8.318342e-07, 8.77929e-07, 1.513856e-06, 
    3.790045e-10, 7.215033e-11, 1.13717e-10, 9.996758e-10, 4.400995e-09, 
    2.788224e-08, 2.636974e-06, 2.608629e-06, 7.195472e-06, 2.310033e-08,
  4.472381e-12, 3.72479e-11, 6.087687e-09, 8.88171e-07, 4.947857e-06, 
    5.613456e-06, 2.051618e-07, 1.412703e-09, 5.92831e-10, 1.225038e-08, 
    1.355667e-07, 6.49749e-07, 2.454346e-06, 1.561531e-06, 7.902311e-08,
  1.382452e-09, 3.793593e-09, 1.718956e-08, 1.632543e-06, 1.069743e-05, 
    2.666123e-05, 2.090467e-06, 2.464479e-09, 2.680076e-09, 4.245166e-09, 
    1.06533e-06, 3.109621e-08, 5.052259e-08, 1.520147e-07, 6.064101e-08,
  2.393472e-06, 5.602843e-07, 3.658427e-06, 2.902347e-05, 3.07831e-05, 
    3.489548e-05, 1.313078e-05, 1.23214e-05, 6.026803e-08, 5.138736e-08, 
    1.854479e-07, 2.525095e-08, 5.494402e-09, 7.434397e-09, 6.983748e-09,
  9.239891e-06, 6.350305e-07, 4.067815e-08, 1.919436e-06, 9.955557e-06, 
    1.464176e-05, 1.392586e-05, 2.011841e-05, 9.109108e-06, 5.683715e-06, 
    1.645974e-10, 7.444739e-10, 4.850559e-10, 2.30554e-09, 1.726585e-07,
  1.265803e-05, 3.197901e-06, 5.674761e-08, 1.37587e-07, 2.117713e-06, 
    6.233494e-06, 1.53336e-05, 6.659538e-06, 5.885702e-06, 1.512714e-09, 
    6.206505e-08, 1.519181e-09, 1.469375e-09, 8.335826e-09, 4.860862e-07,
  4.091115e-06, 1.946622e-06, 5.652788e-07, 1.518216e-06, 3.520153e-06, 
    4.098068e-06, 8.809022e-06, 7.19962e-06, 9.739824e-06, 7.3283e-08, 
    1.563567e-07, 1.918458e-08, 1.81383e-09, 2.486744e-09, 6.71601e-07,
  1.205598e-05, 1.796046e-05, 1.961235e-05, 1.807668e-05, 1.975153e-05, 
    1.831729e-05, 8.263085e-06, 1.21406e-05, 1.628724e-05, 3.423036e-07, 
    3.699906e-07, 1.24476e-07, 5.356267e-09, 4.690015e-09, 7.477786e-09,
  0.0002676636, 0.0002901017, 0.0002133963, 0.0001005956, 8.048004e-05, 
    7.469764e-05, 4.61024e-05, 1.218735e-05, 5.077216e-07, 2.086e-06, 
    1.671815e-06, 8.514283e-07, 1.165121e-07, 8.474293e-08, 1.989168e-09,
  0.0005356273, 0.0006085123, 0.0004804048, 0.000263001, 0.0002437237, 
    0.0001562906, 7.843362e-05, 2.32876e-05, 5.015649e-05, 5.045255e-05, 
    2.779431e-05, 1.200431e-05, 5.79045e-06, 2.572055e-06, 9.796896e-08,
  2.336072e-11, 1.332267e-10, 1.475208e-09, 7.971468e-09, 1.197021e-08, 
    7.775508e-07, 1.939352e-06, 4.053995e-10, 2.581136e-09, 4.516028e-09, 
    3.034936e-08, 1.142535e-07, 7.807292e-06, 4.387162e-06, 5.878919e-08,
  7.48124e-08, 1.558363e-08, 2.992776e-09, 2.463678e-08, 1.588689e-08, 
    4.185864e-07, 3.623899e-06, 6.082076e-07, 6.095159e-08, 1.297338e-07, 
    6.395239e-08, 1.868453e-06, 1.61366e-05, 4.080534e-06, 7.32335e-09,
  4.60961e-07, 1.11924e-06, 1.728335e-07, 3.640563e-08, 4.665239e-07, 
    1.556198e-08, 3.337524e-09, 1.422114e-07, 2.523416e-07, 1.498794e-06, 
    8.201235e-07, 1.818835e-07, 1.592453e-06, 6.959642e-06, 1.799224e-09,
  7.892964e-06, 3.120248e-06, 3.960203e-07, 4.001736e-06, 1.275097e-06, 
    1.846757e-06, 1.366958e-06, 2.431286e-06, 1.43358e-06, 7.833224e-07, 
    8.844353e-08, 7.565117e-08, 1.067149e-08, 2.095029e-09, 4.505469e-09,
  1.040072e-05, 1.766697e-06, 1.826415e-06, 2.300702e-06, 1.160997e-06, 
    6.572977e-07, 2.43446e-06, 4.143651e-06, 1.916769e-06, 5.774329e-06, 
    6.969431e-09, 3.969181e-09, 4.985245e-07, 1.905384e-09, 6.501554e-09,
  1.280254e-05, 6.77014e-06, 1.069471e-05, 2.480844e-05, 2.398083e-05, 
    1.820922e-05, 1.029133e-05, 2.012629e-06, 2.084966e-07, 6.95175e-10, 
    8.697884e-09, 3.535515e-08, 6.340076e-09, 5.267129e-09, 3.807592e-07,
  1.844557e-05, 3.304188e-05, 2.83277e-05, 3.311355e-05, 4.150666e-05, 
    2.756595e-05, 2.128459e-05, 1.14144e-05, 3.513936e-06, 1.924662e-07, 
    3.135469e-08, 2.789166e-08, 8.393967e-09, 1.568174e-08, 7.774474e-07,
  2.227393e-05, 7.812207e-05, 7.06728e-05, 2.718674e-05, 4.3863e-05, 
    5.156526e-05, 8.195244e-05, 7.608953e-05, 3.031092e-05, 2.019361e-06, 
    1.304806e-07, 3.111558e-08, 2.461919e-08, 3.740635e-07, 2.996704e-08,
  0.000149322, 0.0002550232, 0.0002088366, 0.0001423963, 0.0001458691, 
    0.000108883, 6.246952e-05, 6.152664e-05, 2.365229e-05, 9.908304e-06, 
    2.073989e-06, 1.379262e-06, 4.876589e-07, 5.691087e-07, 3.552032e-08,
  0.000150534, 0.0002758645, 0.0002749404, 0.000277181, 0.0003080775, 
    0.0002580194, 0.0001969179, 0.0001724602, 0.0001925706, 9.641856e-05, 
    1.457742e-05, 3.726198e-06, 2.605535e-06, 1.867479e-06, 1.360602e-06,
  9.450686e-09, 5.54682e-07, 3.282409e-06, 5.074091e-06, 7.600357e-07, 
    5.749715e-09, 1.27662e-07, 5.373844e-07, 1.990846e-05, 1.260978e-05, 
    1.043594e-05, 1.183205e-05, 1.567181e-05, 4.106825e-05, 8.55334e-06,
  6.303047e-09, 1.640678e-08, 2.023514e-06, 1.277601e-05, 4.619249e-06, 
    1.396869e-06, 1.7923e-06, 1.34383e-06, 6.021374e-06, 1.610611e-05, 
    1.606131e-05, 2.225955e-05, 4.363661e-05, 6.528523e-05, 5.776587e-06,
  6.345502e-08, 2.935063e-08, 9.793467e-07, 1.504594e-06, 1.036597e-05, 
    1.502061e-06, 8.57789e-08, 1.49595e-06, 5.625991e-06, 2.588787e-05, 
    4.738845e-05, 4.332186e-05, 5.771782e-05, 5.648764e-05, 3.222372e-05,
  1.752609e-06, 2.686554e-07, 3.471987e-06, 7.126307e-06, 8.140365e-06, 
    7.02698e-06, 5.953784e-06, 7.788962e-06, 5.247277e-06, 2.074456e-05, 
    3.467128e-05, 5.420336e-05, 6.418327e-05, 6.110549e-05, 5.933371e-05,
  1.883856e-07, 6.163381e-08, 2.20329e-06, 8.008569e-06, 1.035162e-05, 
    1.074925e-05, 1.222697e-05, 1.780988e-05, 3.277685e-05, 5.40363e-05, 
    1.664901e-05, 1.823669e-05, 4.979853e-05, 1.373985e-05, 2.212445e-05,
  6.673148e-08, 5.353229e-07, 9.469186e-08, 2.036913e-07, 9.422211e-07, 
    4.758429e-06, 5.201528e-06, 1.520905e-05, 5.092992e-05, 5.082522e-05, 
    4.696742e-05, 3.7564e-05, 4.585514e-06, 1.499529e-05, 4.117479e-05,
  2.232384e-06, 2.476016e-06, 7.717012e-08, 1.350128e-08, 3.927705e-08, 
    1.934306e-07, 6.957918e-07, 1.328086e-05, 2.613462e-05, 8.543746e-06, 
    4.739998e-06, 6.01477e-06, 3.861113e-06, 3.407128e-05, 4.443405e-05,
  5.229087e-06, 5.59091e-06, 1.855366e-06, 7.134777e-08, 1.205071e-06, 
    2.125282e-06, 4.799791e-06, 2.60073e-06, 2.44892e-06, 9.247636e-09, 
    1.87527e-09, 1.230259e-07, 1.609163e-06, 4.365091e-05, 1.062541e-06,
  1.077952e-05, 2.3409e-05, 7.961789e-06, 3.495633e-06, 1.011315e-05, 
    1.581987e-05, 1.668469e-05, 1.654367e-05, 4.100437e-07, 8.633959e-07, 
    4.863039e-09, 5.418363e-08, 1.495724e-06, 1.965505e-05, 7.443782e-08,
  1.234623e-05, 3.09336e-05, 1.984491e-05, 4.083708e-06, 2.017186e-05, 
    1.85222e-05, 1.490302e-05, 7.992935e-06, 1.67668e-05, 7.824733e-06, 
    7.747286e-07, 4.944467e-08, 1.590465e-06, 1.990848e-05, 6.619422e-06,
  5.524079e-08, 8.1802e-08, 1.192899e-06, 8.610127e-07, 4.381208e-08, 
    9.035591e-08, 1.439336e-05, 4.153964e-05, 0.0001345487, 0.0001253885, 
    5.719178e-05, 2.0917e-05, 1.746107e-05, 4.75569e-05, 6.8369e-06,
  9.723825e-08, 5.777751e-08, 8.810758e-08, 4.17604e-06, 1.446352e-05, 
    3.759837e-05, 6.307646e-05, 0.0001029211, 0.0001307364, 9.53321e-05, 
    5.282477e-05, 4.125125e-05, 5.4223e-05, 7.498161e-05, 5.57915e-06,
  1.021536e-06, 2.695977e-07, 7.172693e-08, 1.162843e-05, 0.0001169306, 
    8.524293e-05, 8.746482e-05, 0.0001150515, 0.00010802, 4.693525e-05, 
    3.764037e-05, 5.408282e-05, 7.394101e-05, 6.350897e-05, 2.129179e-06,
  9.745263e-06, 1.349048e-06, 1.057283e-05, 9.085342e-05, 0.0001421377, 
    0.0001286652, 8.203692e-05, 7.055254e-05, 4.422781e-05, 2.442423e-05, 
    3.119564e-05, 4.147258e-05, 4.640281e-05, 3.87373e-05, 6.955499e-06,
  1.468843e-05, 1.7731e-05, 5.671635e-05, 0.0001359341, 0.0001365275, 
    8.702772e-05, 5.216577e-05, 1.888187e-05, 1.590323e-05, 1.457675e-05, 
    2.982943e-08, 7.746698e-06, 2.754853e-05, 1.927949e-05, 2.743788e-05,
  1.842558e-05, 7.781951e-05, 0.0001078687, 0.0001356722, 8.322668e-05, 
    2.761485e-05, 8.619838e-06, 4.733053e-06, 1.711044e-06, 3.4976e-08, 
    2.083454e-05, 9.415809e-06, 3.907147e-07, 2.290579e-05, 5.248503e-05,
  4.318983e-05, 9.797992e-05, 8.345194e-05, 6.354467e-05, 1.760762e-05, 
    1.394485e-05, 3.715753e-06, 8.172216e-06, 1.037479e-05, 3.68822e-05, 
    5.580007e-05, 2.945709e-05, 8.638916e-06, 2.414166e-05, 4.417141e-05,
  5.316282e-05, 8.844697e-05, 4.397403e-05, 1.698202e-05, 1.634575e-05, 
    1.570707e-05, 1.439756e-05, 2.428462e-05, 5.237075e-05, 9.271145e-05, 
    7.700498e-05, 4.635829e-05, 1.294368e-05, 7.117417e-05, 1.063055e-05,
  6.270606e-05, 6.867733e-05, 3.178186e-05, 1.848623e-05, 3.34344e-05, 
    6.225704e-05, 6.542214e-05, 5.545767e-05, 6.034915e-05, 9.706626e-05, 
    5.371478e-05, 3.681424e-05, 1.637959e-05, 7.360027e-05, 2.971293e-05,
  6.509609e-05, 7.116485e-05, 3.982392e-05, 2.339654e-05, 4.145318e-05, 
    6.626578e-05, 7.832322e-05, 1.929279e-05, 4.147485e-05, 5.970053e-05, 
    6.202232e-05, 6.844844e-05, 6.328117e-05, 8.790267e-05, 5.624679e-05,
  5.53674e-07, 7.869833e-07, 7.562696e-07, 9.279442e-07, 1.027058e-06, 
    8.116197e-07, 2.520713e-06, 3.810382e-06, 6.204511e-05, 0.0001262, 
    0.0001110451, 6.150819e-05, 3.630948e-05, 7.269032e-05, 5.190857e-05,
  7.864589e-07, 8.461084e-07, 8.763761e-07, 1.102105e-06, 4.787002e-07, 
    7.813761e-07, 7.010502e-06, 2.96619e-05, 8.657316e-05, 8.794806e-05, 
    7.257314e-05, 5.330843e-05, 3.837869e-05, 5.570378e-05, 8.073122e-05,
  7.33242e-07, 7.78358e-07, 5.952172e-07, 4.478575e-07, 1.749239e-05, 
    1.917335e-05, 1.251261e-05, 4.544685e-05, 6.136361e-05, 4.621936e-05, 
    5.218562e-05, 4.817943e-05, 5.281837e-05, 3.794611e-05, 5.213132e-05,
  5.106741e-07, 3.580058e-07, 3.827888e-07, 5.166776e-06, 2.701972e-05, 
    4.538759e-05, 3.85485e-05, 3.121464e-05, 3.104583e-05, 2.906247e-05, 
    3.890718e-05, 4.083158e-05, 5.752595e-05, 3.984258e-05, 2.754401e-05,
  3.265228e-07, 3.132905e-07, 9.699285e-07, 1.932833e-05, 4.944998e-05, 
    5.886666e-05, 4.703858e-05, 1.898929e-05, 1.632508e-05, 1.704374e-05, 
    8.03692e-08, 3.717018e-07, 0.0001053535, 6.858793e-05, 0.0001114069,
  4.227092e-07, 4.506312e-06, 2.872637e-05, 5.868909e-05, 6.647492e-05, 
    5.154382e-05, 1.406586e-05, 2.341455e-06, 3.625747e-06, 5.553872e-06, 
    1.725202e-05, 3.235045e-05, 1.157132e-05, 7.642089e-05, 0.0001348734,
  2.266794e-06, 2.283927e-05, 4.276292e-05, 6.227755e-05, 3.596767e-05, 
    1.062434e-05, 3.009568e-06, 3.351671e-06, 2.514352e-05, 2.646457e-05, 
    4.464473e-05, 7.141053e-05, 7.275352e-05, 9.888847e-05, 8.493467e-05,
  8.721884e-06, 4.222737e-05, 4.574569e-05, 2.300463e-05, 7.762635e-06, 
    3.415887e-06, 8.623575e-07, 7.701201e-06, 7.194866e-05, 2.394775e-05, 
    4.340706e-05, 5.96419e-05, 5.67872e-05, 0.0001348964, 5.505416e-05,
  1.585508e-05, 3.618193e-05, 1.867264e-05, 5.051448e-06, 6.608975e-06, 
    1.356463e-05, 2.36172e-05, 4.143954e-05, 4.84596e-06, 8.286886e-06, 
    1.703997e-05, 1.717562e-05, 4.955971e-05, 0.0001344227, 0.0001121436,
  5.127489e-06, 3.335499e-06, 3.567101e-06, 1.695845e-06, 1.063056e-05, 
    2.637658e-05, 2.985863e-05, 3.344049e-06, 1.475948e-06, 4.12421e-06, 
    4.325415e-06, 1.130218e-05, 6.957199e-05, 0.0001730893, 0.0001206757,
  5.40011e-08, 8.35967e-08, 2.489498e-07, 4.837447e-07, 5.849487e-07, 
    7.73459e-07, 8.512051e-07, 1.181829e-06, 7.977717e-06, 3.921762e-05, 
    7.186188e-05, 5.9126e-05, 0.0001376852, 0.0001938976, 6.51501e-05,
  3.204934e-07, 5.162801e-07, 5.215545e-07, 5.759477e-07, 5.648517e-07, 
    5.259431e-07, 5.112836e-07, 1.664875e-06, 5.557503e-05, 0.0001597622, 
    0.0001683662, 0.0001768056, 0.000226993, 0.0001366438, 6.675239e-05,
  5.143716e-07, 5.822055e-07, 5.8944e-07, 5.338824e-07, 3.952226e-07, 
    3.2487e-07, 6.927056e-07, 3.977662e-05, 0.0001694995, 0.0001672399, 
    0.0001434211, 0.0001495363, 0.0001205771, 7.124506e-05, 1.147138e-05,
  9.287203e-06, 6.264692e-07, 6.934514e-07, 1.102372e-06, 2.405753e-06, 
    1.304156e-05, 5.06154e-05, 0.0001216125, 0.0001261071, 7.685297e-05, 
    8.203028e-05, 4.45584e-05, 2.646924e-05, 3.023935e-05, 1.884939e-05,
  4.425484e-05, 1.805193e-05, 1.924601e-06, 2.716381e-06, 1.097709e-05, 
    5.756675e-05, 8.21698e-05, 5.608047e-05, 2.803972e-05, 1.747141e-05, 
    1.948623e-05, 2.827033e-06, 4.62747e-06, 2.764753e-06, 2.445463e-05,
  7.450481e-05, 6.759191e-05, 2.993852e-05, 6.518714e-05, 7.943947e-05, 
    6.971553e-05, 3.953513e-05, 1.141122e-05, 1.171561e-05, 1.537127e-05, 
    8.448313e-06, 4.142955e-06, 4.785154e-07, 1.099811e-06, 2.991117e-05,
  5.812386e-05, 6.765046e-05, 7.291904e-05, 0.0001230628, 9.855077e-05, 
    4.906836e-05, 1.09042e-05, 1.04343e-05, 3.168381e-05, 1.466373e-05, 
    3.329796e-06, 6.925272e-06, 4.550324e-06, 5.025178e-06, 9.27177e-06,
  3.330898e-05, 5.295205e-05, 7.567881e-05, 6.360515e-05, 5.20469e-05, 
    2.012433e-05, 4.592093e-06, 1.090665e-05, 2.755176e-05, 4.948117e-06, 
    1.169309e-06, 2.37318e-06, 2.755484e-06, 1.726808e-05, 1.035465e-06,
  5.069556e-06, 3.255942e-05, 3.148289e-05, 2.166469e-05, 3.355514e-05, 
    6.068548e-05, 4.003272e-05, 3.300311e-05, 1.659515e-05, 5.283241e-05, 
    8.546017e-06, 6.66969e-07, 2.373023e-06, 8.095567e-06, 1.857798e-06,
  6.381904e-06, 2.595203e-05, 4.708852e-05, 3.845913e-05, 6.400167e-05, 
    6.785095e-05, 7.890425e-05, 7.602323e-05, 0.0001269004, 4.315525e-05, 
    7.353276e-06, 1.374376e-06, 2.826014e-06, 1.220808e-05, 1.71965e-05,
  1.341606e-07, 1.269237e-06, 4.732488e-06, 4.329368e-06, 2.272291e-06, 
    5.716885e-06, 1.518329e-05, 1.865919e-05, 4.045327e-05, 3.243711e-05, 
    1.128364e-05, 6.718663e-06, 6.990438e-07, 1.724466e-07, 1.105054e-08,
  5.223306e-08, 3.316287e-07, 9.352151e-07, 6.067931e-06, 1.025223e-05, 
    1.263122e-05, 2.004925e-05, 2.200298e-05, 6.240248e-05, 5.518176e-05, 
    4.644245e-05, 1.88645e-05, 8.722676e-06, 4.405726e-06, 1.578407e-07,
  6.163911e-06, 4.727282e-06, 3.374649e-07, 1.277941e-06, 2.537369e-05, 
    5.688462e-05, 3.019079e-05, 4.874537e-05, 7.9831e-05, 9.160094e-05, 
    6.344865e-05, 2.772099e-05, 1.470864e-05, 1.444729e-05, 1.496236e-06,
  8.671364e-05, 4.603775e-05, 5.08011e-05, 9.512516e-05, 9.764297e-05, 
    0.0001098216, 9.588574e-05, 7.915038e-05, 7.367547e-05, 7.8803e-05, 
    4.247972e-05, 2.343755e-05, 5.439571e-05, 2.159495e-05, 5.035415e-06,
  0.0001260416, 0.0001290303, 0.0001379562, 0.0001480162, 0.0001804171, 
    0.0002055627, 0.0001865831, 0.0001233829, 9.224638e-05, 2.528236e-05, 
    1.252697e-06, 2.168246e-06, 1.849463e-05, 1.395811e-05, 3.910942e-05,
  5.189545e-05, 8.284647e-05, 0.0001007825, 0.0001557827, 0.0002476658, 
    0.0003173923, 0.0002796837, 0.0002293481, 0.0001469504, 8.566794e-05, 
    0.0001556662, 0.0002159992, 3.375782e-05, 3.983772e-05, 0.0001100337,
  3.160176e-05, 6.242286e-05, 4.310251e-05, 7.866181e-05, 0.0001401963, 
    0.0002111589, 0.0002487279, 0.0003080071, 0.0003303814, 0.0003578714, 
    0.0002424918, 0.0001572381, 4.355011e-05, 0.000164655, 0.0001701216,
  4.869335e-05, 6.890016e-05, 4.69992e-05, 6.206102e-05, 6.856897e-05, 
    0.0001161744, 0.0001623666, 0.0002402203, 0.00031905, 0.000265832, 
    0.0001951389, 0.0001950707, 0.0001991512, 0.0002768273, 5.368099e-05,
  7.547032e-05, 9.531667e-05, 7.328519e-05, 6.040451e-05, 7.636035e-05, 
    0.0001060121, 0.0001076636, 0.0001260267, 0.0001356009, 0.0001349403, 
    0.0001515996, 0.0001409524, 0.0001499486, 0.0001619535, 0.0001281305,
  6.101311e-05, 5.329941e-05, 4.767381e-05, 2.174917e-05, 3.348909e-05, 
    3.950094e-05, 4.51236e-05, 2.381664e-05, 4.683302e-05, 9.331635e-05, 
    9.571343e-05, 5.059444e-05, 2.265983e-05, 3.243266e-05, 5.342124e-05,
  8.159466e-08, 5.863652e-08, 2.875411e-07, 1.408792e-06, 9.661861e-07, 
    3.323382e-06, 8.418045e-06, 2.565159e-05, 0.0001131713, 0.0001479192, 
    0.0001353942, 4.843889e-05, 9.085433e-06, 8.164314e-06, 6.773072e-06,
  9.357263e-07, 1.183509e-06, 4.738497e-08, 5.345569e-07, 2.713508e-06, 
    6.071386e-06, 4.432602e-06, 8.714032e-06, 4.617013e-05, 9.490608e-05, 
    0.0001094506, 6.33528e-05, 2.582369e-05, 2.619709e-05, 9.07297e-07,
  8.860492e-06, 6.003301e-06, 2.672982e-07, 8.340412e-08, 1.771896e-06, 
    1.562612e-06, 1.33254e-06, 7.012813e-06, 2.564979e-05, 5.277699e-05, 
    6.068255e-05, 4.868806e-05, 2.335582e-05, 1.230499e-05, 1.056126e-07,
  6.880204e-05, 6.307175e-06, 3.590796e-06, 6.082933e-06, 4.233833e-06, 
    7.195896e-06, 6.161492e-06, 1.329086e-05, 2.050999e-05, 2.930982e-05, 
    6.285943e-05, 7.522921e-05, 3.882343e-05, 1.725162e-05, 5.667628e-07,
  8.819439e-05, 1.883608e-05, 1.097796e-06, 6.28882e-07, 1.094134e-06, 
    4.491062e-06, 6.822756e-06, 1.989513e-05, 3.276077e-05, 7.844575e-05, 
    7.083223e-05, 0.0001140779, 0.0001711899, 6.633914e-05, 4.716242e-05,
  6.606196e-05, 4.680166e-05, 2.39371e-06, 1.049481e-06, 2.364546e-06, 
    7.40529e-06, 5.925876e-06, 2.515278e-05, 4.314809e-05, 3.28271e-05, 
    3.807255e-05, 8.472426e-05, 9.048064e-05, 0.0001031861, 9.425024e-05,
  8.879861e-05, 8.106463e-05, 2.888836e-05, 7.786139e-06, 6.273059e-06, 
    3.443678e-06, 4.500427e-06, 9.572705e-06, 1.567117e-05, 1.441292e-05, 
    1.178459e-05, 1.165083e-05, 1.747023e-05, 5.021846e-05, 4.731104e-05,
  0.0001336903, 0.0001182649, 7.575854e-05, 3.843968e-05, 1.222947e-05, 
    8.206429e-06, 1.779159e-06, 2.353529e-06, 6.438824e-06, 3.939831e-06, 
    4.338714e-06, 4.929584e-06, 9.577906e-06, 5.542103e-05, 3.601289e-05,
  0.0001987381, 0.000181567, 0.0001325815, 6.840128e-05, 4.360953e-05, 
    2.30183e-05, 7.200475e-06, 7.560963e-06, 1.798388e-06, 4.053024e-06, 
    9.194166e-07, 1.855946e-06, 5.7697e-06, 6.040223e-05, 7.83826e-05,
  0.0001610801, 0.0001934035, 0.0001230273, 8.77233e-05, 6.724723e-05, 
    9.849884e-06, 1.789423e-06, 1.842764e-06, 4.588646e-06, 1.691631e-06, 
    1.371629e-06, 5.070819e-06, 4.984049e-06, 1.991784e-05, 1.980224e-05,
  0.0001003378, 0.0001308022, 0.0001507064, 0.0001076595, 4.421703e-05, 
    0.0001233635, 0.000173133, 0.0001227243, 0.00017845, 9.642072e-05, 
    7.702566e-05, 7.454187e-05, 0.0001184332, 0.0001079409, 7.898247e-05,
  8.140869e-05, 0.0001094508, 0.0001483557, 0.0001306169, 0.0001112884, 
    9.28676e-05, 0.0001701817, 0.0002095444, 0.0001688734, 0.000113771, 
    5.125642e-05, 5.651658e-05, 6.855326e-05, 4.665288e-05, 1.238113e-05,
  0.0002179286, 0.0001289364, 9.508545e-05, 0.000152092, 0.000170685, 
    0.0001460604, 0.0001281391, 0.0002562287, 0.0002241212, 0.000110762, 
    6.908338e-05, 4.664481e-05, 5.832749e-05, 5.779991e-05, 1.598807e-05,
  0.0001968511, 0.0001705326, 0.0001964767, 0.0002034321, 0.0001805044, 
    0.0001938051, 0.000249074, 0.0003005779, 0.0002229272, 0.0001181663, 
    8.603161e-05, 4.576942e-05, 5.616474e-05, 6.293777e-05, 0.0001126166,
  0.0001252893, 0.0001328122, 0.0001559769, 0.000107728, 8.52671e-05, 
    0.0001300111, 0.0001657301, 0.0001928121, 0.0002004733, 0.0001803192, 
    5.176568e-05, 9.219212e-05, 0.0001694632, 8.349506e-05, 0.0001606589,
  5.364791e-05, 8.806206e-05, 6.987576e-05, 6.580906e-05, 5.399428e-05, 
    3.974952e-05, 6.912302e-05, 8.847361e-05, 0.0001512994, 4.080505e-05, 
    8.370527e-05, 0.0001273304, 9.098854e-05, 0.0001161814, 0.0001952349,
  5.159587e-05, 4.863518e-05, 5.729163e-05, 8.981915e-05, 9.319161e-05, 
    4.56859e-05, 3.28015e-05, 5.554888e-05, 4.129649e-05, 1.039871e-08, 
    1.247085e-07, 1.171201e-05, 2.911452e-05, 9.073016e-05, 0.0001053268,
  2.935273e-05, 2.398234e-05, 3.901161e-05, 9.234162e-05, 0.0001299138, 
    8.253751e-05, 5.124774e-05, 4.955806e-05, 4.326805e-05, 2.978936e-06, 
    1.357476e-06, 7.047222e-07, 4.331202e-06, 6.477119e-05, 4.074894e-05,
  3.296059e-05, 2.083013e-05, 2.674062e-05, 7.226147e-05, 0.0001249712, 
    0.0001046382, 6.732252e-05, 0.000122725, 3.183289e-05, 1.731509e-05, 
    1.014669e-05, 3.222158e-06, 1.867824e-06, 4.684436e-05, 0.0001400769,
  1.877396e-05, 2.158267e-05, 5.996456e-05, 5.707342e-05, 0.0001134112, 
    0.0001415814, 0.0001235799, 9.779888e-05, 0.000101853, 6.278003e-05, 
    2.975501e-05, 1.868833e-06, 6.436515e-06, 4.760061e-05, 0.000115788,
  9.038972e-06, 1.049393e-05, 1.917452e-05, 1.804548e-05, 1.339626e-05, 
    2.213513e-05, 3.152455e-05, 3.762235e-05, 0.000144205, 0.0001119388, 
    6.303128e-05, 6.4003e-05, 4.9293e-05, 7.207011e-05, 7.330773e-06,
  1.252024e-10, 3.194753e-10, 3.202221e-06, 6.454572e-06, 3.012134e-06, 
    9.291404e-06, 3.628535e-05, 0.000103514, 0.0001586643, 0.0001176692, 
    7.97414e-05, 8.19979e-05, 4.909745e-05, 5.538762e-05, 1.73436e-05,
  2.642178e-08, 4.121295e-08, 6.572512e-08, 5.518422e-08, 2.343623e-06, 
    1.085023e-05, 3.818534e-05, 0.0001202717, 0.0001570754, 0.000112798, 
    7.939884e-05, 5.941681e-05, 3.598858e-05, 2.58782e-05, 3.589845e-07,
  1.181673e-06, 7.381838e-07, 6.29186e-06, 1.167206e-05, 1.154061e-05, 
    1.833855e-05, 3.219112e-05, 7.173712e-05, 9.320726e-05, 9.862839e-05, 
    0.0001752946, 0.000163342, 9.611608e-05, 4.414696e-05, 6.277334e-06,
  2.405475e-07, 2.357306e-07, 1.823101e-06, 1.080227e-05, 1.181988e-05, 
    2.894946e-05, 3.06162e-05, 4.252488e-05, 6.501711e-05, 0.0001518877, 
    0.0001079319, 0.0001856191, 0.0003044455, 0.0001264557, 0.0001000626,
  2.139491e-08, 1.48065e-07, 3.953596e-07, 2.632034e-06, 8.051563e-06, 
    1.605274e-05, 2.710279e-05, 3.124349e-05, 3.96849e-05, 1.017995e-05, 
    2.201577e-05, 4.087596e-05, 9.251451e-05, 0.0001720403, 0.0001234269,
  6.419479e-07, 3.681714e-07, 7.201276e-07, 1.038183e-06, 2.182024e-06, 
    3.321279e-06, 1.171962e-05, 8.865824e-06, 1.010698e-05, 8.232208e-06, 
    6.505205e-06, 5.814312e-06, 1.464236e-05, 0.0001433903, 9.924499e-05,
  3.437875e-07, 1.348214e-06, 1.822016e-06, 2.454037e-06, 4.609029e-06, 
    5.315752e-06, 4.011411e-06, 4.568148e-06, 1.2312e-05, 7.567079e-06, 
    7.15127e-06, 1.131193e-05, 8.17564e-06, 5.283232e-05, 2.2552e-05,
  6.670743e-07, 8.895105e-07, 1.646861e-06, 4.74643e-06, 2.827342e-05, 
    4.612223e-05, 2.644186e-05, 2.72912e-05, 4.051286e-06, 8.346867e-06, 
    5.315446e-06, 7.034787e-06, 4.998185e-06, 2.200655e-05, 2.968737e-05,
  7.808838e-07, 5.359128e-06, 1.569858e-05, 2.977182e-05, 7.070429e-05, 
    9.853273e-05, 8.995021e-05, 6.464522e-05, 7.418876e-05, 5.190158e-05, 
    2.246099e-05, 1.233932e-05, 1.099687e-05, 1.737645e-05, 4.30085e-05,
  1.581771e-05, 4.530112e-06, 4.487425e-06, 5.029148e-06, 2.923488e-06, 
    6.910195e-06, 1.028672e-05, 3.887905e-06, 1.146209e-05, 2.184889e-05, 
    1.223364e-05, 5.204806e-06, 1.62281e-06, 4.829677e-06, 2.295697e-08,
  1.049197e-05, 1.471346e-05, 1.20781e-05, 2.636578e-05, 1.85993e-05, 
    1.676282e-05, 9.139158e-06, 1.074701e-05, 2.171204e-05, 2.120872e-05, 
    1.189174e-05, 4.380908e-06, 2.197051e-06, 6.873707e-06, 3.903536e-09,
  7.757046e-05, 5.484673e-05, 2.944718e-05, 8.022804e-05, 0.0001143007, 
    5.598349e-05, 1.059012e-05, 1.701628e-05, 3.806667e-05, 2.581825e-05, 
    1.080633e-05, 5.592552e-06, 6.330732e-06, 4.373256e-06, 2.458482e-09,
  0.0001042952, 5.055371e-05, 5.908999e-05, 0.0001019489, 9.827576e-05, 
    7.804231e-05, 7.005998e-05, 9.582059e-05, 0.0001061293, 6.184787e-05, 
    2.532272e-05, 1.587871e-05, 1.485183e-05, 3.607489e-06, 5.934744e-07,
  5.636542e-05, 5.966817e-05, 8.012323e-05, 0.0001052051, 0.0001062837, 
    0.0001228995, 0.0001318004, 0.0001765809, 0.0002118623, 0.0002218103, 
    0.0001829065, 0.0001358029, 0.0001108481, 9.287458e-06, 1.276833e-05,
  2.668548e-05, 5.771417e-05, 8.325378e-05, 0.000104004, 0.0001110292, 
    0.0001373121, 0.000196793, 0.0002702127, 0.0003536216, 0.0003880722, 
    0.0002350085, 0.0001774878, 8.624807e-05, 6.035115e-05, 6.515743e-05,
  3.631327e-05, 4.928075e-05, 5.067228e-05, 5.882952e-05, 7.543588e-05, 
    8.259689e-05, 0.0001410433, 0.0002174242, 0.0002804802, 0.0001615507, 
    8.621944e-05, 8.443488e-05, 8.611417e-05, 0.0001922469, 0.0001330878,
  4.052623e-05, 6.482181e-05, 3.852022e-05, 5.138523e-05, 7.021143e-05, 
    6.558017e-05, 7.085173e-05, 9.457108e-05, 0.0001572577, 7.829578e-05, 
    5.268808e-05, 6.680504e-05, 0.0001053474, 0.0002472528, 6.366413e-05,
  5.536718e-05, 8.343506e-05, 7.135297e-05, 9.276636e-05, 0.0001007531, 
    0.0001017932, 7.754595e-05, 0.0001082879, 5.614027e-05, 3.788027e-05, 
    2.255373e-05, 3.680284e-05, 9.555241e-05, 0.0001724514, 7.324897e-05,
  4.195191e-05, 9.018483e-05, 0.0001236899, 0.0001401487, 0.0001532897, 
    0.0001560325, 0.0001316318, 5.854945e-05, 3.488521e-05, 2.194414e-05, 
    1.59563e-05, 1.490009e-05, 5.6535e-05, 8.604027e-05, 8.764892e-05,
  1.319443e-05, 2.331349e-05, 4.172798e-05, 4.906488e-05, 4.626413e-05, 
    3.764224e-05, 4.074261e-05, 2.860338e-05, 7.666818e-05, 5.447899e-05, 
    1.319877e-05, 1.778029e-06, 3.382937e-07, 7.120517e-06, 1.521186e-07,
  9.079516e-06, 2.670062e-05, 6.412633e-05, 0.0001262194, 0.0001029793, 
    0.0001074227, 6.226479e-05, 7.443557e-05, 0.0001439101, 0.0001357058, 
    8.208905e-05, 1.609616e-05, 1.612784e-06, 5.282241e-06, 8.757985e-07,
  7.73499e-06, 2.059529e-05, 3.809142e-05, 7.583426e-05, 9.668325e-05, 
    0.0001205269, 0.0001204037, 0.0001379049, 0.000200764, 0.0002324134, 
    0.0001972554, 0.0001344544, 6.535488e-05, 1.563079e-05, 8.37773e-07,
  2.543724e-06, 1.571737e-05, 1.44658e-05, 3.561757e-05, 6.086007e-05, 
    8.002656e-05, 0.0001213487, 0.000188425, 0.0002322127, 0.0002540796, 
    0.0003395946, 0.0003000312, 0.0001469453, 0.0001049903, 2.032051e-05,
  3.570765e-07, 1.054265e-05, 6.857739e-06, 1.963882e-05, 3.059925e-05, 
    4.937856e-05, 7.165493e-05, 0.000112236, 0.0002051212, 0.0004132128, 
    0.0005566185, 0.0003326387, 0.0003537901, 0.0001286976, 0.0001161754,
  2.783054e-07, 1.144094e-05, 5.295805e-06, 4.28458e-06, 1.725391e-05, 
    3.319527e-05, 4.699599e-05, 6.113498e-05, 9.76294e-05, 8.975509e-05, 
    8.523802e-05, 0.0001009063, 7.843668e-05, 3.43824e-05, 8.227567e-05,
  3.198346e-06, 1.022561e-05, 1.10349e-05, 6.311105e-06, 1.760597e-05, 
    2.925108e-05, 4.279903e-05, 3.434931e-05, 1.288628e-05, 4.718585e-06, 
    1.167735e-05, 2.106419e-05, 1.049232e-05, 2.033098e-05, 4.214578e-05,
  8.742617e-07, 6.821222e-06, 1.669282e-05, 1.803673e-05, 1.688881e-05, 
    3.015094e-05, 3.729701e-05, 2.658215e-05, 5.807073e-05, 1.275453e-05, 
    2.102191e-05, 1.804691e-05, 3.915924e-06, 3.561561e-05, 3.008251e-05,
  3.218909e-07, 6.569554e-06, 1.507142e-05, 2.715767e-05, 4.2536e-05, 
    7.396917e-05, 7.895535e-05, 9.832844e-05, 1.285198e-05, 2.678084e-05, 
    1.919206e-05, 1.64523e-05, 1.052789e-05, 4.00953e-05, 1.31174e-05,
  1.600211e-07, 2.688183e-06, 2.39225e-05, 2.319378e-05, 3.057891e-05, 
    5.983852e-05, 9.666426e-05, 1.946388e-05, 3.45396e-05, 3.287605e-05, 
    2.377036e-05, 2.550796e-05, 2.235594e-05, 4.232945e-05, 2.329855e-05,
  5.468914e-11, 3.452369e-12, 1.289209e-12, 1.46082e-12, 1.215159e-08, 
    8.853979e-07, 5.183889e-06, 3.266859e-05, 8.687314e-05, 0.0001237987, 
    8.352746e-05, 5.100404e-05, 3.176088e-05, 6.504303e-05, 9.635693e-05,
  1.125878e-14, 8.858763e-11, 1.648613e-10, 5.110799e-10, 4.317327e-09, 
    3.894416e-07, 2.838186e-06, 1.117395e-05, 4.847791e-05, 9.216087e-05, 
    0.0001158012, 9.59363e-05, 8.517325e-05, 9.632137e-05, 0.0002103828,
  4.973348e-11, 2.838504e-09, 2.272803e-08, 1.04315e-07, 3.781794e-07, 
    3.156803e-06, 3.32538e-06, 1.058562e-05, 2.275959e-05, 6.013886e-05, 
    9.342955e-05, 0.0001349958, 0.0001131465, 0.0001373906, 0.0001526842,
  9.936985e-09, 6.836701e-08, 2.892153e-07, 5.392458e-06, 7.899622e-06, 
    1.455111e-05, 1.500603e-05, 1.908313e-05, 2.470365e-05, 8.169714e-05, 
    0.0001553827, 0.0001852504, 0.0001133699, 0.0001699556, 0.0001299939,
  2.433563e-08, 4.07834e-07, 1.666434e-06, 5.989873e-06, 6.585913e-06, 
    1.632783e-05, 2.283361e-05, 2.759859e-05, 5.389082e-05, 0.0001044245, 
    5.522013e-05, 6.509179e-05, 0.0001941699, 0.0001257526, 9.080987e-05,
  2.061052e-08, 9.847821e-07, 1.393776e-06, 4.954711e-06, 1.017514e-05, 
    1.935467e-05, 2.316088e-05, 3.260577e-05, 4.406292e-05, 1.961041e-05, 
    1.663413e-05, 2.769485e-05, 3.106405e-05, 4.735968e-05, 6.433589e-05,
  1.941175e-07, 3.582589e-07, 2.017165e-06, 3.598007e-06, 4.580253e-06, 
    9.243361e-06, 2.121486e-05, 2.416867e-05, 3.176248e-05, 2.664094e-05, 
    2.41216e-05, 1.889577e-05, 1.095004e-05, 3.305018e-05, 5.061977e-05,
  1.50062e-07, 2.533017e-07, 1.551658e-06, 1.510836e-06, 4.930243e-06, 
    7.440978e-06, 1.934395e-05, 2.814163e-05, 5.905468e-05, 2.104368e-05, 
    1.647917e-05, 1.388336e-05, 1.069685e-05, 5.082938e-05, 9.737103e-05,
  1.535155e-07, 1.485925e-07, 6.395917e-07, 2.025176e-06, 9.142485e-06, 
    1.7948e-05, 3.079709e-05, 4.260215e-05, 1.695829e-05, 1.58175e-05, 
    7.629616e-06, 1.394314e-05, 1.716099e-05, 5.191948e-05, 6.012064e-05,
  9.650518e-08, 8.686022e-08, 1.555558e-07, 2.549507e-07, 1.423615e-06, 
    6.740873e-06, 2.047045e-05, 1.502853e-05, 1.42891e-05, 6.50193e-06, 
    4.363009e-06, 9.248497e-06, 1.347795e-05, 3.047114e-05, 2.134466e-05,
  4.651722e-10, 6.020001e-10, 1.608597e-09, 9.750255e-09, 6.075103e-08, 
    1.055812e-07, 5.330954e-08, 3.685112e-09, 2.629774e-10, 3.749033e-08, 
    8.421694e-08, 1.429379e-06, 6.115997e-09, 8.547304e-08, 7.796301e-08,
  3.415915e-09, 4.352328e-09, 2.439916e-08, 2.255556e-07, 3.936763e-07, 
    2.123913e-07, 8.651109e-08, 1.300138e-08, 7.07311e-10, 2.069142e-09, 
    1.225261e-07, 4.408665e-07, 1.030816e-07, 6.428834e-07, 9.268737e-07,
  4.788099e-07, 1.089314e-06, 4.323036e-07, 5.48069e-07, 6.45682e-07, 
    7.026103e-07, 1.51303e-07, 2.080451e-08, 2.371133e-08, 1.353729e-08, 
    2.952018e-09, 2.540221e-07, 1.029971e-06, 3.2342e-06, 3.591186e-06,
  3.214599e-06, 4.861308e-06, 5.318269e-06, 5.684795e-06, 3.404633e-06, 
    4.290373e-06, 1.799517e-06, 6.506129e-07, 2.415476e-07, 6.430685e-07, 
    5.639768e-08, 1.435503e-06, 3.96238e-06, 1.445293e-05, 6.901068e-06,
  4.640053e-06, 4.489496e-06, 1.59187e-06, 1.495161e-06, 2.30302e-06, 
    5.143258e-06, 4.705407e-06, 2.519756e-06, 2.859986e-06, 1.257842e-06, 
    3.815612e-09, 1.345189e-06, 1.500031e-05, 1.925314e-05, 2.452587e-05,
  4.240818e-06, 6.62313e-06, 2.304568e-06, 1.261263e-06, 1.788738e-06, 
    4.124322e-06, 3.167304e-06, 2.377651e-06, 8.010848e-07, 9.797705e-09, 
    1.298123e-06, 4.48869e-06, 5.906141e-06, 3.060562e-05, 2.093995e-05,
  4.388291e-06, 3.341695e-06, 4.670478e-06, 1.244195e-06, 5.341376e-06, 
    4.030687e-06, 3.481623e-06, 9.596192e-07, 7.048651e-09, 9.193035e-08, 
    3.296173e-07, 5.044601e-07, 7.180847e-07, 4.223414e-05, 1.091751e-05,
  9.598914e-08, 4.848881e-06, 1.047017e-05, 5.517887e-06, 2.521952e-06, 
    5.066576e-06, 1.167204e-05, 2.533714e-06, 1.892829e-07, 4.415708e-09, 
    1.131599e-07, 6.875344e-07, 9.543917e-07, 2.934123e-05, 7.493301e-06,
  8.432261e-07, 5.133848e-06, 7.467622e-06, 7.133933e-06, 1.215294e-05, 
    1.314376e-05, 5.889121e-06, 2.965937e-06, 3.109063e-08, 4.731798e-08, 
    3.959872e-07, 3.843098e-07, 4.222267e-06, 1.144066e-05, 4.467717e-06,
  2.214673e-06, 6.333959e-06, 1.025361e-05, 8.192084e-06, 1.150342e-05, 
    1.128544e-05, 6.007292e-06, 1.80443e-06, 2.636218e-07, 3.189181e-07, 
    5.682832e-07, 4.556103e-07, 4.239625e-06, 5.300036e-06, 2.517129e-06,
  6.880104e-10, 6.387124e-10, 9.205846e-10, 4.457008e-10, 3.603709e-09, 
    1.980646e-08, 1.115163e-08, 7.056233e-10, 8.395503e-10, 2.077593e-09, 
    1.380831e-07, 2.334806e-06, 8.180479e-07, 2.129201e-06, 9.329811e-08,
  2.335277e-11, 6.994603e-11, 3.662514e-11, 1.069602e-09, 1.207527e-08, 
    7.280237e-07, 6.121005e-07, 4.865037e-08, 1.199745e-08, 9.230095e-09, 
    2.041076e-09, 5.274394e-08, 2.444665e-07, 3.079651e-07, 3.622345e-09,
  3.142933e-08, 2.044446e-08, 1.31691e-09, 8.762733e-10, 8.198144e-07, 
    1.00654e-06, 5.025717e-07, 1.159253e-06, 7.62795e-08, 4.212903e-08, 
    1.019816e-08, 1.601743e-08, 2.106883e-07, 1.394566e-06, 7.148089e-09,
  3.253008e-07, 3.277964e-08, 4.741394e-08, 3.505793e-07, 3.914074e-07, 
    1.082529e-06, 1.835702e-06, 1.588267e-06, 7.497473e-07, 4.219611e-07, 
    1.859189e-07, 1.008849e-07, 3.319623e-08, 1.07031e-06, 2.943986e-08,
  7.375602e-07, 2.088716e-07, 9.419132e-08, 2.368969e-07, 6.059818e-07, 
    2.620431e-06, 2.103983e-06, 2.208069e-06, 3.958948e-06, 1.182349e-06, 
    1.212882e-08, 1.520185e-08, 1.979642e-08, 8.834858e-07, 1.608894e-07,
  7.074723e-08, 5.134885e-07, 7.287684e-08, 2.040757e-07, 1.264693e-06, 
    2.86705e-06, 4.236898e-06, 4.38238e-06, 2.792178e-06, 6.620262e-09, 
    3.024856e-08, 5.880601e-08, 4.657878e-08, 5.809794e-08, 1.021175e-05,
  2.01182e-09, 5.747453e-08, 7.705039e-08, 1.00219e-07, 1.786292e-06, 
    2.084878e-06, 4.23462e-06, 2.546187e-06, 4.349108e-07, 8.228412e-08, 
    3.938041e-07, 1.008993e-06, 6.067257e-07, 2.615917e-05, 1.027659e-05,
  2.809712e-09, 1.350175e-07, 2.56225e-07, 1.415359e-07, 6.639532e-07, 
    3.754637e-06, 3.692399e-06, 7.947487e-06, 9.650906e-07, 1.704787e-06, 
    7.105044e-06, 1.963326e-05, 1.464405e-05, 6.118472e-05, 3.196482e-06,
  4.765725e-08, 7.251152e-07, 7.281355e-07, 1.761207e-06, 4.218256e-06, 
    5.132645e-06, 5.373092e-06, 8.828988e-06, 9.120718e-07, 9.810851e-06, 
    1.670443e-05, 2.671983e-05, 3.562216e-05, 3.598167e-05, 2.96307e-06,
  1.240612e-06, 8.232509e-07, 1.444493e-06, 1.835753e-07, 3.371256e-07, 
    1.737035e-06, 1.818167e-06, 2.475359e-07, 6.037124e-06, 9.004809e-06, 
    1.218358e-05, 1.410407e-05, 2.601169e-05, 3.574927e-05, 1.470179e-05,
  3.525974e-17, 8.145339e-17, 3.697965e-17, 4.233111e-11, 1.004525e-11, 
    1.752932e-11, 2.580787e-11, 3.858927e-09, 3.27908e-10, 6.585709e-10, 
    1.024746e-08, 1.001483e-06, 2.150123e-06, 1.155091e-05, 4.185094e-09,
  6.762995e-12, 4.364741e-13, 3.317329e-09, 1.586827e-08, 4.645349e-09, 
    3.939878e-09, 4.753907e-08, 1.628838e-07, 2.029421e-09, 6.470958e-09, 
    2.1962e-08, 1.737527e-06, 1.180087e-06, 2.929155e-06, 1.023622e-08,
  1.592965e-07, 6.991439e-08, 8.559224e-09, 1.805992e-10, 3.602411e-07, 
    9.445895e-07, 2.730427e-07, 3.321178e-07, 5.755348e-08, 4.327543e-07, 
    1.618909e-06, 1.878406e-06, 1.643547e-06, 3.10289e-06, 1.11861e-08,
  2.567635e-06, 1.773135e-08, 9.717821e-08, 9.707819e-07, 6.445831e-07, 
    8.329601e-07, 6.787848e-07, 2.884037e-06, 9.405788e-07, 2.537243e-06, 
    6.206335e-06, 5.466643e-06, 3.901329e-06, 2.325876e-06, 2.344436e-06,
  2.959578e-06, 8.199198e-07, 1.712767e-08, 7.066762e-09, 6.294391e-09, 
    2.551052e-07, 1.600745e-06, 2.638412e-06, 2.737639e-06, 1.783324e-07, 
    2.037208e-08, 5.411731e-08, 1.536295e-06, 1.769423e-06, 2.687485e-06,
  2.131263e-07, 6.739896e-08, 7.832115e-09, 1.748274e-08, 1.89588e-07, 
    6.956861e-08, 4.265926e-07, 1.217369e-06, 8.760722e-07, 1.859333e-09, 
    3.333351e-08, 2.753356e-07, 2.821714e-07, 1.157522e-06, 2.664591e-05,
  1.315021e-07, 2.186353e-08, 1.876049e-08, 3.32396e-08, 4.561629e-08, 
    4.048283e-08, 5.263516e-07, 7.356427e-08, 3.590714e-08, 8.596895e-09, 
    4.075871e-08, 1.399415e-07, 1.055044e-06, 5.404333e-05, 3.914207e-05,
  1.919533e-07, 4.592226e-07, 2.021678e-07, 1.333562e-07, 1.542518e-07, 
    3.85682e-07, 5.683918e-07, 2.524505e-06, 2.280141e-07, 1.934746e-07, 
    3.115136e-07, 1.214865e-06, 6.015507e-06, 0.0001163595, 3.836876e-06,
  3.067586e-07, 8.658528e-07, 4.889541e-07, 3.116503e-07, 2.944765e-07, 
    1.835526e-06, 1.432909e-06, 4.086595e-06, 4.461033e-07, 3.59253e-06, 
    5.063059e-06, 5.858848e-06, 2.265259e-05, 4.322045e-05, 6.584776e-06,
  4.173855e-07, 4.882819e-07, 5.349658e-07, 4.025426e-07, 3.154094e-07, 
    2.900939e-07, 2.274165e-07, 2.261192e-07, 2.058281e-06, 6.213299e-06, 
    9.875313e-06, 1.353072e-05, 4.083854e-05, 7.43956e-05, 6.580785e-05,
  3.765449e-10, 2.199587e-09, 4.774977e-09, 1.311091e-09, 2.675772e-09, 
    5.203605e-09, 8.918057e-09, 2.863873e-09, 7.675423e-09, 2.867679e-06, 
    7.857883e-06, 2.20705e-05, 2.421011e-05, 3.641671e-05, 1.013135e-06,
  3.99697e-09, 4.363107e-09, 1.105329e-09, 1.048662e-08, 1.204372e-08, 
    2.36171e-08, 9.740326e-09, 3.326431e-07, 7.075228e-06, 7.860682e-08, 
    2.709718e-06, 1.310767e-05, 1.308842e-05, 4.034581e-05, 8.784025e-07,
  4.107921e-08, 2.260436e-06, 4.225979e-09, 1.242427e-08, 4.285037e-08, 
    1.064232e-06, 5.762378e-07, 3.399936e-06, 2.578107e-07, 1.587153e-06, 
    2.04062e-06, 1.549486e-06, 6.920151e-06, 1.306669e-05, 5.595192e-09,
  1.142563e-07, 2.662626e-07, 2.404072e-07, 1.409723e-06, 3.659424e-06, 
    8.235753e-06, 2.263931e-05, 3.621005e-05, 6.756598e-06, 7.884795e-06, 
    1.385433e-05, 7.577416e-06, 1.947851e-06, 2.713245e-06, 1.980861e-06,
  1.623393e-07, 1.010154e-07, 6.111863e-08, 5.733263e-08, 7.640748e-08, 
    1.1077e-05, 2.786057e-05, 5.46628e-05, 4.815719e-05, 2.471636e-05, 
    8.870391e-08, 4.324478e-06, 2.266266e-05, 1.154735e-05, 7.603747e-06,
  2.217878e-07, 2.324231e-07, 2.466415e-07, 2.49112e-07, 4.623979e-07, 
    5.686318e-07, 1.515116e-05, 4.439536e-05, 4.170046e-05, 1.43001e-06, 
    1.018405e-05, 1.786367e-05, 9.502568e-06, 1.129302e-05, 3.548416e-05,
  1.105655e-07, 2.057391e-07, 4.818057e-07, 6.09992e-07, 8.899768e-07, 
    6.492641e-06, 1.268707e-05, 2.002492e-05, 2.43908e-06, 6.927681e-07, 
    6.616863e-07, 7.533316e-06, 9.040075e-06, 1.58239e-05, 1.810246e-05,
  1.85289e-07, 3.135009e-07, 6.116562e-07, 8.264683e-07, 1.037385e-06, 
    7.520378e-06, 1.094723e-05, 2.581601e-05, 1.037204e-05, 2.061513e-06, 
    2.541492e-06, 1.633168e-05, 1.078763e-05, 1.54331e-05, 8.386345e-06,
  1.822622e-07, 5.466476e-07, 9.310074e-07, 1.001342e-06, 2.461064e-06, 
    6.531657e-06, 7.999815e-06, 2.506637e-05, 2.075108e-06, 1.42713e-05, 
    1.125564e-05, 8.2549e-06, 4.901477e-06, 4.672889e-06, 3.883516e-06,
  1.727559e-07, 5.316681e-07, 1.003295e-06, 1.094516e-06, 9.600114e-07, 
    6.95927e-07, 1.069088e-06, 4.84191e-07, 4.902618e-07, 6.334627e-07, 
    3.815555e-07, 1.979291e-07, 2.193092e-07, 7.472025e-07, 1.191009e-06,
  2.072965e-08, 3.212917e-08, 3.422806e-08, 3.576831e-08, 1.285749e-07, 
    9.375646e-08, 9.41517e-08, 9.856921e-08, 1.416893e-07, 2.565839e-07, 
    2.563589e-06, 1.138854e-05, 1.302532e-05, 2.765957e-05, 2.344235e-05,
  4.201947e-08, 6.828785e-08, 7.328808e-08, 1.104913e-07, 2.255652e-07, 
    2.346235e-07, 1.025865e-07, 1.276547e-07, 1.87212e-07, 3.593153e-07, 
    5.841528e-06, 9.56545e-06, 8.579907e-06, 3.583532e-05, 1.590035e-05,
  9.108388e-08, 1.233911e-07, 9.593669e-08, 1.57446e-07, 2.06249e-07, 
    2.148533e-07, 1.924793e-07, 1.660236e-07, 3.414442e-07, 7.410293e-07, 
    1.366622e-06, 1.993813e-06, 2.169765e-05, 3.585634e-05, 1.908197e-05,
  8.451803e-08, 8.542938e-08, 7.019889e-08, 7.404118e-08, 1.417058e-07, 
    2.02833e-07, 5.778446e-07, 2.426406e-06, 6.067929e-07, 7.684095e-07, 
    6.815065e-06, 1.098927e-05, 7.166021e-06, 1.007369e-05, 2.090774e-05,
  7.36811e-08, 1.871188e-07, 1.187761e-07, 3.529257e-08, 4.690198e-08, 
    1.91627e-07, 8.378374e-07, 3.907716e-06, 1.438227e-05, 1.227991e-05, 
    1.062803e-07, 2.666177e-07, 3.029947e-05, 2.69417e-05, 7.235065e-05,
  1.923757e-07, 1.759732e-07, 1.288496e-07, 1.840538e-08, 2.70542e-08, 
    2.475449e-08, 3.563034e-08, 9.786152e-08, 5.729969e-06, 2.30691e-07, 
    2.332025e-07, 9.354468e-07, 7.242542e-06, 3.790031e-05, 0.0001165958,
  1.577947e-07, 1.173012e-07, 9.214678e-08, 1.404911e-08, 2.802562e-08, 
    3.801329e-08, 2.566164e-06, 1.776227e-07, 8.947113e-07, 1.484001e-07, 
    9.111723e-08, 7.247683e-07, 5.59409e-06, 8.62774e-05, 7.508779e-05,
  1.620504e-07, 1.696147e-07, 7.055271e-08, 3.438655e-08, 1.395433e-08, 
    2.144575e-08, 1.308089e-07, 8.108083e-07, 2.236846e-07, 6.017599e-08, 
    2.429527e-08, 2.495339e-06, 3.064504e-06, 2.698385e-05, 2.21956e-05,
  3.427705e-07, 1.404262e-07, 1.222497e-07, 8.919256e-08, 2.616985e-08, 
    1.66601e-07, 3.006861e-07, 6.314395e-06, 1.944105e-08, 3.869946e-08, 
    1.584494e-08, 2.160349e-08, 4.366441e-08, 8.560684e-06, 3.603134e-06,
  2.316431e-07, 3.156174e-07, 3.463776e-07, 2.722154e-07, 1.217716e-07, 
    2.516201e-08, 1.27305e-08, 2.24784e-08, 1.410736e-08, 1.451515e-08, 
    1.36087e-08, 1.231966e-08, 1.525506e-08, 3.706439e-06, 2.972968e-06,
  4.646727e-08, 3.018044e-08, 3.124423e-08, 3.050046e-08, 4.918075e-08, 
    6.662277e-08, 4.984884e-08, 6.003607e-09, 1.795644e-10, 8.822546e-08, 
    8.746062e-07, 3.047051e-06, 3.911788e-06, 5.794207e-06, 3.851585e-09,
  1.264289e-07, 6.55152e-08, 6.905377e-08, 3.59588e-08, 4.810884e-08, 
    8.353607e-08, 8.390604e-08, 1.378145e-08, 3.308031e-07, 4.712449e-09, 
    1.870271e-06, 1.00696e-05, 1.000534e-05, 1.406797e-05, 1.634336e-09,
  2.449194e-07, 2.438773e-07, 7.204554e-08, 7.112691e-08, 8.245118e-08, 
    1.152676e-07, 5.768873e-08, 1.718923e-08, 1.526025e-08, 8.379188e-09, 
    7.452465e-08, 3.686054e-06, 6.702455e-06, 9.828825e-06, 1.768515e-09,
  2.488284e-07, 2.344962e-07, 1.605688e-07, 1.999981e-07, 1.681941e-07, 
    1.280182e-07, 3.089169e-07, 7.746934e-07, 3.343985e-07, 3.053428e-07, 
    3.230595e-09, 1.506858e-09, 7.55546e-07, 1.698111e-06, 1.374164e-08,
  1.525223e-07, 1.567377e-07, 1.786228e-07, 2.268592e-07, 1.645179e-07, 
    1.030967e-07, 8.514687e-08, 6.091135e-07, 5.33597e-06, 6.105744e-06, 
    2.159723e-09, 2.558746e-09, 4.771126e-07, 4.25991e-07, 2.40052e-07,
  8.671589e-08, 6.769534e-08, 9.44414e-08, 1.234001e-07, 1.127497e-07, 
    7.70147e-08, 5.707183e-08, 3.659552e-08, 1.301966e-07, 1.589426e-09, 
    5.112008e-09, 4.57815e-09, 1.284852e-09, 4.738249e-09, 8.161482e-08,
  1.050092e-07, 7.518965e-08, 5.685655e-08, 5.816274e-08, 6.127988e-08, 
    5.123396e-08, 3.792833e-08, 1.698979e-08, 5.747283e-09, 2.700112e-09, 
    7.188827e-09, 3.693279e-09, 1.460575e-09, 2.335975e-07, 4.831551e-07,
  2.840958e-07, 1.572497e-07, 8.689991e-08, 5.961814e-08, 6.452832e-08, 
    6.447575e-08, 5.541333e-08, 3.813188e-08, 9.964057e-09, 5.736712e-09, 
    3.660093e-09, 4.165125e-09, 7.667125e-09, 4.913706e-08, 4.06188e-07,
  5.293683e-07, 3.664529e-07, 1.994915e-07, 1.413166e-07, 9.482072e-08, 
    1.613898e-07, 3.55413e-07, 1.680977e-06, 1.220608e-09, 3.147197e-09, 
    3.98149e-09, 1.769078e-09, 1.235527e-08, 2.359113e-08, 3.866913e-08,
  5.833627e-07, 6.705537e-07, 5.33783e-07, 4.368153e-07, 2.315847e-07, 
    2.053892e-07, 2.368679e-07, 3.108859e-08, 8.920902e-10, 2.03701e-09, 
    5.980971e-10, 1.370512e-09, 1.607988e-08, 4.367792e-08, 7.708963e-08,
  5.455576e-08, 2.246867e-08, 2.462459e-07, 5.107364e-07, 3.52321e-07, 
    1.505221e-07, 1.792133e-07, 2.325033e-08, 1.724914e-09, 5.7463e-07, 
    1.346664e-06, 2.269662e-06, 2.289461e-06, 2.969328e-05, 2.962663e-05,
  2.351943e-07, 4.945674e-08, 1.260271e-07, 4.229165e-07, 2.931181e-07, 
    3.932017e-07, 8.289997e-08, 4.825293e-08, 1.178325e-08, 2.359905e-09, 
    2.682543e-07, 1.123355e-06, 1.842793e-06, 6.548949e-06, 5.534846e-06,
  3.14763e-07, 9.012604e-08, 9.54681e-08, 2.474302e-07, 2.743839e-07, 
    2.112869e-07, 1.918911e-07, 1.172167e-07, 5.455905e-08, 3.294016e-09, 
    1.507733e-09, 4.16647e-07, 7.399599e-07, 2.244726e-06, 1.679523e-09,
  4.659832e-07, 2.430038e-07, 1.816831e-07, 1.826232e-07, 2.795536e-07, 
    1.574288e-06, 1.262788e-05, 2.015743e-05, 4.399977e-06, 3.225681e-06, 
    4.222808e-09, 6.219527e-10, 2.161341e-08, 1.103055e-09, 5.879168e-10,
  4.648879e-07, 3.873256e-07, 2.386669e-07, 1.979433e-07, 4.3224e-07, 
    4.540162e-06, 1.133301e-05, 1.479869e-05, 1.299428e-05, 2.414783e-05, 
    2.334462e-09, 3.83327e-10, 8.460765e-10, 4.249965e-10, 1.416035e-07,
  3.445583e-07, 3.491743e-07, 3.248645e-07, 3.01467e-07, 1.320868e-06, 
    1.225332e-06, 4.100499e-06, 4.444204e-06, 1.13715e-05, 2.693262e-08, 
    7.637129e-10, 7.010942e-10, 4.743521e-09, 4.933192e-08, 2.306865e-06,
  1.651882e-07, 2.259476e-07, 2.797915e-07, 3.437146e-07, 3.592757e-07, 
    4.347702e-07, 7.088297e-07, 3.610394e-07, 7.594986e-08, 5.13274e-09, 
    2.45177e-09, 4.965508e-09, 1.771233e-08, 1.99336e-08, 1.822447e-07,
  9.356705e-08, 1.377323e-07, 1.983389e-07, 3.387155e-07, 3.998589e-07, 
    3.712561e-07, 3.846671e-07, 2.080554e-06, 6.238716e-07, 4.930822e-09, 
    5.830593e-09, 4.119703e-08, 8.103988e-08, 2.370028e-06, 3.718867e-06,
  8.589721e-08, 1.197666e-07, 2.621386e-07, 1.340154e-06, 1.877672e-06, 
    1.656079e-06, 4.832562e-06, 7.327284e-06, 1.80332e-08, 3.588752e-09, 
    1.917271e-08, 3.133148e-08, 3.07013e-08, 3.529899e-06, 2.396327e-06,
  1.22427e-07, 2.304309e-07, 5.19879e-07, 1.22713e-06, 7.561885e-07, 
    6.632181e-08, 1.01815e-06, 8.021463e-09, 8.539957e-09, 9.879219e-09, 
    3.288661e-08, 5.226436e-08, 7.943783e-09, 3.227383e-09, 3.475609e-07,
  3.763863e-09, 8.628421e-10, 2.125667e-09, 3.315969e-09, 7.592305e-09, 
    1.025056e-08, 8.352155e-09, 6.717614e-09, 1.99736e-06, 7.186248e-06, 
    1.712201e-05, 3.162952e-05, 5.124991e-05, 6.435722e-05, 3.972659e-05,
  1.786307e-08, 1.026219e-08, 5.819758e-09, 4.450043e-09, 1.358542e-08, 
    2.388434e-08, 2.077734e-08, 7.464967e-08, 6.788225e-06, 4.066895e-06, 
    1.314636e-05, 3.335833e-05, 3.793797e-05, 4.910681e-05, 3.087216e-05,
  1.186626e-08, 1.097674e-08, 1.166307e-08, 1.116319e-08, 2.481256e-08, 
    5.008254e-08, 4.849028e-08, 3.960075e-06, 4.302516e-06, 1.463263e-06, 
    4.200982e-06, 1.811442e-05, 1.326571e-05, 2.562317e-05, 3.171305e-05,
  9.157485e-09, 8.25921e-09, 1.130153e-08, 2.233077e-08, 4.998453e-08, 
    7.724567e-08, 1.855521e-06, 9.745847e-06, 1.180225e-05, 9.505737e-06, 
    1.933154e-06, 5.381639e-07, 3.458831e-06, 2.086042e-06, 3.889574e-05,
  1.141215e-08, 9.693794e-09, 1.238127e-08, 2.425968e-08, 4.602844e-08, 
    5.85452e-08, 1.744176e-07, 5.121964e-06, 2.142298e-05, 3.920968e-05, 
    1.987499e-08, 9.079925e-09, 2.725415e-07, 5.924869e-09, 1.805046e-06,
  2.159758e-08, 1.731152e-08, 1.791637e-08, 1.914735e-08, 4.261085e-08, 
    9.252525e-08, 8.521828e-08, 6.93278e-07, 4.855889e-06, 2.491619e-08, 
    1.906886e-08, 1.386348e-08, 1.588326e-08, 6.868625e-08, 5.412874e-06,
  3.089891e-08, 2.611797e-08, 4.322118e-08, 3.887098e-08, 7.716353e-08, 
    1.686275e-07, 1.102241e-07, 5.376675e-08, 9.817204e-08, 2.746098e-08, 
    2.688685e-08, 2.46251e-08, 2.426536e-08, 7.125381e-09, 5.842982e-07,
  7.052347e-08, 4.677011e-08, 9.813541e-08, 7.915284e-08, 1.030969e-07, 
    1.470798e-07, 2.333682e-07, 3.474185e-06, 4.599327e-08, 4.381628e-08, 
    5.574035e-08, 9.274982e-08, 1.047327e-07, 2.464132e-06, 7.905549e-07,
  2.858287e-08, 3.283616e-08, 1.488839e-07, 9.642442e-08, 7.286859e-08, 
    5.09089e-07, 1.98399e-06, 1.850766e-05, 4.473856e-08, 4.859933e-08, 
    5.938553e-08, 5.913801e-08, 3.850073e-08, 5.94873e-09, 2.406602e-08,
  1.82907e-08, 7.538404e-08, 9.682516e-08, 4.967967e-08, 5.788882e-08, 
    3.88357e-08, 2.973343e-06, 3.786399e-08, 3.953107e-08, 2.781778e-08, 
    1.810366e-08, 5.487814e-09, 2.933553e-09, 8.723048e-10, 5.516529e-10,
  3.542403e-10, 2.328998e-10, 8.354291e-10, 1.586958e-09, 1.126027e-09, 
    3.001482e-09, 1.112617e-08, 4.318995e-08, 1.738113e-06, 4.704618e-06, 
    9.223336e-06, 4.070536e-05, 0.0001212035, 0.000134092, 8.628999e-05,
  1.541469e-09, 5.240454e-10, 1.001912e-09, 2.30556e-09, 6.192757e-09, 
    9.636846e-09, 4.292485e-08, 1.145832e-07, 5.102058e-07, 1.623471e-06, 
    6.132329e-06, 3.241728e-05, 7.867518e-05, 7.665592e-05, 2.62896e-05,
  2.982638e-08, 4.177571e-09, 8.780203e-10, 3.826038e-09, 2.594603e-08, 
    4.674334e-08, 8.752787e-08, 5.167489e-07, 1.99973e-06, 8.785781e-08, 
    2.739064e-06, 2.190271e-05, 4.508121e-05, 6.618231e-05, 4.868619e-05,
  4.891646e-09, 1.102379e-09, 2.554657e-09, 8.268402e-09, 5.257885e-08, 
    1.074621e-07, 1.536417e-07, 7.977123e-06, 6.709833e-06, 4.507325e-06, 
    3.574533e-07, 5.250265e-07, 1.863183e-05, 5.552427e-05, 0.0001030591,
  8.042667e-09, 7.007414e-09, 9.476156e-09, 1.450906e-08, 4.178651e-08, 
    1.191406e-07, 1.411656e-07, 3.035814e-07, 7.678649e-06, 6.779193e-06, 
    4.620599e-08, 7.291099e-08, 1.012816e-05, 2.634294e-05, 4.753735e-05,
  2.601517e-08, 2.5821e-08, 1.973982e-08, 1.403908e-08, 3.400077e-08, 
    9.957409e-08, 1.075485e-07, 7.882378e-07, 3.863149e-06, 5.36188e-08, 
    1.427886e-07, 1.19502e-07, 2.828333e-08, 4.789642e-08, 2.218794e-05,
  2.30448e-07, 8.70582e-08, 5.039943e-08, 2.638713e-08, 4.636773e-08, 
    9.92763e-08, 7.262126e-07, 8.861542e-08, 4.537521e-08, 8.574852e-08, 
    1.413821e-07, 1.096947e-07, 1.727481e-08, 9.834906e-07, 7.21591e-06,
  1.959125e-06, 1.119352e-06, 1.321097e-07, 3.749094e-07, 2.325557e-07, 
    1.95689e-07, 6.03059e-07, 1.054618e-06, 3.521335e-08, 7.381688e-08, 
    1.23136e-07, 8.210117e-08, 4.1723e-08, 3.410326e-06, 7.000328e-07,
  1.289835e-05, 2.039432e-05, 1.780986e-06, 2.403428e-06, 2.05003e-06, 
    2.648386e-06, 4.54622e-06, 5.622574e-06, 4.715627e-08, 5.994325e-08, 
    3.441841e-08, 1.967959e-08, 1.532585e-08, 1.261328e-09, 3.994523e-08,
  4.823136e-05, 7.928018e-05, 1.548305e-05, 3.379085e-06, 4.532515e-06, 
    1.236311e-06, 4.621055e-07, 2.825981e-08, 3.892127e-08, 1.994707e-08, 
    7.520129e-09, 5.797258e-09, 1.192049e-09, 3.102782e-11, 4.488149e-09,
  3.499258e-08, 3.285336e-07, 4.106586e-06, 5.56125e-06, 1.641237e-07, 
    4.028656e-10, 3.282221e-10, 2.385652e-09, 1.321532e-08, 4.928917e-08, 
    1.358117e-07, 3.341966e-06, 2.050285e-05, 6.041324e-05, 0.0001182414,
  2.044345e-10, 1.049296e-09, 1.54146e-07, 1.514644e-07, 7.120229e-08, 
    6.36934e-09, 2.767817e-10, 7.645461e-10, 3.781675e-09, 3.419094e-08, 
    1.105436e-07, 2.324889e-06, 2.167801e-05, 7.611843e-05, 0.0001059852,
  2.049748e-07, 1.869889e-08, 5.947608e-10, 1.940336e-08, 3.56989e-07, 
    1.186422e-07, 4.999131e-09, 5.034834e-10, 5.128016e-09, 1.960256e-08, 
    6.148697e-08, 1.551114e-06, 3.548285e-05, 8.350188e-05, 8.906226e-05,
  1.020408e-05, 4.583217e-07, 4.284966e-09, 8.487844e-07, 8.892172e-07, 
    1.587132e-06, 2.040835e-07, 2.006117e-09, 2.729291e-08, 1.359358e-06, 
    4.308388e-08, 9.423471e-08, 1.096277e-05, 3.010842e-05, 7.110343e-05,
  9.37545e-08, 3.935968e-08, 2.85882e-08, 1.619772e-08, 6.279555e-09, 
    5.944337e-09, 2.844732e-09, 5.339765e-10, 8.143621e-08, 1.175396e-06, 
    2.375684e-08, 3.661742e-08, 2.512714e-06, 7.434998e-08, 1.649335e-05,
  6.180127e-07, 2.913043e-06, 1.35443e-06, 8.857512e-07, 1.136441e-06, 
    2.074036e-07, 4.393681e-08, 1.301873e-08, 1.951023e-06, 9.637585e-09, 
    5.389877e-08, 1.645413e-08, 1.627782e-09, 8.060221e-08, 1.446179e-05,
  2.754006e-06, 3.838603e-06, 1.6367e-06, 3.305475e-06, 2.799629e-06, 
    9.183956e-07, 9.992862e-07, 3.172598e-06, 9.675191e-07, 3.653074e-08, 
    6.837477e-08, 9.451031e-09, 3.286811e-09, 5.190388e-08, 1.848552e-06,
  1.988135e-05, 1.353763e-05, 5.01021e-06, 1.279461e-05, 2.014158e-05, 
    9.870134e-06, 1.436964e-05, 3.699058e-05, 4.032168e-07, 6.417992e-08, 
    7.240065e-08, 1.975118e-08, 4.208983e-09, 3.938705e-09, 1.71133e-07,
  4.762342e-05, 6.287866e-05, 3.825705e-05, 3.4891e-05, 4.276731e-05, 
    6.062145e-05, 6.444018e-05, 3.242624e-05, 3.320003e-07, 1.115606e-07, 
    5.500725e-08, 2.127105e-08, 2.822009e-09, 2.820085e-08, 2.784315e-09,
  0.0001088432, 0.000100597, 8.672143e-05, 7.406326e-05, 9.755538e-05, 
    9.437194e-05, 8.119823e-05, 4.83652e-05, 1.067032e-05, 2.10371e-07, 
    5.424534e-08, 2.200862e-08, 2.810038e-09, 8.409219e-09, 8.277831e-13,
  7.203805e-08, 2.670963e-06, 6.979604e-06, 7.246067e-06, 3.854577e-06, 
    4.235636e-07, 1.724613e-08, 8.818923e-09, 1.572017e-06, 1.103844e-06, 
    1.352324e-06, 7.516141e-06, 3.747909e-06, 9.031327e-06, 1.111964e-05,
  1.353178e-10, 2.699251e-10, 1.585289e-07, 1.353022e-05, 1.565857e-05, 
    1.282732e-05, 2.695434e-05, 2.499956e-05, 3.456011e-05, 5.861781e-06, 
    4.275443e-06, 1.317371e-05, 2.985414e-07, 6.701453e-06, 5.309092e-06,
  3.493413e-08, 6.670107e-07, 1.039316e-06, 5.437185e-06, 3.090588e-05, 
    3.339263e-05, 2.798444e-05, 6.354386e-05, 5.261793e-05, 4.346159e-05, 
    3.157074e-05, 2.828217e-05, 5.532161e-06, 2.220511e-05, 5.711475e-06,
  1.041611e-05, 4.092458e-06, 5.556594e-06, 1.919152e-05, 2.911659e-05, 
    3.913826e-05, 4.899446e-05, 6.575637e-05, 0.0001108754, 7.414609e-05, 
    3.56758e-05, 1.040575e-05, 9.514915e-06, 1.650004e-05, 3.338742e-05,
  2.127876e-05, 1.214073e-05, 2.183541e-05, 2.024051e-05, 9.673882e-06, 
    1.771101e-05, 2.912182e-05, 4.868199e-05, 0.0001198964, 0.0001670476, 
    8.356668e-05, 5.090457e-05, 2.466826e-05, 1.347087e-06, 1.966551e-05,
  5.630355e-05, 3.901221e-05, 3.707259e-05, 2.554306e-05, 2.084031e-05, 
    3.168899e-05, 3.623084e-05, 7.461576e-05, 9.557889e-05, 0.0001485737, 
    0.000210531, 0.0002609755, 0.0001110635, 1.37629e-05, 1.968808e-05,
  4.572174e-05, 5.660791e-05, 2.589696e-05, 4.198831e-05, 3.411188e-05, 
    3.034534e-05, 6.082082e-05, 8.458487e-05, 2.548712e-05, 2.09786e-06, 
    3.139091e-05, 0.0001669791, 0.000176959, 2.706684e-05, 7.290827e-06,
  4.923937e-05, 6.327945e-05, 5.35725e-05, 4.87595e-05, 4.858319e-05, 
    4.63371e-05, 9.482273e-05, 0.0001230013, 5.687765e-05, 7.146136e-07, 
    1.267066e-09, 5.413968e-06, 0.0001218636, 0.0001048946, 7.121693e-05,
  7.761458e-05, 0.0001028621, 9.523577e-05, 8.786711e-05, 6.133418e-05, 
    7.581706e-05, 0.0001057394, 0.0001477535, 1.322207e-05, 1.046422e-06, 
    3.376744e-09, 1.812771e-09, 2.808575e-06, 3.88048e-05, 4.436142e-05,
  9.999752e-05, 0.0001180725, 0.000141254, 8.710183e-05, 8.482944e-05, 
    9.227551e-05, 5.495729e-05, 2.463424e-05, 9.551595e-06, 7.416404e-07, 
    9.335148e-09, 3.494433e-09, 8.149533e-09, 2.810853e-06, 2.196643e-06,
  8.757771e-09, 3.823821e-09, 9.770843e-06, 7.256221e-06, 9.710703e-06, 
    3.803447e-05, 5.979094e-05, 6.118381e-05, 9.509616e-05, 8.375035e-05, 
    7.604014e-05, 9.274579e-05, 5.202008e-05, 0.0001057272, 2.996052e-05,
  1.470058e-09, 1.129376e-09, 7.896857e-07, 1.081613e-05, 2.88903e-05, 
    4.665781e-05, 5.916237e-05, 6.105979e-05, 9.028251e-05, 4.348297e-05, 
    8.071591e-05, 8.200323e-05, 0.0001194908, 0.0001404646, 0.0001241714,
  8.658577e-07, 3.557103e-06, 6.45058e-06, 1.660213e-05, 3.515541e-05, 
    6.552543e-05, 5.336802e-05, 8.552454e-05, 4.53779e-05, 2.867561e-05, 
    6.31103e-05, 9.779034e-05, 0.000165575, 0.0002430228, 0.0002202393,
  5.602583e-06, 3.812488e-06, 1.38151e-05, 4.457847e-05, 4.399543e-05, 
    4.501586e-05, 7.260733e-05, 8.76019e-05, 7.230722e-05, 5.837181e-05, 
    4.465884e-05, 4.546782e-05, 7.062606e-05, 0.0001489384, 0.0001021616,
  6.533019e-06, 1.459859e-06, 8.901224e-06, 2.066879e-05, 2.359803e-05, 
    2.992667e-05, 6.257032e-05, 7.084487e-05, 5.843788e-05, 9.296068e-05, 
    2.253302e-06, 1.865967e-05, 0.0001055418, 3.147033e-05, 5.575493e-05,
  3.361986e-06, 7.748913e-06, 9.94646e-06, 2.588412e-05, 2.863134e-05, 
    5.304642e-05, 6.252463e-05, 9.939587e-05, 7.394412e-05, 1.833206e-05, 
    1.201127e-06, 2.08805e-05, 4.755875e-05, 8.479248e-05, 8.407461e-05,
  5.772155e-06, 9.295725e-06, 6.429715e-06, 2.593838e-05, 3.152651e-05, 
    5.544269e-05, 0.0001073483, 8.407836e-05, 9.573998e-05, 2.067779e-05, 
    6.08485e-08, 5.399271e-06, 4.698141e-05, 9.408724e-05, 4.954968e-05,
  1.045492e-05, 1.722842e-05, 2.517707e-05, 2.636706e-05, 3.607451e-05, 
    5.344373e-05, 0.0001381017, 0.0001770935, 0.000159798, 3.796051e-05, 
    1.852681e-07, 4.059068e-07, 9.781526e-05, 0.0001638896, 7.739855e-05,
  1.716888e-05, 3.505008e-05, 2.78363e-05, 3.805285e-05, 5.708894e-05, 
    5.580158e-05, 0.0001074645, 0.0001481925, 8.63059e-05, 2.345957e-05, 
    1.689662e-07, 1.473339e-07, 5.377911e-05, 0.0002467215, 0.0002200048,
  3.42566e-06, 1.826091e-05, 4.539298e-05, 4.383755e-05, 5.309076e-05, 
    4.186644e-05, 2.804197e-05, 1.304089e-05, 2.304906e-05, 5.958047e-06, 
    1.057014e-07, 6.43257e-08, 1.336352e-06, 0.0002052422, 0.0001598557,
  8.120957e-13, 7.344312e-10, 5.325566e-10, 3.584763e-09, 8.26137e-09, 
    5.524064e-08, 4.74704e-07, 1.308531e-06, 1.913134e-05, 2.70035e-05, 
    4.701137e-05, 7.169574e-05, 8.240824e-05, 6.364066e-05, 5.801251e-06,
  1.254091e-11, 1.461052e-09, 3.871489e-08, 5.151383e-08, 2.983618e-07, 
    3.651226e-06, 5.030466e-06, 8.317253e-06, 3.805821e-05, 3.491494e-05, 
    5.594322e-05, 6.779388e-05, 7.150411e-05, 4.488266e-05, 2.241284e-05,
  4.041896e-09, 9.035917e-06, 1.353277e-05, 3.424299e-05, 6.452151e-05, 
    5.970744e-05, 3.397119e-05, 6.387306e-05, 5.231302e-05, 1.795104e-05, 
    2.153556e-05, 5.146486e-05, 5.93563e-05, 4.070826e-05, 6.233079e-05,
  4.902971e-06, 1.61455e-05, 4.392883e-05, 8.680016e-05, 7.309989e-05, 
    0.0001043255, 0.0001237248, 0.0001012702, 8.274683e-05, 6.467182e-05, 
    1.536326e-05, 1.208164e-05, 3.722333e-05, 3.740199e-05, 4.1352e-05,
  3.945512e-06, 3.971411e-05, 6.104983e-05, 7.21679e-05, 4.772696e-05, 
    5.617879e-05, 6.498998e-05, 6.093939e-05, 6.158175e-05, 7.399832e-05, 
    3.72385e-07, 3.522814e-07, 1.367035e-05, 1.483305e-05, 4.501767e-05,
  1.208274e-05, 3.203752e-05, 2.626456e-05, 2.846718e-05, 2.402343e-05, 
    4.073458e-05, 3.905796e-05, 7.334018e-05, 8.015799e-05, 3.985258e-05, 
    1.523433e-05, 9.239156e-06, 8.763155e-07, 9.285816e-07, 8.252853e-06,
  6.221699e-06, 1.403394e-05, 1.429341e-05, 8.410531e-06, 1.698381e-05, 
    1.720797e-05, 9.54175e-05, 6.712458e-05, 5.831342e-05, 7.887995e-06, 
    1.440064e-07, 8.007059e-08, 1.676026e-07, 7.931263e-07, 3.093781e-06,
  2.941e-06, 1.075078e-05, 1.175336e-05, 7.562207e-06, 9.891478e-06, 
    1.811682e-05, 5.971377e-05, 0.0001132665, 0.0001189875, 3.898188e-05, 
    1.500073e-06, 2.61732e-07, 2.437264e-07, 1.896545e-05, 2.132603e-05,
  1.461004e-06, 2.968617e-06, 1.318625e-05, 1.945881e-05, 1.543265e-05, 
    3.108379e-05, 4.090937e-05, 0.0001020598, 0.0001031016, 8.882483e-05, 
    2.266464e-05, 3.15686e-06, 8.751046e-07, 7.541755e-06, 2.177735e-05,
  5.621538e-07, 4.456885e-06, 2.419007e-05, 1.999393e-05, 3.400638e-05, 
    3.570545e-05, 4.034405e-05, 1.027979e-05, 3.730274e-05, 3.981128e-05, 
    2.488233e-05, 1.07116e-05, 1.296311e-06, 1.520756e-06, 4.451761e-06,
  4.643049e-11, 2.189493e-09, 2.145836e-07, 5.792688e-08, 1.019875e-08, 
    2.329483e-07, 7.930478e-07, 3.177056e-09, 8.256908e-09, 6.533613e-07, 
    1.052496e-05, 3.671792e-05, 7.57203e-05, 0.0001005029, 1.512502e-05,
  6.610649e-10, 2.070826e-08, 2.691984e-08, 4.788312e-07, 7.569227e-07, 
    3.683305e-06, 7.396148e-06, 9.260366e-06, 1.662123e-06, 1.242139e-07, 
    4.566815e-06, 2.523771e-05, 7.612888e-05, 7.024456e-05, 3.90991e-05,
  6.529612e-09, 9.884612e-07, 2.114531e-08, 2.723501e-07, 5.429868e-06, 
    1.597601e-05, 2.204951e-05, 2.626834e-05, 1.909344e-05, 5.888442e-06, 
    1.080243e-05, 4.312578e-05, 8.759198e-05, 0.000179414, 0.0001974408,
  5.665972e-09, 8.220224e-07, 1.943282e-06, 7.741944e-06, 1.12289e-05, 
    1.9218e-05, 3.914918e-05, 4.685997e-05, 3.923341e-05, 3.960339e-05, 
    7.16507e-05, 6.345032e-05, 7.68197e-05, 0.00021034, 0.0001791328,
  2.418117e-08, 4.471422e-07, 6.899635e-07, 5.149593e-06, 6.806173e-06, 
    1.89221e-05, 2.717736e-05, 4.239235e-05, 5.235766e-05, 0.0001412941, 
    8.463889e-05, 4.714197e-05, 0.0001419797, 8.239182e-05, 0.0001071141,
  4.440222e-10, 2.914494e-07, 1.840787e-06, 1.422849e-06, 4.201946e-06, 
    1.714531e-05, 3.576504e-05, 2.9489e-05, 8.81461e-05, 9.628351e-05, 
    0.0001247665, 0.0001309142, 8.190547e-05, 6.183796e-05, 7.122788e-05,
  3.291276e-08, 1.26637e-06, 1.741642e-07, 7.019145e-07, 4.604368e-06, 
    1.768213e-05, 5.013137e-05, 4.144044e-05, 3.759212e-05, 1.804018e-05, 
    1.754244e-05, 3.499865e-05, 5.818503e-05, 9.533801e-05, 7.795245e-05,
  2.610404e-08, 1.072369e-06, 1.344715e-06, 5.507663e-07, 3.968596e-06, 
    4.450909e-06, 2.260997e-05, 2.715658e-05, 4.7494e-05, 1.123341e-06, 
    1.55994e-06, 4.041108e-06, 2.286953e-05, 0.0001262901, 0.0001016969,
  1.200391e-09, 1.269891e-07, 2.445253e-06, 3.751615e-06, 8.065328e-06, 
    8.993203e-06, 1.686865e-05, 3.147371e-05, 1.081384e-05, 4.055932e-06, 
    2.107161e-06, 1.510761e-06, 8.046953e-06, 0.0001467643, 0.0001998574,
  8.460475e-10, 1.364526e-07, 1.727572e-06, 4.129639e-06, 8.45069e-06, 
    1.356003e-05, 1.962946e-05, 9.524842e-06, 8.475952e-06, 6.868466e-07, 
    3.005761e-06, 2.591607e-06, 1.151147e-05, 0.0001103599, 0.0001617906,
  4.078667e-13, 3.344979e-14, 7.369402e-12, 5.507e-19, 3.545878e-14, 
    1.045532e-13, 1.331702e-14, 9.560014e-10, 5.165658e-07, 3.638311e-05, 
    5.779487e-05, 6.259017e-05, 3.474365e-05, 2.208255e-05, 1.400303e-05,
  1.713127e-11, 1.04736e-23, 4.185977e-24, 2.364469e-24, 1.256845e-17, 
    1.119479e-15, 1.476837e-14, 1.61566e-08, 1.418725e-06, 1.599888e-05, 
    3.193339e-05, 2.629727e-05, 1.686497e-05, 4.482125e-05, 7.590331e-05,
  1.399422e-10, 1.036525e-11, 4.960373e-14, 1.160434e-12, 1.406547e-10, 
    5.150912e-09, 2.020816e-08, 1.323871e-07, 2.544193e-06, 2.236679e-06, 
    1.257993e-05, 1.816776e-05, 2.107237e-05, 0.0001056507, 0.0002247876,
  8.639293e-11, 5.029789e-12, 1.107685e-12, 2.772003e-08, 1.600239e-08, 
    1.157919e-07, 4.029973e-07, 1.828266e-06, 5.44667e-06, 1.99517e-05, 
    5.590012e-05, 5.915237e-05, 5.316282e-05, 0.0002207053, 0.0001868914,
  6.06182e-11, 5.201496e-13, 1.489361e-13, 8.362434e-08, 2.191171e-07, 
    1.082183e-06, 1.885455e-06, 8.864572e-06, 2.434716e-05, 5.746507e-05, 
    5.663525e-06, 9.23045e-06, 0.0001729746, 0.000187732, 0.0001564098,
  2.020604e-11, 2.377916e-09, 3.547149e-13, 2.191692e-08, 8.169147e-07, 
    2.573602e-06, 5.999043e-06, 1.353903e-05, 3.532223e-05, 1.098374e-05, 
    3.767872e-06, 1.85879e-06, 4.686352e-05, 0.0001235706, 0.0001667552,
  3.027818e-11, 5.075588e-13, 5.571042e-13, 9.897723e-08, 7.852508e-07, 
    1.823123e-06, 6.142936e-06, 1.064379e-05, 9.626811e-06, 1.13456e-06, 
    1.457888e-06, 1.737523e-06, 1.611038e-05, 4.919183e-05, 0.0001234968,
  1.091944e-10, 1.317842e-12, 1.703427e-14, 2.289593e-10, 7.880264e-08, 
    1.595426e-07, 2.28915e-06, 5.962722e-06, 7.77537e-06, 1.872576e-06, 
    4.889732e-06, 2.005397e-06, 3.361507e-07, 3.889026e-05, 7.604437e-05,
  1.234201e-09, 1.451464e-10, 1.527266e-11, 4.266283e-10, 4.211097e-10, 
    3.367663e-08, 1.164183e-06, 7.101853e-06, 2.1878e-07, 1.945964e-06, 
    2.541182e-06, 4.766546e-06, 3.295962e-06, 1.533517e-05, 6.799219e-06,
  2.639789e-09, 1.826941e-09, 8.078938e-10, 1.282467e-09, 2.242375e-10, 
    5.016193e-11, 4.137641e-08, 2.229483e-08, 4.015179e-08, 3.202717e-07, 
    2.150365e-06, 3.198563e-06, 6.940577e-06, 2.350365e-05, 1.26052e-05,
  4.632667e-08, 4.25781e-09, 1.458398e-09, 1.031617e-09, 2.208635e-09, 
    2.067081e-09, 1.206908e-09, 5.260327e-10, 1.465158e-08, 2.308602e-06, 
    1.474863e-05, 2.704209e-05, 4.272881e-05, 2.761275e-05, 2.317251e-05,
  3.58047e-09, 7.141933e-10, 2.493594e-09, 6.659972e-09, 8.395864e-09, 
    5.612348e-09, 2.038813e-11, 3.472353e-12, 1.11047e-09, 1.127346e-08, 
    3.050555e-06, 9.793733e-06, 1.452403e-05, 3.393094e-05, 1.137742e-05,
  1.612636e-08, 2.350659e-09, 4.60902e-09, 1.390862e-08, 3.666118e-08, 
    6.919605e-08, 1.582287e-08, 1.438334e-09, 1.983947e-08, 6.797066e-07, 
    1.220101e-06, 1.107376e-05, 2.507849e-05, 6.257244e-05, 1.716565e-05,
  1.42378e-07, 1.257878e-08, 9.436074e-09, 2.090436e-08, 6.919785e-08, 
    4.623071e-07, 3.051697e-07, 2.236352e-07, 3.460255e-07, 7.724609e-07, 
    1.236271e-06, 4.270946e-06, 2.828936e-05, 6.747998e-05, 2.168937e-05,
  1.279348e-06, 4.973127e-08, 1.511277e-08, 1.699044e-08, 5.17186e-08, 
    8.689211e-08, 1.243441e-06, 1.447822e-06, 1.838767e-06, 7.081884e-06, 
    5.065575e-07, 2.291295e-07, 3.126304e-05, 3.597111e-05, 1.819248e-05,
  3.704004e-06, 5.538943e-07, 1.707779e-07, 1.354754e-08, 2.138041e-08, 
    2.967626e-08, 2.205468e-07, 6.899846e-07, 5.13563e-06, 1.478813e-06, 
    1.2647e-06, 2.889878e-07, 1.376817e-05, 4.825493e-06, 2.470021e-05,
  2.217037e-06, 3.630644e-06, 2.337823e-06, 1.354822e-08, 1.125944e-08, 
    1.922219e-08, 1.71954e-07, 2.069685e-06, 1.661245e-06, 9.403498e-07, 
    6.038402e-08, 1.087235e-08, 2.728955e-06, 3.773881e-06, 2.372754e-05,
  2.038466e-05, 3.431978e-05, 1.618622e-05, 1.219679e-08, 9.601791e-09, 
    1.702677e-08, 3.308246e-07, 1.407102e-06, 1.693225e-07, 1.19626e-08, 
    2.28603e-09, 1.569107e-06, 2.721225e-07, 1.242376e-05, 1.672098e-05,
  2.999458e-05, 7.849782e-05, 4.031268e-05, 9.206721e-09, 7.610747e-09, 
    2.602403e-08, 1.035866e-07, 7.779514e-08, 8.398119e-09, 9.640905e-11, 
    4.686659e-08, 1.351941e-06, 5.807705e-08, 7.514823e-06, 5.733229e-06,
  9.585795e-06, 5.673408e-05, 5.336307e-05, 1.908474e-08, 6.044079e-09, 
    1.528878e-09, 9.350308e-10, 7.896429e-10, 1.480569e-11, 1.332463e-10, 
    2.239005e-09, 5.221584e-09, 4.377083e-10, 2.5748e-06, 3.657799e-07,
  1.178354e-05, 4.793263e-06, 4.703525e-06, 7.558537e-07, 6.155748e-06, 
    2.363363e-05, 4.371726e-05, 5.715968e-05, 0.0001160483, 9.698517e-05, 
    4.889975e-05, 2.595156e-05, 1.159356e-05, 1.207434e-05, 5.763963e-06,
  6.741015e-08, 5.659302e-08, 2.081076e-06, 2.597083e-06, 2.946592e-05, 
    4.454676e-05, 5.451639e-05, 5.945272e-05, 8.71661e-05, 6.476976e-05, 
    3.96396e-05, 1.485666e-05, 4.606805e-06, 3.370348e-06, 4.802964e-07,
  8.867806e-09, 1.951218e-05, 6.321789e-06, 5.466452e-06, 4.224918e-05, 
    4.022059e-05, 1.698089e-05, 1.630744e-05, 2.796477e-05, 2.810591e-05, 
    2.405535e-05, 1.570415e-05, 8.600189e-06, 4.977891e-06, 8.449694e-07,
  3.732287e-05, 2.048403e-06, 1.712286e-06, 4.23948e-05, 5.101265e-05, 
    3.423006e-05, 9.555055e-06, 3.248269e-06, 6.39475e-06, 5.832958e-06, 
    8.066137e-06, 2.388159e-06, 7.577627e-06, 1.719784e-06, 1.170176e-05,
  4.845068e-05, 2.402118e-05, 2.997292e-05, 4.530457e-05, 2.196856e-05, 
    8.899169e-06, 3.685018e-06, 6.574538e-06, 3.935178e-06, 2.496113e-06, 
    7.24757e-09, 4.617585e-10, 7.470548e-10, 3.995608e-08, 1.422519e-05,
  0.0001120036, 0.000125324, 0.0001380295, 8.036834e-05, 3.232761e-05, 
    2.667645e-05, 3.110619e-05, 1.763508e-05, 3.722628e-06, 1.205213e-09, 
    1.312157e-08, 7.874409e-10, 2.067693e-12, 1.90081e-07, 1.584953e-05,
  0.0001607665, 0.0002481373, 0.0002763715, 0.0001060966, 5.699212e-05, 
    5.817432e-05, 3.991175e-05, 6.164624e-06, 1.015918e-06, 5.0347e-10, 
    4.18874e-12, 1.746133e-11, 1.580899e-10, 3.413953e-08, 2.809108e-06,
  9.128867e-05, 0.0002257048, 0.0002633741, 5.918145e-05, 2.780416e-05, 
    2.719065e-05, 7.331688e-06, 2.414455e-06, 8.484009e-07, 3.228509e-11, 
    1.153937e-12, 2.684482e-11, 1.446791e-09, 5.015164e-07, 1.902876e-07,
  4.259677e-05, 8.14778e-05, 0.000150241, 3.009191e-05, 4.537585e-06, 
    4.597132e-06, 6.890119e-07, 1.682161e-07, 5.855357e-08, 5.017462e-13, 
    1.237641e-11, 6.736618e-10, 3.303399e-10, 1.722166e-08, 1.893769e-08,
  1.208604e-05, 3.088643e-05, 9.002872e-05, 7.55577e-06, 2.318797e-06, 
    2.674568e-08, 9.008467e-09, 7.958403e-11, 6.78988e-11, 3.171633e-11, 
    2.829045e-10, 1.440323e-09, 5.110985e-10, 5.74351e-09, 1.294449e-07,
  5.897932e-05, 6.766114e-05, 0.0001352338, 0.0001181412, 0.0001547681, 
    0.000161876, 0.0001669618, 0.0001600127, 0.0002338177, 0.0001777431, 
    0.0001424141, 0.0001711089, 0.0001645255, 9.162596e-05, 0.0001015727,
  5.186186e-06, 4.592095e-05, 0.0001267069, 0.0001651608, 0.0002766512, 
    0.0001971382, 0.0001789373, 0.0001769145, 0.0002697512, 0.000229313, 
    0.000240129, 0.0002347766, 0.000173154, 6.938938e-05, 5.606897e-05,
  8.640268e-05, 0.0001847266, 5.139556e-05, 0.0001211627, 0.000198636, 
    0.0001496383, 0.000102279, 0.0001990858, 0.0002240257, 0.0001693866, 
    0.0001502889, 0.0001552578, 0.0001398335, 8.965662e-05, 6.818349e-05,
  0.0002033577, 0.000203466, 0.0001410112, 0.000129131, 0.0001065008, 
    9.354339e-05, 6.544466e-05, 0.0001166876, 0.0001464355, 7.025803e-05, 
    7.459829e-05, 6.213509e-05, 6.780114e-05, 6.071509e-05, 9.164227e-05,
  8.935698e-05, 0.0001060566, 0.0001258906, 0.0001649451, 0.0001943276, 
    0.0001450324, 0.0001278125, 0.0001298692, 7.853468e-05, 3.497404e-05, 
    3.181155e-06, 3.340355e-06, 2.074947e-05, 1.684325e-05, 6.152633e-05,
  4.082157e-05, 0.0001019166, 0.0001091717, 0.0001403862, 0.0001681964, 
    0.0001197668, 8.057784e-05, 6.495322e-05, 4.224118e-05, 1.418391e-07, 
    1.977163e-07, 2.907165e-07, 7.85799e-07, 5.652358e-07, 7.057e-05,
  7.886235e-05, 0.0001763349, 0.0001756524, 0.000125596, 8.774021e-05, 
    0.0001043963, 0.000106493, 6.249269e-05, 1.804591e-05, 1.300494e-08, 
    2.177143e-09, 1.518551e-09, 2.178185e-09, 5.724116e-06, 2.13824e-05,
  8.652725e-05, 0.0001281948, 0.0001910258, 0.0001312729, 6.739797e-05, 
    7.602462e-05, 7.168364e-05, 2.148541e-05, 9.138446e-07, 2.561484e-09, 
    1.716519e-09, 5.266708e-09, 3.162556e-09, 8.556023e-06, 2.454423e-06,
  5.610986e-05, 8.508746e-05, 0.0001352119, 0.0001028537, 3.647692e-05, 
    3.110327e-05, 1.122999e-05, 3.849352e-06, 1.960226e-09, 8.622164e-10, 
    9.836535e-10, 2.748093e-09, 1.563083e-09, 1.116286e-05, 1.123195e-05,
  2.918831e-05, 5.818615e-05, 9.350461e-05, 2.757777e-05, 2.22693e-05, 
    7.457571e-06, 1.522786e-08, 5.399393e-09, 5.411512e-10, 4.272064e-10, 
    1.07248e-09, 9.008341e-10, 2.858281e-10, 4.574959e-07, 1.013546e-10,
  8.544682e-06, 1.028106e-05, 7.452602e-05, 4.198961e-05, 3.942089e-05, 
    4.777115e-05, 6.129546e-05, 1.727097e-05, 6.798611e-05, 6.037097e-05, 
    4.763028e-05, 3.905063e-05, 6.820951e-05, 7.534054e-05, 2.386716e-05,
  1.473586e-05, 5.059501e-05, 0.0001043825, 0.0001204382, 5.115163e-05, 
    7.046685e-05, 5.42668e-05, 4.799102e-05, 7.787022e-05, 3.939121e-05, 
    2.980948e-05, 3.049267e-05, 4.977803e-05, 5.638e-05, 3.069713e-05,
  0.0001171614, 0.000161612, 9.939473e-05, 6.979934e-05, 0.0001082439, 
    0.0001010614, 0.0001270624, 0.0001509496, 7.521887e-05, 2.620994e-05, 
    2.562007e-05, 3.63555e-05, 6.246312e-05, 6.7633e-05, 3.59539e-05,
  6.451879e-05, 0.000108891, 0.0001739323, 0.0001570487, 8.305829e-05, 
    0.0001607817, 0.0002476791, 0.00026595, 0.0001516896, 6.377497e-05, 
    1.877562e-05, 1.928281e-05, 8.106294e-05, 6.538431e-05, 6.285024e-05,
  1.604747e-05, 6.309336e-05, 0.0001820076, 0.0002172804, 0.0001338628, 
    0.0001801758, 0.0002306749, 0.0002984872, 0.0002465867, 9.27107e-05, 
    6.726971e-07, 1.620374e-07, 2.837753e-05, 7.484583e-05, 0.000122068,
  2.570568e-06, 3.690001e-05, 0.0001137821, 0.0001938359, 0.0001920772, 
    0.000114059, 8.083254e-05, 0.0001098549, 0.0001838694, 8.193407e-05, 
    6.042988e-05, 4.215083e-06, 8.565141e-08, 3.330283e-06, 7.169216e-05,
  9.283347e-06, 1.569934e-05, 3.932556e-05, 5.758779e-05, 6.089915e-05, 
    2.349905e-05, 9.655934e-06, 4.815472e-06, 1.679909e-07, 2.731359e-08, 
    5.65614e-09, 1.284458e-08, 1.429042e-08, 2.742123e-05, 4.002679e-05,
  2.038765e-06, 2.582449e-06, 7.165466e-06, 3.605019e-06, 2.830198e-06, 
    3.983592e-06, 2.13916e-06, 5.576467e-06, 1.516187e-06, 5.973028e-09, 
    1.138259e-09, 2.793843e-09, 8.911513e-09, 1.452065e-05, 2.932819e-05,
  8.00381e-07, 8.319128e-07, 2.883269e-06, 2.999297e-06, 3.4344e-06, 
    1.328012e-05, 1.383614e-05, 1.810565e-05, 4.552393e-08, 2.477533e-09, 
    1.55726e-09, 7.031156e-10, 2.935646e-09, 3.563713e-06, 2.809652e-06,
  1.602919e-07, 8.901387e-07, 2.639979e-06, 2.962128e-06, 2.665763e-06, 
    4.828692e-06, 2.985771e-06, 6.904042e-08, 1.120087e-08, 8.534556e-09, 
    2.375059e-09, 6.721943e-10, 1.018359e-09, 8.095433e-07, 1.236413e-06,
  3.845888e-06, 3.934804e-05, 8.862641e-05, 5.114084e-05, 2.670386e-05, 
    4.049628e-05, 3.770534e-05, 3.124481e-06, 3.593176e-05, 4.055894e-05, 
    5.807437e-05, 8.20948e-05, 7.703985e-05, 5.680852e-05, 5.547231e-06,
  3.412048e-07, 1.289499e-05, 0.0001081697, 0.0001532776, 8.465416e-05, 
    6.345478e-05, 4.340194e-05, 4.257981e-05, 4.720933e-05, 2.963961e-05, 
    4.976652e-05, 4.498349e-05, 5.869887e-05, 4.742798e-05, 5.36862e-06,
  1.216862e-06, 2.872128e-06, 2.772074e-05, 8.258205e-05, 0.000125818, 
    7.932131e-05, 0.0001106184, 9.728234e-05, 5.965645e-05, 2.597372e-05, 
    3.295401e-05, 3.883946e-05, 3.908493e-05, 5.313845e-05, 1.736241e-05,
  7.957316e-07, 2.314297e-06, 3.123375e-05, 8.28441e-05, 6.848488e-05, 
    4.105843e-05, 5.785065e-05, 0.0001096536, 0.0001093368, 5.342282e-05, 
    1.454582e-05, 2.884394e-05, 5.504128e-05, 8.652644e-05, 9.671677e-05,
  3.386449e-06, 3.34391e-07, 7.190926e-06, 3.146609e-05, 2.493392e-05, 
    2.844004e-05, 2.226392e-05, 5.283343e-05, 8.838192e-05, 4.767591e-05, 
    1.082502e-06, 1.787339e-07, 1.283551e-05, 2.721072e-05, 8.782721e-05,
  1.84124e-07, 2.632717e-07, 6.764577e-07, 7.155631e-06, 2.213292e-05, 
    2.900835e-05, 2.531922e-05, 1.521045e-05, 4.311178e-05, 2.207756e-05, 
    2.132655e-05, 1.132599e-06, 1.630335e-07, 7.80663e-06, 2.563972e-05,
  8.067667e-09, 2.781989e-08, 4.255673e-08, 2.265981e-06, 1.173516e-05, 
    1.417931e-05, 1.119358e-05, 6.961068e-06, 2.019651e-07, 9.917209e-09, 
    1.347015e-08, 5.295976e-08, 8.19398e-08, 2.489629e-05, 2.428076e-05,
  5.325606e-08, 1.191915e-08, 2.521813e-07, 8.493578e-08, 6.589211e-07, 
    1.963662e-06, 5.737822e-06, 6.99498e-06, 5.18138e-07, 1.610102e-09, 
    2.425233e-09, 3.469662e-08, 1.2782e-07, 2.687833e-05, 3.859404e-05,
  6.518196e-08, 1.284427e-08, 8.455245e-08, 2.933693e-07, 7.895433e-07, 
    2.955444e-06, 5.150921e-06, 4.455619e-06, 1.48627e-08, 4.57331e-08, 
    2.363537e-09, 5.749247e-09, 6.269206e-08, 2.761858e-06, 6.663323e-06,
  6.330785e-08, 3.525593e-08, 3.743831e-08, 1.704572e-08, 2.589219e-07, 
    1.641639e-07, 5.058868e-07, 1.123304e-07, 2.217281e-08, 6.646646e-08, 
    5.657574e-09, 5.438838e-09, 1.229476e-08, 8.395466e-07, 3.920211e-06,
  4.94221e-08, 1.497278e-08, 1.007355e-06, 1.866292e-06, 4.60639e-07, 
    5.917354e-06, 1.810532e-05, 1.715346e-05, 2.028868e-05, 1.390333e-05, 
    3.923964e-05, 3.625695e-05, 4.715697e-05, 6.72942e-05, 6.878933e-05,
  1.772547e-07, 2.690163e-08, 5.729995e-06, 1.773396e-06, 6.165638e-09, 
    1.284694e-06, 7.501405e-06, 1.691761e-05, 3.969272e-05, 2.680374e-05, 
    2.383824e-05, 2.710779e-05, 4.198213e-05, 7.220513e-05, 8.29355e-05,
  2.038533e-07, 6.196211e-06, 1.277685e-05, 1.273462e-07, 1.564132e-07, 
    9.814637e-08, 4.614504e-07, 9.392303e-07, 1.391115e-05, 3.059559e-05, 
    2.410568e-05, 4.630382e-05, 3.9721e-05, 5.420683e-05, 7.589931e-05,
  4.21256e-07, 3.381579e-06, 1.77062e-06, 5.880674e-06, 9.64293e-07, 
    7.30221e-07, 8.263205e-07, 2.700295e-06, 5.437977e-06, 1.627718e-05, 
    9.723411e-06, 2.595961e-05, 2.534326e-05, 5.624253e-05, 2.218857e-05,
  8.874684e-07, 6.850772e-07, 3.833808e-07, 7.356256e-07, 4.536215e-07, 
    6.329091e-07, 2.966248e-07, 8.313349e-07, 3.910928e-06, 7.036014e-06, 
    3.218319e-07, 6.674209e-07, 3.694637e-06, 1.290737e-05, 2.063192e-05,
  1.38392e-06, 1.635847e-06, 3.447243e-06, 3.032423e-06, 3.200441e-06, 
    7.311844e-07, 5.89471e-07, 1.684238e-07, 8.810354e-07, 6.235278e-09, 
    2.522491e-08, 5.998143e-08, 1.512255e-08, 5.38773e-06, 3.335403e-06,
  3.859019e-06, 2.767862e-06, 8.092145e-06, 1.070491e-05, 5.950378e-06, 
    4.37282e-06, 2.068487e-06, 6.599137e-07, 6.90439e-09, 1.825208e-09, 
    5.219152e-10, 8.082201e-08, 3.284994e-08, 1.473787e-05, 3.440085e-06,
  5.956949e-06, 9.610014e-06, 1.692824e-05, 1.21605e-05, 1.287381e-05, 
    1.220436e-05, 5.20124e-06, 4.424404e-06, 1.180963e-08, 5.177234e-09, 
    2.428674e-10, 8.192622e-08, 3.388059e-08, 1.855267e-05, 6.718014e-06,
  8.193772e-06, 8.021522e-06, 1.766907e-05, 2.56417e-05, 1.666767e-05, 
    9.681154e-06, 8.991249e-06, 1.744894e-05, 2.209026e-08, 9.091773e-09, 
    1.791608e-08, 3.946105e-09, 1.722975e-08, 9.612179e-06, 2.094184e-06,
  1.26842e-06, 1.35145e-06, 6.866372e-06, 3.778995e-06, 2.195534e-06, 
    7.425925e-07, 2.474584e-06, 1.480942e-08, 1.299265e-08, 8.677381e-09, 
    5.726181e-09, 1.206781e-09, 4.157584e-09, 5.466572e-06, 2.82689e-06,
  1.1399e-08, 3.200493e-09, 2.532343e-09, 1.109478e-06, 1.91333e-08, 
    3.627516e-09, 3.13673e-09, 3.259746e-10, 1.926222e-10, 7.67808e-11, 
    2.988609e-09, 9.268573e-08, 1.350692e-09, 1.694547e-07, 9.446994e-07,
  7.492781e-08, 1.952894e-08, 5.527074e-08, 2.055954e-07, 1.560368e-07, 
    1.053421e-06, 3.688158e-07, 4.658276e-07, 6.120302e-06, 3.695019e-06, 
    5.506191e-06, 3.896455e-06, 8.537249e-10, 2.550129e-09, 1.194111e-08,
  1.744991e-07, 1.729428e-07, 3.588672e-07, 1.21876e-06, 2.015731e-06, 
    1.787179e-06, 2.439142e-06, 8.135731e-06, 2.738504e-05, 2.979502e-05, 
    1.715051e-05, 1.338609e-05, 4.785035e-06, 2.974542e-07, 7.591094e-10,
  4.412311e-07, 3.289904e-07, 3.095419e-06, 6.07827e-06, 3.283968e-06, 
    7.424596e-06, 4.775166e-06, 2.4576e-05, 3.799791e-05, 5.748147e-05, 
    1.349392e-05, 1.425917e-05, 1.125185e-05, 7.024385e-10, 2.163165e-10,
  1.662645e-06, 1.943806e-06, 2.887254e-06, 2.033219e-06, 2.560887e-06, 
    4.472903e-06, 6.288518e-06, 9.624882e-06, 3.542979e-05, 5.564016e-05, 
    1.214652e-09, 1.136901e-09, 3.858852e-09, 2.362339e-09, 5.003248e-09,
  2.772424e-06, 5.292679e-06, 2.555453e-06, 2.674249e-06, 5.731684e-06, 
    6.970379e-06, 1.092706e-05, 6.515766e-06, 2.67973e-05, 3.814699e-09, 
    4.02117e-09, 6.963134e-09, 1.180767e-08, 5.425161e-08, 7.404253e-07,
  1.495001e-05, 6.746074e-06, 4.534787e-06, 7.905692e-06, 3.960006e-05, 
    6.094579e-06, 9.406073e-06, 1.994158e-05, 1.474244e-05, 4.855028e-09, 
    2.550831e-09, 7.23495e-09, 1.012522e-08, 1.12714e-08, 1.144741e-07,
  3.051791e-05, 3.3536e-05, 2.463125e-05, 2.258246e-05, 1.842064e-05, 
    2.429853e-05, 1.059181e-05, 3.087858e-05, 3.495025e-05, 1.193297e-06, 
    8.241974e-09, 8.171089e-09, 1.358764e-08, 1.996782e-08, 1.742882e-08,
  6.026265e-05, 0.000101001, 9.402265e-05, 7.428901e-05, 8.861448e-05, 
    8.930112e-05, 3.601406e-05, 4.656701e-05, 1.275131e-06, 5.346888e-06, 
    3.867493e-08, 1.679934e-08, 4.223763e-08, 2.352668e-08, 1.360768e-08,
  1.293248e-05, 4.996263e-05, 7.557716e-05, 6.188956e-05, 0.0001043089, 
    7.951829e-05, 5.3704e-05, 1.341206e-05, 2.613709e-05, 1.263043e-05, 
    9.185074e-07, 3.32205e-08, 4.635507e-09, 1.475583e-08, 1.809148e-09,
  9.067755e-08, 5.318672e-08, 1.316966e-06, 2.325816e-08, 7.626298e-09, 
    1.826668e-09, 2.704381e-09, 1.816289e-09, 4.048932e-09, 7.100166e-08, 
    5.158392e-07, 1.19199e-06, 3.466875e-07, 1.601308e-06, 4.129656e-09,
  1.040406e-07, 6.740706e-08, 4.539529e-08, 2.37399e-08, 1.163507e-08, 
    1.988539e-07, 4.940061e-09, 3.030089e-09, 9.0519e-08, 1.330802e-06, 
    5.700772e-06, 4.493277e-06, 3.623936e-07, 5.803968e-07, 2.890949e-09,
  1.124171e-07, 9.802724e-08, 6.519185e-08, 3.273427e-08, 6.939492e-07, 
    3.619657e-06, 2.017569e-06, 6.40256e-06, 4.739638e-06, 4.236647e-06, 
    3.501958e-06, 9.635919e-06, 4.539514e-06, 4.894758e-06, 1.005385e-09,
  1.232365e-06, 1.238161e-07, 2.703269e-06, 5.136323e-06, 3.85614e-06, 
    8.713097e-06, 1.732021e-05, 1.160092e-05, 1.225271e-05, 8.433145e-06, 
    3.442178e-06, 2.79519e-06, 8.758453e-06, 3.622907e-06, 1.445294e-07,
  1.741396e-05, 1.744734e-07, 3.45838e-07, 1.16728e-06, 1.503206e-06, 
    4.524426e-06, 7.920629e-06, 1.981896e-05, 8.978307e-06, 6.107794e-06, 
    4.216372e-09, 4.687039e-10, 2.548526e-06, 5.597944e-10, 8.158323e-06,
  6.55599e-05, 1.018163e-05, 1.596714e-07, 1.261917e-06, 1.328822e-06, 
    3.274065e-06, 2.251707e-06, 5.127718e-06, 5.231762e-06, 9.408291e-09, 
    4.689351e-09, 1.626072e-09, 1.338507e-10, 5.356454e-09, 3.689572e-07,
  0.0001104204, 4.195141e-05, 8.09386e-06, 9.824445e-06, 1.337628e-05, 
    4.333249e-06, 6.790717e-06, 1.266139e-06, 2.885406e-06, 6.583719e-08, 
    2.804761e-08, 1.150773e-08, 1.46153e-09, 6.315314e-07, 3.81663e-07,
  0.0002154948, 0.0001717493, 4.677657e-05, 1.635529e-05, 2.020414e-05, 
    2.233962e-05, 1.280684e-05, 1.50414e-05, 5.940095e-06, 5.340401e-06, 
    2.326461e-06, 2.737074e-06, 3.267625e-07, 5.238243e-06, 9.671799e-07,
  0.0003042132, 0.0002815814, 0.0001915484, 5.980543e-05, 3.46936e-05, 
    2.943991e-05, 1.417764e-05, 4.035003e-05, 6.176193e-06, 1.364703e-05, 
    7.569554e-06, 7.813494e-06, 6.024281e-06, 2.992741e-06, 5.469735e-06,
  0.0001977597, 0.0002386348, 0.000215636, 0.0001177474, 5.506466e-05, 
    2.72777e-05, 2.869529e-05, 2.224351e-05, 5.762604e-05, 3.611837e-05, 
    1.526471e-05, 1.290745e-05, 7.695326e-06, 4.007871e-06, 9.304985e-07,
  3.163624e-07, 1.009827e-07, 1.827634e-07, 7.045588e-07, 5.344648e-07, 
    1.619663e-06, 3.328036e-06, 1.502196e-07, 1.272031e-06, 8.597918e-06, 
    2.380993e-05, 5.43391e-05, 2.649466e-05, 1.529297e-05, 1.995648e-09,
  2.891491e-08, 2.627917e-08, 5.58915e-08, 5.174577e-06, 5.532242e-06, 
    1.792203e-05, 3.54819e-05, 8.795521e-06, 1.059074e-05, 7.695527e-06, 
    1.595503e-05, 1.857923e-05, 4.191654e-05, 4.089325e-05, 1.840888e-06,
  1.627578e-05, 2.669416e-06, 4.258582e-06, 4.506775e-06, 3.027299e-05, 
    2.740549e-05, 2.53841e-05, 2.569462e-05, 1.531583e-05, 1.047386e-05, 
    9.014741e-06, 2.160439e-05, 9.111949e-05, 5.559034e-05, 8.907924e-06,
  0.0001471946, 8.293759e-06, 3.416628e-05, 3.811961e-05, 5.036279e-05, 
    2.300855e-05, 3.023164e-05, 4.880998e-05, 1.382423e-05, 7.121521e-06, 
    2.007903e-05, 4.753988e-06, 3.07963e-05, 4.832985e-05, 2.891633e-05,
  0.0001694104, 9.011106e-06, 1.25595e-06, 1.274931e-05, 1.515043e-05, 
    1.70186e-05, 4.396669e-05, 3.257777e-05, 1.154692e-05, 7.077198e-06, 
    2.863646e-09, 1.941179e-09, 1.694385e-05, 1.716835e-05, 5.625094e-05,
  8.274047e-05, 7.875622e-05, 2.001374e-05, 3.356933e-05, 3.446548e-05, 
    3.660874e-05, 2.253645e-05, 2.94647e-05, 4.245324e-05, 4.673544e-09, 
    5.033934e-07, 1.324911e-06, 1.533013e-07, 3.675676e-06, 1.77841e-05,
  0.0001038449, 0.0001325583, 9.787439e-05, 0.0001011597, 5.929873e-05, 
    3.400267e-05, 4.339791e-05, 5.063502e-05, 6.596041e-05, 2.389087e-06, 
    2.172977e-06, 7.818269e-08, 3.353682e-08, 2.082838e-06, 1.650322e-06,
  0.0002687288, 0.0002657018, 0.0001495063, 0.0001142743, 7.602994e-05, 
    4.329349e-05, 2.271796e-05, 3.309915e-05, 7.126437e-05, 9.935153e-06, 
    2.049861e-06, 2.047273e-07, 4.807013e-08, 1.317405e-05, 7.349269e-08,
  0.0004901194, 0.000407006, 0.0002617395, 0.000159255, 0.0001334102, 
    8.039565e-05, 2.443226e-05, 2.398943e-05, 2.938082e-08, 2.341172e-06, 
    4.943081e-06, 1.804428e-06, 1.210272e-07, 2.138523e-05, 1.955526e-06,
  0.0004332254, 0.0004504085, 0.0004341766, 0.0002629786, 0.0001723845, 
    7.003068e-05, 1.218509e-05, 3.894173e-09, 2.797574e-08, 8.729062e-07, 
    5.233814e-06, 4.646752e-06, 4.631737e-06, 7.345655e-06, 5.190918e-07,
  2.757499e-05, 5.48928e-06, 1.927221e-05, 5.106808e-06, 5.205455e-07, 
    7.031719e-10, 7.334982e-07, 2.093849e-05, 6.321064e-05, 0.0001063297, 
    5.489909e-05, 7.453468e-05, 3.839457e-05, 3.23779e-05, 2.072193e-08,
  2.466006e-06, 9.841345e-06, 3.10478e-05, 1.2007e-05, 1.031253e-06, 
    1.661159e-08, 5.399841e-09, 2.93841e-05, 4.778456e-05, 8.635782e-05, 
    9.407276e-05, 9.778699e-05, 7.556113e-05, 4.348637e-05, 2.844525e-06,
  8.067283e-05, 5.487179e-05, 1.744846e-05, 1.246341e-05, 1.737982e-05, 
    2.477312e-06, 4.925258e-08, 9.749127e-06, 1.692034e-05, 3.401925e-05, 
    8.884314e-05, 6.031581e-05, 0.0001001593, 5.806564e-05, 6.96395e-06,
  0.0001280791, 2.554083e-05, 4.116317e-05, 5.307064e-05, 2.540551e-05, 
    2.35189e-05, 9.541611e-07, 2.294514e-07, 3.651126e-06, 7.712468e-06, 
    3.584502e-05, 8.602452e-05, 7.32341e-05, 6.274966e-05, 4.822334e-05,
  0.0001369936, 2.718427e-05, 3.623723e-05, 4.564173e-05, 4.709919e-05, 
    3.144641e-05, 1.517926e-05, 7.004846e-06, 9.285537e-08, 4.71213e-07, 
    1.575057e-09, 8.975754e-09, 1.709875e-05, 3.94583e-05, 7.679881e-05,
  3.309409e-05, 6.41156e-05, 3.161934e-05, 5.384972e-05, 5.225618e-05, 
    3.8389e-05, 2.72655e-05, 2.455491e-05, 1.106572e-05, 9.120736e-10, 
    1.253043e-07, 2.808869e-06, 6.61906e-08, 9.494414e-06, 2.6316e-05,
  1.8657e-05, 3.769815e-05, 2.820805e-05, 4.111082e-05, 4.779276e-05, 
    3.25677e-05, 3.622884e-05, 2.585256e-05, 1.152064e-05, 1.432338e-09, 
    3.971653e-10, 1.091245e-09, 3.135812e-09, 2.288838e-05, 3.524714e-05,
  2.084632e-05, 4.767679e-05, 2.574785e-05, 2.505594e-05, 2.874204e-05, 
    3.685924e-05, 2.410536e-05, 2.280819e-05, 1.666394e-05, 3.222263e-10, 
    9.862162e-11, 4.473714e-11, 2.950732e-10, 2.524503e-05, 3.236164e-05,
  5.289846e-05, 5.620514e-05, 4.115612e-05, 2.590812e-05, 3.965754e-05, 
    3.491573e-05, 3.3101e-05, 3.361458e-05, 1.471712e-07, 1.547903e-09, 
    3.449747e-10, 1.302845e-10, 1.997741e-10, 3.959219e-06, 2.964605e-05,
  3.626521e-05, 6.286291e-05, 6.177673e-05, 3.432257e-05, 5.227341e-05, 
    6.663516e-05, 3.244221e-05, 6.539697e-06, 4.284282e-06, 7.938965e-08, 
    4.12272e-10, 2.323786e-08, 1.597035e-09, 3.885244e-08, 5.568792e-06,
  1.275991e-05, 4.591331e-06, 2.238859e-05, 1.41984e-05, 1.799199e-06, 
    3.992328e-09, 5.561807e-06, 6.268801e-05, 0.0003501507, 0.0005753088, 
    0.0004174763, 0.0002737852, 0.0002323795, 0.0001122392, 1.22654e-05,
  6.890366e-08, 4.618837e-06, 3.155084e-05, 3.380409e-05, 1.897626e-05, 
    4.710859e-06, 1.878814e-05, 4.247923e-05, 0.0001989839, 0.0003570759, 
    0.0004106783, 0.0003807534, 0.0002643704, 8.870444e-05, 4.759372e-06,
  1.945563e-05, 1.705357e-05, 2.57693e-05, 2.798228e-05, 3.411091e-05, 
    1.026312e-05, 4.358968e-06, 4.315844e-05, 0.0001040605, 0.0001826478, 
    0.00029884, 0.0003680284, 0.0003435066, 0.0001201492, 4.258181e-06,
  3.243236e-05, 8.697564e-06, 2.980893e-05, 3.894596e-05, 3.539339e-05, 
    2.748213e-05, 2.624939e-05, 3.300346e-05, 6.207499e-05, 5.782631e-05, 
    0.0001691909, 0.0002819342, 0.0002607147, 0.0001191546, 1.624473e-05,
  3.798229e-05, 7.336733e-06, 1.54379e-05, 3.121632e-05, 2.885158e-05, 
    3.157904e-05, 4.36907e-05, 3.015707e-05, 2.307816e-05, 2.218699e-05, 
    1.249873e-06, 4.675285e-05, 0.0003080718, 3.797618e-05, 1.91028e-05,
  2.864654e-05, 3.690719e-05, 2.416614e-05, 3.01994e-05, 3.361526e-05, 
    2.91239e-05, 4.772762e-05, 4.386752e-05, 2.368309e-05, 8.257603e-09, 
    7.019838e-09, 3.906224e-06, 0.0002644728, 0.0001163627, 2.248323e-05,
  2.016242e-05, 2.278147e-05, 5.052837e-06, 7.855804e-06, 1.773952e-05, 
    1.944626e-05, 2.75547e-05, 3.578785e-05, 1.832872e-05, 7.273238e-09, 
    4.338708e-09, 8.999004e-07, 8.128994e-05, 0.0001883956, 6.662332e-05,
  1.870844e-05, 4.329437e-05, 1.935844e-05, 3.661166e-06, 7.782427e-06, 
    1.734734e-05, 2.329881e-05, 5.677233e-05, 2.153488e-05, 4.22045e-09, 
    1.590126e-09, 3.27619e-09, 7.863208e-06, 0.0002828824, 0.0001699569,
  4.078592e-05, 5.192424e-05, 6.813709e-05, 4.035448e-05, 4.161841e-05, 
    3.505038e-05, 3.454395e-05, 5.985233e-05, 2.256145e-07, 3.715951e-09, 
    2.290802e-09, 4.329817e-09, 5.711267e-08, 0.0003498871, 0.0004900266,
  4.93033e-05, 9.765453e-05, 6.351422e-05, 6.227893e-05, 6.846731e-05, 
    6.666403e-05, 3.57824e-05, 5.524921e-06, 8.683227e-09, 5.669688e-10, 
    1.010702e-09, 2.014761e-09, 3.58762e-09, 4.698726e-05, 0.000188386,
  2.283473e-05, 1.026442e-05, 7.979862e-05, 2.005094e-05, 3.287675e-05, 
    3.248595e-05, 5.542632e-05, 7.084962e-05, 0.0001656068, 0.0002121373, 
    0.0001733193, 9.162202e-05, 4.115644e-05, 6.078586e-05, 6.155724e-05,
  3.032718e-06, 2.197028e-06, 4.034919e-05, 6.443969e-05, 7.204451e-05, 
    3.928605e-05, 6.583834e-05, 7.021057e-05, 0.0001086558, 0.0001208923, 
    9.837402e-05, 8.213663e-05, 9.692187e-05, 7.792784e-05, 5.945714e-05,
  2.870924e-05, 1.663613e-05, 2.510802e-05, 4.849209e-05, 5.346251e-05, 
    2.557167e-05, 3.674368e-05, 5.827076e-05, 7.374405e-05, 5.562158e-05, 
    4.199138e-05, 9.094027e-05, 0.0001930144, 0.0001871691, 9.13547e-05,
  7.340557e-05, 7.480364e-06, 4.054791e-05, 5.931079e-05, 4.558142e-05, 
    6.701359e-05, 4.165005e-05, 7.92941e-05, 5.487097e-05, 1.024405e-05, 
    3.620191e-05, 0.0001632152, 0.000233084, 0.000247827, 8.197499e-05,
  5.493747e-05, 5.084454e-06, 2.767701e-05, 4.546201e-05, 6.982486e-05, 
    9.728815e-05, 0.0001106816, 7.294868e-05, 4.395572e-05, 3.361733e-05, 
    1.150846e-07, 2.169321e-05, 0.0004233991, 0.0002121786, 7.132591e-05,
  3.614536e-05, 5.228784e-05, 4.785653e-05, 6.014615e-05, 6.949504e-05, 
    7.492951e-05, 8.812156e-05, 7.634233e-05, 3.661221e-05, 3.050857e-08, 
    4.679184e-08, 2.898812e-05, 0.0002975947, 0.0002867792, 6.527454e-05,
  3.777362e-05, 7.564331e-05, 5.181678e-05, 6.089141e-05, 5.684823e-05, 
    8.753136e-05, 8.828771e-05, 4.362876e-05, 1.323016e-05, 1.196787e-08, 
    1.275315e-08, 2.372306e-05, 0.0002408017, 0.0003589848, 8.237143e-05,
  2.584072e-05, 5.009878e-05, 5.977332e-05, 5.647581e-05, 8.721808e-05, 
    0.0001304608, 9.45386e-05, 7.42102e-05, 3.665536e-06, 8.766914e-09, 
    3.853919e-09, 6.502038e-06, 0.0001250978, 0.0003467414, 0.0001318932,
  2.881236e-05, 4.08194e-05, 5.009777e-05, 6.41528e-05, 6.96795e-05, 
    9.618992e-05, 0.0001281851, 0.0001156378, 2.054504e-06, 7.258351e-09, 
    5.983139e-09, 4.828203e-06, 0.0001030693, 0.0005845965, 0.0002989795,
  3.211343e-05, 3.778443e-05, 3.590569e-05, 4.938252e-05, 4.15841e-05, 
    7.806738e-05, 3.057162e-05, 1.816728e-05, 3.888946e-07, 3.686993e-09, 
    2.833207e-09, 1.29715e-06, 0.0001012965, 0.0004142185, 0.0002106258,
  4.168598e-05, 3.793453e-05, 0.000125387, 5.603021e-05, 4.072995e-05, 
    3.849408e-05, 3.963794e-05, 1.923333e-05, 5.704521e-05, 7.397755e-05, 
    6.337938e-05, 8.306297e-05, 2.577927e-05, 7.698766e-05, 0.0001083159,
  4.375614e-06, 1.497347e-05, 6.267218e-05, 8.440844e-05, 3.818818e-05, 
    3.58321e-05, 5.226476e-05, 5.067282e-05, 6.732581e-05, 4.526409e-05, 
    7.915376e-05, 5.139312e-05, 3.878572e-05, 8.110254e-05, 9.564881e-05,
  5.773301e-05, 4.706292e-05, 1.975626e-05, 7.671712e-05, 7.823648e-05, 
    3.775427e-05, 2.060347e-05, 6.290042e-05, 8.417046e-05, 7.688566e-05, 
    4.812614e-05, 5.645964e-05, 5.555452e-05, 7.244819e-05, 9.272213e-05,
  8.246229e-05, 4.583284e-05, 9.503634e-05, 6.063683e-05, 7.198674e-05, 
    5.082834e-05, 5.017607e-05, 0.0001126487, 9.621459e-05, 8.030519e-05, 
    6.552916e-05, 4.958165e-05, 3.81579e-05, 4.410204e-05, 0.0001181547,
  6.901697e-05, 7.671278e-05, 8.224617e-05, 8.027947e-05, 6.348323e-05, 
    9.853274e-05, 0.000158708, 0.0001067933, 0.0001125024, 7.510377e-05, 
    1.95603e-07, 5.952097e-08, 1.016806e-05, 1.671709e-05, 0.0001254372,
  3.805973e-05, 7.236131e-05, 5.218298e-05, 5.898064e-05, 6.507492e-05, 
    5.508156e-05, 0.0001183317, 0.0002061168, 8.812268e-05, 1.113922e-05, 
    1.831914e-05, 2.212123e-06, 4.267697e-07, 1.311285e-05, 2.631648e-05,
  1.412888e-05, 2.970418e-05, 4.182108e-05, 5.981751e-05, 7.343758e-05, 
    6.831103e-05, 0.0001370327, 0.0001744502, 9.096954e-05, 4.919004e-05, 
    9.642236e-06, 8.97248e-07, 6.014461e-06, 7.781162e-05, 4.047015e-05,
  5.747587e-06, 2.717813e-05, 0.0001197324, 0.0001753482, 0.0001076172, 
    0.0001843312, 0.0002942337, 0.0002366857, 9.270174e-05, 2.514108e-05, 
    8.526725e-07, 1.189073e-05, 8.803127e-06, 0.0001029377, 4.358226e-05,
  9.61774e-06, 1.818461e-05, 0.0001485898, 0.000273199, 0.0002031476, 
    0.0002820691, 0.0004140509, 0.0002525618, 6.468692e-07, 1.486448e-06, 
    4.475851e-07, 1.865333e-05, 2.83697e-05, 8.095355e-05, 2.937209e-05,
  6.343463e-06, 3.222227e-06, 9.576454e-05, 0.000267193, 0.0003255271, 
    0.0004258754, 0.0003383472, 2.893042e-05, 2.192768e-07, 1.026377e-07, 
    2.724069e-06, 3.865862e-05, 8.049179e-05, 7.743922e-05, 6.518176e-05,
  1.86459e-06, 7.1186e-06, 2.003542e-05, 2.229338e-05, 1.128154e-05, 
    5.76307e-06, 6.948232e-06, 3.205968e-06, 3.733868e-05, 4.057703e-05, 
    2.260837e-05, 3.079516e-05, 3.904973e-05, 5.928093e-05, 0.0001490145,
  1.751199e-09, 3.617936e-06, 6.320982e-05, 7.638513e-05, 6.207434e-05, 
    2.86271e-05, 2.404572e-05, 9.233127e-06, 3.21516e-05, 2.626424e-05, 
    1.991228e-05, 1.532095e-05, 3.071431e-05, 2.950388e-05, 8.912253e-05,
  2.452997e-05, 2.706438e-05, 0.0001051817, 0.0001400683, 0.0001390162, 
    5.55933e-05, 3.313554e-05, 4.547029e-05, 4.371603e-05, 3.246712e-05, 
    2.63672e-05, 2.423814e-05, 2.281449e-05, 4.161397e-05, 8.45217e-05,
  4.812211e-05, 3.912982e-05, 5.083896e-05, 0.0001242094, 0.0001294847, 
    8.045625e-05, 6.06491e-05, 4.778984e-05, 5.241573e-05, 3.962079e-05, 
    2.141536e-05, 2.152829e-05, 3.523304e-05, 3.884616e-05, 0.0001342024,
  8.032902e-05, 2.053193e-05, 5.210247e-05, 9.697893e-05, 9.60752e-05, 
    9.47044e-05, 4.766804e-05, 4.293132e-05, 6.213457e-05, 3.804403e-05, 
    1.879631e-07, 3.730547e-07, 2.087695e-05, 1.32844e-05, 0.0001376211,
  9.127339e-06, 2.065262e-05, 1.506322e-05, 2.875426e-05, 4.303195e-05, 
    4.548764e-05, 2.848954e-05, 7.611923e-05, 7.316791e-05, 1.131807e-06, 
    1.224279e-06, 1.375857e-07, 8.682239e-07, 1.035977e-05, 0.0001021084,
  6.40451e-06, 1.205844e-05, 5.294865e-06, 6.884819e-06, 1.285567e-05, 
    1.036684e-05, 2.475617e-05, 7.5911e-05, 0.0001000445, 3.667251e-06, 
    5.597871e-07, 1.904946e-07, 6.859166e-07, 2.062178e-05, 8.88162e-05,
  7.135882e-06, 1.293137e-05, 2.384113e-05, 2.727775e-05, 3.436309e-05, 
    6.293547e-05, 0.0001083195, 0.000160207, 0.0001497662, 1.942418e-05, 
    6.246513e-07, 9.402282e-09, 6.370789e-08, 1.481559e-05, 0.0001004065,
  4.46386e-06, 1.068888e-05, 3.373784e-05, 9.997606e-05, 0.0001503598, 
    0.0001621557, 0.0001823208, 0.0002499173, 0.0001256526, 7.338873e-05, 
    7.157437e-08, 4.058275e-08, 7.243188e-08, 3.218586e-05, 8.363739e-05,
  2.761937e-06, 6.956421e-06, 3.854942e-05, 0.0001025297, 0.0001707001, 
    0.0001818822, 0.0001574194, 8.91435e-05, 4.456904e-05, 2.642956e-05, 
    9.751559e-06, 6.856303e-08, 7.464968e-07, 7.173517e-05, 6.248553e-05,
  1.248248e-06, 9.783492e-07, 1.114779e-06, 3.800443e-07, 9.009747e-09, 
    1.146754e-07, 3.527887e-06, 1.022087e-05, 1.751709e-05, 1.987307e-05, 
    2.289865e-05, 3.088613e-05, 6.30778e-05, 6.456092e-05, 4.722569e-06,
  2.53917e-10, 1.539788e-07, 8.965008e-06, 3.039823e-06, 1.065182e-06, 
    3.1186e-06, 5.01215e-07, 2.375083e-06, 1.646981e-05, 1.599743e-05, 
    1.47945e-05, 2.07939e-05, 4.860928e-05, 4.256435e-05, 2.75532e-05,
  8.511603e-06, 2.079766e-05, 2.53765e-05, 2.393935e-05, 2.36634e-05, 
    2.062789e-05, 9.015687e-06, 1.395377e-05, 3.400436e-05, 3.730266e-05, 
    3.119918e-05, 2.504079e-05, 4.59986e-05, 5.560155e-05, 3.768205e-05,
  2.232133e-05, 6.07495e-06, 8.174244e-06, 3.918309e-05, 1.846274e-05, 
    1.384106e-05, 1.834262e-05, 1.675636e-05, 3.808332e-05, 4.276207e-05, 
    3.979209e-05, 2.194812e-05, 4.555563e-05, 6.145194e-05, 7.398504e-05,
  4.40583e-05, 1.281524e-05, 1.927884e-05, 2.338149e-05, 2.722354e-05, 
    4.02502e-05, 4.785989e-05, 5.080382e-05, 3.799746e-05, 6.346263e-05, 
    6.948114e-07, 4.527554e-09, 2.05532e-05, 1.893614e-05, 6.689087e-05,
  5.802057e-05, 5.168427e-05, 3.621431e-05, 4.960568e-05, 6.209358e-05, 
    5.367196e-05, 0.0001026649, 0.000107992, 5.733979e-05, 1.409864e-06, 
    6.260292e-08, 9.866318e-10, 3.972915e-09, 5.882075e-06, 1.614036e-05,
  5.701508e-05, 6.927171e-05, 3.095895e-05, 6.049987e-05, 7.104286e-05, 
    6.530187e-05, 5.147561e-05, 7.753802e-05, 6.785252e-05, 4.226652e-08, 
    2.662221e-08, 2.720845e-10, 2.903789e-10, 2.190529e-05, 5.077407e-05,
  2.039116e-05, 6.575853e-05, 6.555674e-05, 6.179462e-05, 7.611397e-05, 
    7.478673e-05, 6.557041e-05, 8.878091e-05, 9.14589e-05, 9.631804e-06, 
    7.395418e-09, 7.998006e-11, 3.682441e-10, 5.438564e-05, 5.955675e-05,
  1.259321e-05, 6.077466e-05, 4.171841e-05, 5.570557e-05, 8.177327e-05, 
    7.717167e-05, 3.631058e-05, 6.450846e-05, 7.432376e-06, 1.120383e-07, 
    1.758826e-08, 9.70341e-10, 5.126239e-10, 1.583935e-05, 4.379109e-05,
  3.490705e-05, 2.711627e-05, 3.869822e-05, 3.527936e-05, 6.36234e-05, 
    0.0001032906, 4.428738e-05, 1.173284e-06, 4.171035e-07, 1.785588e-05, 
    2.12298e-05, 8.541339e-08, 4.735728e-09, 2.625622e-05, 4.368535e-05,
  2.429769e-06, 1.888705e-09, 1.062348e-05, 8.545901e-06, 4.086388e-06, 
    3.154407e-05, 5.655986e-05, 1.946004e-05, 9.592054e-08, 2.184561e-07, 
    8.278718e-06, 7.888304e-05, 0.0001632216, 0.0001164112, 2.143622e-05,
  1.87614e-06, 2.855563e-09, 2.308079e-05, 1.173151e-05, 2.095359e-05, 
    2.846182e-05, 3.954206e-05, 7.651516e-06, 2.516252e-06, 2.167456e-06, 
    7.483367e-06, 4.165337e-05, 5.496277e-05, 5.734157e-05, 1.421905e-05,
  2.278531e-05, 1.714287e-05, 7.345059e-06, 5.763931e-06, 3.285001e-05, 
    4.140739e-05, 2.136451e-05, 1.528678e-05, 1.38444e-05, 7.897492e-06, 
    1.738173e-05, 4.688418e-05, 0.000112918, 0.0001313297, 5.820487e-05,
  6.63476e-05, 3.130938e-05, 1.849576e-05, 2.772326e-05, 3.430935e-05, 
    3.210722e-05, 3.134192e-05, 2.271032e-05, 2.456197e-05, 2.020812e-05, 
    3.776532e-05, 5.721883e-05, 0.0001171594, 0.0001558715, 0.0001795269,
  3.834032e-05, 8.791559e-05, 6.892327e-05, 4.91824e-05, 3.558548e-05, 
    2.308067e-05, 1.313988e-05, 2.914103e-05, 3.178395e-05, 3.399749e-05, 
    1.7529e-08, 1.991617e-08, 8.282537e-05, 9.881603e-05, 0.0001344354,
  5.552234e-05, 6.803998e-05, 0.0001175752, 9.296287e-05, 7.286976e-05, 
    6.644881e-05, 6.177019e-05, 6.546475e-05, 5.830799e-05, 6.70173e-08, 
    3.185676e-09, 7.46871e-09, 1.458621e-08, 4.790775e-05, 8.201384e-05,
  4.277108e-05, 4.653511e-05, 5.690691e-05, 0.0001046281, 8.249227e-05, 
    0.0001519154, 0.0001199731, 5.713456e-05, 1.583309e-05, 1.391645e-09, 
    2.952292e-10, 1.671249e-10, 2.676134e-09, 6.627804e-05, 6.690821e-05,
  1.124253e-05, 3.723303e-05, 3.010743e-05, 3.56955e-05, 8.253207e-05, 
    0.0001274403, 0.0001288819, 7.353843e-05, 1.334041e-05, 3.665956e-09, 
    5.110908e-10, 3.534496e-11, 9.301193e-10, 9.802107e-05, 5.115441e-05,
  9.899349e-06, 2.895721e-05, 4.071648e-05, 5.114176e-05, 3.689881e-05, 
    0.0001224665, 9.390837e-05, 8.880765e-05, 1.165893e-06, 1.838726e-09, 
    8.555819e-11, 6.60574e-11, 7.832309e-10, 3.37295e-05, 2.509319e-05,
  6.849636e-06, 9.399635e-06, 2.119217e-05, 2.681743e-05, 5.083354e-05, 
    3.159114e-05, 2.732432e-05, 3.312528e-06, 8.666768e-09, 1.901817e-09, 
    2.189906e-10, 5.532757e-10, 6.305915e-10, 2.572456e-05, 6.04981e-06,
  2.655501e-07, 1.836663e-05, 5.194585e-05, 4.559435e-05, 6.457579e-05, 
    0.0001069289, 0.000128461, 0.0001270226, 0.0001538874, 0.0001381412, 
    0.0001428994, 0.000156899, 9.281894e-05, 3.330484e-05, 4.03442e-06,
  5.760975e-09, 1.730593e-07, 7.592351e-05, 6.394844e-05, 5.351177e-05, 
    9.731677e-05, 0.00019269, 0.0001309456, 8.830513e-05, 9.565493e-05, 
    0.0001280277, 0.0001246258, 7.658312e-05, 2.498917e-05, 6.426707e-06,
  3.567348e-05, 6.155974e-05, 2.064996e-05, 1.594027e-05, 4.762438e-05, 
    8.374404e-05, 9.4804e-05, 4.748108e-05, 4.484698e-05, 5.015857e-05, 
    7.66992e-05, 7.602278e-05, 4.815358e-05, 1.827501e-05, 1.634205e-06,
  2.620074e-05, 2.96589e-05, 5.244428e-05, 6.599819e-05, 6.644978e-05, 
    9.038002e-05, 8.166958e-05, 5.703674e-05, 6.238223e-05, 5.639237e-05, 
    5.382699e-05, 7.149379e-05, 2.370293e-05, 4.05693e-06, 3.291169e-06,
  3.068072e-06, 1.297079e-05, 2.265124e-05, 3.575195e-05, 2.717356e-05, 
    1.283534e-05, 1.597383e-05, 1.94431e-05, 6.513613e-05, 0.0002105778, 
    8.384673e-06, 3.115343e-06, 8.701752e-06, 3.706049e-07, 1.419784e-05,
  2.603367e-06, 1.394536e-05, 1.909663e-05, 1.390128e-05, 1.844566e-05, 
    2.040296e-05, 9.96758e-06, 9.548355e-06, 2.043073e-05, 3.339098e-07, 
    2.771499e-08, 6.86389e-08, 4.525356e-06, 2.250578e-07, 2.331816e-05,
  1.039821e-06, 5.083906e-06, 1.082795e-05, 1.973564e-05, 2.175029e-05, 
    3.853354e-06, 2.184614e-06, 8.519681e-07, 7.531848e-06, 7.520489e-09, 
    1.755708e-09, 3.999689e-09, 4.810108e-08, 1.237984e-05, 2.089432e-05,
  4.071321e-08, 3.211365e-06, 3.205493e-06, 4.809252e-06, 1.777895e-05, 
    6.112707e-06, 2.03554e-06, 2.348322e-06, 4.366077e-06, 8.015958e-08, 
    6.750322e-10, 8.711337e-10, 9.508517e-09, 6.775164e-05, 1.186628e-05,
  6.77042e-09, 9.781429e-07, 2.748214e-06, 1.864611e-06, 5.952735e-06, 
    1.165439e-05, 5.260552e-06, 5.815224e-06, 3.073554e-08, 1.211718e-09, 
    4.4681e-10, 6.130094e-10, 1.708476e-09, 9.513368e-05, 3.453764e-05,
  2.853855e-09, 3.558093e-08, 8.844258e-07, 6.774588e-07, 1.686806e-08, 
    2.127624e-09, 1.033172e-07, 5.923374e-07, 2.855044e-09, 1.358007e-09, 
    8.319213e-10, 9.048235e-10, 1.734374e-09, 3.013623e-05, 1.376485e-06,
  4.765661e-10, 2.280153e-06, 1.643201e-05, 2.78042e-05, 8.134792e-05, 
    0.0001117201, 9.929947e-05, 3.302533e-05, 0.0001051775, 0.0001104139, 
    7.223384e-05, 3.221927e-05, 7.700904e-06, 3.980438e-06, 5.192601e-08,
  9.356308e-10, 2.982479e-10, 8.488097e-07, 3.535692e-05, 6.121161e-05, 
    7.295204e-05, 8.223037e-05, 5.974013e-05, 0.0001036911, 0.0001222901, 
    9.77467e-05, 5.493476e-05, 9.178327e-06, 6.790262e-06, 4.983133e-08,
  3.301184e-06, 4.499685e-06, 5.572845e-06, 2.820022e-05, 5.976035e-05, 
    6.334845e-05, 4.895658e-05, 5.296215e-05, 0.0001156602, 0.0001580442, 
    0.0001296374, 7.301831e-05, 2.765388e-05, 3.752958e-05, 5.777348e-06,
  2.003996e-06, 3.229541e-09, 1.462006e-06, 8.020094e-06, 3.419761e-05, 
    2.670311e-05, 6.178061e-05, 4.608459e-05, 8.619761e-05, 9.603595e-05, 
    7.580377e-05, 6.675841e-05, 1.418029e-05, 4.508505e-05, 4.698465e-05,
  6.480947e-06, 5.931593e-06, 6.654471e-08, 9.14345e-08, 9.802027e-07, 
    1.599649e-05, 1.607068e-05, 2.790723e-05, 3.85495e-05, 0.0001416442, 
    4.991868e-06, 1.690154e-06, 9.951353e-07, 2.03916e-06, 3.416758e-05,
  2.410348e-05, 5.761503e-06, 9.424598e-06, 4.339358e-08, 2.69166e-09, 
    2.147738e-06, 1.393221e-05, 1.350567e-05, 1.487151e-05, 6.778214e-08, 
    2.025938e-08, 4.721713e-08, 1.536675e-09, 6.878319e-08, 2.412923e-05,
  1.5161e-05, 4.460244e-05, 1.892594e-05, 9.874225e-06, 8.520554e-08, 
    9.607602e-10, 5.623146e-07, 7.545451e-07, 3.738343e-08, 6.152627e-10, 
    1.347401e-09, 5.598872e-09, 1.996409e-10, 5.02358e-08, 3.721034e-06,
  1.231613e-05, 2.286303e-05, 5.897618e-05, 2.173832e-05, 1.160944e-05, 
    3.815143e-07, 5.589213e-08, 2.664853e-08, 4.957953e-08, 4.057912e-11, 
    1.07402e-10, 7.593602e-10, 1.251743e-08, 2.230567e-05, 7.272832e-07,
  1.021293e-05, 2.083963e-05, 2.800683e-05, 2.927479e-05, 1.141526e-05, 
    1.006758e-05, 4.002205e-06, 2.54287e-08, 1.888383e-10, 3.036832e-10, 
    6.212851e-12, 1.537891e-10, 1.800901e-09, 1.344138e-05, 3.295909e-08,
  9.575564e-08, 1.165994e-06, 3.547323e-05, 2.716655e-05, 1.503078e-05, 
    8.252779e-06, 1.158713e-05, 8.247988e-09, 2.761268e-11, 1.54865e-09, 
    1.38091e-10, 1.358362e-10, 1.057651e-09, 2.86653e-06, 5.371328e-10,
  7.546693e-09, 1.339825e-06, 2.265106e-05, 4.697411e-05, 8.460467e-05, 
    9.847932e-05, 4.912909e-05, 3.384672e-06, 1.414362e-05, 2.213833e-05, 
    4.927007e-05, 4.044025e-05, 4.582596e-05, 2.825919e-05, 2.291158e-05,
  2.264013e-09, 3.826319e-09, 3.5901e-05, 7.355798e-05, 6.874284e-05, 
    8.563029e-05, 6.37574e-05, 1.699987e-05, 1.75424e-05, 2.952904e-05, 
    4.524266e-05, 2.587554e-05, 2.737138e-05, 2.70611e-05, 3.399177e-06,
  2.072968e-05, 5.870137e-05, 5.613939e-05, 7.990012e-05, 9.407566e-05, 
    8.715755e-05, 3.094308e-05, 3.527416e-05, 3.51317e-05, 3.806252e-05, 
    7.333434e-05, 8.47116e-05, 5.097188e-05, 5.518966e-05, 3.793712e-07,
  1.045056e-05, 4.5536e-05, 0.0001259926, 0.0001032516, 3.037853e-05, 
    3.812745e-05, 2.133859e-05, 1.433862e-05, 6.650413e-05, 2.95249e-05, 
    5.57518e-05, 6.448131e-05, 0.0001027372, 5.107008e-05, 1.414877e-05,
  4.12992e-05, 3.926988e-05, 0.0001060986, 0.000138631, 3.1932e-05, 
    4.397972e-06, 3.121776e-05, 2.930776e-05, 2.447666e-05, 4.323634e-05, 
    2.010402e-08, 1.23076e-08, 6.836747e-05, 3.951766e-05, 4.42747e-05,
  7.427607e-05, 0.0001428104, 9.810214e-05, 0.0001484042, 0.0001027758, 
    3.028577e-05, 6.169995e-06, 1.451495e-05, 1.401762e-05, 8.439278e-10, 
    4.889065e-10, 2.754266e-09, 5.869061e-09, 2.467608e-05, 2.396605e-05,
  6.730469e-05, 0.0001458815, 9.570385e-05, 7.597395e-05, 0.000120356, 
    8.124719e-05, 2.387058e-06, 5.110775e-06, 8.534587e-09, 1.790969e-10, 
    1.250432e-10, 3.435211e-10, 2.642305e-10, 4.145253e-05, 3.473265e-05,
  2.943174e-05, 0.0001004178, 9.937616e-05, 7.67243e-05, 6.925708e-05, 
    8.347438e-05, 2.977311e-05, 3.148464e-05, 7.643732e-08, 1.038836e-10, 
    2.800473e-11, 1.938428e-10, 2.913379e-09, 6.385436e-05, 8.380794e-05,
  2.826839e-06, 6.441661e-05, 7.114788e-05, 0.0001451916, 0.0001589094, 
    0.000106199, 3.260093e-05, 2.791686e-05, 8.882439e-09, 5.848435e-10, 
    8.116507e-12, 1.907345e-10, 3.819203e-09, 4.327474e-05, 5.32086e-05,
  3.703399e-06, 2.504929e-05, 8.94045e-05, 0.0001440842, 0.000318711, 
    7.933084e-05, 1.676352e-05, 2.631395e-06, 5.455704e-09, 3.954831e-10, 
    3.451882e-12, 4.050553e-11, 3.227626e-10, 1.222758e-05, 8.77286e-06,
  2.56224e-09, 3.158882e-09, 3.857077e-07, 3.843867e-06, 1.188258e-05, 
    2.899201e-05, 7.122699e-05, 7.309671e-05, 0.0001135274, 7.533342e-05, 
    4.277288e-05, 4.660709e-05, 7.523915e-05, 9.036809e-05, 2.141615e-05,
  3.230061e-09, 2.196118e-09, 4.279854e-06, 1.541351e-05, 1.215586e-05, 
    3.976217e-05, 9.088478e-05, 0.0001101291, 0.0001273335, 5.591859e-05, 
    5.195573e-05, 4.992796e-05, 7.925354e-05, 8.656692e-05, 4.237042e-05,
  6.63335e-06, 8.307557e-06, 5.721282e-06, 3.24288e-05, 8.27098e-05, 
    7.594278e-05, 8.902234e-05, 0.0001261469, 7.163939e-05, 6.789604e-05, 
    3.502399e-05, 7.801242e-05, 5.574373e-05, 8.818421e-05, 3.428701e-05,
  4.705906e-06, 4.46891e-06, 2.685957e-05, 6.305673e-05, 7.781582e-05, 
    0.0001385871, 0.000103941, 0.0001126525, 6.914557e-05, 0.0001027957, 
    8.734928e-05, 4.105845e-05, 6.711084e-05, 3.465902e-05, 3.119184e-05,
  5.108233e-07, 7.901665e-07, 6.294498e-06, 4.032472e-05, 7.319284e-05, 
    0.0001302665, 0.000130851, 0.0001046906, 9.730157e-05, 9.313121e-05, 
    6.448276e-08, 2.284883e-08, 3.18622e-05, 3.364747e-05, 1.089838e-05,
  2.089302e-08, 7.344847e-06, 7.926196e-06, 4.229057e-05, 6.060703e-05, 
    0.0001083313, 0.0001092963, 0.0001255456, 0.0001494474, 1.007187e-06, 
    5.911077e-08, 1.71867e-09, 1.373878e-09, 2.721466e-05, 2.38944e-05,
  2.462983e-05, 2.997576e-05, 5.713835e-05, 7.158683e-05, 6.807268e-05, 
    4.950984e-05, 0.0001266365, 0.0001965616, 3.832019e-05, 2.761529e-07, 
    1.667018e-10, 9.172561e-11, 1.445675e-09, 3.683605e-05, 3.284495e-05,
  2.489835e-05, 4.585621e-05, 8.149339e-05, 7.428385e-05, 6.95203e-05, 
    6.676037e-05, 0.0001719363, 0.0001345848, 2.522889e-05, 1.772147e-09, 
    3.098606e-11, 1.353336e-11, 7.225966e-10, 7.374419e-05, 0.0001461772,
  2.608575e-05, 4.206656e-05, 9.543464e-05, 6.917753e-05, 5.051225e-05, 
    8.053372e-05, 0.000116776, 0.0001503696, 2.165346e-07, 2.672806e-09, 
    3.818109e-11, 6.975234e-10, 9.81017e-10, 6.371213e-05, 0.0001113991,
  2.478455e-05, 4.339113e-05, 8.707199e-05, 2.83128e-05, 1.540751e-05, 
    2.98923e-05, 2.653167e-05, 1.490502e-05, 1.14638e-06, 1.805288e-09, 
    7.536349e-12, 7.19442e-12, 2.815095e-10, 2.188293e-05, 2.449359e-05,
  6.462088e-08, 6.023177e-06, 4.977039e-05, 7.072562e-05, 7.252484e-05, 
    5.65155e-05, 4.065369e-05, 2.448433e-05, 1.844652e-05, 2.957853e-05, 
    2.95747e-05, 2.932028e-05, 3.557354e-05, 6.65308e-05, 6.585848e-05,
  2.647863e-09, 1.32044e-09, 1.144281e-05, 6.060083e-05, 9.373363e-05, 
    7.198834e-05, 8.44298e-05, 3.027071e-05, 4.384745e-05, 3.746933e-05, 
    5.328534e-05, 4.189762e-05, 4.217768e-05, 9.722854e-05, 0.0001151631,
  2.101744e-05, 1.553095e-05, 1.153765e-05, 1.821641e-05, 7.682535e-05, 
    8.270512e-05, 3.802741e-05, 3.566901e-05, 6.942398e-05, 7.118769e-05, 
    9.319849e-05, 5.262072e-05, 9.161602e-05, 8.241463e-05, 0.0001039471,
  4.422309e-05, 1.607196e-05, 3.236788e-05, 3.6208e-05, 3.191761e-05, 
    4.37626e-05, 4.588869e-05, 6.218808e-05, 9.534484e-05, 0.0001049672, 
    9.19097e-05, 7.531552e-05, 0.0001087155, 7.088787e-05, 6.335203e-05,
  1.133602e-05, 8.59828e-06, 1.298213e-05, 2.119218e-05, 1.295727e-05, 
    3.921786e-05, 5.838638e-05, 6.939682e-05, 0.0001101264, 0.0001048975, 
    7.270938e-08, 1.102263e-05, 7.388139e-05, 0.0001419185, 0.0001056797,
  1.089876e-05, 3.752026e-05, 2.769525e-05, 2.136686e-05, 1.543908e-05, 
    2.875955e-05, 5.412938e-05, 9.668227e-05, 7.329134e-05, 1.735193e-07, 
    2.829658e-05, 1.140427e-05, 4.728472e-07, 1.039653e-05, 2.576715e-05,
  2.309984e-05, 5.014971e-05, 5.043318e-05, 9.390088e-05, 6.906855e-05, 
    7.408864e-05, 0.0001264636, 0.0001025885, 2.884689e-05, 2.539729e-05, 
    1.183791e-05, 2.646145e-09, 2.600478e-09, 4.224602e-06, 1.611051e-05,
  2.127375e-05, 6.764371e-05, 8.5568e-05, 6.524069e-05, 9.744715e-05, 
    0.0001590574, 0.0001199647, 0.0001042821, 6.65297e-05, 1.425308e-05, 
    6.460769e-09, 6.425217e-10, 1.66082e-09, 2.904146e-06, 9.63321e-06,
  6.813743e-06, 2.359056e-05, 3.02513e-05, 8.989753e-06, 1.816003e-05, 
    4.080029e-05, 6.751219e-05, 6.98638e-05, 2.876135e-05, 6.592626e-07, 
    6.555115e-09, 4.363791e-10, 8.027918e-10, 1.183452e-05, 1.186264e-05,
  8.420861e-07, 2.339561e-06, 2.309972e-06, 1.069288e-07, 2.236373e-06, 
    1.037093e-06, 6.128786e-06, 4.414219e-06, 1.009872e-05, 9.905003e-09, 
    9.025453e-10, 1.158573e-11, 5.559234e-11, 5.692696e-06, 3.170728e-07,
  1.963466e-10, 7.622092e-10, 2.017037e-05, 3.873538e-05, 5.680725e-05, 
    8.272536e-05, 0.0001138625, 0.0001124647, 9.651965e-05, 4.394343e-05, 
    3.453101e-05, 3.982391e-05, 1.548745e-05, 1.441348e-05, 1.611994e-05,
  6.812e-12, 5.932966e-10, 5.071623e-06, 1.638141e-05, 4.881233e-05, 
    7.451358e-05, 0.0001277504, 0.0001151155, 8.896291e-05, 4.035986e-05, 
    2.631217e-05, 3.221811e-05, 2.103209e-05, 1.712254e-05, 8.892464e-06,
  7.631686e-06, 9.944869e-07, 6.158257e-09, 7.164449e-08, 1.666795e-05, 
    3.547563e-05, 4.478915e-05, 8.006563e-05, 7.423531e-05, 4.483635e-05, 
    4.765399e-05, 4.258991e-05, 4.237099e-05, 3.529668e-05, 7.360197e-06,
  7.33429e-07, 4.823853e-06, 3.833389e-06, 1.992501e-06, 1.03113e-05, 
    2.689976e-05, 6.619257e-05, 8.228596e-05, 6.608223e-05, 5.985622e-05, 
    6.48203e-05, 5.117041e-05, 4.590129e-05, 3.989312e-05, 9.855308e-06,
  3.56415e-06, 9.125654e-06, 4.008958e-06, 2.833104e-06, 8.302434e-07, 
    1.138402e-05, 5.14843e-05, 7.263081e-05, 8.683444e-05, 8.94464e-05, 
    7.667469e-09, 1.541143e-08, 1.188738e-05, 1.268841e-05, 1.64493e-05,
  9.412572e-07, 8.013387e-06, 1.237408e-05, 7.555494e-06, 4.070849e-06, 
    5.731793e-06, 2.353491e-05, 3.747517e-05, 7.224937e-05, 6.315262e-09, 
    4.324686e-08, 7.615297e-09, 5.446855e-10, 6.380789e-06, 2.489246e-05,
  5.635226e-08, 1.010695e-06, 2.230551e-06, 1.004318e-05, 1.860174e-05, 
    2.096691e-05, 3.19122e-05, 3.293742e-05, 1.440631e-05, 1.46001e-08, 
    3.487693e-09, 1.618738e-10, 2.707398e-10, 1.114601e-05, 4.059028e-05,
  1.682272e-07, 2.438893e-07, 2.40848e-07, 3.566638e-06, 1.906984e-06, 
    2.271237e-05, 5.089196e-05, 8.380727e-05, 2.586121e-05, 1.824045e-08, 
    3.454074e-10, 3.566458e-10, 9.23504e-10, 4.770951e-05, 3.830922e-05,
  1.89289e-07, 1.346135e-07, 1.346827e-07, 6.519299e-09, 2.380253e-07, 
    1.108805e-06, 2.444735e-05, 7.213731e-05, 1.292009e-08, 1.769321e-07, 
    6.69423e-10, 2.972231e-10, 4.263881e-10, 7.990918e-06, 1.163664e-05,
  8.252248e-08, 1.132589e-07, 6.487376e-08, 1.720206e-08, 1.539128e-09, 
    1.562971e-09, 9.751986e-07, 1.433457e-07, 6.671776e-09, 1.16777e-09, 
    4.038459e-10, 3.612028e-10, 1.631466e-10, 2.051265e-08, 1.966437e-09,
  1.391447e-09, 3.423825e-10, 2.274349e-10, 8.291865e-09, 6.454948e-06, 
    3.846123e-05, 3.300021e-05, 2.896928e-05, 4.158099e-05, 2.507706e-05, 
    4.405038e-05, 7.944302e-05, 0.0001149876, 0.0001009065, 0.0001135299,
  1.264464e-09, 1.455167e-10, 8.255215e-09, 1.306761e-08, 3.966582e-08, 
    1.615238e-05, 4.605452e-05, 5.288007e-05, 6.292082e-05, 4.495048e-05, 
    3.919098e-05, 6.140223e-05, 0.0001208825, 9.015761e-05, 9.058322e-05,
  2.092374e-06, 2.825384e-06, 2.229693e-06, 4.005937e-09, 2.376682e-09, 
    5.825581e-07, 5.46415e-06, 5.601931e-05, 6.659922e-05, 2.820831e-05, 
    7.033833e-05, 6.642681e-05, 7.345473e-05, 6.214056e-05, 4.804511e-05,
  1.707747e-05, 1.671673e-05, 2.440226e-05, 1.825473e-05, 2.434672e-06, 
    1.06982e-07, 9.217089e-07, 1.481315e-05, 4.845682e-05, 7.414154e-05, 
    0.0001104711, 7.325302e-05, 8.293357e-05, 5.982421e-05, 4.007214e-05,
  1.72729e-05, 6.377177e-06, 1.809943e-05, 1.759522e-05, 1.825137e-06, 
    2.077228e-07, 4.774816e-07, 5.294953e-06, 2.583816e-05, 4.401457e-05, 
    2.378597e-08, 5.37282e-08, 3.69929e-05, 5.161521e-05, 6.619738e-05,
  2.276424e-06, 2.485695e-05, 2.080542e-05, 3.032913e-05, 2.128494e-05, 
    1.34432e-06, 4.667201e-07, 1.980624e-06, 2.752371e-06, 6.146854e-10, 
    7.373356e-09, 6.726393e-09, 3.80955e-09, 1.774603e-06, 7.490947e-05,
  5.498278e-08, 2.226895e-05, 2.439635e-05, 5.466183e-05, 5.418675e-05, 
    2.519155e-05, 3.088765e-06, 3.51171e-07, 2.728064e-06, 9.855902e-10, 
    1.448791e-09, 8.543644e-10, 1.373253e-09, 1.506846e-05, 5.763028e-05,
  1.067673e-07, 6.575893e-06, 3.75393e-05, 6.177629e-05, 7.223434e-05, 
    7.937873e-05, 2.316276e-05, 1.331037e-06, 1.078415e-06, 7.222111e-10, 
    1.17977e-09, 4.777008e-10, 1.090911e-09, 1.493891e-05, 4.217476e-05,
  1.750043e-07, 1.508405e-05, 2.390616e-05, 3.785199e-05, 7.915492e-05, 
    0.0001096249, 6.800691e-05, 3.489292e-05, 4.690521e-10, 6.091441e-10, 
    4.831501e-10, 2.288441e-10, 3.78853e-10, 6.73899e-06, 1.160103e-05,
  1.518392e-06, 5.773174e-06, 5.329995e-06, 1.413496e-05, 3.874595e-05, 
    7.249061e-05, 5.632718e-05, 3.924272e-06, 5.501703e-07, 1.187113e-10, 
    2.371148e-10, 1.84352e-11, 1.234771e-11, 3.805964e-07, 1.000518e-06,
  2.455569e-09, 2.070613e-09, 6.992028e-09, 3.101525e-08, 2.147909e-07, 
    7.683242e-07, 4.405994e-07, 1.359521e-07, 4.627766e-07, 3.393608e-06, 
    5.184629e-06, 1.611665e-05, 1.154062e-05, 2.349922e-05, 4.395814e-05,
  5.476398e-10, 8.90697e-10, 1.577087e-08, 6.931666e-08, 1.995185e-06, 
    6.297563e-06, 3.116056e-06, 1.188453e-06, 4.21339e-06, 3.902923e-06, 
    6.158269e-06, 2.987284e-06, 5.68561e-06, 2.302362e-05, 6.590345e-05,
  1.980864e-09, 4.497856e-07, 2.528522e-08, 5.44616e-08, 4.369344e-06, 
    1.002356e-05, 2.923312e-06, 2.723192e-06, 6.317539e-06, 6.675432e-06, 
    9.29441e-06, 4.717665e-06, 1.922281e-05, 2.397224e-05, 5.338459e-05,
  8.035238e-06, 7.289806e-07, 8.33676e-06, 2.515518e-05, 1.280629e-05, 
    2.06216e-05, 2.247542e-05, 1.302645e-05, 1.961202e-05, 1.37823e-05, 
    1.714467e-05, 2.874658e-05, 3.76086e-05, 4.029976e-05, 6.954592e-05,
  3.669858e-06, 3.545049e-06, 1.175001e-05, 1.059666e-05, 9.400772e-06, 
    1.80377e-05, 2.62831e-05, 3.073605e-05, 1.826727e-05, 2.452617e-05, 
    3.206501e-09, 2.040567e-09, 3.338332e-06, 1.373926e-05, 4.443333e-05,
  1.015775e-05, 2.851107e-05, 4.537664e-05, 7.684743e-05, 5.731824e-05, 
    4.850736e-05, 4.633157e-05, 5.896272e-05, 4.761825e-05, 2.220756e-10, 
    1.611796e-09, 1.684903e-09, 1.139465e-09, 2.274566e-07, 2.612917e-05,
  6.342888e-06, 3.207459e-05, 7.518185e-05, 9.776085e-05, 0.0001098622, 
    0.0001263249, 8.768843e-05, 6.567479e-05, 2.713071e-05, 2.196099e-10, 
    1.317241e-09, 1.100982e-09, 1.011547e-09, 5.65425e-08, 6.320373e-06,
  1.775754e-05, 1.316504e-05, 3.962931e-05, 7.86177e-05, 0.0001435927, 
    0.0001699993, 0.0001623195, 0.0001163555, 5.460323e-05, 1.421226e-09, 
    1.323201e-09, 1.08365e-09, 5.047276e-10, 6.334453e-09, 8.136729e-06,
  2.103651e-05, 5.919117e-06, 1.556733e-05, 6.517996e-05, 0.0001437155, 
    0.0001381126, 0.0002887129, 0.0002685459, 1.604399e-08, 2.412989e-08, 
    2.299808e-09, 9.396715e-10, 7.119541e-10, 4.498039e-08, 2.70966e-07,
  6.592118e-05, 2.748935e-05, 1.015222e-05, 2.14977e-05, 0.0001076066, 
    0.0001213593, 0.0001614359, 0.0002362481, 0.0001377816, 5.058936e-06, 
    8.185822e-09, 2.303191e-09, 1.222266e-09, 2.451433e-09, 1.856798e-08,
  3.983935e-09, 4.315915e-10, 1.328648e-07, 2.972561e-08, 2.989149e-09, 
    2.718694e-08, 5.49525e-08, 6.22265e-08, 5.147955e-08, 6.969408e-08, 
    1.841621e-06, 4.903711e-06, 1.860761e-05, 3.666874e-05, 3.689212e-06,
  3.578343e-06, 5.062197e-09, 6.516827e-06, 2.532686e-06, 4.049403e-08, 
    6.753814e-09, 1.137286e-08, 3.465671e-08, 4.229831e-08, 3.630777e-08, 
    8.064452e-07, 1.488475e-06, 3.686778e-06, 1.870177e-05, 2.213129e-06,
  0.000113934, 8.09848e-05, 1.487582e-05, 9.223203e-06, 1.158782e-05, 
    4.561966e-06, 8.431874e-08, 4.664363e-08, 3.230058e-08, 1.811886e-08, 
    8.998249e-08, 2.26723e-06, 8.667263e-06, 9.45819e-06, 8.937412e-07,
  0.0001789005, 2.476539e-05, 5.578064e-05, 5.385076e-05, 2.404789e-05, 
    1.264408e-05, 1.010177e-05, 7.367121e-06, 5.0973e-06, 2.483785e-08, 
    9.105555e-08, 2.562962e-06, 1.965858e-05, 1.39377e-05, 1.32966e-05,
  0.0002058946, 4.423958e-05, 2.511416e-05, 5.783288e-05, 3.703886e-05, 
    2.734143e-05, 1.484104e-05, 1.64728e-05, 1.621555e-05, 3.698755e-06, 
    4.581669e-09, 1.143781e-09, 5.850174e-06, 1.146608e-06, 2.936777e-05,
  0.0001286424, 7.186491e-05, 4.082702e-05, 7.002655e-05, 7.252984e-05, 
    3.891498e-05, 1.779542e-05, 1.335274e-05, 1.205926e-05, 2.9852e-10, 
    2.173069e-07, 5.082479e-08, 2.020269e-10, 3.701404e-07, 2.211559e-05,
  0.0001463796, 0.0001041009, 4.477886e-05, 5.334864e-05, 4.701426e-05, 
    6.394889e-05, 3.918557e-05, 2.386566e-05, 6.28814e-06, 8.984531e-10, 
    3.450556e-08, 1.506895e-08, 8.782404e-10, 1.847282e-06, 1.040781e-05,
  0.0002006774, 0.0002710466, 0.0001363297, 7.936213e-05, 6.380224e-05, 
    6.368548e-05, 6.472582e-05, 6.972447e-05, 4.247336e-05, 7.671667e-08, 
    4.064979e-07, 8.043537e-07, 8.327109e-09, 1.102806e-05, 9.505169e-07,
  0.00022794, 0.000144242, 0.0001094573, 6.917767e-05, 5.852782e-05, 
    8.973281e-05, 9.646195e-05, 0.0001081766, 4.907352e-06, 4.957198e-06, 
    1.297386e-06, 4.913829e-07, 3.239659e-07, 9.258476e-06, 5.050972e-07,
  0.0001707622, 0.0001620093, 9.280356e-05, 6.814372e-05, 6.533716e-05, 
    6.679428e-05, 8.521262e-05, 8.105121e-05, 9.796026e-05, 1.298417e-05, 
    2.179139e-06, 5.334847e-07, 1.023008e-06, 2.163299e-05, 3.949202e-06,
  1.27727e-05, 2.212364e-07, 7.052549e-06, 3.580031e-06, 1.675887e-06, 
    1.510805e-06, 2.564803e-06, 2.817928e-07, 2.454373e-06, 5.214563e-06, 
    3.434116e-06, 1.09676e-06, 1.595239e-06, 9.729078e-06, 3.597083e-09,
  1.219881e-06, 7.730628e-08, 1.977685e-05, 1.708646e-05, 4.025929e-06, 
    5.019032e-06, 2.122433e-06, 1.992613e-06, 4.83685e-06, 4.815607e-06, 
    2.025221e-06, 2.94449e-06, 2.244635e-06, 1.454496e-05, 3.653051e-09,
  6.81241e-05, 5.874838e-05, 3.024432e-05, 3.222253e-05, 4.851455e-05, 
    2.231321e-05, 7.094917e-06, 6.270136e-06, 1.284771e-05, 5.551941e-06, 
    8.413864e-06, 8.254525e-06, 1.387273e-05, 1.31698e-05, 1.71841e-08,
  9.624912e-05, 2.709775e-05, 4.489881e-05, 7.155127e-05, 5.790088e-05, 
    3.309591e-05, 4.756723e-05, 2.931747e-05, 3.529742e-05, 2.127132e-05, 
    1.753947e-05, 1.594744e-05, 2.866719e-05, 3.587435e-05, 9.987552e-06,
  0.0001199347, 2.282189e-05, 2.94799e-05, 4.530543e-05, 4.648935e-05, 
    4.49713e-05, 5.568933e-05, 5.299475e-05, 3.521601e-05, 3.359685e-05, 
    3.583797e-09, 2.015074e-09, 1.015136e-05, 2.037326e-06, 6.362569e-06,
  4.766346e-05, 7.860074e-05, 4.791178e-05, 6.50158e-05, 6.771117e-05, 
    4.477712e-05, 4.561124e-05, 5.110235e-05, 6.167532e-05, 5.178649e-06, 
    1.483552e-06, 2.333825e-07, 9.707367e-09, 2.191514e-07, 1.29578e-05,
  4.548253e-05, 7.704039e-05, 8.087381e-05, 7.645959e-05, 0.0001111455, 
    0.0001071054, 0.0001203129, 7.530895e-05, 9.876255e-05, 8.18247e-06, 
    6.478742e-08, 6.741408e-08, 7.008069e-09, 4.467833e-05, 4.481178e-05,
  8.862195e-05, 0.0001140955, 0.0001312168, 0.0002356293, 0.0002820762, 
    0.0002594815, 0.0002722181, 0.000233145, 0.0001695029, 1.288128e-05, 
    1.183465e-06, 2.146739e-06, 5.651575e-09, 0.0001551729, 3.542356e-05,
  6.821426e-05, 9.978915e-05, 0.0001173193, 0.0002704782, 0.0003258206, 
    0.0002577285, 0.0002298205, 0.0002207865, 3.13332e-05, 2.507568e-06, 
    7.494057e-07, 4.563098e-06, 1.437724e-06, 0.0001354733, 7.397845e-05,
  0.0001115187, 0.0001260116, 0.0001738722, 0.0001898175, 0.0001953198, 
    0.0001169784, 7.33199e-05, 7.053446e-06, 1.401024e-06, 2.267754e-06, 
    2.08645e-06, 2.22512e-06, 2.810876e-06, 8.066009e-05, 0.0001087681,
  4.069883e-06, 7.686271e-06, 2.684748e-05, 2.244104e-05, 3.778204e-06, 
    8.230524e-08, 2.727804e-06, 1.076822e-05, 1.995132e-05, 3.041947e-05, 
    0.0001127303, 0.0002033257, 0.0002281171, 0.0002225487, 0.0001335148,
  5.252407e-11, 1.245117e-09, 4.929449e-05, 4.49472e-05, 2.125741e-05, 
    1.104593e-05, 3.55649e-06, 1.42613e-05, 4.025577e-05, 5.840639e-05, 
    0.0001178414, 0.0001330163, 0.0001898053, 0.0001617508, 0.0002219969,
  4.594411e-06, 7.438099e-06, 1.275538e-05, 2.475293e-05, 2.405568e-05, 
    4.030415e-05, 9.062461e-06, 1.737229e-05, 5.39515e-05, 7.548447e-05, 
    0.0001485108, 0.0002060467, 0.0001238074, 8.510028e-05, 8.48909e-05,
  1.945655e-06, 9.518178e-06, 2.221719e-05, 3.735705e-05, 1.719074e-05, 
    3.941286e-05, 5.712434e-05, 3.665235e-05, 5.045743e-05, 9.864776e-05, 
    0.0003086454, 0.0003535168, 0.0001806129, 7.914157e-05, 1.63544e-05,
  1.582619e-06, 5.701973e-06, 1.449412e-05, 3.22802e-05, 3.180526e-05, 
    6.964971e-05, 4.350532e-05, 4.935711e-05, 7.353729e-05, 0.0002040064, 
    7.106087e-05, 8.812228e-05, 0.0002737844, 0.0001381718, 6.872986e-05,
  3.174603e-07, 6.873533e-06, 8.202104e-06, 1.119177e-05, 2.982687e-05, 
    7.565879e-05, 9.202954e-05, 9.566679e-05, 0.0001541075, 0.000115532, 
    0.0001126046, 3.322979e-05, 2.098797e-05, 5.448141e-05, 9.985156e-05,
  2.240969e-06, 5.592378e-06, 6.338516e-06, 5.548532e-06, 1.834748e-05, 
    7.455752e-05, 0.0001569974, 0.000196475, 0.0001972904, 0.0001304041, 
    6.162488e-05, 3.393473e-05, 8.856078e-06, 7.678827e-05, 7.962488e-05,
  1.462877e-07, 3.904782e-06, 7.047698e-06, 2.501054e-06, 2.717554e-06, 
    1.508272e-05, 5.374444e-05, 8.546097e-05, 0.0001266828, 4.760557e-05, 
    2.807545e-05, 2.275422e-05, 9.813725e-06, 0.0001269124, 0.0001052761,
  1.071934e-07, 1.650933e-06, 5.847614e-06, 5.62369e-06, 7.603382e-06, 
    1.242676e-05, 1.806938e-05, 5.144836e-05, 1.027766e-05, 2.676764e-06, 
    4.108186e-06, 3.39751e-06, 1.377631e-06, 3.044339e-05, 2.903408e-05,
  2.410634e-08, 2.322573e-07, 2.633455e-06, 2.251406e-06, 2.997727e-06, 
    1.053797e-05, 2.539154e-05, 1.335552e-05, 5.129229e-06, 5.921755e-06, 
    6.438674e-06, 6.977141e-06, 5.472457e-06, 1.76037e-05, 1.267434e-05,
  3.42148e-10, 2.630707e-08, 5.074775e-06, 1.706196e-08, 1.239189e-10, 
    4.589214e-09, 2.567928e-08, 1.432644e-07, 8.98067e-06, 6.062321e-05, 
    8.864115e-05, 4.375606e-05, 5.548522e-05, 2.002376e-05, 3.804459e-05,
  2.658667e-10, 7.414225e-10, 1.901785e-07, 2.456841e-07, 1.122435e-10, 
    2.846571e-10, 2.57069e-10, 1.883945e-08, 7.174604e-06, 3.745304e-05, 
    5.227117e-05, 7.631821e-05, 5.2772e-05, 1.005501e-05, 7.166964e-05,
  3.364801e-08, 4.608986e-06, 1.931559e-07, 2.06331e-08, 3.131968e-09, 
    4.134391e-10, 7.299081e-10, 9.44374e-10, 2.349617e-07, 4.119066e-06, 
    1.175278e-05, 2.868391e-05, 8.794463e-06, 7.814398e-06, 2.999536e-05,
  5.571938e-06, 2.126589e-06, 1.888567e-06, 2.067065e-07, 7.320278e-09, 
    6.665035e-08, 6.542514e-08, 1.553353e-08, 6.249314e-08, 1.76816e-06, 
    8.002963e-06, 2.568986e-05, 8.473636e-06, 1.865344e-05, 2.283937e-06,
  5.924164e-06, 2.129174e-06, 1.389143e-06, 2.00014e-06, 6.74073e-08, 
    3.352933e-08, 5.690687e-08, 2.802356e-08, 5.965816e-08, 4.267566e-07, 
    1.665056e-07, 2.386713e-06, 3.367479e-05, 2.381243e-05, 1.262644e-05,
  6.012397e-06, 1.056558e-05, 7.245774e-06, 7.417572e-06, 1.002294e-05, 
    5.849525e-07, 9.95818e-08, 4.206516e-08, 2.901207e-08, 6.841741e-10, 
    6.238379e-07, 8.48733e-07, 2.293941e-06, 2.044766e-05, 1.110363e-05,
  2.254446e-06, 3.904897e-06, 7.94789e-06, 2.131411e-05, 8.812574e-06, 
    5.523403e-06, 2.29253e-06, 1.496629e-08, 2.381666e-09, 6.829627e-10, 
    7.768743e-11, 5.093611e-08, 6.216648e-08, 1.916333e-05, 7.28506e-06,
  4.690459e-07, 4.969176e-06, 6.80531e-06, 1.313653e-05, 1.895024e-05, 
    1.352094e-05, 9.376418e-06, 2.597892e-06, 2.898031e-07, 1.526525e-08, 
    1.071942e-10, 5.583691e-08, 4.975565e-09, 3.823233e-06, 2.847044e-07,
  5.312643e-09, 2.920149e-06, 1.01329e-05, 1.653681e-05, 2.3886e-05, 
    2.712146e-05, 2.433377e-05, 8.394274e-06, 5.397034e-07, 4.477388e-08, 
    1.552922e-10, 5.276156e-11, 4.541735e-10, 2.279429e-07, 9.853537e-08,
  2.304867e-09, 1.025705e-06, 7.528827e-07, 5.254128e-06, 7.732968e-06, 
    7.813996e-06, 5.038486e-06, 4.95943e-06, 9.202379e-06, 2.761235e-06, 
    3.703631e-09, 2.531488e-10, 2.718223e-10, 4.185721e-08, 2.311985e-07,
  1.474495e-08, 7.062823e-10, 1.214536e-07, 3.73901e-08, 5.466985e-09, 
    4.342602e-09, 4.220151e-08, 2.513999e-09, 3.88559e-06, 5.694023e-06, 
    2.913841e-06, 1.525893e-05, 3.561222e-05, 5.800033e-05, 6.898292e-05,
  7.225304e-09, 8.361821e-10, 2.535342e-07, 3.461591e-06, 3.463225e-06, 
    9.389344e-06, 7.281005e-06, 1.629099e-05, 4.016278e-05, 3.466381e-05, 
    2.662944e-05, 2.993438e-05, 4.090583e-05, 4.889726e-05, 3.187199e-05,
  1.064632e-08, 7.061775e-10, 8.831537e-10, 2.677437e-08, 8.041149e-06, 
    1.884891e-05, 2.283239e-05, 4.482896e-05, 8.418602e-05, 7.812343e-05, 
    0.0001027016, 9.684481e-05, 7.393828e-05, 4.401116e-05, 2.56086e-05,
  1.257029e-08, 1.056412e-09, 6.545884e-09, 5.753487e-08, 2.11103e-07, 
    5.792025e-06, 1.427713e-05, 3.766819e-05, 7.714239e-05, 0.0001189085, 
    0.0001885312, 0.0001674088, 0.0001050262, 4.433459e-05, 2.638237e-05,
  1.739748e-08, 2.987589e-09, 3.062416e-10, 5.346139e-10, 7.715085e-09, 
    3.547395e-07, 3.302372e-06, 1.811837e-05, 5.493061e-05, 0.0001280529, 
    2.107915e-08, 2.682471e-07, 2.498685e-05, 5.046109e-06, 2.696072e-06,
  2.818099e-08, 4.895222e-09, 4.487768e-10, 9.560714e-10, 7.158733e-07, 
    1.811398e-06, 1.044735e-05, 3.963681e-05, 6.796471e-05, 2.604366e-09, 
    5.420804e-09, 1.510187e-08, 6.398893e-09, 2.409627e-06, 1.193999e-07,
  3.229606e-08, 3.920752e-09, 4.518667e-10, 1.110705e-08, 1.595e-06, 
    2.639462e-06, 1.779096e-05, 4.925095e-05, 6.586926e-05, 3.510605e-09, 
    9.079709e-09, 7.939221e-09, 3.971186e-09, 3.456878e-05, 2.7436e-05,
  2.624127e-08, 5.139102e-08, 3.405769e-07, 1.104945e-06, 1.081481e-06, 
    1.348838e-05, 3.463104e-05, 7.061559e-05, 8.509629e-05, 1.675633e-07, 
    5.712791e-07, 3.714282e-07, 2.262347e-08, 1.841121e-05, 1.8133e-05,
  2.419152e-08, 7.852763e-07, 1.625724e-06, 4.605889e-06, 9.9926e-06, 
    1.968935e-05, 2.863704e-05, 7.12995e-05, 1.653457e-06, 9.760352e-06, 
    8.936984e-06, 7.866566e-06, 4.517526e-06, 1.358262e-05, 8.719368e-06,
  9.778664e-08, 5.222017e-07, 2.347413e-06, 1.778647e-06, 7.561016e-06, 
    8.689338e-06, 7.331603e-06, 7.74162e-08, 3.262531e-06, 1.558437e-05, 
    1.62321e-05, 1.43456e-05, 1.066977e-05, 8.451787e-06, 8.159582e-06,
  3.018147e-07, 8.097534e-08, 5.219933e-08, 3.866038e-08, 2.404889e-08, 
    1.125792e-08, 4.167074e-09, 6.152716e-09, 7.46464e-09, 2.05459e-06, 
    5.974042e-06, 2.263402e-05, 7.387954e-05, 0.0001034884, 2.091442e-05,
  1.846141e-07, 1.60651e-08, 2.142328e-08, 2.078325e-08, 1.217925e-08, 
    4.892816e-09, 1.088398e-08, 1.427963e-08, 4.536022e-07, 1.554433e-06, 
    3.818047e-06, 2.455966e-05, 7.064139e-05, 6.868879e-05, 8.729377e-05,
  9.315464e-08, 2.354439e-08, 3.884868e-09, 1.414481e-08, 4.435688e-07, 
    3.488569e-08, 1.444135e-08, 8.77654e-09, 2.625118e-06, 7.121403e-06, 
    1.650279e-05, 6.642901e-05, 6.211206e-05, 0.0001031768, 0.0001279489,
  2.930415e-07, 2.013763e-07, 2.726804e-06, 1.62723e-06, 2.474782e-07, 
    3.137123e-07, 2.417778e-06, 1.013077e-06, 4.606017e-06, 1.282229e-05, 
    4.99653e-05, 6.765841e-05, 8.363418e-05, 8.854543e-05, 1.610938e-05,
  2.273405e-06, 6.360911e-08, 4.035454e-08, 1.707038e-06, 3.303043e-08, 
    3.055051e-07, 5.604753e-07, 2.832878e-06, 8.62398e-06, 1.611226e-05, 
    8.448824e-07, 1.658051e-07, 2.292512e-05, 1.642693e-05, 1.948219e-05,
  4.306691e-06, 2.390364e-06, 6.90434e-08, 7.101147e-06, 6.468517e-06, 
    7.4934e-08, 8.116942e-07, 4.447159e-07, 9.987251e-06, 6.335825e-07, 
    2.230768e-08, 1.1795e-08, 7.256159e-09, 8.478525e-06, 5.023196e-05,
  5.16716e-06, 9.487757e-06, 4.310634e-06, 9.645987e-06, 3.896777e-06, 
    7.622044e-08, 1.510209e-08, 2.340399e-07, 1.52453e-08, 5.283785e-10, 
    1.740938e-09, 1.110008e-09, 2.206842e-10, 2.659844e-05, 4.669164e-05,
  5.179725e-06, 1.60747e-05, 6.988997e-06, 7.829252e-06, 1.233524e-05, 
    6.406269e-06, 1.022941e-06, 1.951532e-06, 1.134612e-08, 4.543456e-10, 
    2.126326e-09, 2.693872e-09, 9.834198e-10, 2.468508e-05, 2.091869e-05,
  3.071686e-06, 1.325239e-05, 1.438956e-05, 1.480933e-05, 5.275471e-06, 
    2.561664e-05, 1.905067e-05, 2.657346e-05, 4.699087e-09, 1.357772e-09, 
    9.692014e-09, 3.250527e-09, 1.15716e-09, 1.155341e-05, 6.508295e-06,
  1.061173e-06, 1.614971e-06, 4.190169e-06, 2.175318e-06, 1.949487e-06, 
    8.591335e-07, 1.215967e-05, 3.528826e-06, 3.114626e-07, 1.834565e-08, 
    2.864278e-09, 1.755063e-09, 1.170402e-09, 1.064141e-05, 6.208952e-06,
  4.696128e-09, 6.721645e-09, 1.8736e-08, 2.107922e-08, 1.932736e-08, 
    1.928382e-08, 1.649075e-07, 3.205243e-07, 5.579413e-06, 2.128679e-05, 
    2.451997e-05, 3.389309e-05, 6.608019e-05, 4.864841e-05, 8.79202e-05,
  7.782253e-09, 8.804207e-09, 2.497866e-08, 1.979488e-08, 4.771649e-08, 
    3.595083e-06, 8.30702e-06, 9.491542e-06, 3.170624e-05, 3.117471e-05, 
    4.156799e-05, 3.844957e-05, 5.303674e-05, 8.467022e-05, 5.660327e-05,
  1.42024e-08, 2.5507e-08, 1.874391e-08, 2.561851e-08, 3.864267e-06, 
    1.090312e-05, 1.852715e-05, 3.602214e-05, 7.778978e-05, 6.41744e-05, 
    5.434835e-05, 5.430124e-05, 9.27898e-05, 9.380114e-05, 2.544749e-05,
  3.72232e-08, 1.319834e-07, 1.210011e-06, 1.249637e-05, 1.58667e-05, 
    2.553519e-05, 2.135099e-05, 3.13497e-05, 5.990144e-05, 0.0001011179, 
    7.956832e-05, 6.775036e-05, 9.507698e-05, 6.245058e-05, 3.143004e-05,
  7.672051e-08, 1.033518e-07, 1.019278e-07, 8.088358e-08, 1.351642e-06, 
    1.265045e-05, 1.668147e-05, 2.951457e-05, 5.004222e-05, 6.258155e-05, 
    5.195077e-06, 3.568339e-08, 1.957398e-05, 1.893448e-05, 3.874025e-05,
  4.322294e-08, 6.694621e-08, 5.843402e-08, 7.996659e-08, 1.884886e-06, 
    1.096063e-05, 1.499284e-05, 1.003748e-05, 4.242879e-05, 8.080141e-09, 
    1.55777e-08, 5.851296e-08, 4.464471e-08, 5.432696e-08, 6.76703e-06,
  2.43739e-08, 1.100976e-06, 1.801591e-07, 3.949471e-06, 8.534244e-06, 
    1.422026e-05, 2.141668e-05, 1.92227e-05, 1.432547e-05, 2.937919e-09, 
    1.563334e-08, 1.018602e-07, 2.21802e-07, 1.434277e-07, 1.610004e-06,
  1.858695e-08, 1.407421e-06, 9.979882e-07, 3.492079e-07, 5.581826e-06, 
    1.758696e-05, 3.194125e-05, 4.456911e-05, 2.804311e-05, 1.083376e-09, 
    7.940771e-09, 1.234321e-07, 2.944342e-07, 1.744171e-07, 2.138958e-05,
  1.2374e-08, 5.923092e-06, 5.065908e-06, 7.449406e-06, 2.393067e-05, 
    4.942725e-05, 5.97429e-05, 8.325076e-05, 7.315634e-07, 1.334374e-08, 
    6.803837e-09, 9.636648e-08, 1.717062e-07, 2.31045e-06, 1.473709e-05,
  1.879121e-07, 8.01012e-06, 1.869559e-05, 1.861588e-05, 3.150646e-05, 
    2.878649e-05, 2.691049e-05, 4.048352e-08, 9.576911e-07, 1.201396e-06, 
    1.015818e-08, 1.20245e-07, 1.207073e-07, 2.217042e-08, 5.560554e-09,
  3.0086e-09, 3.097631e-09, 3.979252e-09, 2.249823e-08, 5.009494e-08, 
    4.4424e-08, 2.733818e-08, 2.397091e-08, 1.281516e-07, 1.667952e-06, 
    5.699859e-06, 9.217387e-06, 1.522558e-05, 2.980461e-05, 6.486044e-05,
  5.040149e-09, 8.996954e-09, 2.130506e-08, 1.886005e-08, 6.359853e-08, 
    6.039031e-08, 3.025566e-08, 1.151228e-08, 1.897471e-06, 5.237808e-06, 
    1.48025e-05, 3.687357e-05, 2.767569e-05, 3.563195e-05, 6.36945e-05,
  1.548565e-08, 3.943992e-08, 4.280153e-08, 5.815351e-08, 5.210126e-07, 
    3.525586e-07, 6.939981e-08, 6.13962e-06, 1.598417e-05, 3.631172e-05, 
    3.740552e-05, 6.299677e-05, 8.274549e-05, 5.616732e-05, 3.508369e-05,
  1.688129e-08, 2.469378e-08, 8.016796e-08, 3.162095e-06, 9.289743e-07, 
    8.774451e-06, 1.92491e-05, 3.203647e-05, 6.467765e-05, 0.0001072567, 
    0.0001257699, 9.14401e-05, 7.043084e-05, 6.155379e-05, 1.159061e-05,
  2.469958e-08, 2.161377e-08, 2.181601e-08, 9.17892e-07, 6.104281e-07, 
    1.107595e-05, 2.742278e-05, 6.425401e-05, 0.0001589457, 0.0001308368, 
    1.351944e-05, 1.585612e-05, 7.522805e-05, 1.837858e-05, 9.001396e-06,
  4.524922e-08, 1.174015e-06, 4.02595e-08, 3.284473e-06, 8.671415e-06, 
    1.95971e-05, 3.295745e-05, 9.305616e-05, 0.0001471088, 1.579457e-08, 
    8.445996e-07, 6.986372e-07, 3.974634e-08, 6.72055e-06, 5.109406e-05,
  5.77272e-08, 8.313018e-08, 1.341422e-07, 2.799762e-06, 6.769134e-06, 
    1.485825e-05, 2.810712e-05, 7.229526e-05, 0.000136447, 6.211438e-08, 
    1.062544e-09, 2.404838e-09, 9.400013e-09, 4.258457e-05, 8.499675e-05,
  3.317907e-08, 1.191489e-06, 4.953871e-06, 5.975921e-07, 3.748849e-06, 
    1.609767e-05, 3.006911e-05, 9.00657e-05, 0.0001957479, 2.078153e-09, 
    1.451424e-09, 1.3506e-08, 1.120077e-08, 0.0001117691, 4.756813e-05,
  2.972197e-08, 3.011215e-06, 2.369235e-06, 1.303658e-06, 3.83969e-06, 
    1.624826e-05, 3.228167e-05, 5.928702e-05, 3.168502e-07, 4.093521e-07, 
    6.181365e-07, 4.488548e-07, 5.227114e-07, 4.06669e-05, 3.494239e-05,
  3.544149e-08, 6.645497e-08, 1.370881e-07, 9.349599e-09, 9.004854e-07, 
    7.497682e-06, 1.873236e-05, 2.03955e-06, 5.139896e-07, 1.372461e-06, 
    2.547524e-06, 6.72656e-06, 6.480989e-06, 5.57252e-05, 3.038734e-05,
  6.052608e-08, 3.05783e-09, 2.79047e-07, 5.833113e-07, 3.927244e-06, 
    2.075087e-06, 3.535682e-07, 1.519196e-08, 1.74619e-08, 2.983993e-06, 
    1.474083e-05, 2.993631e-05, 4.048131e-05, 5.640273e-05, 1.153857e-05,
  6.331761e-08, 6.509049e-09, 6.783865e-07, 7.765663e-06, 3.509307e-06, 
    1.418913e-05, 3.185029e-06, 1.053818e-06, 4.373137e-07, 2.686045e-06, 
    6.113429e-06, 1.597847e-05, 2.806905e-05, 5.008371e-05, 6.492413e-06,
  3.624093e-07, 5.876185e-07, 2.272873e-06, 9.049614e-06, 8.679813e-06, 
    1.992606e-05, 9.008028e-06, 7.310169e-06, 1.939562e-05, 1.882187e-05, 
    2.515391e-05, 3.228745e-05, 5.866793e-05, 3.644982e-05, 2.471258e-05,
  1.799747e-06, 9.073482e-07, 1.145833e-05, 1.626973e-05, 2.707771e-05, 
    4.055774e-05, 3.284866e-05, 3.618521e-05, 4.131539e-05, 4.490646e-05, 
    5.81227e-05, 6.25746e-05, 7.527932e-05, 9.249704e-05, 4.709646e-05,
  1.573229e-05, 5.695685e-06, 5.327276e-06, 8.457607e-06, 2.118059e-05, 
    1.55661e-05, 1.334698e-05, 2.592889e-05, 3.340708e-05, 3.767723e-05, 
    1.954181e-08, 1.230498e-08, 6.804513e-05, 7.335033e-05, 6.949635e-05,
  3.55561e-05, 3.77746e-05, 1.567834e-05, 6.580332e-06, 2.845658e-05, 
    3.545411e-05, 2.075927e-05, 9.255609e-06, 2.563834e-05, 4.635969e-08, 
    4.581917e-08, 4.540254e-07, 3.091185e-08, 2.208187e-05, 8.41498e-05,
  4.868166e-05, 3.981912e-05, 1.470134e-05, 2.941698e-05, 6.666039e-05, 
    4.687261e-05, 2.721529e-05, 7.397223e-06, 3.010611e-05, 9.446611e-09, 
    1.203455e-09, 4.650321e-08, 3.30567e-09, 2.579515e-05, 7.805176e-05,
  1.909225e-05, 2.376359e-05, 1.546931e-05, 2.077794e-05, 5.626214e-05, 
    6.104075e-05, 5.437439e-05, 5.536031e-05, 6.768199e-05, 4.716856e-08, 
    9.673606e-10, 2.579001e-07, 2.270019e-09, 7.331705e-06, 1.517856e-05,
  7.029906e-06, 1.733916e-05, 1.844441e-05, 4.196631e-05, 3.807559e-05, 
    6.671864e-05, 7.521153e-05, 7.051695e-05, 4.483702e-09, 1.00981e-08, 
    6.64934e-08, 5.938537e-07, 4.903532e-07, 2.036717e-06, 2.091389e-07,
  7.052175e-06, 2.254015e-05, 4.236258e-05, 3.306243e-05, 2.658997e-05, 
    2.288277e-05, 2.28951e-05, 3.809405e-09, 1.01132e-08, 7.813978e-08, 
    4.181884e-09, 1.071959e-07, 1.671994e-06, 8.957441e-06, 2.778123e-06,
  2.286751e-09, 5.054627e-09, 5.373691e-07, 3.374471e-07, 8.737885e-06, 
    2.459526e-05, 3.606257e-05, 9.671558e-06, 2.216814e-05, 7.925325e-05, 
    8.948505e-05, 9.982426e-05, 6.075292e-05, 2.886554e-05, 5.511933e-07,
  4.079659e-10, 1.003159e-09, 2.211821e-07, 1.211369e-05, 2.348708e-05, 
    6.542032e-05, 9.059497e-05, 6.647939e-05, 6.971313e-05, 2.560698e-05, 
    2.7572e-05, 3.641554e-05, 4.956369e-05, 4.626059e-05, 2.720509e-06,
  3.546027e-07, 4.901069e-06, 7.805092e-06, 3.53527e-05, 5.728475e-05, 
    9.572943e-05, 0.0001671218, 0.0001361701, 0.0001147521, 7.077234e-05, 
    3.650299e-05, 3.012993e-05, 2.68917e-05, 4.310251e-05, 1.385089e-06,
  6.082577e-06, 7.01709e-06, 2.851409e-05, 6.43642e-05, 6.069968e-05, 
    0.0001591885, 0.0001195235, 0.0002018267, 0.000183118, 0.0002229248, 
    0.0001097331, 6.911641e-05, 6.49643e-05, 6.054645e-05, 1.902681e-05,
  3.479682e-06, 1.199464e-05, 1.56275e-05, 3.860615e-05, 4.782608e-05, 
    0.000103948, 0.0001013981, 0.000142856, 0.0001651339, 0.0001794637, 
    1.117412e-05, 4.672872e-06, 5.750754e-05, 4.819972e-05, 7.949422e-05,
  1.337011e-05, 3.214165e-05, 4.051721e-05, 6.024518e-05, 6.590541e-05, 
    3.792181e-05, 5.551221e-05, 0.0001215868, 0.0001328381, 2.087369e-05, 
    5.152797e-05, 4.349742e-05, 2.591649e-06, 2.24191e-05, 9.741514e-05,
  2.814955e-05, 5.902399e-05, 4.083973e-05, 6.098324e-05, 5.603157e-05, 
    7.52784e-05, 0.0001218169, 0.000110857, 0.0001135615, 1.356739e-05, 
    1.58149e-05, 1.285201e-05, 3.730632e-06, 1.22468e-05, 8.893609e-05,
  1.960325e-05, 6.974221e-05, 6.376803e-05, 6.217338e-05, 7.915907e-05, 
    8.306018e-05, 0.0001481024, 0.0001696348, 0.0001104243, 1.168689e-05, 
    2.209482e-06, 3.251011e-06, 2.334566e-06, 9.338331e-06, 3.969179e-05,
  1.066865e-05, 7.205335e-05, 5.17124e-05, 9.218753e-05, 0.000107577, 
    0.0001341442, 0.0001426657, 0.0001308634, 5.869969e-05, 4.246152e-05, 
    1.230056e-05, 8.926059e-07, 3.273031e-07, 2.191174e-05, 3.359984e-05,
  8.333879e-06, 2.699963e-05, 6.572282e-05, 6.602644e-05, 9.847971e-05, 
    9.880973e-05, 0.0001107234, 2.877121e-05, 5.50959e-05, 4.252942e-05, 
    2.781025e-05, 4.994136e-06, 7.657005e-07, 1.183299e-05, 2.408782e-05,
  6.006847e-06, 3.002052e-08, 1.939039e-05, 2.737321e-07, 1.838267e-05, 
    1.502043e-05, 7.00633e-05, 7.022951e-05, 6.544013e-05, 2.663259e-05, 
    1.359804e-05, 6.088284e-06, 7.290044e-06, 2.885992e-05, 1.267802e-05,
  1.02078e-06, 3.76249e-09, 7.861484e-06, 6.7279e-06, 2.082762e-06, 
    1.936454e-05, 5.818964e-05, 8.335122e-05, 9.105267e-05, 5.425736e-05, 
    3.001396e-05, 1.910901e-05, 2.349211e-05, 4.225258e-05, 1.541603e-05,
  8.312666e-06, 1.294385e-05, 5.037656e-06, 5.136892e-06, 1.265985e-05, 
    1.245777e-05, 1.13281e-05, 6.106936e-05, 9.839624e-05, 8.176846e-05, 
    6.547062e-05, 7.469975e-05, 4.998676e-05, 6.111682e-05, 1.601455e-05,
  5.680766e-05, 3.317638e-05, 5.336512e-05, 8.225496e-05, 4.351037e-05, 
    4.547275e-05, 5.133383e-05, 5.220075e-05, 7.787671e-05, 0.000176565, 
    0.0001183182, 9.71421e-05, 7.358415e-05, 8.025074e-05, 6.053859e-05,
  2.257952e-05, 6.491531e-05, 7.348043e-05, 9.107085e-05, 8.840241e-05, 
    6.666413e-05, 5.89613e-05, 8.094909e-05, 0.000112763, 8.179484e-05, 
    1.866049e-05, 1.929878e-05, 0.0001278991, 5.835216e-05, 0.0001102779,
  2.133214e-05, 4.362122e-05, 7.316918e-05, 0.0001182596, 0.000117395, 
    0.0001045663, 0.0001261663, 0.0001150471, 0.0001177963, 1.537372e-06, 
    9.618971e-06, 4.738519e-05, 3.512255e-05, 3.198632e-05, 0.0001402819,
  8.478083e-05, 3.824431e-05, 2.316403e-05, 4.794717e-05, 5.332005e-05, 
    9.029663e-05, 0.0002077403, 0.0003053559, 0.000232551, 2.372538e-07, 
    9.830333e-08, 1.969586e-07, 6.929634e-06, 9.154445e-05, 0.0001428416,
  9.66833e-05, 0.0001061879, 5.054245e-05, 2.575038e-05, 4.116762e-05, 
    8.660198e-05, 0.0001676761, 0.00024811, 0.0002737354, 2.61392e-05, 
    2.343616e-07, 1.582781e-08, 2.746457e-08, 0.0001473815, 7.217233e-05,
  0.0001073967, 0.0001384814, 0.0001519768, 0.0001021299, 3.758644e-05, 
    5.469987e-05, 0.0001255445, 0.0001666294, 7.621132e-06, 8.128513e-06, 
    2.109532e-06, 1.617586e-08, 1.63218e-08, 9.351371e-05, 6.90223e-05,
  5.81824e-05, 0.0001013174, 0.0001662481, 0.0001544534, 0.0001041694, 
    2.452312e-05, 2.350423e-05, 8.090637e-06, 6.540409e-07, 2.252817e-07, 
    3.379992e-09, 1.972152e-09, 5.36298e-09, 4.868908e-05, 4.176082e-05,
  1.345242e-06, 4.356832e-05, 0.0002080021, 0.0001010268, 6.772423e-05, 
    4.428759e-05, 7.480547e-05, 5.04905e-05, 8.223236e-05, 7.637057e-05, 
    6.374936e-05, 5.306797e-05, 6.21568e-05, 5.361962e-05, 2.516666e-06,
  2.382022e-09, 7.258544e-09, 0.0001421051, 0.0001667653, 9.349361e-05, 
    4.722744e-05, 7.917275e-05, 0.0001100738, 0.0001773902, 0.0001579767, 
    0.0001001902, 6.073543e-05, 7.513812e-05, 8.08156e-05, 3.981684e-06,
  1.806016e-05, 4.869649e-05, 3.556829e-05, 5.045435e-05, 5.387796e-05, 
    3.309427e-05, 3.450374e-05, 0.0001363256, 0.0002175556, 0.0002419878, 
    0.0002695106, 0.0002153674, 0.0001537346, 0.0001028569, 4.674688e-06,
  2.971061e-05, 4.67463e-05, 8.094938e-05, 5.899477e-05, 6.023009e-05, 
    4.342108e-05, 6.371404e-05, 0.0001060124, 0.0002503384, 0.0002745695, 
    0.0002762042, 0.0002219915, 0.0001993403, 0.0001114542, 2.024661e-05,
  2.647972e-05, 4.963576e-05, 6.799494e-05, 9.735557e-05, 8.70084e-05, 
    9.900725e-05, 7.578587e-05, 0.0001353374, 0.0002913148, 0.0003423443, 
    7.391773e-05, 0.0001032916, 0.000187919, 8.307192e-05, 6.638636e-05,
  2.95431e-05, 4.682337e-05, 7.944253e-05, 6.147089e-05, 6.208384e-05, 
    8.04076e-05, 9.975508e-05, 0.0001419255, 0.0002329042, 8.049529e-05, 
    2.421584e-05, 0.000145062, 0.0001135921, 9.401108e-05, 0.0001556795,
  3.850868e-05, 6.113938e-05, 6.249754e-05, 5.14294e-05, 8.632272e-05, 
    0.0001263028, 0.0002236392, 0.0001178773, 0.0001689158, 7.89336e-05, 
    1.357101e-05, 2.787296e-05, 4.492868e-05, 0.0001259628, 0.0001480645,
  1.640823e-05, 5.142438e-05, 7.876991e-05, 3.796461e-05, 2.639885e-05, 
    7.866124e-05, 0.0001577125, 5.015704e-05, 9.530417e-05, 7.893301e-05, 
    6.174722e-06, 1.132727e-06, 1.485159e-06, 9.49542e-05, 0.0001147888,
  6.991142e-06, 4.084467e-05, 4.539041e-05, 7.231813e-05, 8.80945e-05, 
    7.276228e-05, 7.895573e-05, 7.022212e-05, 1.595756e-05, 6.051387e-05, 
    5.909284e-06, 6.057741e-07, 1.899965e-07, 7.452151e-05, 0.0001392125,
  1.93757e-06, 1.720797e-05, 7.875512e-05, 8.028997e-05, 0.0001239583, 
    7.257875e-05, 0.0001320247, 3.75713e-06, 1.933491e-05, 2.452489e-05, 
    1.164001e-05, 2.12208e-06, 8.898028e-07, 5.247103e-05, 8.571074e-05,
  6.598026e-09, 1.855035e-05, 7.585465e-05, 6.495179e-05, 6.2769e-05, 
    8.515309e-05, 0.0001453637, 0.0001260331, 0.0002394615, 9.470432e-05, 
    3.677572e-05, 2.978806e-05, 2.341463e-05, 2.655481e-05, 2.93962e-08,
  8.564318e-10, 5.737273e-10, 2.679285e-05, 4.696202e-05, 3.340849e-05, 
    6.332574e-05, 9.056455e-05, 9.250198e-05, 9.008014e-05, 6.921407e-05, 
    8.263323e-05, 7.101188e-05, 1.947407e-05, 2.39535e-05, 9.134021e-07,
  2.494589e-08, 8.283134e-07, 3.48336e-07, 2.227606e-07, 2.60959e-05, 
    5.428147e-05, 6.002724e-05, 6.3119e-05, 0.0001933975, 0.0001778772, 
    0.0001811184, 0.0001080292, 5.299054e-05, 3.568924e-05, 9.11827e-06,
  3.551751e-07, 1.809886e-07, 3.339486e-06, 1.21774e-05, 2.62788e-05, 
    8.137663e-05, 7.141045e-05, 0.0001342493, 0.0001774273, 0.0002320847, 
    0.0002599071, 0.0002394385, 8.166925e-05, 0.0001064003, 2.672502e-05,
  2.652624e-08, 2.720869e-10, 2.283207e-06, 2.781265e-06, 8.535336e-06, 
    4.744171e-05, 7.543866e-05, 0.0001143301, 0.0001265935, 0.0003034768, 
    0.0003239375, 0.0001812823, 0.0003812136, 0.0001271545, 0.0001250948,
  2.168036e-09, 3.282699e-07, 3.097881e-07, 1.567841e-06, 3.738766e-06, 
    3.361787e-05, 7.386872e-05, 9.398832e-05, 4.234273e-05, 2.099679e-05, 
    6.219994e-05, 0.0002133908, 0.0002456641, 0.0002880594, 0.000158212,
  7.224884e-10, 6.481377e-08, 2.142061e-08, 1.161814e-06, 3.401718e-06, 
    8.606905e-06, 6.619278e-05, 5.428774e-05, 2.311524e-05, 3.792688e-06, 
    1.727975e-05, 4.727567e-05, 5.457664e-05, 0.0003247143, 0.0002243865,
  4.746324e-09, 3.115028e-09, 1.684098e-08, 6.021542e-07, 1.807553e-06, 
    4.411838e-06, 2.176507e-05, 3.702371e-05, 2.498571e-05, 4.126134e-06, 
    3.221131e-06, 2.432985e-06, 1.430448e-06, 0.0002106306, 0.0002290739,
  1.27365e-08, 4.305599e-09, 7.290961e-08, 1.347497e-06, 6.124491e-06, 
    1.045507e-05, 1.314022e-05, 2.041762e-05, 8.505757e-07, 1.510402e-05, 
    1.695614e-06, 7.578883e-08, 1.564226e-05, 0.0002004279, 0.0002886049,
  9.854514e-09, 8.47296e-09, 6.315489e-09, 2.362941e-09, 2.325287e-07, 
    2.762304e-06, 8.194679e-06, 1.193838e-07, 4.459014e-06, 3.031341e-06, 
    1.514712e-06, 4.623869e-08, 5.308577e-07, 9.939889e-05, 0.0001499433,
  2.524086e-13, 1.036652e-11, 9.396563e-09, 9.896355e-09, 7.088509e-13, 
    3.626345e-09, 5.35469e-07, 1.399769e-05, 3.788997e-05, 7.061035e-05, 
    8.001738e-05, 8.598515e-05, 6.721442e-05, 6.850914e-05, 7.324151e-05,
  1.219304e-10, 1.527645e-11, 4.690257e-07, 6.557219e-07, 1.574095e-13, 
    4.379096e-09, 3.371886e-08, 6.913857e-07, 1.393839e-05, 3.226657e-05, 
    3.996018e-05, 5.205124e-05, 6.096672e-05, 6.808758e-05, 5.934109e-05,
  1.0225e-08, 8.787248e-09, 1.285802e-09, 4.194917e-10, 3.444091e-09, 
    2.968947e-07, 1.513299e-08, 4.314496e-07, 5.400714e-06, 1.430959e-05, 
    1.760568e-05, 2.616427e-05, 5.152117e-05, 5.445731e-05, 2.893139e-05,
  4.118912e-08, 3.112264e-08, 2.019218e-08, 2.940398e-08, 2.635764e-08, 
    6.443587e-06, 3.843915e-06, 2.866053e-06, 7.841733e-06, 1.33166e-05, 
    4.447102e-06, 5.790667e-06, 1.029373e-05, 2.422511e-05, 1.755441e-06,
  9.169765e-07, 7.841629e-08, 3.376893e-08, 1.685541e-08, 1.356747e-09, 
    1.000616e-08, 1.84813e-07, 5.354978e-06, 9.23837e-06, 6.244908e-06, 
    1.495777e-10, 1.221778e-09, 1.933423e-06, 2.607621e-06, 1.515906e-05,
  1.431953e-07, 1.230139e-07, 7.992268e-08, 2.823237e-08, 1.042299e-08, 
    9.234745e-09, 7.670647e-06, 6.055538e-07, 2.516451e-06, 1.643568e-10, 
    2.69148e-11, 2.273236e-10, 5.469143e-08, 2.761838e-05, 4.53076e-05,
  1.538973e-07, 1.886325e-07, 2.602087e-07, 1.811533e-07, 6.977712e-08, 
    1.501235e-08, 7.019898e-07, 1.077092e-07, 1.618668e-08, 3.51329e-10, 
    3.134872e-12, 1.994492e-10, 4.973882e-06, 2.562521e-05, 4.706395e-05,
  1.641744e-07, 2.305913e-07, 4.622759e-07, 2.118229e-07, 1.102876e-07, 
    4.506695e-08, 9.183473e-08, 1.131287e-06, 4.437708e-09, 5.004436e-11, 
    5.888458e-12, 5.589701e-12, 5.182227e-08, 1.772405e-05, 9.189676e-06,
  7.567416e-07, 6.500245e-07, 9.013307e-07, 1.813434e-06, 4.907843e-06, 
    1.836741e-06, 1.348868e-06, 9.592725e-07, 4.866988e-10, 1.001319e-10, 
    1.795072e-09, 2.038429e-11, 1.435813e-08, 2.339526e-06, 9.132803e-08,
  1.571502e-06, 2.037279e-06, 1.668057e-06, 7.177413e-07, 3.380567e-07, 
    2.776136e-07, 5.791362e-07, 1.341217e-08, 5.884492e-10, 2.052845e-10, 
    2.59295e-09, 1.902631e-10, 1.071872e-09, 1.066109e-06, 7.346405e-08,
  8.663909e-09, 1.410897e-08, 9.426977e-09, 1.921347e-09, 7.785175e-10, 
    3.146569e-10, 4.91573e-11, 4.028577e-11, 2.735978e-10, 1.339666e-09, 
    6.18341e-09, 4.477961e-08, 9.80684e-08, 3.180803e-06, 2.080691e-05,
  1.137808e-08, 1.695191e-08, 1.993995e-08, 8.313846e-09, 3.571603e-09, 
    6.411248e-09, 6.691906e-09, 1.076159e-09, 3.026418e-07, 9.998082e-09, 
    3.238219e-08, 8.749683e-09, 9.216755e-09, 5.185557e-07, 7.72563e-06,
  6.701569e-08, 6.973158e-08, 4.038677e-08, 1.764012e-08, 1.261116e-08, 
    9.891139e-09, 3.349284e-09, 4.237133e-09, 2.547625e-06, 5.518665e-07, 
    5.3108e-08, 1.85909e-08, 3.381945e-09, 1.191351e-08, 7.387174e-09,
  8.874001e-08, 8.828329e-08, 5.41641e-08, 2.891395e-08, 2.606008e-08, 
    2.907939e-08, 2.630248e-08, 1.16483e-06, 4.65504e-06, 1.198262e-06, 
    1.848294e-08, 1.004985e-08, 2.328783e-10, 1.987674e-11, 4.075376e-10,
  1.152221e-07, 1.098962e-07, 7.80776e-08, 5.566528e-08, 3.594676e-08, 
    2.927107e-08, 3.673947e-08, 2.706214e-07, 9.257764e-06, 1.151636e-05, 
    2.656239e-10, 7.513009e-15, 3.564253e-12, 1.98567e-13, 3.587807e-09,
  1.382293e-07, 1.687206e-07, 2.461108e-07, 1.139172e-06, 8.3941e-07, 
    3.282339e-08, 1.240368e-07, 1.134188e-06, 1.001977e-05, 2.469173e-10, 
    1.260038e-11, 4.288628e-12, 2.947903e-13, 5.728617e-14, 9.598418e-12,
  8.364719e-08, 1.077799e-07, 9.267763e-07, 1.14887e-05, 3.238441e-06, 
    6.230166e-08, 3.158116e-08, 1.38458e-08, 4.593165e-06, 2.834526e-10, 
    3.98542e-11, 2.339687e-11, 1.261674e-22, 2.431266e-13, 4.08459e-11,
  1.223474e-07, 1.120629e-06, 3.666588e-07, 3.537471e-07, 2.48995e-07, 
    8.94907e-08, 5.424894e-08, 8.947623e-07, 2.040761e-06, 2.763191e-10, 
    1.063507e-10, 5.974684e-12, 1.515486e-22, 2.646481e-14, 2.102024e-11,
  3.724742e-07, 2.364254e-05, 2.441246e-05, 8.049507e-06, 2.446744e-06, 
    9.360957e-07, 6.780461e-08, 2.394467e-06, 1.974432e-09, 3.225477e-10, 
    1.774958e-10, 5.079546e-11, 2.420603e-23, 6.195467e-24, 9.913922e-12,
  4.954406e-07, 7.038624e-06, 3.446457e-05, 2.363122e-05, 3.650783e-06, 
    2.644904e-06, 8.311146e-08, 7.391193e-08, 1.113351e-08, 4.482534e-10, 
    3.450126e-10, 2.064396e-10, 5.034284e-11, 1.476548e-12, 4.45075e-10,
  1.229996e-08, 1.288771e-08, 9.123451e-09, 2.163159e-09, 1.603837e-09, 
    9.040938e-11, 3.05545e-12, 1.338673e-12, 1.368017e-11, 2.625749e-10, 
    3.270743e-10, 8.524556e-10, 1.099404e-10, 2.437246e-09, 2.711587e-10,
  1.346718e-08, 2.419974e-08, 2.54862e-08, 8.02793e-09, 1.83098e-09, 
    4.790096e-10, 7.411783e-11, 2.596086e-13, 1.295894e-07, 5.545652e-10, 
    2.613472e-10, 5.022064e-12, 3.856474e-10, 1.191442e-08, 1.286661e-10,
  1.081241e-08, 2.173472e-08, 4.771621e-08, 4.816048e-08, 1.295437e-08, 
    1.399914e-09, 8.183811e-11, 5.927934e-09, 1.28447e-06, 4.203486e-06, 
    4.948876e-09, 1.895622e-12, 1.984616e-10, 2.139414e-10, 6.593414e-11,
  2.24558e-08, 4.884672e-08, 4.801698e-08, 6.725433e-08, 4.283055e-08, 
    1.975446e-08, 1.644648e-09, 1.416038e-07, 1.247697e-06, 3.115725e-06, 
    2.229886e-06, 8.489407e-10, 4.849774e-10, 1.043003e-10, 7.807941e-11,
  1.410723e-07, 9.799092e-08, 7.32231e-08, 8.227152e-08, 6.777954e-08, 
    4.462577e-08, 1.258536e-08, 2.116732e-07, 1.687542e-08, 1.630967e-06, 
    1.342033e-10, 7.533649e-11, 1.196298e-09, 7.61619e-11, 1.000004e-11,
  4.106707e-07, 2.885425e-07, 1.790028e-07, 1.096655e-07, 8.220643e-08, 
    5.998977e-08, 3.538049e-08, 8.128796e-09, 3.040205e-07, 1.062462e-10, 
    5.034143e-10, 2.685504e-11, 4.774261e-11, 6.412437e-10, 2.782499e-11,
  5.36977e-07, 3.687761e-07, 2.440999e-07, 1.514894e-07, 1.396469e-07, 
    7.138647e-08, 2.598981e-07, 1.894151e-08, 5.440565e-10, 2.421845e-09, 
    3.80446e-10, 1.079878e-10, 8.592765e-11, 7.977973e-11, 1.393641e-11,
  3.018528e-07, 1.601905e-06, 1.108269e-05, 4.828401e-06, 2.4144e-06, 
    5.378457e-06, 3.121033e-06, 6.346132e-07, 8.036628e-09, 1.91009e-09, 
    2.383903e-10, 1.352061e-10, 1.512141e-10, 2.713192e-11, 1.867782e-08,
  1.377041e-07, 1.9436e-07, 7.356867e-07, 1.997743e-05, 1.971857e-05, 
    3.966844e-05, 1.542003e-05, 6.266683e-06, 1.106125e-08, 1.331029e-09, 
    1.705938e-10, 8.495075e-11, 1.00323e-10, 1.730245e-11, 4.960404e-12,
  2.540711e-07, 9.772224e-08, 5.683874e-08, 9.687732e-08, 1.247966e-05, 
    1.189298e-05, 9.639395e-06, 3.297749e-08, 2.158213e-08, 3.561752e-09, 
    4.733641e-10, 6.698177e-11, 5.925049e-11, 3.450936e-11, 7.995035e-12,
  3.415849e-08, 1.082177e-09, 1.163056e-08, 2.004692e-09, 2.444066e-09, 
    9.937472e-11, 3.649909e-11, 4.306925e-11, 3.358708e-11, 1.627775e-12, 
    4.046661e-09, 7.49144e-07, 9.694693e-07, 2.184963e-08, 1.44021e-09,
  6.513353e-08, 4.490222e-09, 8.432776e-09, 6.818709e-09, 7.332451e-09, 
    2.690233e-08, 1.707267e-08, 1.21037e-10, 3.280301e-10, 1.112141e-10, 
    5.482374e-12, 5.072903e-10, 4.184146e-07, 4.805367e-09, 9.004008e-11,
  7.105579e-08, 2.630576e-08, 2.756028e-08, 3.134744e-08, 1.313228e-07, 
    1.385623e-06, 1.916901e-08, 1.510739e-06, 1.608066e-05, 4.545405e-07, 
    3.556734e-07, 2.497337e-10, 5.467832e-07, 1.865385e-08, 1.403721e-11,
  1.111258e-07, 8.493348e-08, 3.358666e-08, 1.224982e-05, 5.58954e-06, 
    8.224863e-06, 3.949316e-06, 7.427714e-06, 3.042261e-05, 3.21575e-05, 
    3.629042e-05, 6.286872e-06, 4.63726e-06, 1.263163e-08, 7.408316e-11,
  1.38837e-07, 1.317674e-07, 4.924814e-08, 5.542049e-07, 1.69564e-06, 
    4.560682e-06, 1.081923e-05, 9.433395e-06, 1.018499e-05, 2.552725e-05, 
    6.898385e-09, 6.36301e-10, 1.740229e-06, 2.645092e-09, 7.557113e-08,
  1.301692e-07, 1.365378e-07, 1.160851e-07, 2.980636e-06, 2.714081e-06, 
    4.580269e-06, 1.685543e-05, 2.146994e-05, 1.416613e-06, 4.080313e-09, 
    2.492372e-09, 1.058396e-09, 5.347026e-09, 7.781732e-08, 6.77703e-08,
  7.032815e-08, 2.853883e-06, 1.87393e-07, 4.138838e-06, 7.975505e-06, 
    9.288364e-06, 6.02776e-06, 2.3793e-07, 4.201997e-09, 3.809173e-09, 
    4.206087e-09, 4.709848e-09, 6.154915e-10, 5.971458e-10, 1.762501e-06,
  2.870702e-08, 6.634316e-08, 1.068719e-07, 1.131233e-06, 1.620001e-05, 
    1.634325e-05, 2.504021e-05, 4.439311e-08, 7.486157e-09, 4.135927e-09, 
    3.732845e-09, 2.892417e-09, 3.642342e-09, 6.375486e-10, 1.864617e-06,
  2.936519e-09, 1.366285e-08, 5.415894e-08, 2.248621e-07, 1.095367e-06, 
    1.25132e-05, 1.172695e-05, 1.075505e-07, 2.336319e-09, 3.200194e-09, 
    3.842435e-09, 2.562789e-09, 4.987484e-09, 2.573819e-08, 3.919621e-08,
  2.456799e-12, 1.18657e-10, 4.664006e-09, 5.133659e-09, 8.726365e-09, 
    1.087951e-09, 1.95231e-09, 5.852944e-10, 2.250507e-09, 2.884039e-09, 
    3.376834e-09, 2.803789e-09, 2.485441e-09, 6.116199e-09, 3.073693e-09,
  6.894401e-08, 4.618102e-08, 1.810831e-08, 1.288085e-09, 3.960093e-10, 
    3.65958e-10, 6.684112e-10, 5.622159e-10, 5.927405e-10, 2.110663e-10, 
    5.428226e-11, 7.613754e-09, 4.238687e-10, 1.004279e-08, 4.162293e-09,
  6.60944e-08, 5.072555e-08, 3.206006e-08, 8.788151e-07, 1.994342e-06, 
    9.872805e-07, 9.146541e-08, 8.645545e-08, 1.297352e-07, 1.291282e-08, 
    8.459761e-10, 8.989511e-10, 5.66585e-09, 1.125517e-07, 2.402461e-10,
  7.447448e-08, 4.870834e-08, 9.584461e-07, 1.375453e-06, 7.288515e-06, 
    1.548651e-05, 3.037068e-06, 2.59912e-06, 2.625321e-05, 2.577725e-05, 
    1.387781e-06, 1.792097e-06, 9.076409e-07, 1.016936e-06, 1.093715e-10,
  5.160669e-08, 3.750878e-08, 9.96211e-06, 6.906792e-05, 3.465337e-05, 
    7.465061e-05, 5.401966e-05, 2.952413e-05, 4.238244e-05, 6.992249e-05, 
    1.685797e-05, 3.040004e-06, 8.402117e-06, 1.976769e-06, 3.076851e-09,
  2.101534e-08, 1.45753e-08, 1.737657e-08, 2.841901e-06, 2.905195e-05, 
    9.34987e-05, 8.92039e-05, 6.763321e-05, 8.081878e-05, 3.211433e-05, 
    2.745526e-08, 7.240748e-09, 2.616668e-06, 4.652558e-07, 3.298654e-06,
  6.283389e-09, 8.192687e-07, 3.918731e-06, 9.865276e-06, 2.561571e-05, 
    9.523108e-05, 0.0001416434, 7.660086e-05, 1.538611e-05, 2.738118e-08, 
    6.668582e-09, 3.116652e-09, 3.458095e-08, 4.815387e-06, 2.253237e-05,
  3.215881e-05, 5.13184e-05, 6.60279e-05, 4.753546e-05, 3.230859e-05, 
    2.890422e-05, 3.818781e-05, 5.57477e-07, 6.548117e-08, 4.125153e-09, 
    3.821304e-09, 3.544781e-09, 4.600696e-09, 1.692758e-05, 4.136005e-05,
  5.408253e-05, 0.0001170368, 0.0001340249, 0.0002112986, 0.0001200673, 
    6.456544e-05, 8.89848e-06, 1.740008e-06, 1.655256e-06, 6.526087e-09, 
    3.279516e-09, 4.411413e-09, 3.615064e-09, 3.142018e-05, 8.469154e-05,
  1.576425e-05, 5.275855e-05, 7.280143e-05, 8.64832e-05, 0.0001405011, 
    8.290106e-05, 2.01522e-05, 1.074019e-05, 4.975961e-07, 3.1968e-07, 
    1.832449e-08, 8.203812e-09, 2.960403e-09, 6.637937e-06, 1.776068e-05,
  4.129086e-09, 1.975146e-07, 5.991118e-07, 4.170211e-06, 6.953108e-06, 
    8.236627e-06, 1.595338e-05, 2.883988e-05, 5.839006e-05, 3.334114e-05, 
    4.123079e-06, 3.880398e-08, 6.684238e-08, 2.243854e-06, 2.552983e-06,
  6.677834e-08, 8.155627e-08, 4.105505e-06, 3.793198e-06, 2.843015e-06, 
    7.380129e-06, 1.01654e-06, 1.172908e-06, 4.794034e-06, 1.74854e-05, 
    8.8197e-06, 6.961112e-10, 4.360354e-10, 6.702487e-09, 2.943518e-09,
  2.417295e-09, 2.400569e-08, 7.002962e-08, 2.651687e-06, 2.378695e-05, 
    2.93036e-05, 1.614742e-05, 1.102777e-05, 3.344892e-05, 3.40687e-05, 
    2.001935e-05, 9.062877e-08, 4.543223e-09, 1.429996e-09, 8.938209e-10,
  1.499612e-08, 2.209016e-09, 5.785263e-08, 7.124219e-08, 1.92845e-05, 
    3.312356e-05, 3.846742e-05, 4.328634e-05, 3.988941e-05, 6.208855e-05, 
    7.04189e-05, 3.103534e-05, 3.47358e-06, 5.594952e-09, 6.354005e-10,
  1.873014e-10, 5.082276e-09, 8.107563e-09, 5.314175e-07, 1.315103e-05, 
    3.147934e-05, 6.002972e-05, 7.536897e-05, 7.736733e-05, 8.000795e-05, 
    0.0001156981, 6.609307e-05, 1.935963e-05, 2.875574e-07, 2.909646e-09,
  7.031868e-10, 1.586262e-08, 2.673123e-09, 8.461805e-09, 2.993716e-08, 
    8.648426e-06, 3.71584e-05, 9.274256e-05, 0.0001066491, 7.698388e-05, 
    6.447198e-09, 8.651127e-07, 4.573619e-05, 2.421646e-05, 1.696004e-07,
  4.181264e-06, 1.272041e-05, 4.051868e-05, 1.78327e-05, 7.335007e-06, 
    2.196336e-05, 6.204024e-05, 7.073189e-05, 1.494141e-05, 9.963072e-08, 
    9.290726e-09, 5.399166e-09, 8.556667e-09, 7.194786e-06, 3.478289e-05,
  9.732526e-05, 0.0001113471, 9.325798e-05, 6.977341e-05, 5.597011e-05, 
    4.769568e-05, 3.779218e-05, 1.714541e-05, 2.8576e-06, 2.835853e-09, 
    1.168349e-09, 3.926024e-09, 1.37978e-08, 5.560832e-05, 7.251689e-05,
  6.655106e-05, 0.0001188712, 0.0001211612, 0.0001106525, 0.0001372924, 
    0.0001307053, 8.129112e-05, 1.69959e-05, 4.087509e-06, 1.032614e-08, 
    1.538473e-08, 3.667161e-08, 6.561156e-07, 4.162157e-05, 0.0001014708,
  1.120247e-05, 5.30393e-05, 4.42579e-05, 4.081527e-05, 6.879046e-05, 
    7.402193e-05, 5.746265e-05, 1.514509e-05, 1.30902e-08, 4.66623e-07, 
    6.752418e-07, 7.440309e-07, 1.079927e-06, 4.22685e-05, 8.803829e-05,
  4.665005e-09, 1.709079e-05, 2.188395e-05, 2.407993e-05, 1.858292e-05, 
    2.147694e-05, 5.602308e-06, 8.409286e-08, 4.287081e-08, 2.345639e-08, 
    3.330519e-07, 1.754067e-08, 1.835002e-07, 2.123743e-05, 1.491506e-05,
  2.720754e-10, 2.383303e-10, 9.152854e-09, 6.936704e-07, 7.087067e-06, 
    3.110655e-05, 1.816895e-05, 6.950441e-06, 1.298215e-05, 2.46467e-05, 
    4.172883e-05, 4.378509e-05, 1.123644e-05, 4.678576e-06, 1.125667e-09,
  1.688458e-11, 1.098536e-10, 7.591696e-09, 1.760795e-06, 1.930317e-05, 
    4.436534e-05, 5.351344e-05, 3.22982e-05, 5.858856e-05, 3.903569e-05, 
    3.664767e-05, 3.846915e-05, 1.60827e-05, 1.395923e-05, 1.215605e-09,
  9.85991e-10, 1.384189e-11, 2.118634e-10, 2.34836e-06, 4.479293e-05, 
    5.577663e-05, 6.453026e-05, 6.254314e-05, 9.033173e-05, 4.614816e-05, 
    4.054391e-05, 6.769574e-05, 6.551506e-05, 4.913336e-05, 2.516406e-09,
  1.645409e-08, 1.691463e-09, 4.022491e-09, 2.491109e-05, 9.774516e-05, 
    0.0001224396, 9.620901e-05, 0.0001021525, 0.0001487392, 6.408097e-05, 
    1.469504e-05, 3.174568e-05, 4.840818e-05, 0.0001440598, 8.210457e-07,
  1.414744e-08, 7.651537e-09, 3.606763e-09, 2.124762e-05, 5.441138e-05, 
    0.0001033372, 0.0001148424, 0.0001960713, 0.0001126202, 3.417232e-05, 
    4.852953e-07, 3.773658e-08, 2.006991e-05, 4.253096e-05, 6.714448e-05,
  7.603158e-05, 6.158256e-05, 5.871107e-05, 6.226049e-05, 9.905338e-05, 
    3.117965e-05, 4.437577e-05, 2.418957e-05, 2.997194e-05, 5.831279e-07, 
    3.473352e-08, 8.744248e-09, 9.814909e-08, 7.093002e-06, 0.000100196,
  0.000108233, 5.66412e-05, 5.838238e-05, 2.98199e-05, 4.573653e-05, 
    6.226116e-05, 3.908355e-05, 5.571951e-05, 1.681636e-05, 7.697807e-09, 
    3.596015e-09, 3.22614e-09, 1.052435e-08, 2.819867e-05, 0.0001644898,
  6.70615e-05, 7.447326e-05, 8.692651e-05, 7.293934e-05, 8.99958e-05, 
    5.673772e-05, 4.322211e-05, 1.330097e-05, 1.043711e-05, 9.445567e-09, 
    7.198209e-09, 8.247551e-09, 1.169785e-08, 6.229823e-05, 0.0001321756,
  1.797053e-05, 4.735409e-05, 5.683929e-05, 5.837762e-05, 4.262866e-05, 
    5.588492e-05, 9.138296e-06, 1.596708e-05, 2.964003e-08, 5.696185e-09, 
    5.718426e-09, 3.323535e-09, 1.680904e-08, 2.869539e-05, 0.0001274158,
  3.62102e-09, 5.956872e-06, 3.042019e-05, 2.009573e-05, 2.482235e-05, 
    7.609246e-06, 7.578489e-06, 3.848546e-08, 5.089456e-08, 2.149283e-09, 
    2.78417e-09, 4.125708e-09, 3.52822e-09, 2.350822e-05, 1.941727e-05,
  4.109282e-07, 1.688198e-07, 1.039422e-06, 6.711313e-06, 2.411221e-05, 
    3.055717e-05, 2.976981e-05, 2.95313e-05, 5.000931e-05, 6.850515e-05, 
    9.408637e-05, 0.0001137076, 5.378735e-05, 4.956443e-05, 5.331302e-08,
  7.967458e-09, 4.398204e-09, 2.544209e-07, 5.54879e-06, 5.532514e-05, 
    8.984758e-05, 0.0001104246, 9.550626e-05, 0.0001129032, 0.0001128567, 
    0.0001072493, 0.0001424238, 8.290575e-05, 7.78195e-05, 1.233122e-07,
  1.01301e-06, 2.647231e-06, 3.516152e-06, 4.143488e-08, 2.87275e-05, 
    0.0001235749, 0.0001458355, 0.0001282065, 0.0001941852, 0.0001584078, 
    0.0001730594, 0.0001442282, 0.0001044599, 0.0001045338, 7.970103e-09,
  2.392474e-05, 7.71209e-07, 6.624368e-07, 3.93604e-05, 6.081126e-05, 
    0.0001404647, 0.0002153219, 0.0001785102, 0.0002030693, 0.0001455799, 
    0.00010446, 0.0001890372, 0.0001161924, 0.0001578293, 7.109516e-06,
  3.560613e-05, 8.808918e-05, 0.0001373714, 0.0002058832, 0.0001423961, 
    0.0001141839, 0.0001255984, 5.854027e-05, 3.306773e-05, 6.530558e-05, 
    1.950031e-06, 5.826975e-08, 0.0001029639, 0.0001178707, 0.0001098718,
  0.0001343689, 0.0001090615, 8.516629e-05, 6.417969e-05, 8.886509e-05, 
    0.0001167638, 3.299675e-05, 3.158437e-05, 1.880135e-05, 4.793168e-08, 
    1.05697e-08, 7.945219e-09, 1.926835e-08, 2.742774e-05, 0.0001369072,
  0.0001993777, 9.557379e-05, 4.619489e-05, 4.292053e-05, 4.968307e-05, 
    6.051105e-05, 2.470707e-05, 2.794525e-05, 1.636653e-05, 6.261044e-09, 
    3.342904e-09, 2.440261e-09, 3.399599e-09, 1.165113e-05, 0.000102215,
  0.0001091031, 0.0001111622, 8.877822e-05, 0.0001008079, 9.828564e-05, 
    3.316116e-05, 1.264647e-05, 8.378502e-06, 8.373341e-06, 2.372105e-09, 
    2.471283e-09, 9.823714e-10, 1.54775e-09, 4.131919e-05, 3.799151e-05,
  6.589435e-05, 6.839907e-05, 5.587685e-05, 9.67114e-05, 8.424208e-05, 
    8.364222e-05, 2.142045e-05, 2.783432e-05, 9.537638e-10, 1.718729e-09, 
    8.153261e-09, 7.660467e-10, 3.935651e-12, 1.981185e-06, 2.690925e-06,
  5.368743e-06, 3.11855e-05, 1.566745e-05, 3.442014e-05, 2.945939e-05, 
    1.306228e-05, 6.454539e-07, 8.714859e-09, 1.865718e-11, 2.524799e-13, 
    6.878515e-16, 2.024607e-13, 1.477154e-11, 2.192624e-09, 1.533369e-09,
  2.606593e-06, 3.672203e-06, 8.375851e-06, 8.696124e-06, 5.788743e-07, 
    4.059887e-07, 4.205121e-06, 4.178971e-06, 1.153609e-05, 2.049971e-07, 
    3.426173e-08, 2.436085e-08, 3.525478e-08, 9.28671e-06, 8.368977e-09,
  1.983251e-07, 2.256169e-06, 1.440567e-05, 1.991139e-05, 5.094232e-06, 
    1.09254e-05, 2.470202e-05, 1.447993e-05, 2.53464e-05, 1.117623e-05, 
    3.120202e-06, 8.740827e-07, 7.350593e-06, 1.60629e-05, 1.465515e-08,
  0.0001246483, 0.0001066192, 3.457722e-05, 2.706312e-05, 6.005719e-05, 
    5.217944e-05, 0.0001169775, 0.0001114317, 8.902849e-05, 6.897836e-05, 
    4.835955e-05, 3.065503e-05, 2.739217e-05, 6.161817e-05, 9.331005e-07,
  0.0003852844, 0.0002493172, 0.0001688146, 0.0001228331, 0.0001494007, 
    0.0002293223, 0.0001749187, 0.0001990887, 0.0002356576, 0.000210423, 
    0.000159739, 5.591522e-05, 0.0001114746, 0.0001407465, 1.753393e-05,
  0.0004182215, 0.0003595522, 0.0002806697, 7.588937e-05, 2.264163e-05, 
    1.821239e-05, 2.221239e-05, 2.877553e-05, 0.0001123919, 0.0001728928, 
    5.32178e-06, 1.281782e-05, 0.0001012318, 9.236644e-05, 0.0001208451,
  0.0002001581, 0.0001085173, 0.0001079457, 8.458358e-05, 8.651739e-06, 
    3.469665e-05, 3.673987e-05, 9.029527e-05, 0.0002200945, 0.0001302592, 
    0.0001112334, 3.134812e-05, 3.363266e-06, 4.849795e-05, 0.0001845678,
  0.0001684984, 0.0001241803, 8.309398e-05, 4.258789e-05, 2.84368e-05, 
    1.414849e-05, 1.156589e-05, 1.970667e-05, 1.886227e-05, 3.899459e-05, 
    2.222263e-05, 1.334641e-05, 2.741759e-06, 0.0001943299, 0.0001184237,
  6.726961e-05, 7.839652e-05, 5.426651e-05, 3.527642e-05, 3.870946e-05, 
    1.586895e-05, 2.531823e-06, 5.915497e-06, 7.998156e-07, 7.999935e-07, 
    1.60768e-06, 3.543512e-06, 1.003254e-05, 0.0003253595, 9.55448e-05,
  1.609698e-05, 3.540167e-05, 3.335774e-05, 3.291985e-05, 2.185477e-05, 
    1.297581e-05, 4.955054e-06, 1.163085e-05, 4.288154e-09, 5.111439e-07, 
    5.055607e-08, 2.205697e-07, 2.014261e-06, 9.355823e-05, 6.286599e-05,
  1.004386e-08, 7.250999e-07, 5.21456e-06, 7.058725e-07, 9.287047e-08, 
    4.967642e-09, 1.193801e-08, 1.711052e-12, 1.919822e-12, 9.669785e-10, 
    5.887999e-08, 2.514209e-08, 2.938654e-08, 3.046235e-05, 8.997542e-06,
  2.383487e-06, 6.072154e-07, 3.584481e-06, 3.829133e-06, 8.3781e-08, 
    5.897859e-10, 1.703714e-10, 1.695547e-09, 1.169853e-08, 1.525631e-07, 
    2.318826e-08, 1.286748e-08, 4.608971e-09, 7.603731e-09, 5.100524e-09,
  5.320212e-07, 1.136557e-06, 5.143085e-06, 8.62817e-06, 1.160277e-06, 
    1.832888e-08, 4.840303e-10, 2.396905e-10, 5.197412e-09, 4.789088e-08, 
    3.051701e-07, 2.520845e-07, 1.050022e-08, 1.530473e-07, 5.540933e-09,
  0.0001292993, 0.0001816518, 3.22006e-05, 5.698187e-06, 7.712234e-06, 
    3.928337e-07, 8.810733e-08, 5.681092e-08, 5.805668e-07, 1.444226e-06, 
    8.594375e-06, 1.75008e-05, 1.488979e-05, 1.392269e-05, 1.710344e-07,
  0.0003025707, 0.0002314809, 0.0001886052, 5.606593e-05, 3.982992e-05, 
    0.0001740333, 7.828642e-05, 1.505936e-05, 1.403555e-05, 7.036736e-06, 
    2.136001e-05, 3.723717e-05, 3.950323e-05, 6.542598e-05, 1.10492e-05,
  0.0002362627, 0.0001173358, 0.0001230968, 0.000117523, 0.0001216831, 
    0.0001317436, 9.63477e-05, 0.0001255521, 9.317105e-05, 4.118333e-05, 
    1.274211e-08, 1.528978e-07, 0.0001560855, 4.219846e-05, 9.897839e-05,
  1.289756e-05, 4.873696e-06, 1.701354e-06, 2.317421e-06, 1.579313e-05, 
    3.748331e-05, 3.92096e-05, 3.622952e-05, 9.488926e-06, 8.686148e-08, 
    7.440291e-08, 2.457542e-08, 4.141069e-09, 2.342164e-05, 8.386325e-05,
  9.566831e-06, 7.966967e-07, 9.765442e-08, 1.177005e-07, 2.530456e-06, 
    9.462485e-06, 1.525463e-05, 3.390815e-06, 3.039673e-06, 5.791383e-06, 
    2.068635e-08, 3.767783e-08, 3.118449e-08, 6.326203e-05, 7.997889e-05,
  4.638771e-07, 1.024293e-05, 1.798729e-06, 6.647014e-07, 6.130289e-07, 
    3.084631e-06, 1.239245e-06, 2.531162e-07, 1.366858e-05, 1.983652e-05, 
    1.430585e-05, 7.559715e-06, 5.216646e-07, 0.0001124252, 5.960075e-05,
  2.654386e-08, 2.749524e-07, 1.116752e-06, 1.572395e-06, 2.730649e-06, 
    1.343619e-06, 1.509968e-07, 3.298014e-07, 8.313654e-09, 4.944121e-06, 
    4.329044e-06, 5.091379e-06, 1.122033e-05, 2.652792e-05, 0.0001278435,
  5.010904e-11, 1.559505e-10, 7.055875e-10, 1.337734e-10, 1.791659e-09, 
    1.142375e-09, 5.920553e-10, 2.766576e-11, 1.026399e-09, 7.596623e-09, 
    2.416961e-08, 9.011925e-08, 7.114754e-06, 0.0002833403, 0.0001394829,
  1.999554e-06, 1.615772e-06, 1.165198e-06, 2.360733e-08, 4.973828e-11, 
    2.257434e-09, 1.950672e-09, 1.666051e-09, 1.455963e-09, 1.079556e-06, 
    7.759231e-06, 1.41736e-05, 3.416712e-07, 1.003695e-06, 8.219887e-08,
  1.155465e-08, 6.806709e-06, 8.173414e-05, 1.187723e-05, 3.275522e-06, 
    2.353666e-09, 1.213398e-09, 1.034377e-09, 9.232826e-08, 2.217958e-06, 
    8.396076e-06, 1.467976e-05, 6.880414e-06, 3.416294e-06, 3.135584e-07,
  8.272329e-05, 0.0001414362, 0.0001080863, 0.0001042496, 5.368864e-05, 
    1.820579e-05, 5.273639e-08, 7.656104e-09, 1.551842e-06, 1.844072e-05, 
    1.330869e-05, 2.39096e-05, 2.877575e-05, 4.299105e-05, 2.149638e-06,
  5.341707e-05, 6.307293e-05, 0.0001283322, 0.0001542147, 0.0001456262, 
    0.0001044752, 1.858876e-05, 4.925137e-06, 1.650278e-05, 2.940918e-05, 
    5.21298e-05, 8.6138e-05, 6.320085e-05, 0.0001165498, 2.948671e-05,
  2.765175e-05, 3.126363e-05, 7.656065e-05, 0.0001244268, 0.0001112009, 
    8.040192e-05, 3.728298e-05, 4.358051e-05, 2.589563e-05, 1.433012e-05, 
    3.19919e-08, 9.312142e-07, 8.437712e-05, 6.000794e-05, 7.391425e-05,
  7.476541e-06, 3.578363e-05, 6.558208e-05, 8.45435e-05, 8.199021e-05, 
    5.596177e-05, 3.0053e-05, 9.789312e-06, 1.662695e-06, 1.698971e-08, 
    1.022303e-07, 1.735912e-08, 9.13793e-08, 5.443127e-05, 0.0001077355,
  9.449392e-06, 1.267072e-05, 2.049619e-05, 5.691028e-05, 5.442571e-05, 
    2.639825e-05, 9.154241e-06, 5.710285e-07, 2.009502e-08, 1.210249e-08, 
    1.3683e-08, 1.223286e-05, 3.588081e-05, 8.659922e-05, 0.0001269483,
  4.426839e-06, 6.429141e-07, 3.159552e-07, 2.56546e-06, 1.696691e-05, 
    2.647087e-05, 3.358916e-06, 5.979811e-07, 1.135132e-09, 1.858992e-09, 
    4.740098e-09, 2.821043e-08, 6.659536e-08, 0.0001612073, 9.869895e-05,
  7.208397e-06, 8.265992e-06, 4.448011e-07, 1.507615e-07, 2.299395e-07, 
    1.087649e-06, 9.234975e-07, 1.301774e-07, 4.555695e-10, 1.615919e-09, 
    2.254783e-09, 1.642704e-09, 1.776328e-09, 9.535934e-05, 5.45007e-05,
  1.214241e-05, 5.945155e-06, 2.129291e-06, 3.809882e-10, 4.647337e-11, 
    1.197081e-10, 9.502117e-11, 1.940612e-10, 1.801275e-10, 8.390166e-10, 
    1.533484e-09, 1.743336e-09, 2.735476e-09, 6.300335e-05, 5.805005e-05,
  9.948257e-09, 4.510981e-06, 7.881462e-05, 4.536341e-05, 8.342415e-09, 
    9.567001e-09, 9.790138e-09, 9.774938e-09, 1.875915e-06, 2.054969e-05, 
    4.200899e-05, 2.467909e-05, 4.288235e-05, 7.478268e-05, 7.443284e-05,
  1.617768e-08, 5.852237e-08, 0.0001622648, 0.0001003545, 1.674889e-07, 
    2.375776e-08, 3.66915e-09, 1.406626e-08, 8.037371e-07, 1.185606e-05, 
    4.545067e-05, 3.898993e-05, 4.874564e-05, 6.912673e-05, 6.621177e-05,
  8.156796e-05, 0.0001986789, 0.0002083184, 5.219229e-05, 7.00829e-08, 
    3.426744e-07, 2.795226e-08, 1.205101e-06, 6.240013e-06, 4.395131e-05, 
    4.675372e-05, 5.715976e-05, 0.0001203388, 8.165876e-05, 7.682729e-05,
  9.127131e-05, 0.000170164, 0.0001407128, 8.702859e-05, 3.182935e-05, 
    1.553307e-05, 7.499538e-06, 6.396021e-06, 5.256498e-05, 5.733405e-05, 
    5.738288e-05, 8.50279e-05, 9.775128e-05, 0.0001289447, 9.899979e-05,
  4.536643e-05, 8.119406e-05, 7.351011e-05, 7.973118e-05, 3.917746e-05, 
    1.805644e-05, 5.030869e-05, 6.344242e-05, 5.808632e-05, 2.205018e-05, 
    6.610744e-09, 2.582759e-08, 7.301927e-05, 8.658742e-05, 5.772943e-05,
  3.583498e-05, 3.488241e-05, 2.319551e-05, 8.261991e-06, 3.48094e-06, 
    8.660459e-06, 1.313811e-05, 2.357752e-05, 2.524878e-05, 3.138149e-09, 
    2.73494e-09, 7.747742e-09, 3.311144e-08, 5.090349e-05, 4.226878e-05,
  4.396091e-05, 3.341311e-05, 1.168387e-05, 1.011618e-06, 2.050161e-07, 
    3.934842e-09, 5.775477e-06, 8.855534e-07, 4.721865e-06, 3.595935e-09, 
    4.353988e-08, 1.172342e-08, 2.775457e-08, 5.624688e-05, 8.37179e-05,
  1.985547e-05, 2.987817e-05, 3.637497e-05, 1.751063e-06, 2.002779e-09, 
    3.86528e-08, 1.110743e-07, 1.531955e-05, 4.636427e-06, 7.719795e-09, 
    3.796938e-08, 3.123007e-08, 9.04187e-09, 5.778613e-05, 2.694126e-05,
  3.645585e-05, 5.816614e-05, 5.554518e-05, 3.010371e-05, 1.542886e-05, 
    7.937268e-07, 7.363572e-07, 1.217904e-05, 1.52959e-10, 5.636314e-10, 
    1.021655e-09, 3.996468e-09, 1.911332e-08, 2.059363e-05, 3.691601e-06,
  9.043815e-06, 2.459401e-05, 6.676246e-05, 1.620646e-05, 1.064851e-05, 
    4.43577e-06, 2.771798e-09, 2.430479e-10, 7.585158e-11, 2.74262e-11, 
    3.086622e-11, 1.01117e-10, 6.380317e-10, 9.752419e-09, 3.322545e-10,
  4.027357e-09, 1.471717e-05, 5.708466e-05, 4.538682e-05, 9.460891e-06, 
    1.228157e-06, 6.96766e-06, 3.457309e-08, 1.314059e-06, 8.901417e-06, 
    3.058144e-05, 3.983215e-05, 6.570932e-05, 0.0001122336, 0.0001007451,
  4.412285e-09, 5.173407e-09, 0.0001040497, 0.0001299454, 3.221821e-05, 
    2.807785e-05, 8.139092e-06, 5.278921e-07, 5.848212e-06, 1.362159e-05, 
    3.035192e-05, 3.665353e-05, 0.0001051577, 0.0001316184, 0.0001512021,
  3.195214e-05, 5.104087e-05, 3.873921e-05, 3.371805e-05, 6.585605e-05, 
    6.398412e-05, 1.274554e-05, 4.114728e-06, 6.353529e-06, 2.729521e-05, 
    7.712047e-05, 0.0001054675, 0.0001280756, 0.0001207714, 0.0001064115,
  5.949746e-05, 4.55642e-05, 4.278235e-05, 4.919932e-05, 7.425356e-05, 
    8.109985e-05, 7.87578e-05, 4.343997e-05, 4.306527e-05, 6.572211e-05, 
    0.0001169308, 0.0001079637, 0.0001495908, 0.0001306176, 0.0001301148,
  1.715141e-05, 6.596286e-05, 2.337596e-05, 5.132795e-06, 5.224863e-06, 
    3.055408e-05, 8.086865e-05, 8.44039e-05, 0.000139749, 0.0001896451, 
    5.253376e-07, 2.928212e-08, 0.0001277312, 0.0001288546, 6.331159e-05,
  2.984475e-05, 7.51711e-05, 9.535539e-05, 5.639043e-05, 1.53571e-05, 
    1.349123e-05, 3.359862e-05, 4.267212e-05, 4.315897e-05, 1.80541e-07, 
    5.51149e-09, 1.230843e-08, 1.206074e-08, 6.589215e-05, 0.0001030414,
  2.175864e-05, 6.227987e-05, 0.0001018781, 0.0001173427, 6.800544e-05, 
    5.657547e-05, 2.997962e-05, 3.051176e-05, 1.135437e-08, 3.052713e-09, 
    5.692407e-10, 4.421935e-10, 5.226101e-09, 9.359934e-05, 3.760897e-05,
  2.131105e-05, 5.833207e-05, 0.0001166678, 0.0001122584, 0.0001154702, 
    3.574476e-05, 1.185127e-05, 1.107779e-05, 4.074705e-06, 7.129948e-10, 
    1.407445e-10, 2.626526e-10, 2.903141e-09, 0.0001214383, 6.19261e-05,
  1.88323e-05, 4.240788e-05, 7.51546e-05, 7.096222e-05, 5.791664e-05, 
    3.94482e-05, 1.172699e-06, 1.36729e-05, 7.078991e-09, 4.802124e-10, 
    4.72219e-11, 6.281325e-10, 3.211065e-09, 5.097052e-05, 2.992831e-05,
  1.817391e-06, 6.107883e-05, 0.0001076023, 5.374888e-05, 2.602059e-05, 
    1.173137e-05, 1.385826e-06, 8.636623e-09, 4.490971e-09, 9.034123e-11, 
    3.706379e-10, 2.168419e-09, 4.73185e-09, 2.168074e-05, 5.583163e-06,
  1.863406e-09, 3.00958e-07, 3.063989e-05, 2.371191e-05, 1.745892e-05, 
    2.111572e-05, 6.004716e-05, 7.02074e-05, 0.0001352645, 0.0001419692, 
    0.0001200004, 7.791913e-05, 6.426781e-05, 0.0001709095, 0.0001094238,
  9.052322e-09, 4.584803e-09, 3.977111e-05, 5.240594e-05, 6.456846e-05, 
    0.0001006792, 0.0001294142, 7.758407e-05, 7.046657e-05, 0.0001198759, 
    0.0001303284, 0.0001245704, 0.0001453303, 0.000130712, 0.0001698839,
  0.0001203492, 0.0001067632, 5.014445e-05, 5.838899e-05, 0.0001515469, 
    0.0001182761, 9.237459e-05, 0.0001041304, 0.0001023151, 0.0001161767, 
    0.0001378475, 0.0001630138, 0.0001813352, 0.0002225541, 0.0002063842,
  0.000227841, 0.0001571693, 8.995061e-05, 9.312668e-05, 7.75152e-05, 
    8.009955e-05, 9.239672e-05, 9.69411e-05, 0.0001329038, 9.196162e-05, 
    0.0002019584, 0.0002047934, 0.000121422, 0.0001983168, 0.0001915129,
  0.0001378211, 0.000102211, 5.111704e-05, 3.47092e-05, 2.512227e-05, 
    3.246142e-05, 3.601087e-05, 2.886962e-05, 3.918989e-05, 0.0001060761, 
    9.122514e-06, 3.318161e-06, 0.0001959687, 0.0002063575, 0.0001967935,
  4.309391e-05, 8.840001e-05, 5.78136e-05, 5.980842e-05, 6.225178e-05, 
    4.283003e-05, 3.830249e-05, 3.263972e-05, 3.922802e-05, 2.062306e-07, 
    1.67284e-05, 7.748647e-06, 2.270153e-05, 8.809387e-05, 0.0001739462,
  2.213984e-05, 2.66833e-05, 3.113175e-05, 4.822406e-05, 5.159971e-05, 
    5.592216e-05, 3.998907e-05, 2.116777e-05, 1.189356e-05, 7.856132e-06, 
    2.142724e-07, 9.302525e-08, 4.099221e-05, 0.0001930402, 0.0002058536,
  7.486916e-06, 2.07446e-05, 2.368882e-05, 1.349722e-05, 2.496596e-05, 
    2.19292e-05, 3.06773e-05, 2.713157e-05, 5.402468e-05, 1.087277e-08, 
    2.206216e-09, 9.812287e-09, 7.13036e-08, 0.0002619068, 0.0002427167,
  1.25522e-05, 1.97214e-05, 2.550428e-05, 3.649389e-05, 2.640088e-05, 
    2.652453e-05, 3.569138e-05, 6.528271e-05, 1.232672e-06, 2.304847e-08, 
    2.255939e-09, 1.885627e-09, 1.426046e-08, 0.000137328, 0.0001109027,
  1.927274e-05, 3.471785e-05, 5.539418e-05, 2.77575e-05, 4.443512e-05, 
    5.280308e-05, 1.911337e-05, 1.217056e-06, 6.819796e-08, 1.673542e-08, 
    1.003141e-08, 4.082529e-09, 5.034182e-09, 6.448651e-05, 6.374294e-05,
  3.349431e-08, 8.408936e-06, 1.55757e-05, 1.304717e-06, 2.545365e-07, 
    8.211357e-07, 8.399841e-06, 4.544647e-07, 5.120073e-06, 1.651782e-05, 
    2.798667e-05, 4.331776e-05, 5.949521e-05, 0.0001296076, 0.0001508379,
  3.573564e-10, 2.559752e-09, 3.574258e-05, 6.911185e-05, 7.986864e-05, 
    9.048518e-05, 6.171924e-05, 4.228414e-05, 5.808122e-05, 5.876671e-05, 
    9.138228e-05, 9.995006e-05, 0.0001555377, 0.0001805561, 0.0002575334,
  2.428595e-05, 4.576213e-05, 6.115834e-05, 7.107091e-05, 8.184528e-05, 
    9.167319e-05, 8.869545e-05, 8.351982e-05, 0.0001311471, 0.0001219753, 
    0.0001282492, 0.0001052842, 0.0001497917, 0.0001922345, 0.0001350333,
  8.735356e-06, 1.578924e-05, 1.498722e-05, 3.10496e-05, 4.651869e-05, 
    3.323812e-05, 4.794627e-05, 4.709858e-05, 6.061834e-05, 0.0001084146, 
    0.0001653461, 0.0001279215, 0.00019491, 0.0003805652, 0.000160575,
  2.37456e-06, 6.162166e-06, 4.941936e-06, 5.131164e-06, 1.303789e-05, 
    3.109681e-05, 2.587424e-05, 2.514765e-05, 0.000117919, 0.0002935523, 
    1.641056e-05, 8.068623e-06, 0.0004246505, 0.0004142613, 9.738301e-05,
  1.121284e-06, 1.76005e-05, 8.009841e-06, 5.970845e-06, 1.087352e-05, 
    3.735454e-05, 4.890522e-05, 4.439875e-05, 0.0001001412, 1.478713e-05, 
    4.80523e-05, 1.034318e-05, 9.275062e-05, 0.0001403924, 8.907478e-05,
  1.108701e-06, 1.292878e-05, 1.172936e-05, 6.931848e-06, 2.165036e-05, 
    3.976295e-05, 4.822269e-05, 4.064335e-05, 1.992573e-05, 1.434729e-05, 
    8.469833e-07, 2.619985e-07, 8.731266e-05, 0.00015458, 7.038478e-05,
  2.111166e-07, 1.191351e-05, 1.838639e-05, 9.78993e-06, 1.705247e-05, 
    2.379367e-05, 1.820315e-05, 1.754514e-05, 1.688395e-05, 1.919736e-07, 
    1.511404e-08, 3.546223e-08, 4.794027e-07, 0.0001546867, 7.876709e-06,
  1.064977e-06, 1.412615e-05, 1.864701e-05, 1.169286e-05, 2.048645e-05, 
    5.476188e-06, 2.386039e-05, 3.088327e-05, 1.886337e-07, 3.005236e-07, 
    3.723413e-09, 1.353342e-08, 5.000656e-08, 4.942604e-05, 2.645893e-05,
  5.787792e-09, 9.937539e-07, 1.053269e-05, 6.644577e-06, 1.260885e-05, 
    9.932824e-06, 7.006064e-06, 1.316924e-08, 2.326781e-09, 3.616175e-08, 
    4.492951e-09, 6.844462e-09, 7.898357e-09, 4.03688e-07, 2.132786e-05,
  4.397051e-11, 1.627576e-10, 3.542528e-06, 4.075416e-07, 3.397285e-07, 
    5.02857e-07, 8.888994e-08, 9.607824e-07, 1.923907e-07, 3.028482e-05, 
    3.946747e-05, 9.473244e-05, 0.00013303, 0.0001581467, 0.0001690998,
  4.130295e-11, 6.966399e-10, 5.849967e-08, 1.741411e-06, 1.612187e-06, 
    3.479919e-06, 5.921889e-06, 3.913033e-06, 2.682707e-05, 3.876899e-05, 
    5.898925e-05, 7.621464e-05, 0.0001432937, 0.0001022527, 0.0001632067,
  2.259356e-07, 7.807129e-07, 1.562859e-08, 2.866609e-08, 1.450135e-07, 
    3.924384e-06, 4.574523e-06, 3.019883e-05, 3.775901e-05, 3.631943e-05, 
    4.006057e-05, 4.361794e-05, 5.513944e-05, 5.095072e-05, 7.385164e-05,
  5.732808e-07, 7.090503e-07, 9.164151e-07, 2.421782e-06, 1.491986e-06, 
    5.071014e-06, 5.455285e-06, 9.938615e-06, 2.037812e-05, 3.051992e-05, 
    0.0001260183, 8.128969e-05, 4.925638e-05, 7.12459e-05, 6.603132e-05,
  4.72266e-07, 7.778722e-07, 1.765081e-07, 6.632602e-07, 1.492049e-07, 
    2.813586e-06, 4.573509e-06, 6.3875e-06, 1.759327e-05, 5.089491e-05, 
    6.927789e-06, 1.40461e-05, 0.0002324812, 9.166114e-05, 0.0001014819,
  6.24137e-06, 1.710128e-05, 2.410679e-05, 1.30582e-05, 2.273623e-06, 
    5.660521e-06, 7.003074e-06, 7.912969e-06, 1.489378e-05, 6.062772e-07, 
    6.081736e-06, 2.334293e-05, 7.152332e-05, 8.721395e-05, 8.984016e-05,
  1.278355e-05, 2.947647e-05, 1.341266e-05, 5.255579e-05, 9.879814e-06, 
    1.264564e-06, 4.972149e-06, 1.025199e-06, 5.588067e-07, 5.455052e-08, 
    1.416436e-08, 6.205777e-06, 5.764823e-05, 6.852986e-05, 9.500264e-05,
  8.231923e-06, 3.786419e-05, 6.353132e-05, 6.92898e-05, 8.329601e-05, 
    1.388288e-05, 8.977049e-06, 3.657871e-06, 3.475912e-07, 2.315682e-09, 
    2.5995e-09, 2.195175e-08, 1.428213e-05, 0.0002061284, 5.101542e-05,
  1.264436e-05, 5.436488e-05, 9.830701e-05, 0.0001222467, 0.0001038349, 
    5.016231e-05, 1.280938e-05, 5.668928e-06, 8.914508e-08, 5.142169e-10, 
    5.16635e-10, 1.467715e-09, 3.398373e-08, 0.000114328, 7.821454e-05,
  5.337894e-06, 5.776265e-05, 9.180363e-05, 7.818325e-05, 9.216226e-05, 
    5.203304e-05, 3.98523e-07, 1.046672e-08, 2.564891e-10, 1.041159e-09, 
    8.662928e-10, 4.852955e-09, 5.732087e-09, 1.427069e-06, 4.18176e-06,
  6.579132e-11, 1.072632e-11, 3.351167e-08, 2.474516e-10, 1.018463e-12, 
    1.962747e-17, 6.18232e-25, 2.368455e-12, 2.09546e-09, 1.126549e-05, 
    4.255722e-05, 8.814743e-05, 0.0002273071, 0.000124848, 0.0001057748,
  2.017625e-09, 2.353209e-11, 6.646777e-09, 2.555958e-09, 2.079e-12, 
    6.056034e-17, 1.006477e-23, 9.684073e-11, 2.438662e-06, 1.751539e-05, 
    4.648188e-05, 7.4729e-05, 0.0001096546, 5.598676e-05, 5.997433e-05,
  2.894144e-08, 1.295566e-06, 5.60792e-09, 1.09746e-09, 1.059352e-09, 
    6.513827e-09, 3.863725e-14, 1.897393e-11, 1.766388e-07, 1.617867e-05, 
    1.62057e-05, 3.071926e-05, 3.389887e-05, 2.612291e-05, 2.247631e-05,
  9.277197e-06, 5.583742e-06, 2.354713e-05, 1.774639e-05, 9.822482e-06, 
    4.841051e-06, 3.48499e-10, 8.640756e-09, 1.326413e-06, 9.757046e-06, 
    8.7699e-06, 1.422159e-05, 6.872608e-06, 2.183597e-05, 2.674528e-05,
  2.174045e-05, 6.729248e-06, 7.506697e-06, 1.320553e-05, 8.836997e-07, 
    7.393197e-06, 5.834775e-07, 6.191088e-07, 2.255289e-06, 6.886323e-06, 
    1.962121e-08, 5.917015e-07, 1.200034e-05, 3.891717e-05, 1.560568e-05,
  2.05395e-05, 2.85232e-05, 2.604832e-05, 2.912967e-05, 2.870133e-05, 
    1.080022e-05, 1.121393e-05, 5.484422e-06, 3.599138e-07, 1.707637e-08, 
    3.155539e-09, 8.284453e-09, 7.113297e-07, 2.592802e-05, 4.993394e-05,
  3.747478e-05, 4.11073e-05, 4.023448e-05, 5.211886e-05, 6.287428e-05, 
    6.007999e-05, 3.804587e-05, 1.312904e-06, 3.612497e-09, 2.978472e-11, 
    2.738402e-10, 1.021892e-09, 2.515795e-06, 4.976883e-05, 4.656085e-05,
  2.222221e-05, 5.33415e-05, 4.751474e-05, 2.633038e-05, 4.980923e-05, 
    5.858104e-05, 8.089647e-05, 3.046507e-05, 7.644423e-09, 7.646619e-11, 
    9.247964e-11, 3.039833e-08, 9.8283e-08, 4.515413e-05, 2.027957e-05,
  2.022058e-05, 3.135971e-05, 5.279567e-05, 4.863464e-05, 7.016835e-05, 
    9.933609e-05, 0.0001132086, 7.702078e-05, 1.66828e-09, 3.246237e-10, 
    3.113478e-10, 2.875405e-10, 3.391892e-09, 7.820952e-06, 1.081447e-06,
  1.528857e-05, 2.849168e-05, 5.174898e-05, 6.783025e-05, 9.185798e-05, 
    9.405431e-05, 0.0001276786, 9.433074e-07, 2.321406e-06, 3.409e-07, 
    6.84769e-10, 7.043379e-10, 1.582032e-07, 1.109814e-06, 1.520423e-07,
  4.263055e-10, 6.506926e-10, 1.032961e-09, 3.462152e-11, 6.009452e-12, 
    5.109035e-12, 6.431365e-14, 2.046797e-12, 3.191681e-10, 4.200569e-08, 
    2.152314e-06, 4.660501e-05, 6.736217e-05, 4.949588e-05, 3.203789e-05,
  3.385629e-11, 1.825688e-11, 1.097396e-10, 2.400162e-11, 7.585904e-12, 
    1.283323e-09, 1.677323e-09, 1.044497e-09, 3.275138e-08, 2.684581e-06, 
    1.190962e-05, 4.971427e-05, 6.673852e-05, 4.694196e-05, 1.935167e-05,
  1.219665e-10, 1.179731e-10, 2.447423e-09, 7.863574e-11, 1.139512e-09, 
    6.204033e-08, 1.728998e-09, 7.986036e-09, 7.576907e-07, 2.086411e-05, 
    3.993194e-05, 0.0001013791, 0.0001339354, 8.107151e-05, 5.437406e-06,
  3.405848e-10, 2.582435e-10, 1.30213e-08, 3.483822e-07, 7.889398e-07, 
    1.944507e-06, 2.807354e-06, 2.458409e-07, 8.630611e-07, 1.580106e-05, 
    6.25433e-05, 0.0001180881, 0.0001423452, 8.184079e-05, 2.548689e-05,
  9.722565e-10, 5.364411e-10, 4.087591e-10, 1.754054e-09, 5.574278e-09, 
    2.692001e-07, 9.647241e-07, 3.888778e-07, 2.727346e-06, 1.2667e-05, 
    2.091912e-09, 6.446705e-09, 5.955929e-05, 4.268654e-05, 9.216847e-06,
  3.480691e-09, 6.598311e-09, 1.745369e-09, 7.835252e-09, 1.887459e-08, 
    4.450806e-08, 2.988149e-06, 3.888476e-06, 8.665312e-06, 3.680272e-11, 
    3.125509e-10, 3.6738e-10, 2.677438e-10, 4.133382e-06, 6.082523e-05,
  1.182965e-09, 1.554752e-08, 8.346504e-09, 3.88956e-08, 1.079903e-06, 
    2.845157e-07, 4.008353e-06, 8.850503e-07, 7.102803e-08, 1.107828e-12, 
    5.366165e-12, 7.686902e-13, 9.260024e-11, 8.083038e-08, 2.293705e-05,
  6.929732e-10, 7.034738e-07, 1.05154e-06, 2.963478e-08, 1.87976e-06, 
    1.301915e-05, 1.810332e-05, 2.790993e-05, 4.414397e-06, 2.405286e-11, 
    2.747227e-11, 1.113371e-11, 3.968018e-11, 7.519174e-06, 9.466102e-06,
  1.087265e-08, 7.737308e-06, 7.919148e-06, 1.434689e-05, 3.280764e-05, 
    5.72836e-05, 6.60453e-05, 0.000109021, 2.552993e-09, 3.571178e-10, 
    2.72556e-10, 1.443895e-10, 1.518211e-10, 1.211043e-05, 2.337741e-05,
  5.867338e-07, 4.154565e-06, 1.122445e-05, 1.58102e-05, 6.297487e-05, 
    0.0001031597, 0.0001004682, 4.022234e-08, 5.998947e-09, 2.700534e-09, 
    9.91498e-10, 4.137872e-10, 2.637388e-10, 1.165841e-05, 1.209093e-05,
  3.795335e-12, 7.979963e-12, 8.336133e-12, 7.653007e-12, 3.034857e-12, 
    3.677883e-13, 4.42332e-14, 1.818183e-11, 8.317651e-09, 3.474777e-08, 
    2.511241e-06, 2.022519e-05, 5.195385e-05, 7.531927e-05, 1.614392e-05,
  7.985347e-12, 4.30156e-12, 2.907433e-12, 2.236381e-12, 1.130422e-12, 
    6.010002e-13, 1.518801e-12, 6.975387e-12, 4.525282e-09, 3.847756e-08, 
    2.511121e-06, 2.194008e-05, 4.999799e-05, 7.051919e-05, 1.348652e-05,
  2.324109e-12, 3.130186e-13, 3.696779e-12, 3.260629e-10, 1.917973e-11, 
    1.382287e-10, 9.177e-11, 6.949766e-09, 3.080362e-08, 3.447819e-06, 
    2.61002e-05, 5.177481e-05, 0.000147752, 0.0001906761, 3.75644e-05,
  1.181184e-12, 6.114129e-13, 1.047296e-10, 1.307337e-09, 2.59816e-10, 
    8.830906e-09, 2.460456e-07, 2.336243e-06, 5.406053e-06, 3.511621e-05, 
    7.545208e-05, 9.645645e-05, 0.0002148537, 0.000227908, 0.0001019639,
  3.912111e-12, 1.170984e-11, 3.629004e-11, 8.60419e-10, 6.637892e-10, 
    1.951945e-08, 8.382455e-07, 8.141634e-06, 3.512158e-05, 6.417798e-05, 
    1.094851e-07, 9.055617e-09, 2.608145e-05, 8.263459e-05, 0.0001149703,
  1.476998e-11, 1.303238e-09, 4.072744e-09, 1.085399e-08, 3.026972e-09, 
    8.479785e-08, 4.176666e-06, 3.080803e-05, 2.815647e-05, 4.697866e-08, 
    3.105148e-07, 1.661609e-07, 4.744146e-07, 1.773564e-05, 0.000245858,
  3.000268e-11, 8.004616e-09, 8.239321e-09, 7.405557e-09, 1.69244e-08, 
    1.579612e-08, 2.640656e-06, 9.574423e-06, 1.918876e-05, 5.499086e-08, 
    2.328251e-10, 1.315864e-08, 1.224449e-07, 5.669893e-06, 0.0001283122,
  9.51477e-19, 2.997476e-12, 2.151643e-08, 7.663314e-09, 2.276077e-08, 
    8.589627e-07, 1.269625e-06, 3.254273e-05, 2.660718e-05, 2.546051e-09, 
    3.006839e-10, 3.103706e-10, 1.563975e-09, 1.644106e-06, 4.0646e-05,
  7.776634e-12, 2.152671e-09, 2.034289e-08, 1.972041e-07, 1.293596e-06, 
    4.843592e-06, 7.283855e-06, 2.740978e-05, 2.860844e-09, 6.50038e-10, 
    6.854356e-09, 2.124805e-10, 6.507026e-10, 6.69547e-07, 1.220347e-07,
  4.333472e-12, 4.026693e-11, 4.115062e-09, 2.002141e-07, 3.44147e-07, 
    4.026223e-06, 4.486884e-06, 1.983147e-07, 9.730002e-09, 3.237945e-09, 
    2.169513e-09, 1.517338e-09, 7.078138e-10, 3.753053e-07, 3.422295e-09,
  6.736112e-11, 6.094388e-11, 6.25635e-09, 5.807179e-09, 3.889703e-09, 
    1.568882e-09, 1.589669e-09, 1.403383e-09, 3.18309e-09, 1.513249e-08, 
    6.514418e-08, 4.37985e-06, 3.906674e-05, 4.354905e-05, 2.069575e-05,
  7.267111e-12, 4.766651e-11, 7.242213e-09, 1.564986e-08, 3.717046e-10, 
    4.562255e-10, 3.175511e-10, 1.59309e-10, 8.034664e-08, 4.672299e-06, 
    3.012596e-05, 7.14511e-05, 8.762305e-05, 7.944661e-05, 3.976661e-05,
  2.393356e-13, 1.065417e-10, 1.44064e-09, 5.197821e-10, 7.62836e-10, 
    1.92872e-08, 4.772557e-09, 4.606413e-07, 1.321808e-05, 5.151643e-05, 
    9.707242e-05, 0.0001581769, 0.0001560696, 0.0001404551, 3.837466e-05,
  3.010928e-17, 4.842993e-12, 1.398313e-09, 2.045714e-08, 7.436884e-09, 
    2.426762e-06, 3.263938e-06, 8.317266e-06, 3.429888e-05, 1.940078e-05, 
    0.0001195923, 0.0001053701, 5.915453e-05, 0.0001165215, 4.661691e-05,
  1.021055e-27, 6.370844e-21, 3.81494e-31, 1.720222e-14, 1.112522e-09, 
    1.647471e-07, 3.422213e-06, 8.949168e-06, 1.275328e-05, 4.010646e-05, 
    4.991917e-06, 1.553297e-06, 2.180205e-05, 6.002116e-05, 3.212444e-05,
  5.843328e-13, 5.501379e-11, 5.02657e-28, 2.717405e-12, 1.893065e-09, 
    1.172849e-07, 2.939315e-06, 6.691857e-06, 2.321973e-05, 1.147669e-07, 
    7.55007e-07, 1.564355e-06, 3.706173e-06, 1.110786e-05, 7.471351e-05,
  2.001684e-25, 5.475313e-12, 5.177416e-12, 5.782605e-11, 1.547804e-09, 
    2.672511e-08, 2.268081e-06, 2.328732e-06, 1.835023e-06, 1.020213e-10, 
    1.872374e-10, 9.832648e-09, 2.067222e-06, 8.574244e-06, 8.128773e-05,
  9.205302e-11, 2.848686e-09, 2.248181e-09, 4.813946e-12, 1.23237e-10, 
    4.24436e-08, 2.341831e-07, 4.099862e-06, 3.489824e-06, 1.594169e-10, 
    1.429304e-10, 2.793474e-10, 6.341987e-08, 2.378464e-05, 5.560655e-05,
  2.283686e-17, 1.059146e-15, 1.796594e-10, 1.033473e-11, 1.580973e-09, 
    2.008255e-09, 3.081244e-08, 1.772704e-07, 1.933254e-10, 3.651242e-15, 
    4.684723e-11, 5.784576e-12, 3.882819e-11, 2.320349e-05, 1.926766e-05,
  3.312165e-24, 1.147698e-25, 3.047046e-16, 1.368524e-11, 1.791086e-13, 
    6.40325e-21, 1.232743e-15, 6.153782e-11, 2.101426e-12, 8.764229e-21, 
    2.747259e-25, 3.199307e-24, 2.530549e-10, 5.536263e-06, 7.827185e-06,
  1.100109e-26, 3.056691e-14, 3.792614e-27, 2.435274e-25, 1.00826e-15, 
    4.703702e-13, 2.381785e-09, 1.661029e-08, 5.573575e-06, 1.212563e-05, 
    1.850675e-05, 4.93925e-05, 6.089411e-05, 2.26557e-05, 9.531234e-06,
  5.009908e-30, 9.446241e-28, 2.199125e-26, 4.086246e-25, 3.05711e-24, 
    1.153466e-11, 2.184015e-07, 1.209766e-05, 5.807679e-05, 0.0001037567, 
    0.000155959, 0.0001888986, 0.0001476302, 6.111799e-05, 3.504128e-05,
  8.381903e-18, 3.160909e-13, 2.147411e-13, 7.246453e-19, 9.241303e-13, 
    2.675068e-10, 7.544664e-09, 2.369001e-05, 6.894807e-05, 0.0001068502, 
    0.0002476397, 0.0003969482, 0.0003743272, 0.0001696869, 0.0001775945,
  3.298511e-11, 6.169951e-11, 8.512193e-11, 3.354077e-12, 3.493024e-11, 
    7.181252e-09, 1.096991e-07, 2.528463e-06, 1.556145e-05, 3.535343e-05, 
    0.0002805293, 0.0002422579, 0.000264582, 0.0001954523, 0.0001420895,
  2.747857e-09, 2.117392e-10, 2.081673e-09, 1.673148e-15, 1.718279e-12, 
    1.120665e-10, 3.050843e-08, 4.198999e-07, 2.49743e-06, 1.034385e-05, 
    2.59998e-07, 7.23505e-07, 0.0001644318, 0.000126497, 5.412302e-05,
  1.545294e-10, 9.047925e-11, 1.706063e-11, 1.854134e-10, 4.896791e-11, 
    3.004699e-12, 4.516852e-09, 1.901066e-07, 2.301953e-10, 1.263156e-09, 
    2.664232e-09, 4.513507e-09, 1.572524e-06, 3.464511e-05, 6.690656e-05,
  4.085283e-10, 2.253678e-09, 3.101928e-10, 1.242073e-09, 1.69322e-10, 
    2.151629e-10, 3.555003e-10, 4.348625e-10, 6.616977e-12, 6.146685e-11, 
    5.401483e-10, 1.00508e-09, 3.126409e-09, 5.122093e-05, 4.781574e-05,
  6.042132e-10, 2.540835e-09, 5.4908e-10, 3.934844e-10, 4.902836e-10, 
    1.172236e-08, 1.427084e-08, 8.383921e-10, 1.227551e-14, 5.99024e-13, 
    1.060909e-14, 5.791247e-11, 1.384856e-09, 5.19726e-05, 2.880053e-05,
  3.457872e-10, 1.71474e-10, 1.079928e-09, 1.817095e-10, 7.836845e-09, 
    6.823339e-09, 8.953976e-09, 1.99156e-10, 1.676769e-12, 3.856215e-23, 
    6.383576e-24, 1.877855e-11, 4.873836e-10, 7.159417e-06, 5.919795e-06,
  4.4187e-11, 9.022091e-11, 3.475822e-10, 1.822081e-09, 1.171374e-10, 
    2.694582e-10, 1.108552e-10, 1.881517e-11, 2.172558e-22, 1.090627e-22, 
    5.324559e-23, 6.614863e-16, 2.066964e-12, 5.186503e-08, 2.47474e-06,
  1.316198e-17, 2.476667e-24, 3.239826e-24, 1.917978e-24, 1.039176e-15, 
    3.395631e-14, 7.01592e-14, 6.871353e-11, 3.867853e-05, 5.472031e-05, 
    2.503976e-05, 4.644398e-05, 4.563001e-05, 4.44379e-05, 4.0682e-05,
  2.798725e-24, 1.273983e-14, 5.843587e-12, 3.19214e-11, 1.95065e-10, 
    1.078921e-09, 9.33155e-14, 1.457303e-09, 1.744296e-05, 5.39771e-05, 
    8.74573e-05, 0.0001282187, 7.202328e-05, 7.457532e-05, 4.33747e-05,
  4.080299e-14, 1.453982e-11, 2.222401e-10, 5.994102e-10, 8.424694e-10, 
    6.594506e-10, 2.29526e-11, 1.456403e-10, 9.922086e-07, 6.117547e-06, 
    3.197326e-05, 0.0002898317, 0.0004716108, 0.0003869609, 0.000157401,
  5.893986e-11, 1.845501e-10, 1.702427e-09, 4.662059e-10, 6.002734e-10, 
    1.016284e-08, 3.080234e-09, 1.593853e-09, 2.58123e-07, 7.173452e-06, 
    3.952597e-05, 9.640388e-05, 0.0004337089, 0.0005934973, 0.000299152,
  5.216856e-10, 1.639926e-09, 1.595974e-09, 1.244911e-09, 1.62668e-09, 
    2.338039e-08, 4.51168e-09, 9.089623e-10, 5.588305e-10, 8.084246e-07, 
    4.009934e-08, 1.158411e-07, 0.0002121001, 5.430634e-05, 4.626514e-05,
  1.573335e-09, 1.587463e-10, 6.650247e-11, 4.478412e-10, 1.984824e-09, 
    6.8769e-09, 2.144674e-09, 9.222155e-09, 8.13907e-09, 1.074965e-09, 
    3.878053e-09, 3.121436e-08, 2.206014e-05, 0.0001098122, 5.137482e-05,
  2.382254e-09, 1.368877e-09, 3.025888e-11, 6.191632e-11, 7.088202e-10, 
    9.36684e-09, 4.680459e-09, 1.09905e-08, 6.967219e-08, 1.172761e-09, 
    5.194391e-10, 4.791431e-09, 5.354359e-08, 9.704018e-05, 9.714944e-05,
  1.779018e-14, 1.423966e-12, 1.38189e-09, 3.938333e-10, 3.68325e-09, 
    3.334558e-08, 1.621769e-07, 3.698421e-07, 5.437936e-07, 2.4562e-09, 
    1.26471e-09, 1.3841e-09, 4.667615e-09, 5.334932e-05, 7.108897e-05,
  1.180578e-12, 3.556534e-12, 4.254708e-11, 7.061527e-09, 2.607532e-07, 
    1.042543e-07, 9.36771e-07, 1.422895e-06, 6.075273e-08, 7.442609e-09, 
    6.324477e-09, 4.178196e-09, 3.848164e-09, 6.582931e-06, 1.102727e-05,
  9.286263e-12, 1.72015e-10, 3.834663e-08, 4.140878e-10, 2.010639e-09, 
    7.779862e-08, 1.966243e-07, 2.504263e-09, 3.313664e-09, 5.87532e-09, 
    3.129626e-09, 4.555976e-09, 1.029676e-08, 1.88086e-08, 2.220922e-07,
  4.954569e-23, 6.791285e-13, 1.58792e-11, 3.662628e-12, 3.183438e-14, 
    1.941263e-13, 5.411054e-11, 3.707169e-11, 1.006398e-08, 8.511864e-06, 
    4.894169e-05, 7.812415e-05, 4.448559e-05, 6.858917e-05, 4.275967e-05,
  4.649208e-14, 4.908221e-23, 4.587443e-12, 2.449684e-12, 1.19105e-12, 
    1.897514e-12, 2.201588e-12, 3.343321e-10, 2.798113e-08, 3.357784e-06, 
    1.501712e-05, 3.003288e-05, 7.006763e-05, 9.447504e-05, 6.633958e-05,
  1.505894e-10, 1.164369e-10, 3.159305e-10, 6.23291e-13, 5.245327e-12, 
    2.829114e-11, 5.644019e-10, 4.641533e-09, 1.302756e-07, 3.12123e-06, 
    1.784848e-05, 2.047135e-05, 2.554896e-05, 6.36645e-05, 6.468446e-05,
  4.280851e-10, 1.936952e-10, 2.764761e-11, 3.709091e-11, 2.442573e-11, 
    2.694676e-08, 8.087576e-08, 3.265715e-07, 2.180999e-06, 2.303712e-05, 
    5.77421e-05, 5.957633e-05, 3.909772e-05, 8.57355e-05, 5.523936e-05,
  1.421826e-09, 2.213684e-10, 6.389228e-11, 4.723263e-11, 2.042852e-10, 
    3.840221e-08, 5.630241e-07, 4.650851e-06, 3.06813e-05, 9.187087e-05, 
    4.140684e-06, 3.214867e-06, 4.908376e-05, 3.498845e-05, 3.401139e-05,
  9.351189e-10, 1.84131e-10, 8.093694e-11, 3.30464e-11, 1.352662e-09, 
    6.578124e-07, 4.071812e-06, 1.381154e-05, 5.172201e-05, 3.966013e-06, 
    3.517353e-06, 1.290364e-06, 1.747051e-05, 9.860931e-05, 8.915678e-05,
  4.287309e-10, 3.308618e-10, 8.167657e-11, 2.460295e-11, 1.156158e-07, 
    5.410303e-08, 1.899593e-06, 4.019668e-06, 5.235996e-06, 3.069144e-07, 
    2.751574e-08, 9.53959e-09, 1.159505e-06, 7.290262e-05, 8.300713e-05,
  6.200604e-10, 8.221988e-11, 7.464448e-11, 2.63425e-10, 1.205968e-08, 
    4.251352e-07, 1.697907e-06, 6.574906e-06, 5.95235e-06, 1.708422e-09, 
    3.329871e-09, 1.073856e-08, 1.761423e-07, 3.572909e-05, 1.971753e-05,
  4.304039e-10, 9.563147e-11, 3.292698e-09, 1.430249e-08, 5.11776e-07, 
    3.643738e-06, 6.509129e-06, 9.644516e-06, 6.091693e-08, 5.482057e-10, 
    2.04931e-09, 7.581164e-09, 1.834714e-08, 1.378907e-05, 8.362004e-06,
  2.83605e-11, 1.688007e-09, 1.30942e-07, 3.463329e-08, 1.210323e-06, 
    5.592937e-06, 4.219953e-06, 1.264912e-08, 4.313774e-11, 8.169844e-11, 
    3.190356e-09, 6.949976e-09, 6.28872e-09, 2.213769e-06, 1.077062e-06,
  8.693668e-08, 4.01407e-08, 2.428901e-08, 9.942156e-09, 5.62471e-09, 
    5.398793e-09, 2.679917e-09, 1.365058e-09, 1.122155e-09, 2.86408e-06, 
    2.128927e-05, 6.964961e-05, 0.0001041564, 6.653164e-05, 3.263311e-05,
  6.912445e-08, 2.265464e-08, 8.398989e-09, 7.396516e-09, 9.389549e-09, 
    7.265577e-09, 2.587487e-09, 1.186741e-09, 2.567926e-08, 1.569852e-06, 
    6.767847e-06, 2.402559e-05, 3.695551e-05, 2.648884e-05, 5.844769e-07,
  6.686759e-08, 2.170425e-08, 1.47766e-08, 1.493032e-08, 6.815098e-08, 
    1.974146e-07, 2.017424e-07, 6.426193e-08, 2.443048e-08, 4.221943e-07, 
    5.299105e-06, 7.300678e-06, 2.827715e-06, 2.580416e-06, 2.441636e-08,
  4.837869e-08, 2.53875e-08, 2.605195e-08, 1.971363e-08, 2.122023e-07, 
    2.988196e-06, 3.297667e-06, 7.532508e-07, 1.019492e-06, 5.815084e-06, 
    1.526533e-05, 8.039872e-06, 2.18405e-06, 2.894909e-06, 3.775609e-07,
  1.289502e-08, 1.6789e-08, 6.912908e-09, 3.472451e-09, 2.223331e-08, 
    9.088786e-07, 3.071542e-06, 2.853214e-06, 1.438806e-05, 4.688022e-05, 
    5.867099e-06, 4.980237e-06, 1.098552e-05, 5.220816e-06, 3.763521e-06,
  1.0021e-08, 5.725413e-09, 8.52601e-10, 3.220338e-11, 6.197946e-11, 
    5.457139e-08, 7.812734e-07, 3.411317e-06, 1.118108e-05, 9.787422e-07, 
    1.951664e-07, 2.323587e-07, 1.947251e-06, 1.331149e-05, 9.374654e-06,
  1.797253e-09, 1.271535e-10, 2.180076e-11, 4.085879e-13, 5.907468e-10, 
    8.262132e-10, 9.734091e-07, 6.216377e-07, 3.752784e-07, 4.699567e-08, 
    2.716506e-08, 1.401344e-08, 1.608362e-08, 7.323577e-06, 2.273723e-06,
  2.528264e-09, 4.933224e-10, 5.817666e-12, 1.32487e-13, 4.899993e-10, 
    4.006158e-07, 9.025229e-08, 1.738917e-07, 1.457618e-07, 1.889719e-09, 
    1.376116e-08, 8.97804e-10, 3.552966e-10, 5.449216e-06, 1.256772e-06,
  7.507657e-10, 1.703023e-09, 4.299415e-11, 1.604505e-11, 3.511901e-10, 
    2.595892e-09, 1.047826e-07, 2.258034e-08, 6.386969e-12, 1.940687e-10, 
    2.990992e-09, 7.851643e-10, 1.563373e-09, 1.92131e-06, 3.120394e-07,
  2.934995e-10, 2.244217e-10, 1.470406e-10, 3.395212e-11, 2.074373e-10, 
    1.533923e-11, 1.633307e-11, 8.141952e-14, 1.731853e-11, 8.350226e-11, 
    1.612522e-11, 1.009819e-09, 3.227279e-07, 3.541046e-06, 1.375688e-07,
  5.294471e-07, 3.322646e-07, 2.93589e-07, 3.190987e-07, 2.681501e-07, 
    1.887274e-07, 1.43397e-07, 1.73839e-07, 1.974272e-07, 2.656286e-07, 
    2.294016e-07, 1.570257e-07, 6.14389e-06, 3.281864e-05, 1.478877e-06,
  4.002321e-07, 2.38254e-07, 2.447825e-07, 2.825781e-07, 2.213392e-07, 
    1.265697e-07, 8.680852e-08, 8.807641e-08, 7.728871e-08, 8.30596e-08, 
    9.619093e-07, 7.19742e-06, 2.868155e-05, 7.611199e-05, 3.621207e-05,
  2.841967e-07, 1.995111e-07, 1.300899e-07, 1.425237e-07, 6.951119e-07, 
    3.453665e-06, 3.796536e-08, 1.508864e-08, 2.333808e-08, 9.315153e-06, 
    1.752282e-05, 2.716104e-05, 4.922694e-05, 7.713047e-05, 8.545465e-05,
  2.095088e-07, 1.667542e-07, 3.137146e-07, 4.45707e-07, 2.655422e-06, 
    4.182346e-06, 1.1929e-06, 2.322731e-07, 8.174928e-07, 9.636414e-06, 
    3.155692e-05, 5.085107e-05, 1.240037e-05, 2.766418e-05, 8.446592e-06,
  5.998366e-08, 2.982846e-08, 2.840594e-08, 1.969661e-08, 1.359609e-08, 
    5.365138e-09, 1.363544e-06, 9.627216e-07, 4.520073e-06, 2.346716e-05, 
    2.023406e-07, 5.49327e-08, 9.759729e-06, 1.883668e-06, 2.064389e-05,
  9.786063e-09, 1.414085e-08, 1.055307e-09, 1.197921e-09, 4.770001e-10, 
    7.329436e-07, 2.555102e-06, 4.550211e-06, 1.607947e-05, 1.390869e-06, 
    6.300735e-09, 1.360934e-06, 1.393589e-06, 1.626615e-06, 5.834137e-06,
  1.039697e-08, 6.05839e-09, 1.372346e-09, 3.623952e-10, 1.627515e-07, 
    3.26529e-08, 2.446271e-06, 9.346326e-06, 2.865642e-05, 8.062383e-06, 
    2.49976e-06, 2.182122e-06, 1.054055e-05, 4.843134e-05, 1.246881e-05,
  5.49236e-09, 3.49038e-09, 3.183574e-08, 5.825058e-08, 5.626337e-08, 
    8.430866e-07, 7.565745e-06, 2.510331e-05, 6.277447e-05, 1.403683e-05, 
    2.198398e-06, 2.658889e-06, 5.447243e-06, 8.614395e-05, 4.63943e-05,
  1.597789e-09, 1.201608e-08, 7.5409e-07, 1.581986e-06, 4.293228e-06, 
    1.020859e-05, 2.39587e-05, 7.130259e-05, 1.847135e-05, 2.489359e-06, 
    1.238201e-06, 5.674527e-06, 1.657629e-05, 9.573624e-05, 6.326042e-05,
  1.433562e-09, 1.745232e-06, 5.188913e-06, 2.091083e-06, 9.848046e-06, 
    1.757786e-05, 2.775199e-05, 1.272397e-05, 1.243761e-06, 1.321096e-06, 
    3.250851e-06, 7.271613e-06, 1.63337e-05, 8.34976e-05, 4.341723e-05,
  7.078611e-09, 4.555794e-08, 1.229792e-07, 2.664804e-08, 1.812506e-08, 
    5.528896e-08, 3.261062e-08, 3.809682e-08, 1.516057e-08, 1.382568e-07, 
    2.748758e-06, 3.014393e-06, 2.143373e-05, 4.358103e-05, 6.694426e-07,
  2.468517e-11, 1.747354e-09, 5.211986e-08, 1.85613e-08, 2.615195e-08, 
    5.247138e-09, 3.500223e-09, 5.430917e-09, 7.992039e-09, 1.765184e-07, 
    1.671099e-06, 7.83436e-06, 2.67109e-05, 4.143881e-05, 6.967781e-12,
  9.163875e-09, 6.984608e-07, 1.563332e-08, 4.909243e-09, 5.073029e-08, 
    2.882701e-06, 1.738788e-09, 9.20354e-09, 1.396316e-06, 2.866863e-06, 
    1.935005e-05, 1.480681e-05, 3.549154e-05, 5.921024e-05, 1.157801e-10,
  2.120627e-06, 1.825046e-06, 1.666943e-06, 2.030295e-07, 3.399203e-07, 
    2.608971e-06, 6.435522e-07, 5.896524e-07, 1.572509e-06, 1.244367e-05, 
    3.161471e-05, 2.681101e-05, 7.889596e-06, 1.207007e-05, 2.387914e-08,
  2.130046e-07, 2.35927e-09, 1.129164e-10, 4.142838e-12, 1.163206e-10, 
    9.655042e-08, 1.522357e-06, 6.099775e-06, 2.260292e-05, 9.319049e-05, 
    1.18429e-05, 8.434458e-08, 4.177831e-06, 3.399858e-06, 1.597726e-06,
  6.923315e-09, 1.020563e-10, 3.375445e-10, 1.769602e-11, 7.809627e-10, 
    9.687616e-08, 2.909484e-06, 1.833139e-05, 6.025811e-05, 1.845223e-05, 
    3.725831e-06, 9.279611e-06, 7.548659e-06, 1.49626e-05, 1.737866e-05,
  3.215076e-09, 4.941799e-10, 1.71237e-09, 6.318256e-10, 4.023782e-07, 
    1.253605e-06, 9.959147e-06, 2.071649e-05, 2.246223e-05, 5.27238e-06, 
    5.860648e-07, 9.102283e-09, 2.714408e-06, 1.390989e-05, 1.017284e-05,
  4.758271e-12, 1.135279e-08, 2.647222e-07, 1.174839e-07, 4.032077e-07, 
    4.927203e-06, 8.598401e-06, 1.100398e-05, 4.311617e-06, 2.164527e-08, 
    2.310082e-07, 3.220204e-07, 2.979801e-07, 9.006287e-06, 6.642597e-07,
  1.132578e-09, 1.662427e-07, 2.348376e-06, 8.982542e-07, 5.470442e-07, 
    1.001871e-06, 1.573121e-06, 1.715778e-06, 1.70801e-08, 2.681104e-07, 
    4.795419e-07, 1.130903e-06, 2.911364e-06, 6.655634e-06, 7.987645e-07,
  6.355032e-10, 8.31809e-08, 1.116576e-06, 7.029611e-08, 4.145583e-07, 
    1.852123e-07, 5.667486e-08, 3.865595e-10, 3.516276e-09, 5.458228e-07, 
    7.287968e-07, 2.072772e-06, 4.057973e-06, 8.143304e-06, 1.341908e-05,
  2.140007e-14, 1.227383e-10, 3.223853e-07, 3.582287e-09, 7.350494e-14, 
    3.986027e-12, 8.998779e-11, 2.290776e-10, 3.470657e-10, 5.276307e-09, 
    1.069268e-07, 2.489104e-05, 8.579288e-05, 1.762909e-05, 2.062502e-07,
  4.932013e-11, 2.790239e-09, 1.619954e-09, 5.410433e-09, 7.078385e-09, 
    2.456092e-11, 2.350247e-10, 8.783336e-10, 3.99156e-09, 8.983886e-08, 
    4.546333e-06, 1.181793e-05, 5.465539e-05, 1.59016e-05, 3.062768e-08,
  1.472059e-09, 1.930343e-07, 3.096337e-10, 7.922816e-10, 2.252566e-08, 
    9.955116e-08, 7.222081e-08, 1.842469e-08, 1.175713e-07, 1.887157e-06, 
    5.239775e-06, 6.355875e-06, 5.784985e-06, 4.349743e-06, 3.091539e-08,
  2.229121e-08, 3.928735e-07, 3.249285e-09, 3.262274e-10, 7.657697e-08, 
    2.792544e-06, 2.552702e-06, 1.120626e-06, 4.229968e-06, 3.073978e-05, 
    7.230735e-05, 6.152242e-05, 2.011137e-05, 1.570388e-05, 9.12259e-08,
  4.682756e-06, 1.179827e-07, 3.815447e-10, 2.29997e-10, 3.831929e-09, 
    7.888565e-07, 6.191918e-06, 1.108886e-05, 4.157799e-05, 0.0001334345, 
    1.179826e-05, 1.757404e-06, 2.316036e-05, 8.276437e-06, 5.894631e-07,
  3.224685e-05, 9.665621e-07, 2.121551e-10, 3.574158e-10, 2.525129e-08, 
    1.16106e-06, 8.355658e-06, 1.668416e-05, 5.705006e-05, 5.372696e-06, 
    1.859825e-06, 2.413298e-06, 3.327021e-06, 1.285046e-05, 1.239109e-05,
  2.860001e-05, 1.176846e-06, 1.927117e-10, 4.22426e-09, 4.023427e-07, 
    5.900994e-07, 4.895639e-06, 7.019407e-06, 1.155428e-05, 1.484357e-06, 
    1.31506e-06, 2.498754e-06, 2.257052e-06, 2.133013e-05, 1.29e-05,
  1.273647e-08, 2.219859e-09, 1.026346e-11, 3.134789e-10, 3.416847e-09, 
    1.470137e-08, 9.916886e-07, 7.641684e-06, 8.060522e-06, 7.132969e-07, 
    7.566518e-07, 1.23757e-06, 1.17763e-06, 1.622399e-05, 1.014235e-05,
  7.447775e-11, 1.642144e-10, 2.465921e-15, 5.096457e-12, 1.77043e-10, 
    1.472583e-08, 1.913351e-06, 8.071543e-06, 1.78992e-07, 2.266232e-07, 
    1.186826e-07, 3.499267e-07, 3.521464e-07, 8.258467e-06, 7.543642e-06,
  9.731159e-12, 3.353586e-14, 5.094577e-17, 1.464693e-13, 1.017109e-11, 
    8.756228e-10, 6.925217e-07, 1.829632e-08, 6.659185e-09, 5.636105e-08, 
    2.553087e-17, 7.353744e-10, 3.868776e-09, 4.957649e-07, 2.278869e-06,
  4.622751e-13, 2.695586e-11, 1.644468e-11, 1.132515e-10, 1.844983e-10, 
    1.570658e-13, 2.095795e-12, 1.417032e-16, 1.490548e-11, 1.696022e-08, 
    1.010347e-07, 2.606194e-05, 3.548403e-05, 3.823488e-06, 4.003634e-07,
  4.576856e-12, 2.799129e-10, 2.221009e-13, 1.601054e-13, 1.498051e-11, 
    1.474338e-10, 1.991025e-10, 8.096714e-11, 5.301442e-09, 2.43469e-06, 
    1.448652e-05, 3.758689e-05, 3.935237e-05, 9.690407e-06, 1.850491e-06,
  7.052844e-09, 1.335849e-08, 3.522011e-09, 8.144584e-10, 9.308953e-07, 
    1.542307e-08, 7.325835e-09, 1.989692e-09, 3.176647e-08, 5.14661e-06, 
    1.370554e-05, 3.027106e-05, 5.224042e-05, 1.32678e-05, 1.992541e-08,
  2.742704e-06, 3.752571e-06, 5.454785e-06, 7.781964e-06, 9.045458e-06, 
    1.899335e-06, 5.164861e-07, 2.339455e-08, 4.212235e-07, 5.514103e-06, 
    5.64048e-06, 2.501859e-06, 1.33775e-07, 1.40064e-06, 1.641844e-08,
  1.09732e-06, 2.258477e-08, 7.385468e-09, 6.676777e-09, 4.565955e-09, 
    7.926965e-07, 3.511203e-06, 2.356581e-06, 1.252928e-05, 3.826373e-05, 
    1.679252e-07, 4.093653e-09, 4.541376e-10, 2.264677e-07, 6.594528e-08,
  1.884267e-08, 8.929265e-09, 2.682611e-09, 3.492683e-09, 4.010181e-08, 
    8.359642e-07, 2.766346e-06, 2.860191e-06, 6.159183e-06, 4.5295e-08, 
    2.80257e-10, 3.676012e-10, 5.874568e-08, 2.013259e-07, 1.341345e-07,
  7.331445e-09, 7.440074e-10, 1.011972e-09, 3.572161e-10, 3.871217e-08, 
    4.333291e-07, 2.802513e-06, 3.363407e-07, 2.278748e-07, 4.305473e-10, 
    1.984996e-12, 6.363049e-16, 1.075726e-09, 4.210372e-07, 2.686116e-07,
  1.660328e-09, 6.029699e-10, 5.433566e-10, 3.077506e-09, 9.290481e-10, 
    9.99511e-08, 3.751048e-07, 1.810918e-07, 3.388489e-08, 5.03969e-12, 
    5.322308e-27, 0, 1.060616e-12, 9.123909e-08, 1.143055e-08,
  6.255631e-11, 2.761648e-10, 3.384063e-10, 5.957503e-10, 3.785216e-11, 
    4.276616e-09, 2.827402e-08, 1.908668e-07, 8.418666e-10, 2.264253e-14, 0, 
    3.448609e-29, 1.493596e-11, 5.267881e-08, 1.408127e-07,
  6.180252e-10, 6.128582e-10, 4.737204e-10, 2.942974e-10, 1.479431e-10, 
    2.356201e-10, 7.189589e-10, 3.062586e-09, 9.880843e-13, 2.767634e-28, 0, 
    2.122946e-19, 2.449796e-10, 3.622717e-08, 4.442565e-09,
  3.347145e-15, 3.319433e-15, 6.500629e-12, 6.098038e-11, 4.634153e-10, 
    1.547893e-10, 8.575018e-11, 6.852333e-12, 2.71647e-11, 3.526552e-11, 
    7.968244e-10, 4.527062e-09, 9.427712e-07, 1.049573e-08, 2.326571e-09,
  3.611288e-26, 4.316472e-14, 5.329208e-16, 1.474598e-25, 1.700452e-11, 
    7.760463e-12, 7.418597e-14, 8.502353e-13, 8.103957e-13, 2.263017e-10, 
    3.558976e-08, 8.559897e-06, 1.049382e-05, 5.147428e-07, 2.270406e-09,
  3.173451e-14, 5.794493e-14, 3.748917e-15, 2.776416e-12, 1.017087e-10, 
    4.515768e-09, 9.226634e-11, 3.285153e-10, 7.328307e-11, 4.236558e-08, 
    1.441867e-05, 3.478479e-05, 4.099186e-05, 7.804475e-06, 3.063986e-10,
  1.778905e-12, 4.224956e-12, 2.67738e-12, 1.682391e-09, 4.33484e-08, 
    1.84801e-07, 3.359198e-08, 6.412242e-10, 1.206148e-08, 8.697273e-06, 
    2.29346e-05, 3.054285e-05, 5.026023e-05, 1.201358e-05, 3.132347e-10,
  4.540342e-12, 1.528362e-11, 2.04681e-11, 1.018721e-11, 3.403917e-13, 
    3.489135e-09, 4.143168e-11, 4.382056e-09, 1.724351e-07, 4.39013e-06, 
    7.15263e-08, 1.952138e-09, 4.529659e-06, 1.622177e-06, 2.213687e-06,
  5.843172e-11, 2.4981e-11, 3.711715e-11, 1.345956e-11, 5.87916e-14, 
    5.186573e-12, 1.03604e-11, 7.801174e-10, 4.621223e-08, 7.407474e-08, 
    1.069569e-10, 7.366267e-11, 1.241408e-09, 2.244475e-07, 1.871205e-05,
  5.024984e-09, 7.180659e-10, 2.42605e-11, 1.143592e-12, 7.213159e-13, 
    2.649119e-14, 5.268769e-15, 1.607142e-12, 3.936284e-11, 3.234342e-15, 
    4.105484e-26, 1.939789e-17, 1.829866e-11, 1.080509e-07, 1.768828e-05,
  4.312818e-09, 8.112815e-10, 1.426215e-10, 1.523821e-11, 4.165799e-12, 
    2.463266e-12, 2.205348e-12, 1.423891e-17, 3.284922e-26, 1.364511e-26, 
    1.5377e-27, 6.73814e-27, 1.525196e-26, 2.952853e-07, 8.104568e-08,
  5.863466e-10, 1.898885e-10, 4.880626e-09, 8.994928e-10, 1.228159e-11, 
    4.33492e-12, 2.793039e-11, 8.710168e-13, 7.028409e-26, 1.547793e-26, 
    7.240655e-33, 2.83613e-32, 9.043968e-29, 1.645732e-14, 8.118455e-12,
  5.639749e-10, 1.275513e-09, 8.75369e-09, 8.778683e-11, 7.048754e-11, 
    6.901014e-13, 2.114989e-10, 6.453651e-12, 2.240058e-25, 2.755519e-26, 
    7.538078e-28, 0, 0, 6.4044e-17, 1.496435e-16,
  2.103561e-10, 4.384533e-10, 1.351608e-09, 8.962371e-10, 8.491612e-10, 
    3.98646e-10, 1.096805e-10, 1.714327e-11, 3.09869e-11, 1.08497e-10, 
    2.303865e-09, 1.228429e-08, 4.255041e-07, 5.031141e-07, 5.546633e-10,
  2.158343e-11, 1.845118e-10, 8.668563e-10, 4.885265e-10, 2.856482e-10, 
    7.296505e-11, 1.834012e-25, 5.05907e-25, 2.350095e-13, 3.619619e-12, 
    9.173488e-11, 5.868542e-07, 2.079264e-06, 5.433163e-07, 2.636416e-10,
  3.15153e-13, 1.421586e-11, 2.79853e-11, 3.373272e-10, 5.561573e-11, 
    9.447766e-11, 8.244638e-12, 1.054922e-13, 1.057331e-16, 1.982059e-11, 
    6.469213e-08, 8.103372e-07, 3.036728e-06, 5.51592e-06, 1.512136e-11,
  2.894967e-11, 3.729492e-09, 3.265004e-10, 4.555101e-10, 6.020051e-08, 
    7.9045e-07, 3.903825e-10, 1.671768e-09, 8.527755e-11, 2.247869e-07, 
    3.346224e-07, 4.618476e-07, 5.674185e-06, 1.002981e-05, 2.343067e-09,
  3.920269e-09, 2.048501e-09, 5.2479e-10, 4.656404e-11, 5.482634e-11, 
    1.218183e-09, 1.525685e-08, 1.117387e-08, 5.703435e-09, 1.781289e-07, 
    3.111802e-12, 1.320652e-10, 2.064171e-06, 7.499271e-07, 9.323317e-06,
  4.282854e-09, 3.575459e-09, 2.134463e-09, 7.159448e-11, 6.927788e-10, 
    7.744487e-10, 6.559787e-10, 3.384797e-09, 4.632519e-10, 4.142525e-10, 
    2.733655e-13, 6.001808e-11, 3.203995e-10, 2.663026e-08, 5.631599e-06,
  1.896377e-06, 3.254071e-07, 2.930813e-07, 3.24671e-09, 1.274533e-09, 
    2.955375e-09, 6.717576e-09, 1.306778e-09, 3.788641e-09, 9.544638e-12, 
    1.000204e-22, 9.331937e-23, 4.796724e-11, 1.723557e-09, 1.21711e-05,
  5.869078e-10, 4.96665e-09, 1.301219e-06, 1.778453e-06, 2.255582e-06, 
    1.805566e-06, 3.634202e-06, 2.000046e-09, 1.007522e-10, 4.39241e-10, 
    4.959858e-10, 8.494887e-15, 1.326639e-09, 4.253907e-08, 6.642737e-06,
  5.444152e-10, 4.424106e-09, 5.92674e-06, 1.047088e-05, 1.183598e-05, 
    2.359784e-05, 1.828751e-05, 6.390364e-07, 4.798733e-10, 1.866609e-09, 
    2.362918e-09, 9.517058e-10, 5.691029e-10, 1.515948e-06, 9.487968e-09,
  7.524085e-10, 1.988847e-09, 8.457273e-07, 2.21508e-06, 7.971524e-06, 
    2.067819e-06, 5.967909e-08, 1.539967e-09, 2.407436e-09, 5.584148e-09, 
    4.820798e-09, 7.861279e-10, 5.710404e-10, 3.08098e-10, 2.207267e-10,
  3.564946e-25, 3.044225e-25, 2.250963e-12, 6.322966e-12, 2.681247e-13, 
    1.488991e-11, 1.89362e-12, 2.254034e-11, 2.22766e-11, 3.687482e-11, 
    5.241794e-11, 1.827096e-07, 4.629964e-06, 6.928636e-07, 3.476383e-11,
  5.165464e-26, 6.173746e-26, 5.691812e-26, 4.77689e-13, 5.309178e-13, 
    1.047682e-12, 2.073238e-12, 3.323126e-10, 2.572371e-11, 5.566977e-10, 
    2.598902e-08, 5.003796e-06, 2.119889e-05, 8.101282e-06, 5.381701e-08,
  1.319669e-16, 2.528558e-15, 3.090623e-12, 8.745346e-10, 7.171598e-11, 
    8.823556e-12, 3.434031e-11, 6.573777e-07, 4.718222e-06, 9.638434e-06, 
    3.265225e-05, 5.544756e-05, 7.580568e-05, 2.841163e-05, 1.312354e-07,
  8.179084e-11, 2.37881e-11, 1.670171e-07, 6.796536e-06, 3.495658e-07, 
    5.002375e-06, 1.096815e-05, 4.290183e-05, 4.099185e-05, 3.852727e-05, 
    2.538198e-05, 2.971664e-05, 6.35294e-05, 5.154067e-05, 1.119214e-08,
  1.616766e-08, 1.289947e-09, 9.844856e-07, 2.238228e-06, 1.631196e-06, 
    5.457769e-06, 1.751656e-05, 6.157428e-05, 4.80205e-05, 7.925242e-06, 
    1.39262e-09, 2.757175e-11, 2.390683e-06, 2.440383e-06, 6.559915e-07,
  4.466731e-10, 5.977494e-07, 8.101632e-07, 1.08374e-08, 2.925506e-09, 
    4.978427e-07, 1.893435e-05, 4.73563e-06, 3.431232e-06, 6.488541e-10, 
    6.577123e-10, 4.023751e-10, 1.230062e-10, 3.208454e-07, 6.007638e-06,
  2.452458e-09, 2.027749e-07, 1.485386e-06, 3.551841e-07, 1.347474e-09, 
    3.56377e-10, 1.038807e-09, 2.485837e-09, 1.793098e-08, 3.003019e-10, 
    1.350798e-08, 6.945904e-09, 3.28333e-09, 1.447693e-09, 1.861167e-05,
  2.942226e-10, 2.329934e-07, 9.958398e-06, 9.328235e-06, 1.103891e-05, 
    5.248934e-06, 2.178464e-06, 1.113302e-08, 5.714147e-10, 1.721034e-09, 
    2.695308e-09, 4.520998e-09, 1.229803e-08, 4.688046e-06, 1.421677e-05,
  1.829651e-13, 7.387827e-09, 8.526849e-06, 1.991479e-05, 3.765968e-05, 
    5.808404e-05, 3.428751e-05, 2.65932e-07, 2.014104e-09, 8.182359e-10, 
    3.678978e-09, 8.600695e-09, 1.043587e-08, 2.441623e-06, 7.007982e-09,
  2.37746e-12, 1.060896e-11, 3.17314e-10, 1.509977e-08, 2.769082e-06, 
    7.03567e-06, 2.963444e-06, 1.262889e-09, 2.823947e-09, 3.52393e-09, 
    2.752192e-09, 5.916017e-09, 2.388615e-08, 4.617002e-09, 5.669258e-09,
  9.61832e-28, 4.977441e-27, 5.595328e-26, 1.291873e-13, 7.879465e-13, 
    4.334672e-12, 2.144756e-13, 1.269888e-12, 3.701087e-11, 2.146263e-09, 
    1.163075e-09, 1.521615e-06, 2.639651e-06, 6.620321e-07, 4.045186e-10,
  2.20034e-27, 2.063177e-26, 6.193652e-17, 4.83398e-12, 7.223233e-11, 
    1.237383e-10, 9.851398e-14, 2.787063e-09, 9.950389e-09, 1.251204e-08, 
    6.272306e-07, 6.156895e-06, 1.221183e-05, 1.026191e-05, 7.712069e-09,
  7.422979e-18, 3.27237e-15, 8.537673e-10, 8.442232e-09, 1.033329e-06, 
    3.512518e-06, 5.479117e-08, 1.580727e-06, 6.246071e-06, 1.393833e-05, 
    4.615288e-05, 9.009321e-05, 0.0001379193, 8.802087e-05, 4.329557e-08,
  7.430126e-13, 3.025804e-10, 6.305794e-10, 5.365778e-09, 1.055921e-06, 
    5.530364e-06, 1.265277e-05, 2.721595e-05, 1.584277e-05, 4.912135e-05, 
    4.910902e-05, 5.17052e-05, 0.0001726327, 0.0001336785, 5.005222e-07,
  2.336426e-11, 9.571609e-10, 1.009931e-07, 7.812284e-09, 1.349917e-08, 
    3.83841e-07, 7.05225e-06, 2.189613e-05, 2.499702e-05, 2.995583e-05, 
    3.853764e-09, 8.917755e-09, 9.785605e-06, 3.119364e-05, 3.289762e-05,
  7.93998e-08, 1.034511e-06, 1.345922e-06, 5.059727e-07, 1.473753e-08, 
    2.007839e-07, 6.110725e-06, 2.862955e-06, 3.055113e-06, 7.917292e-10, 
    8.175956e-09, 2.916999e-09, 2.562669e-08, 2.864105e-06, 7.583937e-05,
  1.757662e-06, 2.173262e-06, 3.798631e-06, 8.604064e-06, 4.024499e-06, 
    1.319228e-06, 4.395937e-08, 1.19036e-08, 1.131316e-08, 3.985635e-09, 
    5.260178e-09, 3.397777e-09, 8.829152e-10, 7.044883e-07, 5.143695e-05,
  1.21825e-09, 2.042255e-07, 3.516e-06, 1.342708e-05, 2.601198e-05, 
    3.418823e-06, 5.068748e-06, 7.596014e-09, 4.934656e-09, 1.893287e-09, 
    9.485716e-09, 3.114449e-09, 1.041085e-09, 1.484323e-05, 1.458628e-05,
  2.314226e-11, 5.375519e-10, 1.105676e-06, 2.429891e-05, 2.540874e-05, 
    3.506579e-05, 2.615419e-05, 2.400711e-09, 2.904149e-09, 1.272096e-09, 
    2.683222e-09, 1.852648e-09, 9.854556e-10, 2.67467e-06, 1.219144e-08,
  5.689454e-14, 6.711888e-15, 2.548464e-10, 5.525881e-09, 1.520844e-06, 
    3.846494e-06, 2.555402e-08, 5.122775e-09, 1.606316e-09, 3.919279e-10, 
    1.619215e-09, 2.075345e-09, 2.756366e-10, 6.113257e-10, 1.51584e-09,
  1.11404e-11, 1.198523e-10, 6.599798e-11, 1.318929e-10, 1.87729e-11, 
    3.353225e-10, 6.05118e-10, 1.23857e-09, 5.746845e-07, 1.049517e-08, 
    9.338819e-07, 9.771272e-06, 6.934667e-06, 6.375106e-06, 1.586378e-08,
  9.946203e-13, 5.016075e-10, 4.412399e-08, 1.283946e-08, 4.811731e-09, 
    1.267879e-09, 4.446321e-06, 6.214758e-06, 6.018054e-06, 9.481424e-06, 
    9.01245e-06, 3.627695e-05, 0.0001332117, 0.0001329748, 2.747772e-06,
  1.105449e-10, 2.156004e-08, 1.254185e-08, 2.30491e-05, 8.577151e-05, 
    5.594046e-05, 5.191254e-05, 3.82541e-05, 3.700362e-05, 2.488329e-05, 
    4.263677e-05, 6.593118e-05, 8.961043e-05, 0.0001805167, 1.96026e-05,
  4.232237e-10, 4.127644e-09, 2.270183e-07, 2.152934e-05, 4.03275e-05, 
    8.579312e-05, 0.0001102865, 6.70419e-05, 2.93709e-05, 1.861338e-05, 
    4.059285e-05, 3.922437e-05, 3.513046e-05, 0.0001301377, 3.7878e-05,
  1.65463e-07, 3.701077e-06, 1.840192e-05, 5.395023e-05, 4.958992e-05, 
    7.062019e-05, 9.722137e-05, 4.274406e-05, 1.589002e-05, 2.212215e-05, 
    1.981112e-08, 1.672668e-08, 3.288133e-05, 2.776907e-05, 3.549757e-05,
  1.247691e-05, 1.634706e-05, 6.27245e-05, 3.408813e-05, 2.549759e-05, 
    5.708384e-05, 6.732201e-05, 5.405805e-06, 1.102527e-06, 3.875587e-09, 
    1.827972e-09, 5.368249e-09, 1.255934e-08, 3.723997e-05, 0.0001174912,
  4.583668e-05, 5.835532e-05, 0.000140168, 7.331397e-05, 5.483251e-05, 
    4.426052e-05, 5.109913e-05, 8.1677e-07, 3.649342e-09, 2.005534e-09, 
    1.573691e-09, 1.999682e-09, 3.905048e-09, 2.887103e-05, 0.0001067724,
  1.068086e-05, 5.60669e-05, 0.000115196, 0.0001281376, 7.691334e-05, 
    7.202801e-05, 5.41448e-05, 2.192552e-06, 7.034813e-09, 2.523145e-09, 
    2.108284e-09, 1.556419e-09, 1.916926e-09, 2.314452e-05, 3.641516e-05,
  5.998576e-09, 2.201964e-05, 4.895372e-05, 8.166653e-05, 6.584293e-05, 
    5.378679e-05, 1.386095e-05, 5.829811e-06, 1.033589e-08, 3.434124e-09, 
    2.762018e-09, 2.725917e-09, 2.35359e-09, 1.215493e-08, 9.24638e-09,
  3.171355e-09, 6.4553e-07, 1.385842e-05, 1.886227e-05, 2.754878e-05, 
    7.721595e-06, 1.909026e-07, 8.974659e-09, 6.867319e-09, 7.273019e-09, 
    1.180595e-08, 4.834869e-09, 1.147566e-08, 7.193914e-09, 8.027797e-09 ;

 sftlf =
  0.0008770345, 0.4596241, 0.9892928, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.01035247, 0.004304647, 0.6546783, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.8534847, 0.8118016, 0.9951549, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1,
  0.9894952, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0.4452189, 0.3028796, 0.7140614, 1, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.9903189, 0.3150955, 0.0007410151, 0, 0.02645395, 
    0.9012984, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.681631, 0, 0, 0, 0.004980796, 0.7708192, 1,
  1, 1, 1, 1, 1, 1, 1, 1, 0.5536854, 0, 0, 0, 0.004666397, 0.9395298, 1,
  1, 1, 1, 1, 1, 1, 1, 0.9995009, 0.3626226, 0, 0, 0, 0, 0.8367797, 1,
  1, 1, 1, 1, 1, 0.8451425, 0.7016711, 0.3953246, 0, 0, 0, 0, 0.006316811, 
    0.8673657, 1 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0.2038203, 25.08469, 362.922, 581.3585, 583.7158, 677.0037, 892.3406, 
    840.3151, 1394.918, 1845.667, 2078.668, 2048.803, 1746.472, 1895.031, 
    903.5963,
  0.04938461, 3.284697, 202.5217, 654.3141, 903.2668, 1076.606, 1196.302, 
    1163.293, 1639.916, 1906.256, 1988.945, 1916.741, 1695.228, 1807.269, 
    774.2457,
  790.1076, 1114.346, 653.3495, 780.126, 1392.106, 1491.591, 1273.753, 
    1344.373, 1825.463, 2046.944, 2142.644, 2067.535, 1930.862, 1770.506, 
    591.146,
  1359.809, 1341.669, 1435.043, 1594.124, 1615.893, 1763.274, 1677.539, 
    1645.991, 1875.931, 2003.645, 2040.039, 1879.801, 1919.839, 1717.029, 
    1138.974,
  1205.389, 1290.31, 1192.454, 1271.409, 1283.839, 1439.06, 1538.882, 
    1587.552, 1685.139, 1482.705, 108.3495, 67.86669, 940.4369, 898.4109, 
    1612.947,
  1168.617, 1342.769, 1106.133, 1029.211, 1110.353, 1151.071, 1218.088, 
    1182.275, 1031.226, 58.02261, 0, 0, 7.641389, 710.6758, 2161.482,
  1244.873, 1316.863, 1112.963, 998.5415, 1017.03, 1014.576, 1020.14, 
    838.6226, 484.287, 0, 0, 0, 0, 1273.715, 2180.106,
  896.0552, 1198.27, 1151.006, 981.8504, 1010.922, 1103.887, 1045.003, 
    880.1057, 498.0692, 0, 0, 0, 0, 1386.297, 1186.975,
  625.923, 1015.673, 1096.604, 994.0698, 1069.039, 1288.357, 1166.806, 
    927.0013, 34.64387, 0, 0, 0, 0, 678.2806, 439.0615,
  346.5426, 755.811, 896.7624, 677.1516, 656.058, 642.5463, 557.833, 
    41.91994, 0, 0, 0, 0, 0, 191.3587, 93.07086 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
