netcdf atmos_daily.00010101-00010701.ps.tile5 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float ps(time, grid_yt, grid_xt) ;
		ps:_FillValue = 1.e+20f ;
		ps:missing_value = 1.e+20f ;
		ps:units = "Pa" ;
		ps:long_name = "Surface Air Pressure" ;
		ps:cell_methods = "time: mean" ;
		ps:cell_measures = "area: area" ;
		ps:time_avg_info = "average_T1,average_T2,average_DT" ;
		ps:standard_name = "surface_air_pressure" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:07 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile5.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile5.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 ps =
  101521.8, 101399.9, 101303.7, 101201.7, 101124.1, 101047, 100976.4, 
    100929.4, 100926.2, 100938.1, 100960.8, 100985, 101004.7, 101022.2, 
    101046.4,
  101744.7, 101621.1, 101529.4, 101423.5, 101336.7, 101258.5, 101202.7, 
    101161.3, 101123.4, 101093.9, 101073.3, 101071.7, 101082.5, 101093.4, 
    101111.7,
  101941.7, 101823.5, 101732.9, 101633.7, 101547.1, 101460.5, 101383.3, 
    101315.8, 101268.2, 101234.2, 101216.1, 101199.9, 101192.6, 101188.6, 
    101188.9,
  102112, 102008.3, 101920.9, 101827.6, 101742.7, 101658.9, 101586.7, 
    101517.5, 101452.9, 101397, 101352.3, 101319.4, 101298.3, 101285.3, 
    101278.1,
  102267.6, 102173.3, 102085, 101997.2, 101914.9, 101831.6, 101755.5, 101682, 
    101621.1, 101564.5, 101514.2, 101468.6, 101430.2, 101399.9, 101378.7,
  102411.3, 102316.8, 102231.9, 102145.8, 102066.3, 101990.2, 101919.2, 
    101849.1, 101779.2, 101717.2, 101659.2, 101608.2, 101563.2, 101525.9, 
    101493.7,
  102546.1, 102450.9, 102365.6, 102278.9, 102198.4, 102122, 102051.5, 
    101986.5, 101921.2, 101857, 101799.5, 101742.3, 101691.6, 101644.1, 
    101603.9,
  102665.9, 102568.7, 102486.9, 102400.9, 102320.7, 102242.5, 102169.6, 
    102104.6, 102043.7, 101983.3, 101923.4, 101862.2, 101807.8, 101756.8, 
    101712,
  102765.3, 102671, 102590.1, 102504.3, 102427.4, 102350.6, 102276.4, 
    102203.4, 102140.8, 102082.3, 102027.8, 101971.4, 101915, 101857.3, 
    101806.8,
  102840.9, 102755.9, 102672.7, 102592.3, 102513.8, 102438.4, 102368.5, 
    102298.5, 102230.7, 102165.1, 102109.4, 102055, 102003.4, 101947.4, 
    101893.3,
  101974.9, 101830.8, 101693, 101542.4, 101395.2, 101227.3, 101115.4, 
    101031.4, 101081.8, 101064.5, 101013.1, 101013.2, 101051.6, 101085.8, 
    101110.7,
  102136, 101998.8, 101871.9, 101731.1, 101602.6, 101471.7, 101352.3, 
    101216.6, 101116.3, 101072.2, 101086.2, 101083.6, 101079.4, 101085.4, 
    101104.6,
  102291.4, 102162.4, 102043.6, 101905.1, 101770.4, 101627.7, 101494.4, 
    101382, 101271.6, 101179.1, 101108.7, 101076, 101070.2, 101087.4, 101116.7,
  102424.8, 102305.8, 102201.3, 102081, 101958.3, 101829.6, 101691, 101557.4, 
    101449.4, 101361.6, 101281.2, 101218.6, 101178.3, 101151, 101140.6,
  102551, 102440.5, 102330.5, 102222.8, 102112.5, 101994.6, 101873.8, 
    101735.2, 101606.8, 101518, 101445.5, 101360.6, 101306.6, 101251, 101233.8,
  102658.5, 102558.3, 102451.6, 102350, 102247.3, 102141.5, 102038, 101930.7, 
    101816.1, 101708.4, 101620.2, 101522.5, 101431.2, 101347.8, 101297.7,
  102759.2, 102657.4, 102555.9, 102457.7, 102357.5, 102264.3, 102162.5, 
    102063.8, 101965.4, 101854.9, 101753.8, 101672, 101573.9, 101486.1, 
    101417.8,
  102846.6, 102745.3, 102646.2, 102550.8, 102455.4, 102362.7, 102272.8, 
    102185.5, 102099.1, 102009.5, 101904.8, 101792.5, 101689, 101586.5, 
    101513.5,
  102917.5, 102819.9, 102722.9, 102627.7, 102536.1, 102450, 102358.6, 
    102272.6, 102188.2, 102110.6, 102025.4, 101935.4, 101844.3, 101746, 
    101660.4,
  102975.5, 102880.2, 102786.3, 102693, 102602.8, 102519.6, 102437.9, 
    102356.7, 102278.5, 102201.3, 102125.6, 102042.4, 101959.2, 101878.2, 
    101794.5,
  101901.9, 101755.2, 101618.6, 101469.5, 101337.2, 101216.8, 101145.4, 
    101129.2, 101142.3, 101131.8, 101145.3, 101162.5, 101178.7, 101191.9, 
    101186.4,
  102041.9, 101903.6, 101778.4, 101639.5, 101492.5, 101361.8, 101250.5, 
    101178.1, 101147.1, 101159, 101173, 101179.5, 101191.4, 101197.1, 101204.9,
  102170.3, 102036.7, 101906.9, 101764.6, 101628.3, 101492.2, 101376.6, 
    101275.6, 101211.2, 101172.3, 101173.4, 101183.7, 101201.1, 101221.4, 
    101230.5,
  102286.4, 102166.1, 102046, 101916.1, 101777.3, 101638.3, 101509.1, 
    101380.7, 101285.1, 101228.9, 101185.8, 101185.2, 101210.3, 101221, 
    101222.4,
  102396.5, 102281.4, 102164.6, 102043.9, 101919.1, 101790, 101654.6, 
    101518.1, 101402.9, 101322, 101260.5, 101212.2, 101202.5, 101211.3, 
    101234.2,
  102495.1, 102389.2, 102276.7, 102167.7, 102049.5, 101935.2, 101818.4, 
    101697, 101586.6, 101453.8, 101344.8, 101280.2, 101258.3, 101254.1, 
    101267.2,
  102581.9, 102479.9, 102378.7, 102272.9, 102167.2, 102060.3, 101953.2, 
    101834.8, 101706.3, 101591.8, 101482.5, 101376.1, 101317.6, 101298.9, 
    101303.7,
  102658, 102555.7, 102467.9, 102365.1, 102268.3, 102167.3, 102072.9, 
    101976.3, 101863.6, 101727.1, 101609.3, 101514.2, 101442.6, 101406.6, 
    101383.3,
  102718.8, 102621.3, 102538, 102447.9, 102355.8, 102260.4, 102170.3, 
    102070.5, 101975.9, 101875.3, 101757.1, 101656.9, 101575.5, 101526.4, 
    101499.1,
  102766.2, 102671.8, 102591.3, 102509.5, 102431.4, 102340.3, 102259.8, 
    102176, 102084.1, 101983.9, 101888.5, 101795.8, 101717, 101664.6, 101616.2,
  101349.5, 101229, 101117, 101028.3, 100964.8, 100924, 100886.8, 100883.7, 
    100881.1, 100886, 100894.3, 100907.1, 100917.2, 100939.6, 100956.3,
  101484.5, 101381.4, 101276.6, 101164.2, 101057.7, 101003.1, 100985.3, 
    100963.5, 100955.3, 100964.5, 100967.5, 100972.9, 100981.2, 100992.6, 
    101008.2,
  101599.9, 101497.7, 101396.8, 101296.4, 101194.3, 101081.3, 101033.8, 
    101024.9, 101017.3, 101020.7, 101026.9, 101038.5, 101044.1, 101055.1, 
    101064.1,
  101727.6, 101617.5, 101506.9, 101408.5, 101303.3, 101184.7, 101081.3, 
    101059.1, 101064.6, 101072.8, 101073.4, 101088.1, 101095.9, 101105.7, 
    101114.8,
  101842.6, 101725.5, 101615.7, 101518.8, 101413.3, 101288.5, 101158.4, 
    101091.2, 101080.2, 101098.7, 101104.6, 101123.8, 101136.2, 101147.3, 
    101151.8,
  101948.6, 101830.1, 101720.9, 101623.3, 101528.6, 101413.8, 101256.2, 
    101132.4, 101102.1, 101108.5, 101128.8, 101151.1, 101167.6, 101176.8, 
    101180.7,
  102044.9, 101928.1, 101819.3, 101713.3, 101627.5, 101532.3, 101387.4, 
    101228.7, 101146.5, 101122.7, 101135.8, 101156.8, 101174.4, 101187.3, 
    101204.2,
  102124.9, 102012.1, 101912.5, 101804.6, 101714.5, 101623.7, 101513.8, 
    101359, 101235.8, 101168.4, 101160.1, 101167.6, 101197.9, 101213.2, 
    101234.5,
  102188, 102088, 101993.3, 101887, 101794, 101710.9, 101607.3, 101473.5, 
    101327.7, 101232.5, 101202.8, 101175.6, 101203.3, 101211.1, 101262.8,
  102233.5, 102148.3, 102063.3, 101962.9, 101874.3, 101795.4, 101709.8, 
    101587.4, 101447.7, 101316.1, 101253.9, 101222.7, 101233.7, 101257, 
    101307.8,
  100321.4, 100312, 100310.2, 100320.1, 100340.7, 100371.2, 100418.4, 
    100475.1, 100525.3, 100579.8, 100632, 100688.9, 100743.7, 100780, 100823.6,
  100420.4, 100398.1, 100390.2, 100394.5, 100412.5, 100437.9, 100470.4, 
    100515.2, 100569, 100626.3, 100676.5, 100728.8, 100773.8, 100818.2, 
    100867.7,
  100524.2, 100486.4, 100462.1, 100449, 100450.9, 100468.7, 100502.2, 
    100547.8, 100603, 100657.2, 100706.5, 100757.6, 100804.1, 100853.4, 
    100900.1,
  100639.9, 100584.2, 100549, 100524.8, 100516.2, 100521, 100548.8, 100592.4, 
    100643.7, 100694.4, 100742.4, 100795, 100839.4, 100884.4, 100937.8,
  100760, 100700.1, 100643.5, 100603.8, 100581.3, 100574.2, 100591, 100630.4, 
    100679.3, 100729.7, 100778.9, 100831.8, 100874, 100918.5, 100964.8,
  100882.9, 100815.9, 100751.6, 100704.9, 100661.7, 100638.6, 100639.8, 
    100667.8, 100713.2, 100765.1, 100815.2, 100870, 100910.4, 100956.5, 
    100999.8,
  101000.2, 100933.9, 100858.1, 100804.9, 100754.2, 100716.4, 100700, 
    100704.6, 100744.8, 100793.3, 100843.9, 100897.3, 100942.3, 100994, 
    101038.8,
  101088.9, 101033.2, 100964.8, 100906.5, 100850.5, 100801.1, 100759.4, 
    100747.5, 100777.2, 100816.4, 100866.5, 100916.3, 100969.1, 101025.1, 
    101074,
  101165.6, 101109.5, 101053.3, 100994.7, 100949.1, 100891.3, 100834.6, 
    100793.4, 100797.5, 100835.4, 100886.4, 100934.6, 100990.7, 101051, 
    101103.6,
  101213.2, 101171.4, 101121.2, 101074, 101023.9, 100982.5, 100919, 100861.7, 
    100827.3, 100855.3, 100896.1, 100944, 101006.6, 101066, 101125.7,
  99621.78, 99614.84, 99642.65, 99678.5, 99723.67, 99785.69, 99864.3, 
    99950.99, 100049.5, 100142.4, 100229.4, 100313.9, 100397.4, 100480.3, 
    100559.8,
  99740.27, 99733.27, 99768.73, 99796.49, 99843.06, 99894.59, 99963.13, 
    100044.2, 100136.1, 100222.7, 100303.8, 100379.6, 100460.3, 100540.5, 
    100619,
  99819.14, 99814.03, 99851.73, 99883.59, 99939.66, 99993.05, 100063.8, 
    100140.5, 100224.9, 100307.5, 100386.1, 100460.5, 100534.1, 100605.6, 
    100679.1,
  99897.23, 99894.93, 99934.61, 99971.49, 100030.4, 100080.9, 100150.7, 
    100224.1, 100304.8, 100384.7, 100463.2, 100533.6, 100601.9, 100670, 
    100741.6,
  99952.72, 99950.85, 99999.04, 100042.4, 100100.7, 100155.7, 100225, 100299, 
    100376.5, 100458.1, 100535.5, 100610.4, 100676, 100739.3, 100804.6,
  99995.22, 99985.03, 100045.1, 100092.4, 100155.1, 100215.1, 100286.2, 
    100361.4, 100442.7, 100521.2, 100600.7, 100673.2, 100739.5, 100803.2, 
    100866.7,
  100020.9, 100017.9, 100068.2, 100121.2, 100192, 100257.6, 100332.4, 
    100412.2, 100497.2, 100577.3, 100655.1, 100728.8, 100795.8, 100863.1, 
    100929.9,
  100030.7, 100052.2, 100069.8, 100138.6, 100210.1, 100283.3, 100364.6, 
    100448, 100537.5, 100620.8, 100699.5, 100777.8, 100843.1, 100915.9, 
    100980.7,
  100056.3, 100087.3, 100082, 100153.2, 100218, 100296.6, 100381.9, 100470.7, 
    100562.5, 100650.9, 100734.6, 100818.1, 100882.4, 100959, 101028.8,
  100129.3, 100111.1, 100101.6, 100161.2, 100224.1, 100309.4, 100388.4, 
    100484.4, 100579, 100671.4, 100761.6, 100846.2, 100915.4, 100994, 101070.1,
  99025.85, 99083.84, 99188.75, 99287.48, 99404.54, 99518.75, 99645.55, 
    99760.05, 99882.01, 100014.6, 100160.6, 100311.1, 100450.9, 100581, 
    100695.1,
  99001.58, 99067.72, 99172.98, 99274.4, 99392.2, 99506.98, 99630.13, 
    99754.21, 99901.95, 100022.1, 100202, 100348.6, 100497.8, 100626.6, 
    100741.4,
  98965.44, 99047.81, 99177.09, 99295.95, 99425.41, 99536.67, 99657.81, 
    99801.32, 99940.22, 100069.4, 100263.6, 100417.2, 100570.6, 100693, 
    100803.8,
  98925.18, 99012.45, 99146.87, 99275.12, 99415.62, 99539.31, 99664.34, 
    99824.21, 99944.7, 100104.5, 100300.2, 100471.6, 100627.4, 100749.2, 
    100859.4,
  98891.56, 98974.27, 99118.34, 99274.74, 99418.96, 99564.96, 99694.42, 
    99865.17, 99976.3, 100154.3, 100344, 100537.7, 100689.8, 100813.2, 100922,
  98869.16, 98945.1, 99092.12, 99264.93, 99418.08, 99584.61, 99731.81, 
    99901.15, 100008.9, 100193.7, 100387.4, 100594, 100744.6, 100874.5, 
    100983.1,
  98886, 98928.76, 99079.99, 99263.64, 99434.17, 99611.59, 99779.66, 
    99940.01, 100066.3, 100245.3, 100441.3, 100652.8, 100803.2, 100941.7, 
    101047.6,
  98921.39, 98937.13, 99071.52, 99262.02, 99446.52, 99638.86, 99821.97, 
    99980.97, 100129.1, 100302.3, 100501.1, 100706.1, 100861.7, 101002.8, 
    101109.7,
  98950.84, 98968.2, 99063.2, 99267.09, 99461.66, 99671.73, 99865.55, 
    100028.4, 100197.8, 100370, 100566.7, 100762, 100924.2, 101064.5, 101175.9,
  98971.48, 98999.24, 99072.41, 99275.41, 99478.88, 99701.1, 99910.74, 
    100077, 100265.6, 100440.4, 100633.5, 100823.9, 100985.8, 101129.6, 
    101241.3,
  99910.26, 100030.7, 100132.3, 100242.1, 100371.6, 100498, 100611.4, 
    100724.8, 100857, 100991.2, 101112.3, 101221.9, 101312.6, 101382.7, 
    101438.4,
  99906.72, 100014, 100107, 100219.1, 100354.4, 100480.8, 100607.2, 100734.6, 
    100869.5, 101011, 101139.8, 101258.1, 101352.1, 101426.8, 101485.3,
  99900.82, 100025.6, 100135.4, 100239, 100375.2, 100514.1, 100648.2, 
    100776.8, 100925.3, 101066.2, 101199.9, 101315.5, 101407.9, 101481.2, 
    101540.4,
  99899.69, 100023.2, 100126.8, 100233.9, 100369.7, 100516.3, 100650.9, 
    100786.4, 100947.2, 101094.9, 101239.4, 101358.5, 101454.2, 101529.8, 
    101590.4,
  99905.12, 100029.1, 100134.6, 100258, 100384.7, 100535.2, 100670.6, 
    100822.9, 100982, 101139.1, 101290.1, 101407.9, 101504.6, 101580, 101641.2,
  99903.31, 100037.6, 100141.3, 100273.9, 100390.4, 100546.2, 100683, 
    100848.5, 101006.3, 101176, 101330.5, 101454.4, 101555.3, 101634.4, 
    101697.9,
  99897.23, 100041.4, 100157.7, 100294.4, 100414.3, 100565.2, 100709.8, 
    100882.7, 101037.5, 101216.7, 101376.3, 101503.6, 101605.3, 101684.5, 
    101747.2,
  99887.65, 100037, 100168.5, 100304.1, 100439, 100578.3, 100737.9, 100911.4, 
    101070, 101252.9, 101416.2, 101548.1, 101652.7, 101733.4, 101797.7,
  99880.62, 100026.9, 100177, 100315.6, 100467.4, 100596.9, 100770.5, 
    100941.3, 101106.2, 101288, 101456.1, 101594.3, 101700.3, 101782.5, 
    101848.5,
  99872.12, 100015.6, 100181.4, 100328.5, 100490.9, 100615.9, 100797.1, 
    100968.9, 101140.4, 101321.2, 101495.4, 101638.9, 101747, 101834, 101900.8,
  100635.4, 100677.1, 100743.2, 100833.7, 100936.6, 101050.7, 101185.8, 
    101330.3, 101474, 101609.7, 101726.8, 101818.9, 101885.2, 101928, 101954.8,
  100640.6, 100665.7, 100726.5, 100813.3, 100914.4, 101022.8, 101147, 
    101295.4, 101451.8, 101601.8, 101726.4, 101825.6, 101897.5, 101948.2, 
    101980.1,
  100614.5, 100652.3, 100721.4, 100805.4, 100925.5, 101031.7, 101157.9, 
    101304.8, 101464.5, 101614.6, 101738.7, 101838, 101915, 101969.1, 102001.6,
  100602.3, 100639.7, 100705.3, 100777.8, 100898.9, 101009.8, 101136, 101287, 
    101454.3, 101610.4, 101741.2, 101846.4, 101927.6, 101984.8, 102021.7,
  100586.5, 100615.9, 100679.7, 100761.4, 100868.8, 101000.5, 101136.6, 
    101281.8, 101457, 101614.8, 101749.4, 101855.5, 101940.6, 102000.7, 
    102037.5,
  100571.1, 100593.6, 100652.3, 100746.5, 100839.6, 100976.8, 101114.9, 
    101265.2, 101449.1, 101611.5, 101754.2, 101864.6, 101954.9, 102017.4, 
    102059.7,
  100560.1, 100581.7, 100630.7, 100737.1, 100814.5, 100961.4, 101103, 
    101257.9, 101443.8, 101611.1, 101760.8, 101874.9, 101968.1, 102031.5, 
    102077.8,
  100547.5, 100584.3, 100619.8, 100738.5, 100793.3, 100940.5, 101086, 
    101247.5, 101433.6, 101605.9, 101762.3, 101883.1, 101977.9, 102043.8, 
    102094.7,
  100545.1, 100589.1, 100621.8, 100745, 100781.3, 100927.7, 101071.1, 
    101245.4, 101426.8, 101601.5, 101761.4, 101885.8, 101983.4, 102051.2, 
    102105.9,
  100541, 100594.8, 100632.7, 100739.7, 100783.3, 100909.6, 101053.2, 101241, 
    101418.3, 101593.3, 101756.5, 101885.4, 101988.7, 102063.5, 102120.8,
  100838.3, 100891.8, 100950.2, 100997.4, 101060.1, 101132.4, 101159.9, 
    101199, 101280.6, 101364, 101448.7, 101546.3, 101628.6, 101688, 101731.6,
  100803.8, 100884.1, 100945.6, 100998.4, 101062.3, 101133.3, 101173.8, 
    101207.3, 101242.7, 101336.4, 101424.6, 101521.3, 101611, 101677.8, 
    101730.3,
  100784.3, 100864.3, 100927.7, 100983.9, 101047, 101123.9, 101166.3, 
    101212.8, 101248.3, 101322.5, 101418.6, 101512.4, 101602.3, 101672.5, 
    101733.2,
  100747.9, 100834.2, 100911.6, 100980, 101045.2, 101129.7, 101171.3, 101221, 
    101261.4, 101306.3, 101409.8, 101505.6, 101593.8, 101664.4, 101731.6,
  100711, 100796.3, 100886.4, 100961.2, 101030.3, 101121.2, 101172.9, 
    101217.1, 101260.7, 101303.8, 101397.6, 101496.8, 101585.5, 101661, 
    101728.5,
  100673.1, 100751.9, 100845.4, 100930.1, 101014.9, 101104.3, 101175.7, 
    101218.2, 101255.6, 101294, 101382.5, 101487.9, 101580.4, 101659.9, 
    101729.6,
  100629.9, 100701.2, 100797.7, 100883.3, 100984.6, 101074.1, 101168, 
    101213.8, 101259.8, 101296.7, 101370.4, 101477, 101574.8, 101658.1, 
    101729.7,
  100585.8, 100647.7, 100738.1, 100826.2, 100938.6, 101032.7, 101148.4, 
    101208.5, 101257.7, 101293.1, 101359.2, 101466, 101567.9, 101655.5, 
    101731.1,
  100531.9, 100594.1, 100676, 100762, 100878.1, 100987.7, 101112.9, 101198.4, 
    101254.1, 101289.2, 101352.7, 101453.9, 101560.5, 101650.9, 101730.4,
  100476, 100543.8, 100603.9, 100696, 100809.8, 100935.5, 101067.3, 101177.3, 
    101240.4, 101288.9, 101345.4, 101443, 101551.7, 101646.6, 101733.5,
  99674.96, 99832.32, 100002, 100155.5, 100298.9, 100454.1, 100617.4, 
    100789.7, 100943.5, 101082.7, 101204.8, 101307.4, 101395.8, 101464.6, 
    101522.9,
  99588.38, 99738.71, 99901.54, 100068.2, 100212.6, 100371.3, 100538.4, 
    100719.6, 100886.2, 101037.5, 101171.3, 101287.1, 101380.9, 101457, 
    101523.9,
  99531.98, 99685.85, 99845.46, 100012.6, 100161.2, 100322.7, 100493, 
    100679.1, 100853.6, 101017.7, 101156.1, 101278.8, 101381.3, 101462.3, 
    101534.9,
  99479.94, 99629.88, 99785.97, 99945.34, 100092.8, 100258.7, 100427.9, 
    100626.8, 100810.5, 100989.7, 101137.4, 101269.4, 101378.9, 101462.6, 
    101537.9,
  99437.95, 99595.29, 99741.33, 99904.73, 100043.8, 100212.9, 100379, 
    100585.1, 100776.4, 100967.6, 101121.3, 101262.1, 101376.3, 101464.4, 
    101545.2,
  99410.56, 99568.59, 99708.43, 99869.02, 100001.1, 100172.1, 100325.6, 
    100536.5, 100735.5, 100939.2, 101104.4, 101254.3, 101374.4, 101469.1, 
    101546.8,
  99397.16, 99557.21, 99691.72, 99854.77, 99976.8, 100150.7, 100289.6, 
    100501, 100699.1, 100915, 101091.7, 101250.6, 101372.8, 101471.9, 101549.7,
  99399.55, 99555.68, 99689.25, 99849.36, 99968.65, 100140.6, 100265.8, 
    100468.2, 100664.1, 100889, 101076.4, 101244.1, 101372.4, 101476, 101557.6,
  99414.16, 99564.43, 99697.37, 99857.33, 99976.94, 100138.4, 100259.7, 
    100447.4, 100638.2, 100866.5, 101064.6, 101237.1, 101371.2, 101478.3, 
    101565.5,
  99445.56, 99587.29, 99717.41, 99870.59, 99997.66, 100146, 100266.7, 100438, 
    100625.2, 100846.9, 101050.8, 101228.4, 101370.7, 101482.7, 101570.8,
  100985.5, 101127.1, 101258.7, 101361.5, 101442.4, 101504.3, 101551.5, 
    101593.2, 101625.9, 101655.4, 101683.1, 101707.9, 101722.2, 101744.2, 
    101788.6,
  100875.4, 101031.4, 101163.4, 101277.9, 101375.2, 101450.2, 101506, 
    101554.2, 101593.8, 101628.8, 101661.2, 101689.6, 101713.8, 101745.5, 
    101788.1,
  100780.4, 100945.9, 101082.2, 101215.6, 101311.1, 101394.4, 101458.4, 
    101514.4, 101565, 101609.7, 101648.1, 101685.1, 101714.7, 101748, 101803,
  100688.8, 100856.5, 101002.2, 101145.4, 101249.2, 101350.4, 101421.2, 
    101485.7, 101541, 101591.1, 101634.1, 101674.7, 101709.2, 101751.2, 
    101806.5,
  100596.8, 100772.8, 100929.3, 101076.7, 101192.4, 101299.6, 101378.5, 
    101451, 101512.1, 101568.4, 101616, 101663.5, 101700.2, 101755.5, 101814.6,
  100513.7, 100694.7, 100858, 101008.4, 101136.6, 101247.6, 101338.2, 
    101413.1, 101481.9, 101545.5, 101597.2, 101650.8, 101695.5, 101755, 
    101821.6,
  100439.2, 100623, 100790.6, 100945.4, 101081.2, 101198.6, 101297.3, 
    101376.8, 101454.5, 101522.7, 101582.4, 101639.3, 101688.7, 101761.3, 
    101829.6,
  100373.8, 100558.2, 100728.7, 100886.5, 101028, 101151.8, 101257.2, 
    101343.7, 101427.4, 101499.4, 101567.6, 101628.5, 101684.6, 101763.3, 
    101836.9,
  100314.4, 100500.4, 100672.8, 100833.2, 100979.5, 101108.2, 101218.4, 
    101312.5, 101402.2, 101478.4, 101554.4, 101622.4, 101681.9, 101768.7, 
    101844.1,
  100261.2, 100447.3, 100621.6, 100784, 100934.5, 101066.2, 101183.1, 
    101284.5, 101379.9, 101459.8, 101546.4, 101617.4, 101681.2, 101775.2, 
    101852.3,
  102335.7, 102386.5, 102441.4, 102478.7, 102500.6, 102510.2, 102503.8, 
    102487.6, 102461.6, 102421, 102379, 102326.7, 102281.7, 102223.9, 102176.1,
  102278.4, 102343.1, 102409.6, 102457.4, 102488.3, 102509.5, 102511, 
    102500.9, 102478.6, 102445, 102406.2, 102356.4, 102308.1, 102260, 102198.3,
  102214.3, 102285.6, 102348.5, 102407.6, 102452, 102482.6, 102499, 102497.3, 
    102487.1, 102456.9, 102425.1, 102378.2, 102330.6, 102283.1, 102234.6,
  102142.4, 102233.4, 102307.9, 102381.6, 102426.1, 102464.8, 102490.7, 
    102495.9, 102491.3, 102468.7, 102441.7, 102398.3, 102355.9, 102301.5, 
    102260.5,
  102065.3, 102162.6, 102240.7, 102332.1, 102380.2, 102426.2, 102462.3, 
    102477.7, 102484.3, 102469.1, 102446.6, 102409.9, 102370.1, 102319.7, 
    102279.4,
  101977.5, 102087.2, 102174.2, 102278.4, 102336.9, 102390.9, 102434.4, 
    102459.3, 102471.5, 102463.8, 102449.3, 102416.4, 102383.2, 102330.5, 
    102297,
  101880.7, 102007.1, 102097.3, 102212.5, 102283.3, 102346.2, 102398.4, 
    102431.9, 102452.3, 102454.1, 102441.3, 102417.2, 102389, 102342.1, 
    102310.7,
  101784.6, 101913.2, 102018.8, 102139.5, 102224.9, 102298.1, 102357.8, 
    102400.5, 102426, 102436, 102430.3, 102411.1, 102389.6, 102346.9, 102322.8,
  101678.1, 101818.2, 101932.6, 102061.7, 102159, 102240.8, 102309.9, 
    102363.9, 102393.6, 102412.1, 102411.6, 102398.7, 102384.4, 102346, 
    102327.6,
  101570.4, 101721.4, 101842.4, 101979.5, 102086.1, 102180.8, 102257, 102319, 
    102357.5, 102382.3, 102391.6, 102382.6, 102370.5, 102342.4, 102324.6,
  101662.4, 101764.6, 101855.4, 101943.4, 102010.6, 102064.3, 102102.4, 
    102133.2, 102151, 102154.7, 102149.5, 102127.1, 102103.3, 102074.3, 102051,
  101713.7, 101824.4, 101918.2, 102003.2, 102062.2, 102118.5, 102155, 
    102185.9, 102200.6, 102206, 102200.7, 102182.9, 102154.1, 102116.6, 102081,
  101780.3, 101884.8, 101977.3, 102059.3, 102119.3, 102167.8, 102206.1, 
    102231.7, 102251.1, 102254.3, 102249.7, 102229.9, 102203.8, 102163.2, 
    102125.6,
  101831.3, 101934.7, 102037, 102108.2, 102175.5, 102217.4, 102257.3, 
    102280.9, 102300.3, 102305.2, 102298.8, 102281.6, 102255, 102216.5, 
    102170.2,
  101877.3, 101975.9, 102081.7, 102157.5, 102224.2, 102265.4, 102303.4, 
    102327.1, 102343.4, 102348.1, 102344.7, 102328.6, 102304.3, 102268.9, 
    102220.4,
  101917.2, 102013.6, 102118.6, 102197.8, 102264, 102312.2, 102344.3, 
    102372.1, 102387.6, 102391.7, 102385, 102368.3, 102345.6, 102307.8, 
    102269.3,
  101960.4, 102050, 102148.4, 102233.3, 102301, 102348, 102384.9, 102409.3, 
    102427.1, 102434, 102426.6, 102411.4, 102384.8, 102346, 102306.8,
  102006.7, 102087.9, 102177.6, 102262.6, 102333.7, 102381.7, 102418.1, 
    102445.3, 102461.2, 102470, 102464, 102447, 102424, 102383.9, 102338.9,
  102055.3, 102127.4, 102206.5, 102287.5, 102356.8, 102411.2, 102453.4, 
    102475.8, 102493.2, 102501.5, 102498.1, 102481, 102457.8, 102422.3, 
    102377.6,
  102101.8, 102160.6, 102233.5, 102307, 102372.5, 102435.4, 102473.4, 102506, 
    102518.2, 102532.9, 102533.1, 102512.9, 102489, 102451.9, 102411.4,
  100257.5, 100406.7, 100533.8, 100669.5, 100797.9, 100920.6, 101041.6, 
    101146.7, 101241.2, 101321.8, 101396.9, 101459.1, 101514.2, 101554.9, 
    101582.7,
  100273.7, 100416.8, 100554.2, 100689.6, 100829.6, 100970.2, 101087.2, 
    101191, 101278.4, 101356.3, 101427.5, 101488.7, 101538.4, 101573.9, 
    101598.5,
  100323.2, 100458, 100603.6, 100744, 100893.5, 101034.1, 101151.5, 101252.7, 
    101340.9, 101416.4, 101482.1, 101533.4, 101574.4, 101602.4, 101620.9,
  100370.4, 100484.5, 100641, 100791.1, 100952.4, 101096.1, 101210.8, 101311, 
    101396.8, 101471, 101530.5, 101579.7, 101614.5, 101638.7, 101653.2,
  100419.4, 100530, 100711.2, 100862.6, 101030.6, 101169.4, 101279.8, 
    101387.9, 101470.4, 101546.8, 101602, 101644.2, 101671.8, 101686.1, 
    101693.1,
  100469.7, 100606.9, 100786.4, 100939.8, 101104.8, 101241.2, 101355.7, 
    101466.1, 101547.2, 101619.3, 101668.2, 101704.6, 101728, 101741.1, 101742,
  100533.4, 100700.9, 100864.4, 101024.8, 101183.9, 101316.9, 101440.8, 
    101542.5, 101625.1, 101689.3, 101735.4, 101767.7, 101786.4, 101795.5, 
    101793.9,
  100613.5, 100795.4, 100944.4, 101105.7, 101258.5, 101395, 101518, 101613, 
    101695.9, 101755.3, 101798.3, 101828.2, 101846, 101853.5, 101852.7,
  100704.2, 100883.5, 101031.8, 101188.8, 101343.1, 101479.8, 101597.8, 
    101691.7, 101769.7, 101828.2, 101868.9, 101898.3, 101912.8, 101917.6, 
    101916.4,
  100814.1, 100970.9, 101122.3, 101276.9, 101426.1, 101561.7, 101672.7, 
    101767.6, 101841.5, 101898.4, 101939, 101966.7, 101981.4, 101985, 101981.5,
  100157.8, 100286.2, 100425.9, 100547.6, 100669.6, 100794.1, 100904.2, 
    101005.8, 101100.5, 101188.1, 101261.4, 101318.9, 101370.2, 101412, 
    101450.5,
  100070.7, 100209.8, 100340.3, 100469.3, 100602.7, 100723.1, 100835, 
    100938.7, 101037.8, 101128.4, 101212.4, 101282.5, 101343.2, 101393.5, 
    101431.7,
  99998.38, 100136.4, 100270.3, 100414.2, 100542.9, 100664.6, 100781.2, 
    100890.6, 100996.2, 101093.3, 101181.4, 101259.9, 101330.3, 101389.8, 
    101437.9,
  99933.31, 100069.3, 100205.8, 100344.2, 100469.1, 100597.8, 100718.8, 
    100831, 100942, 101048.1, 101145.3, 101232, 101310.7, 101379.1, 101434.7,
  99883.5, 100018.1, 100153.1, 100289.8, 100416.8, 100555.5, 100676.1, 
    100798.8, 100917.9, 101027.2, 101129.2, 101222.7, 101309.3, 101382.4, 
    101445.3,
  99853.61, 99983.83, 100119, 100247.7, 100384.7, 100524.6, 100649.8, 
    100777.8, 100898.3, 101010.3, 101120.3, 101222, 101314, 101389.8, 101458,
  99850.94, 99963.91, 100098.1, 100227.9, 100372.6, 100509, 100644, 100779.8, 
    100899.7, 101018.9, 101132.9, 101237.3, 101329.2, 101408.6, 101476.7,
  99857.66, 99966.39, 100106.6, 100236.9, 100379.2, 100518.9, 100668.8, 
    100798.8, 100921.4, 101043.7, 101156.3, 101262.3, 101357.8, 101436.9, 
    101503.5,
  99891.05, 99999.82, 100138.2, 100272.1, 100417.3, 100565.1, 100713.2, 
    100836.7, 100967.5, 101086.3, 101203.1, 101307.8, 101401.2, 101475.8, 
    101538.7,
  99947.07, 100062.5, 100206.1, 100333.4, 100487.4, 100635.7, 100775.1, 
    100902.9, 101034.9, 101150, 101266, 101364.4, 101451, 101524.5, 101586.4,
  102125.8, 102176, 102229.2, 102266.2, 102297.7, 102312.1, 102312.7, 
    102315.8, 102300.8, 102274.4, 102243, 102202.3, 102163, 102113.9, 102066.6,
  102026.9, 102095.4, 102162.7, 102209.4, 102246.7, 102270.6, 102284.5, 
    102291.2, 102283.2, 102266.7, 102236.8, 102203, 102169.9, 102124.8, 
    102086.5,
  101929.4, 102004.7, 102081.7, 102140, 102190.6, 102227.6, 102250.3, 102264, 
    102265.9, 102255.7, 102233.4, 102203.6, 102169.9, 102130.3, 102092.5,
  101817.5, 101910.8, 101999.4, 102071, 102132.3, 102178.9, 102210.5, 
    102230.7, 102238.6, 102237.4, 102220.3, 102197.5, 102167.1, 102134.9, 
    102094,
  101699.2, 101799.1, 101903.7, 101992.8, 102060.9, 102119.4, 102162.7, 
    102190.8, 102207.7, 102214.7, 102205.3, 102190.3, 102162.6, 102134.3, 
    102093.9,
  101559.8, 101685.7, 101797.2, 101904.8, 101985.2, 102053.7, 102108.7, 
    102146.9, 102170.7, 102185.9, 102183.1, 102177, 102153.6, 102133, 102087,
  101414.5, 101558.3, 101681.9, 101808.9, 101903.3, 101985, 102047.7, 
    102098.1, 102129.6, 102153.3, 102156.2, 102160.8, 102143, 102126.6, 
    102079.4,
  101260.7, 101422.4, 101563.2, 101704.1, 101813.6, 101911, 101981.5, 
    102042.9, 102083.8, 102114.8, 102124.9, 102136, 102128.2, 102113.6, 
    102075.3,
  101108.8, 101280.4, 101437.2, 101592.4, 101721.5, 101830, 101914.6, 
    101984.1, 102038.1, 102076.5, 102094.5, 102109.8, 102111.5, 102098.8, 
    102066.6,
  100958.1, 101138.3, 101310.3, 101478.6, 101622, 101746.5, 101843.8, 
    101922.7, 101988, 102034.9, 102064.2, 102085.2, 102093.1, 102080.4, 
    102052.9,
  102964.2, 102956.5, 102937.3, 102905.3, 102861.5, 102810.6, 102757.1, 
    102693, 102629.4, 102564.8, 102496.2, 102418.9, 102350.4, 102292.1, 
    102208.7,
  102982.3, 102981.3, 102958.1, 102935.7, 102897.8, 102852.7, 102800.8, 
    102742.7, 102678.1, 102610.3, 102540.8, 102466.1, 102390.2, 102317.4, 
    102246.6,
  102992.9, 102991.4, 102971.4, 102952.1, 102921.2, 102881.5, 102830.5, 
    102772, 102713.7, 102648.6, 102574.3, 102500.7, 102421, 102356.1, 102278,
  102988.5, 102993.3, 102982.5, 102963.2, 102940.8, 102905.6, 102860.5, 
    102807.9, 102748.9, 102684.4, 102611.4, 102536.8, 102456.2, 102388, 
    102305.3,
  102985.7, 102988.9, 102983.8, 102967.2, 102948.7, 102917.4, 102879.9, 
    102833.7, 102775.4, 102713.3, 102645.4, 102570.4, 102490.1, 102414.4, 
    102331.3,
  102964.1, 102974.3, 102977, 102967.9, 102947.9, 102923.2, 102886.4, 
    102851.3, 102802.5, 102740.1, 102672.7, 102602.7, 102522.3, 102446.6, 
    102361.9,
  102928.4, 102945.4, 102958.9, 102956.1, 102941.7, 102920.6, 102891.1, 
    102856, 102814.3, 102757.1, 102694.5, 102628.1, 102549.5, 102476.6, 
    102389.6,
  102887.8, 102905.6, 102930.8, 102932.5, 102927.5, 102918.8, 102890.3, 
    102856.9, 102821.1, 102765.8, 102710.8, 102644.5, 102573.3, 102498.8, 
    102419.2,
  102832.8, 102863.5, 102889.6, 102905.4, 102903.9, 102902.4, 102880, 
    102854.9, 102818.4, 102768.6, 102721, 102659.8, 102589.6, 102514.2, 
    102438.9,
  102769.3, 102813.6, 102841.3, 102863.5, 102870, 102875.5, 102863, 102843.5, 
    102809.4, 102764.3, 102722.1, 102667.7, 102601.4, 102526.5, 102458.3,
  102773.9, 102753.1, 102734.4, 102691.6, 102646.6, 102594.8, 102534.4, 
    102473.3, 102403.7, 102329.3, 102252.9, 102180.6, 102107.4, 102040, 
    101968.2,
  102832.9, 102813.8, 102792.7, 102754.1, 102704.7, 102651.7, 102592.2, 
    102527.9, 102458.7, 102385.4, 102310.7, 102232.4, 102159.3, 102078.4, 
    102006.8,
  102887.4, 102868.9, 102843.4, 102809.1, 102760.1, 102707.9, 102645.7, 
    102580.6, 102511.2, 102436.8, 102360.3, 102279.8, 102204.1, 102130, 
    102048.9,
  102940.6, 102925.1, 102894.8, 102859.3, 102812.3, 102755.8, 102698.9, 
    102634, 102563.5, 102486, 102411.4, 102331.6, 102251.3, 102170.2, 102095.7,
  102988.2, 102973, 102944.3, 102903.6, 102860.3, 102805.6, 102743, 102680.9, 
    102613.9, 102534.8, 102458.7, 102378.1, 102296, 102212.7, 102132.8,
  103022.1, 103004.7, 102980.2, 102939.8, 102901.1, 102851.9, 102784.5, 
    102727, 102662.9, 102579.6, 102502.6, 102424.7, 102340.8, 102257.8, 
    102173.3,
  103038.3, 103028.5, 103014.2, 102969.6, 102930.2, 102883.2, 102825.8, 
    102763.8, 102703.9, 102625.1, 102543.7, 102466.5, 102382.8, 102296.4, 
    102211.3,
  103048.3, 103033.9, 103029.1, 102993.2, 102953, 102910.1, 102859.7, 
    102799.2, 102738.8, 102665.3, 102581.9, 102505.1, 102422.1, 102337.2, 
    102247.9,
  103042.4, 103042.5, 103033.8, 103006.9, 102969.2, 102927.7, 102881.1, 
    102821.7, 102766.1, 102694.9, 102618.7, 102541.7, 102457.5, 102371.2, 
    102281.9,
  103031.3, 103033.7, 103025.8, 103000.9, 102978.6, 102939.9, 102894, 
    102835.5, 102784.4, 102719.2, 102648.9, 102573.8, 102491.9, 102405.5, 
    102313.6,
  102566.4, 102546.8, 102530.4, 102492.8, 102452.3, 102399.5, 102342, 
    102276.5, 102208.3, 102135.5, 102059.3, 101985.7, 101912.6, 101839.9, 
    101766.8,
  102621.3, 102604.5, 102584.9, 102549.2, 102510.2, 102459.7, 102400, 102335, 
    102269.3, 102198.9, 102126.1, 102043.3, 101967.9, 101887.8, 101811.2,
  102663.1, 102654.2, 102637, 102606.1, 102562.6, 102515.1, 102461.4, 
    102395.4, 102327, 102254.8, 102181.4, 102099.2, 102022.8, 101945.6, 
    101864.5,
  102714.8, 102708.7, 102688.1, 102662, 102622.1, 102568.9, 102515.2, 
    102453.2, 102385.8, 102313.1, 102242.5, 102162, 102077.6, 101996.7, 
    101914.3,
  102762.1, 102756.5, 102737.8, 102710.7, 102676.5, 102622.9, 102568.5, 
    102506.8, 102440.3, 102368, 102295.9, 102217.9, 102131.7, 102049.8, 
    101963.4,
  102811.9, 102808.7, 102786, 102760.9, 102720.9, 102676.7, 102618.3, 
    102560.3, 102492.1, 102422.4, 102348.7, 102274.4, 102188.6, 102102.5, 
    102016.1,
  102852.9, 102853.3, 102841.6, 102809.1, 102763.2, 102719.4, 102665.3, 
    102606.4, 102543, 102472.8, 102399.3, 102323.5, 102241.3, 102152.9, 
    102064.6,
  102890.2, 102896.7, 102883.1, 102853.3, 102814.6, 102759.6, 102711.9, 
    102653.1, 102587.2, 102518.5, 102445.2, 102369.9, 102291.1, 102206.1, 
    102114,
  102924.1, 102928.4, 102912.6, 102882.9, 102846, 102798.8, 102747.9, 
    102696.1, 102627.1, 102560.1, 102488.3, 102412.5, 102333.2, 102251.8, 
    102160.4,
  102939.1, 102945.4, 102936, 102904.9, 102862.3, 102817.5, 102773.6, 
    102725.6, 102659.6, 102594.5, 102523.1, 102451.3, 102374.2, 102294.4, 
    102208,
  102605.1, 102565, 102530.5, 102484.3, 102438.2, 102383.1, 102329.6, 
    102267.6, 102204.9, 102136.7, 102064.5, 101994.6, 101928.9, 101856.5, 
    101787.6,
  102692.7, 102649.4, 102612.4, 102565, 102517.8, 102463, 102404.8, 102341.6, 
    102275.3, 102205.5, 102133.2, 102059.8, 101987.1, 101914.9, 101839.7,
  102776.1, 102728, 102691.7, 102642.3, 102591.1, 102535.4, 102477, 102414.4, 
    102345.4, 102274.3, 102199.3, 102120, 102042.5, 101970, 101890.4,
  102851.2, 102805.3, 102767.3, 102718, 102667.3, 102609, 102548.4, 102483.1, 
    102413.1, 102338.6, 102262.3, 102185.4, 102101.8, 102023.3, 101942.7,
  102919.5, 102879.2, 102839.6, 102786.3, 102737.1, 102676.5, 102615.6, 
    102549.6, 102479.1, 102406.1, 102324.7, 102244.7, 102160.9, 102076.2, 
    101993.7,
  102984, 102947.8, 102911, 102855.4, 102802, 102742.6, 102677.8, 102611.1, 
    102537.4, 102465.1, 102385.1, 102305.2, 102219.3, 102131.8, 102045.8,
  103036.7, 103012.4, 102972.8, 102918, 102861.3, 102801, 102737.5, 102671.1, 
    102595.7, 102523.3, 102442.4, 102357.8, 102275.1, 102183.3, 102095,
  103080.8, 103066.6, 103014.9, 102974.6, 102913.7, 102853.7, 102790.8, 
    102725.6, 102648.4, 102574.6, 102496.2, 102410.4, 102327.1, 102236, 
    102142.9,
  103122.5, 103113.8, 103058.5, 103011.2, 102958.2, 102895.7, 102836.7, 
    102774.7, 102698.4, 102624.3, 102545.2, 102460.3, 102373.8, 102282, 
    102188.4,
  103156.7, 103146.9, 103096.3, 103041, 102987.4, 102932.9, 102872.7, 
    102814.9, 102741.8, 102667.2, 102590.1, 102504.6, 102419.5, 102328.2, 
    102231.6,
  102472.3, 102403.6, 102354.7, 102295, 102245.8, 102191.4, 102138.9, 
    102084.2, 102028.8, 101970.5, 101910.8, 101847.7, 101786.1, 101729.7, 
    101671.6,
  102579.9, 102503, 102462.6, 102401.3, 102347.6, 102285.6, 102227.4, 
    102168.1, 102107.5, 102044.5, 101979.8, 101916.9, 101850.4, 101787.3, 
    101722.3,
  102690, 102625.3, 102569.7, 102498, 102439.1, 102373.9, 102310.5, 102247.6, 
    102182.5, 102117.3, 102048.8, 101976.4, 101904.6, 101837.9, 101770.3,
  102797.2, 102724.9, 102665.7, 102594.2, 102530.3, 102461.7, 102391.7, 
    102325.2, 102255.3, 102184.2, 102112.9, 102038.9, 101963, 101891.5, 
    101818.2,
  102894.5, 102817.2, 102756.7, 102683.6, 102610.8, 102538.9, 102464.5, 
    102391.1, 102321.2, 102246.3, 102172, 102095.3, 102016.9, 101937.8, 
    101862.9,
  102982.8, 102902.1, 102835.5, 102760.6, 102684.6, 102610.5, 102534.1, 
    102455.9, 102379.2, 102303.3, 102225.9, 102148.2, 102067.9, 101986.2, 
    101905.1,
  103062.3, 102974.9, 102905.2, 102831.2, 102751.5, 102674.6, 102593.8, 
    102513.5, 102435.4, 102357.4, 102275.6, 102197.3, 102114, 102031.8, 
    101946.5,
  103129.6, 103046.5, 102965.7, 102890.2, 102813.4, 102730.9, 102650.3, 
    102567.5, 102486.2, 102405.8, 102324.1, 102243, 102158.7, 102074.7, 
    101987.4,
  103183.3, 103104.6, 103022.9, 102941, 102865.2, 102783.4, 102699.2, 
    102617.5, 102532, 102452.3, 102367.4, 102285.3, 102199, 102114.5, 102024.3,
  103225.7, 103147.7, 103071.8, 102986.8, 102908.4, 102826.9, 102744, 
    102657.9, 102574.7, 102491.5, 102406.7, 102322.2, 102235.6, 102149.9, 
    102060.1,
  101780.5, 101676.6, 101601.5, 101511.7, 101430.7, 101349.4, 101281.5, 
    101223, 101170.9, 101123.8, 101081.4, 101047.6, 101016.9, 100996.1, 100979,
  101909.5, 101806.4, 101724.5, 101634.1, 101559.1, 101481.8, 101408.4, 
    101344.2, 101290, 101242.5, 101198, 101163.7, 101134.5, 101109.1, 101077.2,
  102016.3, 101916.3, 101841.7, 101756.4, 101678.7, 101603, 101533.2, 
    101465.4, 101402.2, 101349.4, 101299.8, 101253.3, 101212.4, 101178.8, 
    101144.5,
  102116.8, 102025.8, 101948.6, 101864.8, 101787.5, 101713.8, 101644.8, 
    101581.2, 101517.6, 101459.4, 101411.9, 101366.9, 101324.6, 101284.8, 
    101243.4,
  102210.6, 102122.3, 102044.7, 101967.3, 101893.6, 101818, 101750.3, 
    101682.5, 101623, 101565.7, 101511.7, 101464.8, 101418.3, 101374.8, 
    101333.4,
  102286.4, 102200.8, 102133, 102054, 101985, 101914, 101848.5, 101777.7, 
    101717.6, 101660.2, 101607.4, 101558.8, 101513.6, 101465.9, 101423,
  102344.9, 102260.8, 102200.9, 102130.3, 102060.9, 101992.2, 101931.1, 
    101866.8, 101804.1, 101743.4, 101690.2, 101638.2, 101590.1, 101544.8, 
    101497.8,
  102388.8, 102310.3, 102247.8, 102187.6, 102125.8, 102058.4, 101998, 
    101939.9, 101878.6, 101817, 101760.6, 101708.7, 101657.3, 101614.3, 
    101566.3,
  102424.1, 102350.3, 102286.9, 102226.9, 102174.9, 102112.7, 102052.5, 
    101996.2, 101946, 101883.5, 101825.9, 101771.9, 101721.5, 101670.9, 
    101624.6,
  102442.8, 102379.8, 102318.8, 102261.1, 102208.7, 102156, 102098.4, 102041, 
    101990.7, 101940.3, 101882.9, 101828.8, 101776.4, 101726.7, 101679.6,
  100283.5, 100115.8, 99980.13, 99873.84, 99808.82, 99779.18, 99788.09, 
    99825.4, 99899.98, 99981.16, 100063.3, 100147, 100237, 100316.7, 100389.4,
  100544.1, 100351.7, 100182.6, 100063.4, 99987.12, 99941.91, 99932.08, 
    99948.16, 99985.48, 100038.1, 100106.5, 100176.1, 100244, 100311.4, 
    100386.1,
  100759.2, 100583.9, 100417.3, 100284.8, 100183.3, 100118, 100080.1, 
    100070.8, 100088.5, 100123.2, 100171.6, 100231.5, 100292.5, 100358.7, 
    100412.8,
  100971.2, 100799.4, 100634.5, 100496.6, 100382.4, 100301.6, 100246.7, 
    100218, 100212.4, 100225.2, 100254, 100296.2, 100342.3, 100390.5, 100428.8,
  101155.8, 101003, 100853.7, 100706.9, 100586.3, 100490.2, 100415.9, 
    100368.5, 100341.9, 100332.8, 100345.2, 100371.6, 100402.4, 100438.9, 
    100466,
  101321.3, 101182.6, 101050.7, 100914.8, 100793.8, 100690.1, 100607.6, 
    100544.6, 100501.5, 100481.8, 100461.7, 100471.4, 100473.6, 100495.1, 
    100524.1,
  101466.6, 101346.9, 101226.2, 101104.2, 100990.5, 100893.9, 100801.6, 
    100731.1, 100673.2, 100628, 100599.5, 100577.7, 100574.8, 100586.3, 
    100596.5,
  101593.4, 101491.3, 101389.5, 101281.8, 101176, 101086.5, 101003.8, 100927, 
    100858.8, 100805.7, 100756.9, 100721.8, 100700.3, 100679.8, 100681.4,
  101698.7, 101615.9, 101532.1, 101439.3, 101348.3, 101259.4, 101179.6, 
    101111.4, 101038.6, 100971.6, 100912.7, 100869.5, 100826.7, 100798.1, 
    100778.2,
  101787.1, 101723.3, 101653.4, 101577.2, 101498.3, 101418.2, 101346.5, 
    101278.9, 101213.9, 101150.8, 101081.8, 101026.8, 100976, 100924.3, 
    100893.9,
  99239.94, 99106.39, 98976.13, 98908.66, 98916, 99004.28, 99149.05, 
    99308.64, 99460.3, 99612.25, 99755.87, 99909.23, 100059.5, 100198, 
    100333.6,
  99472.12, 99351.17, 99237.37, 99159.33, 99140.77, 99186.63, 99286.77, 
    99399.8, 99521.18, 99654.73, 99790.68, 99921.97, 100058.9, 100193.9, 
    100320.2,
  99647.51, 99548.17, 99446.13, 99379.7, 99352.2, 99367.82, 99426.62, 
    99511.07, 99615.12, 99727.48, 99845.3, 99963.38, 100085.1, 100207.5, 
    100319.6,
  99836.74, 99746.1, 99669.46, 99598.59, 99561.44, 99560.56, 99588.05, 
    99646.25, 99728.57, 99821.37, 99918.26, 100021.7, 100128.9, 100237.3, 
    100339.4,
  100014.1, 99924.09, 99849.92, 99793.36, 99760.34, 99746.39, 99759.04, 
    99791.22, 99847.35, 99924.56, 100010.4, 100102.8, 100193.5, 100285, 
    100373.5,
  100179.4, 100095.2, 100021.7, 99969.9, 99936.5, 99921.51, 99920.74, 
    99944.42, 99984.23, 100040, 100110.5, 100186, 100262.2, 100342.5, 100421.9,
  100361.9, 100261.9, 100183.6, 100131, 100098.9, 100079.5, 100079.9, 
    100091.1, 100118.9, 100160.3, 100213.5, 100271.2, 100335, 100399.5, 
    100462.8,
  100538.3, 100427.5, 100339.8, 100270.2, 100223.8, 100200.5, 100191.4, 
    100203.3, 100226.9, 100265, 100307.7, 100350.6, 100393.2, 100446.2, 
    100511.2,
  100716, 100592.6, 100495.6, 100418.6, 100365.5, 100327, 100312.6, 100305, 
    100324.7, 100352.4, 100382.9, 100421.4, 100466.2, 100508.1, 100545.6,
  100893.4, 100768.2, 100660.4, 100568.8, 100503.9, 100454.3, 100423.9, 
    100409.2, 100413.6, 100428.5, 100457.5, 100483.1, 100508, 100548, 100610,
  98815.48, 98837.43, 98978.4, 99158.55, 99340.85, 99525.2, 99702.79, 
    99866.32, 100022.6, 100163.3, 100292.2, 100402.8, 100501, 100588.5, 
    100671.1,
  98722.72, 98779.41, 98902.57, 99061.95, 99235.39, 99419.53, 99601.48, 
    99772.55, 99931.46, 100071.7, 100208.4, 100329.7, 100439, 100531.5, 100618,
  98755.77, 98809.16, 98878.83, 99009.23, 99172.17, 99345.77, 99518.6, 
    99688.24, 99846.84, 99994.74, 100129.2, 100254.1, 100368.6, 100470.4, 
    100557.4,
  98873.05, 98888.24, 98917.41, 99016.77, 99149.37, 99306.07, 99464.54, 
    99625.24, 99780.9, 99929.13, 100067.5, 100196.9, 100316.3, 100424.3, 
    100520.4,
  99030.79, 99012.87, 99002.64, 99073.94, 99166.38, 99297.02, 99441.38, 
    99587.09, 99730.08, 99873.79, 100008.2, 100136.4, 100259.8, 100369.8, 
    100469.5,
  99216.84, 99170.84, 99130.32, 99162.54, 99219.65, 99321.73, 99431.87, 
    99563.14, 99698.22, 99834.31, 99962.36, 100091.3, 100209.8, 100328.2, 
    100431.9,
  99391.59, 99334.39, 99283.72, 99279.73, 99306.61, 99376.32, 99460.14, 
    99569.12, 99680.84, 99806.58, 99934.06, 100056.3, 100177.1, 100295, 
    100399.9,
  99561.52, 99486.81, 99430.15, 99415.5, 99419.67, 99450.6, 99509.92, 
    99585.48, 99686.23, 99801.88, 99917.88, 100039.4, 100153.8, 100266.6, 
    100376.1,
  99707.2, 99627.76, 99571.66, 99527.7, 99521.64, 99543.96, 99584.78, 
    99641.05, 99712.23, 99804.64, 99912.27, 100025.2, 100135.7, 100250.7, 
    100362.4,
  99821.81, 99743.55, 99699.54, 99648.24, 99629.1, 99629.73, 99647.62, 
    99698.94, 99752.51, 99824.27, 99911.09, 100012.3, 100127.6, 100240.9, 
    100351.3,
  99360.69, 99476.41, 99628.99, 99772.44, 99907.95, 100021.2, 100139.3, 
    100273.8, 100394.1, 100513.3, 100618.3, 100721.2, 100809.4, 100893, 
    100970.4,
  99265.9, 99404.89, 99571, 99709.34, 99849.44, 99973.93, 100088.8, 100205, 
    100328.7, 100453.8, 100566, 100671.8, 100766.9, 100856.5, 100935.8,
  99156.69, 99308.26, 99481.34, 99623.45, 99772.56, 99905.09, 100024.6, 
    100137.2, 100254.1, 100375, 100496, 100607.5, 100709, 100803.9, 100893.1,
  99052.49, 99215.6, 99403.35, 99551.77, 99709.86, 99847.7, 99979.52, 100097, 
    100210.8, 100330.4, 100452.1, 100571.9, 100678.8, 100779.7, 100869.5,
  98954.83, 99117.78, 99312.71, 99468.3, 99633.53, 99776.38, 99915.59, 
    100039.4, 100155.6, 100272.3, 100393.5, 100517.3, 100629, 100735.1, 
    100830.9,
  98882.98, 99037.22, 99232.18, 99392.95, 99562.77, 99709.91, 99853.41, 
    99984.23, 100105.9, 100223.5, 100338.8, 100467.2, 100587.5, 100696.5, 
    100797,
  98829.94, 98981.65, 99158.2, 99327.3, 99494.68, 99644.88, 99792.95, 
    99926.35, 100051.2, 100173.2, 100288.2, 100414.1, 100540.1, 100655.3, 
    100758.8,
  98813.05, 98954.38, 99107.75, 99271.51, 99435.15, 99587.71, 99736.43, 
    99870.67, 100003, 100122.7, 100242.9, 100367.3, 100496.6, 100617.8, 
    100728.9,
  98830.83, 98951.23, 99075.89, 99237.38, 99388.59, 99540.62, 99686.56, 
    99822.06, 99953.02, 100077.4, 100197, 100320.5, 100452, 100581.1, 100693,
  98868.53, 98976.36, 99072.47, 99218.87, 99359.75, 99505.48, 99643.02, 
    99778.3, 99908.82, 100038.4, 100156, 100282.1, 100414, 100548, 100667,
  98373.07, 98536.88, 98771.48, 98990.34, 99228.7, 99471.94, 99688.7, 
    99898.83, 100094.8, 100272.4, 100437.1, 100580, 100704.5, 100814.8, 
    100913.1,
  98201.23, 98413.18, 98666.7, 98878.38, 99104.61, 99337.87, 99562.52, 
    99787.38, 99990.47, 100182.4, 100345.9, 100498.5, 100634.3, 100756.9, 
    100864.2,
  98124.15, 98329.88, 98549.55, 98761.41, 98979.51, 99212.51, 99448.45, 
    99671.38, 99883.2, 100080.3, 100259, 100421.3, 100565.3, 100695.9, 
    100813.6,
  98100.84, 98284.3, 98487.5, 98687.49, 98900.06, 99118.78, 99354.12, 
    99584.99, 99801.94, 100005.6, 100192.2, 100361.7, 100514.4, 100654.1, 
    100778.8,
  98116.43, 98266.78, 98445.11, 98636.09, 98837.34, 99050.64, 99282.23, 
    99507.66, 99730.87, 99935.45, 100126.6, 100304, 100465.7, 100611.8, 
    100742.4,
  98157.18, 98284.88, 98434.4, 98622.02, 98807.05, 99010.48, 99231.41, 
    99455.69, 99668.92, 99878.58, 100075.3, 100259.8, 100426.4, 100577.2, 
    100712.7,
  98229.59, 98330.51, 98466.28, 98632.95, 98802.4, 98994.26, 99201.31, 
    99419.87, 99632.89, 99842.3, 100036, 100223.7, 100394.6, 100550.4, 
    100686.7,
  98317.43, 98405.56, 98524.59, 98669.22, 98823.48, 99002.47, 99194.17, 
    99402.98, 99615.71, 99817.89, 100013, 100198.4, 100374.6, 100531.7, 
    100671.6,
  98404.75, 98491.44, 98598.99, 98725.88, 98870.6, 99030.97, 99208.37, 
    99407.7, 99612.05, 99810.18, 100001.7, 100189.1, 100362.4, 100521, 
    100660.8,
  98499.93, 98588.55, 98686.44, 98801.48, 98935.23, 99082.09, 99248.97, 
    99435.98, 99625.09, 99819.07, 100007.5, 100189.6, 100359.3, 100522.1, 
    100661.6,
  99714.02, 99826.65, 99967.52, 100122.3, 100279.9, 100421.8, 100556, 
    100681.7, 100793.8, 100902.7, 100996.3, 101086.8, 101160.8, 101232.5, 
    101286.2,
  99542.69, 99682.01, 99832.13, 99982.09, 100142, 100297.4, 100444, 100585.4, 
    100712, 100822.1, 100925.9, 101021.1, 101104.7, 101177.5, 101247.7,
  99329.68, 99473.45, 99637.69, 99802.36, 99974.28, 100148, 100301.7, 
    100454.1, 100591, 100721, 100833.1, 100938.3, 101035.2, 101120, 101199.1,
  99142.63, 99292.3, 99467.23, 99645.04, 99831.05, 100007.9, 100188.9, 
    100351.3, 100503.4, 100645.1, 100771.2, 100883.2, 100988.7, 101079.8, 
    101163.7,
  98973.48, 99106.91, 99271.64, 99459.49, 99660.29, 99854.73, 100043.3, 
    100228, 100393.7, 100544.4, 100682.5, 100809.5, 100921.2, 101024.8, 
    101113.4,
  98821.55, 98940.23, 99103.81, 99285, 99494.13, 99699.75, 99905.71, 
    100097.3, 100283.1, 100450.6, 100601.6, 100737.2, 100859.1, 100970, 
    101066.4,
  98674.25, 98781.97, 98944.98, 99124.33, 99331.04, 99550.62, 99767.02, 
    99975.03, 100170.6, 100351.6, 100514.7, 100661.6, 100795.4, 100912.9, 
    101017.9,
  98544, 98647.82, 98809.55, 98984.59, 99192.62, 99412.3, 99640.42, 99858.33, 
    100066.9, 100258.2, 100436.4, 100591.8, 100732.7, 100860.3, 100971.4,
  98436.44, 98544.32, 98694.6, 98867.3, 99066.79, 99289.1, 99524.9, 99750.3, 
    99968.59, 100170.4, 100356.8, 100522.9, 100672.3, 100807.1, 100925.7,
  98371.3, 98479.74, 98611.76, 98776.59, 98972.52, 99190.64, 99424, 99656.55, 
    99881.61, 100091.2, 100285, 100461.3, 100618, 100757.4, 100885.6,
  100129.8, 100279.2, 100430.9, 100571, 100713.7, 100848.9, 100976.5, 
    101088.8, 101192, 101287.2, 101369.7, 101440.1, 101499.2, 101547.4, 
    101589.5,
  100094.7, 100258.5, 100410.7, 100555.8, 100701.8, 100834.9, 100961.9, 
    101078.2, 101186.3, 101282.8, 101366.5, 101440.4, 101502.5, 101555.7, 
    101597.6,
  100078.7, 100236.2, 100387.5, 100538.6, 100687.6, 100830, 100958.6, 
    101077.4, 101185.2, 101280.6, 101365.4, 101440.9, 101504.7, 101558, 
    101604.4,
  100054.3, 100213.1, 100365.5, 100522.1, 100677.5, 100823.6, 100954.4, 
    101074.5, 101182.2, 101279.5, 101367.1, 101441.4, 101510.2, 101566.5, 
    101611.9,
  100042.1, 100191.2, 100343.4, 100501, 100660.6, 100810.5, 100946.3, 
    101067.7, 101174.6, 101272.5, 101359.2, 101436.5, 101505.5, 101564.9, 
    101611.7,
  100043.9, 100173.2, 100326.5, 100483.3, 100643.8, 100795.3, 100933.6, 
    101057.1, 101166.6, 101264.9, 101352.8, 101431.8, 101501.9, 101562.2, 
    101609.6,
  100042.5, 100161.3, 100309.7, 100464.2, 100623.8, 100777.4, 100918.2, 
    101041.8, 101153.8, 101254.5, 101343.2, 101423.3, 101493.5, 101554.9, 
    101606.9,
  100035.3, 100148, 100294.4, 100443.2, 100603.5, 100757.2, 100898, 101024.8, 
    101138.1, 101239.9, 101333, 101413.6, 101484.2, 101545.5, 101601.5,
  100019.4, 100133.3, 100273.9, 100420.1, 100577.8, 100732, 100876.8, 
    101004.8, 101121.4, 101224.8, 101318.8, 101403.3, 101473.9, 101537.8, 
    101592.5,
  99999.88, 100117.5, 100251.8, 100395.7, 100550.2, 100705.7, 100851.8, 
    100982.6, 101101.5, 101207.7, 101303.6, 101389.5, 101463.4, 101527.1, 
    101586.5,
  100840.7, 100939, 101043, 101116.8, 101194, 101253.4, 101311.9, 101357.3, 
    101450.5, 101522.1, 101596.2, 101658.3, 101716, 101758.3, 101793.6,
  100788.3, 100888.7, 100990.3, 101078.6, 101163.6, 101227.7, 101298.3, 
    101348.3, 101429.9, 101523, 101595.9, 101667, 101725.2, 101772.6, 101811.9,
  100746.9, 100848.1, 100957.3, 101046.9, 101138.6, 101206.2, 101286.2, 
    101352.5, 101419.2, 101522.6, 101603.1, 101683.8, 101741.6, 101795.7, 
    101835.7,
  100699.6, 100809.3, 100921.9, 101013.9, 101110.9, 101189.1, 101269.2, 
    101351.5, 101416.3, 101525.3, 101612.5, 101696.1, 101757.1, 101812.3, 
    101851.2,
  100654.4, 100768.1, 100888.6, 100985.8, 101080.2, 101169.9, 101249.8, 
    101341.3, 101418.6, 101521.3, 101616.7, 101704, 101771.1, 101827.8, 
    101873.9,
  100602.1, 100727.9, 100847.4, 100952.7, 101049.9, 101149.2, 101235.7, 
    101332.1, 101422.6, 101513.9, 101619.8, 101708.6, 101782.1, 101841.5, 
    101891.2,
  100553, 100688.2, 100811.8, 100922.7, 101021.6, 101126.2, 101218.6, 
    101320.4, 101417.8, 101507.9, 101619.9, 101710.7, 101791.3, 101856.6, 
    101908.6,
  100505.1, 100651.6, 100775.3, 100894.2, 100996.2, 101106.4, 101203.8, 
    101308.3, 101410.1, 101506.9, 101617, 101713, 101798.7, 101866.9, 101920.5,
  100469.5, 100624, 100746.9, 100870, 100975.1, 101087.6, 101189.4, 101296.8, 
    101402.6, 101506, 101616.2, 101717.6, 101807.1, 101880.1, 101935.1,
  100444, 100597.2, 100723.5, 100853.5, 100962.6, 101073.8, 101179.5, 101289, 
    101399, 101506.9, 101619, 101725.5, 101816.7, 101889.4, 101946.9,
  100785.8, 100925.1, 101057.9, 101177.8, 101293.7, 101402.5, 101503.9, 
    101599, 101690.7, 101772, 101840.4, 101890.8, 101932.1, 101958.3, 101971.2,
  100807.1, 100950.6, 101082.4, 101196.8, 101313.7, 101417, 101516.5, 
    101613.6, 101711.9, 101797.5, 101864.9, 101922, 101956.6, 101982.9, 
    101998.6,
  100860.7, 101002, 101122.3, 101233.2, 101338.8, 101438.7, 101536.4, 
    101631.1, 101734.1, 101818.8, 101888.8, 101944.5, 101984.6, 102015.8, 
    102034,
  100913.6, 101061.7, 101178.8, 101287, 101385.4, 101473.6, 101569.7, 
    101662.5, 101760.6, 101846.9, 101917, 101974, 102015.4, 102046.8, 102069.2,
  100975.2, 101121.1, 101235.6, 101339.3, 101432.1, 101510.5, 101599.3, 
    101687.8, 101780.8, 101868.6, 101940.9, 102001.2, 102043.3, 102081.1, 
    102099.7,
  101048.6, 101185.5, 101297, 101396.4, 101485.4, 101558.1, 101639.8, 
    101726.1, 101809.7, 101899.4, 101970.1, 102036.2, 102086.6, 102120.8, 
    102137.2,
  101126.1, 101245.7, 101350.4, 101444.2, 101527.1, 101603.9, 101683.1, 
    101766.8, 101847.8, 101928.9, 102004.3, 102066.6, 102115.1, 102151.2, 
    102169.5,
  101204.9, 101315.1, 101418.2, 101503, 101583, 101661, 101734.5, 101817, 
    101890.1, 101965.6, 102036.9, 102098.4, 102143.5, 102180.7, 102201.4,
  101283.8, 101387.4, 101484, 101568.3, 101642.2, 101718.1, 101790.3, 
    101867.7, 101931.4, 102001, 102066, 102127.5, 102172.2, 102212.1, 102234.1,
  101359.1, 101459.1, 101555.8, 101636.9, 101704.7, 101779, 101846.9, 
    101914.8, 101972.6, 102038.1, 102093.6, 102153.1, 102196.5, 102233.7, 
    102258.1,
  100919.5, 100992.4, 101088.6, 101179.8, 101322.8, 101459.8, 101577.7, 
    101681.4, 101766.7, 101837, 101890.5, 101935.5, 101968.1, 101990, 102001.7,
  100883.1, 100981.6, 101089.4, 101173.6, 101311.5, 101450.8, 101579.4, 
    101695.9, 101789.9, 101866.1, 101919.2, 101963, 101993.8, 102017.2, 
    102030.6,
  100904.9, 100995.9, 101096, 101177, 101314.5, 101457.2, 101591.8, 101716.1, 
    101817.1, 101894.6, 101952, 101998.6, 102030.9, 102052.4, 102063.5,
  100911.7, 101019, 101117.3, 101194.2, 101316.5, 101458.3, 101606.6, 
    101741.1, 101847.5, 101929, 101987.9, 102033.7, 102062, 102082.8, 102093.7,
  100931.4, 101058.3, 101133.5, 101222.5, 101332.7, 101472.7, 101623.2, 
    101759.3, 101871.4, 101957.1, 102019.8, 102066.1, 102093.7, 102117.5, 
    102123.4,
  100956.2, 101105.5, 101151.1, 101253.1, 101356.4, 101493.9, 101646.6, 
    101785.4, 101905.4, 101993.3, 102062, 102109.8, 102137.2, 102154.6, 
    102159.5,
  100984, 101136.2, 101187.5, 101295.5, 101399.4, 101526.8, 101680, 101821.7, 
    101941.1, 102032.7, 102104, 102147.1, 102173.8, 102188.1, 102194,
  101009.4, 101145.5, 101217.2, 101340.4, 101434.2, 101559, 101714.5, 
    101855.4, 101979.5, 102073.2, 102142.4, 102188.6, 102215.5, 102228, 
    102235.9,
  101041.4, 101164.6, 101272, 101402.2, 101484.1, 101606, 101748.4, 101888.4, 
    102019.1, 102113.6, 102185.1, 102229.9, 102256.5, 102271.6, 102274.6,
  101083.6, 101207.9, 101334.8, 101467.4, 101546.3, 101663.8, 101783.8, 
    101923.2, 102056.1, 102152.3, 102226.6, 102271.6, 102298.5, 102309, 
    102311.8,
  101162.8, 101251.9, 101360.6, 101456, 101545.6, 101625.2, 101701.3, 
    101770.8, 101842.1, 101906.7, 101964.8, 102007.7, 102041.2, 102071.7, 
    102081.4,
  101101, 101202.7, 101316.2, 101410.5, 101508, 101593.7, 101675.9, 101752.4, 
    101832.3, 101894.2, 101967.6, 102012.6, 102053.7, 102084.6, 102096.8,
  101079.6, 101171.7, 101279.6, 101370.3, 101476, 101561.4, 101650.4, 
    101738.6, 101832, 101903.2, 101975, 102027.2, 102069.2, 102100.8, 102116.2,
  101038.5, 101127.6, 101230.2, 101326.1, 101440.9, 101530, 101635.6, 
    101734.5, 101831.9, 101914.1, 101984.3, 102044.8, 102087.5, 102117.7, 
    102134.6,
  101003, 101091.1, 101193.6, 101286.4, 101402.4, 101499, 101621.5, 101733.4, 
    101832.1, 101918.1, 101991.3, 102056.1, 102101.2, 102134.7, 102152.1,
  100971.3, 101061.7, 101160.4, 101252.6, 101370.2, 101480.6, 101621.5, 
    101732.5, 101836.1, 101923, 102002.2, 102068.7, 102119.9, 102153.5, 
    102173.7,
  100972, 101069.5, 101155.3, 101248, 101363.3, 101481.6, 101629.5, 101737.1, 
    101848, 101931.7, 102017.5, 102083.9, 102138.3, 102177.8, 102198.2,
  100981.2, 101101.5, 101168.2, 101268.7, 101371.8, 101492.4, 101635, 
    101740.7, 101858.5, 101943.4, 102034.5, 102102, 102161.5, 102200, 102224.1,
  101000.6, 101127, 101176.7, 101290.4, 101369.4, 101512, 101639.7, 101753.1, 
    101870.4, 101964.1, 102054.6, 102125, 102185, 102226.3, 102253.3,
  101042.4, 101143.5, 101179.4, 101306.1, 101395.6, 101537.3, 101647.8, 
    101783.2, 101889.4, 101991.9, 102081.1, 102152.9, 102212.8, 102255.9, 
    102282.4,
  101282.7, 101343.4, 101435.7, 101513.9, 101594.4, 101665.6, 101722.2, 
    101764.9, 101795.1, 101823.4, 101844.4, 101872.4, 101897.8, 101915.7, 
    101923.2,
  101338, 101404.8, 101487.2, 101557.8, 101632.8, 101691.8, 101746.2, 
    101789.2, 101822.2, 101851.5, 101865.1, 101883.9, 101911.9, 101927.9, 
    101939.2,
  101383.4, 101454.1, 101535.3, 101602.2, 101672.8, 101728.7, 101776, 101810, 
    101838.7, 101865.8, 101880.4, 101894.1, 101922.7, 101941.4, 101952.2,
  101441.5, 101516.7, 101594.9, 101660.2, 101724.5, 101773, 101817.9, 
    101851.4, 101869.9, 101890.9, 101907.1, 101914.7, 101932.8, 101952, 
    101963.3,
  101492.4, 101573.6, 101640.8, 101703.3, 101763.5, 101810.9, 101853.8, 
    101881.5, 101898.7, 101915.4, 101925.1, 101934.1, 101942.7, 101970.3, 
    101978.9,
  101554.7, 101625.3, 101690.6, 101752.1, 101804.7, 101852, 101885.2, 
    101914.4, 101927.1, 101938.9, 101941.6, 101943.5, 101955, 101976.5, 
    101990.6,
  101604, 101666, 101729, 101783.9, 101835.4, 101881.2, 101913.2, 101939.2, 
    101948.5, 101957.8, 101955.7, 101959.4, 101959.1, 101982.8, 102002.7,
  101636.5, 101695.6, 101754.5, 101808.2, 101860.8, 101900.4, 101931.9, 
    101954.1, 101964.6, 101970.8, 101963.4, 101965, 101967.1, 101990.8, 
    102014.1,
  101649.2, 101707.4, 101767.7, 101816, 101867.6, 101908, 101938.7, 101961, 
    101970.8, 101978.2, 101973.3, 101975.6, 101980.8, 102001.4, 102029.6,
  101645.9, 101707.4, 101771.4, 101818.6, 101864.1, 101905.5, 101937.6, 
    101954, 101975.9, 101982.5, 101978.7, 101978.3, 101992.8, 102012.2, 
    102051.6,
  100369.9, 100477.3, 100571.7, 100690.5, 100813, 100931.9, 101053.3, 101177, 
    101292.6, 101394.7, 101478.6, 101555.3, 101618.2, 101664.9, 101695.9,
  100370.8, 100492, 100548.4, 100665.2, 100787.7, 100908.7, 101044.3, 
    101174.4, 101298.1, 101398.2, 101486.3, 101563.2, 101624.8, 101672, 
    101709.8,
  100402.9, 100508.3, 100576.9, 100649.1, 100781, 100903.4, 101046.6, 
    101175.2, 101305.1, 101412.2, 101504.1, 101580.4, 101641.2, 101686.3, 
    101716.8,
  100408.5, 100502.4, 100593, 100642, 100782.9, 100899.7, 101051.9, 101188.9, 
    101325.5, 101431.2, 101524.5, 101595.9, 101651.1, 101695.2, 101730.1,
  100391.6, 100484.1, 100594.8, 100662.4, 100789.9, 100904.1, 101058.6, 
    101199.1, 101338.2, 101445.5, 101537.5, 101606.6, 101665, 101711.3, 
    101744.1,
  100378.1, 100468.6, 100594.6, 100676.4, 100803.4, 100919.8, 101073.2, 
    101217, 101356.6, 101463.2, 101555.3, 101626.7, 101685.8, 101728.6, 
    101765.7,
  100395.8, 100477.7, 100609.4, 100706.3, 100835, 100951.4, 101096.6, 
    101242.6, 101376.3, 101484, 101572.5, 101642, 101700.5, 101748.4, 101785.1,
  100459.1, 100519.6, 100646.3, 100755.4, 100881, 100993, 101131.9, 101273.9, 
    101402.5, 101506.9, 101590.2, 101659.7, 101718.6, 101765.6, 101798.9,
  100555.7, 100597.6, 100709.5, 100825, 100939.2, 101049.2, 101178.8, 
    101309.2, 101431.1, 101533, 101614.6, 101678.2, 101729.9, 101779.2, 
    101822.4,
  100662.8, 100699.2, 100799.8, 100903.6, 101017.4, 101117.3, 101238.8, 
    101351.5, 101467.3, 101562.1, 101639.9, 101696.2, 101750.4, 101808.7, 
    101847,
  100042.4, 100106, 100234.5, 100358.1, 100474.5, 100575.4, 100689.3, 
    100798.2, 100898.6, 101005.9, 101115.8, 101210.6, 101303.5, 101381.6, 
    101444.5,
  100047.9, 100120.9, 100224, 100342.9, 100463.7, 100546.3, 100653.5, 
    100762.9, 100870.3, 100977.2, 101100.6, 101203.1, 101298.2, 101379.3, 
    101448.6,
  100086.7, 100141, 100239.2, 100337.5, 100453.9, 100541.1, 100640.2, 
    100735.2, 100850, 100956.7, 101088.6, 101197.8, 101293.5, 101378, 101449,
  100118.1, 100167.2, 100267.2, 100353, 100460.7, 100550.1, 100638.3, 
    100704.4, 100836.9, 100935.5, 101080, 101194.6, 101302.5, 101387.3, 
    101461.6,
  100152.4, 100202.5, 100292.8, 100370.5, 100464.4, 100549.9, 100641.9, 
    100693.7, 100819.1, 100914.4, 101063.7, 101185.5, 101299.6, 101389, 
    101465.9,
  100193.9, 100245.7, 100328.9, 100393, 100473.3, 100570.5, 100648.5, 
    100686.1, 100804, 100897.5, 101045, 101176.7, 101299.4, 101395.3, 101475.3,
  100243.9, 100296.6, 100364.6, 100411.2, 100493.8, 100591.6, 100644.7, 
    100693, 100802.7, 100890.7, 101036.8, 101171.4, 101299.4, 101404, 101488.9,
  100302.7, 100351.1, 100406.9, 100439.1, 100510.6, 100605.8, 100658.4, 
    100703.8, 100808.1, 100898.3, 101036.4, 101173.9, 101305.4, 101415.4, 
    101502.7,
  100358.2, 100407.4, 100449, 100470.4, 100530.1, 100630.1, 100685.2, 
    100725.4, 100815.8, 100917.8, 101047, 101185, 101316.5, 101428.8, 101516.6,
  100413, 100459.6, 100497.8, 100506.1, 100546.9, 100644.6, 100686.7, 
    100752.8, 100834.5, 100947.1, 101070.4, 101207.8, 101335.1, 101446.4, 
    101534.4,
  99976.87, 100116.6, 100273.3, 100417.9, 100567.3, 100709.6, 100840.6, 
    100952.7, 101052.4, 101137.4, 101215.1, 101277.9, 101329.3, 101374.1, 
    101425.6,
  99970.72, 100107.2, 100257.7, 100400.2, 100548.8, 100690, 100822.7, 
    100940.8, 101043.9, 101131.8, 101208.6, 101273.2, 101333.3, 101382.1, 
    101433.3,
  99984.36, 100097.4, 100235.7, 100375.8, 100521.4, 100664.6, 100799, 
    100919.3, 101024.1, 101116.5, 101196.8, 101265.5, 101323.4, 101381.5, 
    101434.2,
  99994.31, 100102.4, 100238.1, 100373.4, 100511.4, 100654, 100791, 100915.9, 
    101026.6, 101122, 101204.9, 101276.1, 101337.4, 101393.6, 101447.7,
  100009, 100111.1, 100234.5, 100366.6, 100501.5, 100643.9, 100780, 100904.2, 
    101017.8, 101112.9, 101199, 101270.9, 101337.2, 101395.4, 101452.1,
  100030.1, 100123, 100240.2, 100363.5, 100494.7, 100635.2, 100771.2, 
    100898.4, 101013.1, 101109.6, 101194.4, 101269.8, 101341.8, 101403.3, 
    101460.7,
  100052.6, 100139.1, 100250.1, 100362.4, 100491.4, 100628.8, 100764.2, 
    100889.2, 101004.9, 101098.8, 101186.1, 101266.1, 101344.5, 101403.8, 
    101468.9,
  100077, 100156.7, 100261.3, 100368.2, 100494.5, 100626.2, 100756.2, 
    100880.8, 100992.8, 101091.9, 101178.7, 101263.6, 101345.3, 101409, 
    101480.7,
  100101.5, 100164.9, 100269.2, 100370.6, 100498.5, 100626.2, 100751.7, 
    100869.5, 100978.7, 101077.1, 101162, 101256.6, 101340, 101416.7, 101486.8,
  100115, 100172, 100274.5, 100374.8, 100502.3, 100624.7, 100744.9, 100854.7, 
    100962.4, 101059.5, 101142.6, 101244.7, 101332.8, 101417.1, 101492.1,
  99974.81, 100039.3, 100173.5, 100275.8, 100380.6, 100498.8, 100643.4, 
    100789.4, 100913.9, 101033.4, 101144.8, 101244.3, 101336.3, 101416, 
    101487.7,
  99968.98, 100041.8, 100174, 100275, 100375.8, 100497.8, 100653.5, 100796.7, 
    100923.8, 101042.2, 101156, 101259.7, 101351.9, 101435.9, 101507.2,
  100006.6, 100075.8, 100202.8, 100309, 100407.1, 100514.7, 100681.4, 100815, 
    100947, 101066.4, 101182.8, 101286, 101375.3, 101461.4, 101531.2,
  100025.8, 100102.7, 100225, 100332.3, 100428.5, 100526.3, 100704.9, 
    100833.8, 100969.8, 101090, 101208.2, 101315.5, 101405.6, 101493.5, 
    101560.7,
  100048, 100139.1, 100262, 100368.3, 100465.7, 100554.4, 100734.7, 100862.6, 
    101001.5, 101119.2, 101237.7, 101345.9, 101435.7, 101518.1, 101587.5,
  100078.4, 100177.5, 100307.6, 100403.3, 100509.4, 100590.3, 100762.6, 
    100892.5, 101031.2, 101151.1, 101271.3, 101375.6, 101467.2, 101549.1, 
    101620.1,
  100122, 100226.8, 100364.4, 100455.1, 100560.1, 100642.3, 100797.8, 
    100925.9, 101065.8, 101187.1, 101311.3, 101413.2, 101506.4, 101584.9, 
    101650.2,
  100182.5, 100291.3, 100426.4, 100522.5, 100616.3, 100700, 100834.2, 
    100957.7, 101098.4, 101223.8, 101353.3, 101454.3, 101546.3, 101618.2, 
    101683.6,
  100264.1, 100368.2, 100493.8, 100579.5, 100666.9, 100758.9, 100879.4, 
    100994.5, 101131.5, 101259.8, 101394.1, 101494, 101583.1, 101651, 101720.8,
  100360.8, 100451.9, 100566.1, 100627.2, 100719.7, 100818.7, 100929.5, 
    101039.2, 101162.7, 101301.3, 101427, 101531.1, 101620, 101694.7, 101756.2,
  99790.18, 100000.1, 100208.2, 100399.4, 100568.8, 100720.6, 100849.3, 
    100961.7, 101064, 101158.9, 101260, 101361.1, 101452.3, 101534.9, 101612.1,
  99735.1, 99942.41, 100153.5, 100340.6, 100517.5, 100673.2, 100803.9, 
    100919.6, 101029.5, 101130.6, 101237.3, 101345.1, 101442.6, 101529.5, 
    101611.8,
  99698.41, 99950.58, 100157.7, 100343.6, 100525.1, 100674, 100807.4, 
    100929.3, 101040.8, 101147.8, 101253.3, 101362.5, 101460.9, 101554.8, 
    101634.5,
  99700.39, 99953.24, 100144.6, 100333.3, 100504.5, 100652.7, 100785.6, 
    100909.4, 101026.4, 101139.9, 101250.4, 101361.9, 101469.1, 101566.5, 
    101650.9,
  99731.79, 99970.95, 100147.2, 100340.3, 100503.8, 100652.9, 100789.9, 
    100918.6, 101039, 101154.7, 101270.1, 101384, 101495.5, 101596.2, 101680.2,
  99779.57, 99996.38, 100166, 100343.6, 100505.1, 100655.4, 100792.5, 
    100926.2, 101043.4, 101170.2, 101288.2, 101404.7, 101521.9, 101626.4, 
    101710.8,
  99826.61, 100027.8, 100183.7, 100356.6, 100511.7, 100672, 100812.4, 
    100947.7, 101071.5, 101202.2, 101312.8, 101440.6, 101560.8, 101665.1, 
    101748.7,
  99888.21, 100068.2, 100207, 100374.7, 100542.9, 100695.9, 100837.3, 
    100976.1, 101104.5, 101235.4, 101346.4, 101482.9, 101600, 101706.3, 
    101791.4,
  99968.35, 100128.1, 100248.7, 100419, 100578.5, 100725.9, 100878.4, 
    101022.5, 101158.9, 101264.3, 101396.9, 101533.7, 101649, 101756.7, 
    101837.3,
  100061.9, 100207.9, 100329.8, 100489.8, 100633.5, 100785.1, 100932.9, 
    101082, 101194.1, 101318.1, 101453.9, 101587.7, 101704.6, 101808.2, 
    101886.1,
  101851.5, 101946.1, 102028, 102099.4, 102160.3, 102220.8, 102262.5, 
    102295.8, 102329.1, 102333.7, 102336.2, 102330.2, 102329.4, 102315.5, 
    102305.4,
  101806, 101907, 101987.3, 102061.6, 102128.8, 102186, 102237.1, 102272, 
    102305.9, 102316.3, 102321, 102319.9, 102325.7, 102312.2, 102306.4,
  101747.8, 101852.7, 101930.4, 102011.8, 102078.6, 102143.5, 102202.5, 
    102241.4, 102275.2, 102293.7, 102310.9, 102315.7, 102322.3, 102317.1, 
    102304.5,
  101697.7, 101808.2, 101890.6, 101973.3, 102045, 102115.1, 102175.2, 
    102217.1, 102260, 102283.8, 102295.5, 102313.1, 102313.2, 102313.2, 
    102301.1,
  101641.7, 101763.3, 101846.2, 101935.1, 102003.5, 102081, 102139.5, 
    102185.8, 102233.8, 102263.2, 102285.5, 102301.5, 102307.3, 102311.9, 
    102298.8,
  101595, 101720.8, 101807.6, 101901.4, 101972.6, 102048.7, 102112.8, 102161, 
    102206.4, 102248.2, 102267.1, 102288.8, 102297.1, 102307.3, 102298.2,
  101549.8, 101679.5, 101769.2, 101872.1, 101945.1, 102019.1, 102082.3, 
    102132, 102176.9, 102226, 102252, 102274.9, 102288.5, 102301.6, 102302,
  101513.5, 101640.1, 101739, 101845.8, 101919.9, 101993.7, 102055.2, 
    102101.6, 102148.8, 102198.9, 102232.3, 102254.2, 102277, 102296, 102306.7,
  101478.8, 101608, 101712.2, 101824.1, 101892.4, 101961.9, 102019, 102070.1, 
    102114.2, 102172.1, 102208.1, 102236.7, 102269.1, 102295.6, 102316.1,
  101455.8, 101584.1, 101695.5, 101799.6, 101863.5, 101926, 101986.2, 
    102035.9, 102086.8, 102141.7, 102183.3, 102225.1, 102260.5, 102296.2, 
    102327.1,
  102467, 102580.4, 102671.8, 102746.8, 102799, 102834.9, 102857.6, 102861.4, 
    102855.2, 102836.5, 102812, 102774.6, 102733.2, 102678.1, 102618.5,
  102462, 102579.7, 102676.5, 102752.9, 102812.5, 102856.5, 102882.7, 
    102887.5, 102884.4, 102866.3, 102845.4, 102812.2, 102766.9, 102714.9, 
    102651.5,
  102467.5, 102584.5, 102684.4, 102766.5, 102831.5, 102878.7, 102905.6, 
    102918.4, 102911.4, 102895.8, 102869.9, 102840.6, 102796.8, 102744.6, 
    102681,
  102469.1, 102588.9, 102692.5, 102777.9, 102846.4, 102896.7, 102928.5, 
    102944.2, 102938.3, 102923.5, 102897.1, 102868.7, 102825, 102772, 102709,
  102476, 102596, 102701.9, 102789.3, 102859.7, 102907.9, 102942.3, 102960.3, 
    102960.5, 102943.1, 102920.5, 102889.3, 102846.9, 102795.1, 102734.2,
  102481.9, 102602.8, 102710.6, 102800.1, 102871.3, 102920.2, 102957.1, 
    102972.5, 102977.8, 102963.9, 102942.2, 102911.3, 102871.2, 102819.5, 
    102757.7,
  102489, 102610, 102719.6, 102810.5, 102880.7, 102932, 102968.3, 102986, 
    102992, 102978.9, 102962.2, 102924.6, 102890.8, 102840.6, 102780.2,
  102492.1, 102614.3, 102724.2, 102817.1, 102886.6, 102940.2, 102979.6, 
    102998.6, 103006.5, 102995, 102977, 102943.6, 102906.6, 102860.4, 102804.8,
  102496.8, 102616.9, 102728, 102820.4, 102892.7, 102950.5, 102989, 103010.7, 
    103016.9, 103007.9, 102989.4, 102962, 102924.4, 102873.8, 102825.7,
  102498.4, 102617.4, 102729.2, 102819.2, 102894.2, 102953.1, 102996.8, 
    103017.4, 103026.6, 103018.6, 103002.2, 102974.6, 102937.5, 102887.6, 
    102843.7,
  102432, 102544.9, 102642.5, 102723.1, 102781.9, 102825.4, 102850.3, 
    102860.3, 102850.7, 102826.4, 102790.8, 102747.9, 102699.2, 102657.7, 
    102615.1,
  102412.9, 102533.9, 102637.6, 102726.3, 102796.8, 102845.8, 102879, 
    102888.6, 102884.3, 102865.6, 102836.7, 102795.4, 102739.9, 102696.5, 
    102649.9,
  102400.6, 102527.5, 102636.6, 102733.7, 102808.1, 102864.5, 102896.5, 
    102904.5, 102906.5, 102893.1, 102869.5, 102840.7, 102781.1, 102730.4, 
    102684.6,
  102379.2, 102513.1, 102630, 102730.3, 102811.7, 102876.6, 102910.5, 
    102932.3, 102938.6, 102930.5, 102904.7, 102876, 102828.5, 102769.2, 
    102716.1,
  102353.7, 102495.5, 102619.3, 102725.2, 102815.2, 102885.1, 102927.4, 
    102954.2, 102960.6, 102958.1, 102941.5, 102911.2, 102859.9, 102810.6, 
    102749,
  102325.9, 102473.3, 102606.2, 102718, 102816.9, 102890.3, 102938.7, 
    102971.8, 102985.1, 102980.6, 102966, 102942.6, 102903.8, 102846.7, 
    102783.3,
  102293.1, 102449.6, 102591.7, 102708.9, 102813.4, 102892.3, 102946.6, 
    102986.4, 103007.3, 103010.4, 102994.6, 102966.6, 102931.2, 102881.1, 
    102817.9,
  102257.5, 102424, 102573.4, 102697.5, 102808.1, 102890.3, 102950.5, 102996, 
    103020.3, 103017.5, 103009.5, 102986.7, 102959.8, 102917.5, 102852.6,
  102222.2, 102396.7, 102553.3, 102684.5, 102799.3, 102884.8, 102952.1, 
    103000.6, 103031.3, 103038.9, 103034.7, 103013.4, 102984.5, 102936.9, 
    102886.2,
  102183, 102367.6, 102530, 102668.5, 102786.9, 102877.7, 102950, 103000.6, 
    103037.6, 103045.9, 103047.3, 103029.6, 102999.4, 102963.7, 102915.5,
  102203.5, 102308, 102399.6, 102475.2, 102538.3, 102584, 102620.5, 102642.7, 
    102641.9, 102638.6, 102619.5, 102597, 102568.6, 102538.4, 102501,
  102207.9, 102316.6, 102410.7, 102492, 102563.1, 102620.6, 102661.4, 
    102685.2, 102688.4, 102680.3, 102664.8, 102639.9, 102607.9, 102574.2, 
    102534,
  102216.5, 102331.3, 102428.2, 102512.6, 102588.6, 102648.3, 102689.5, 
    102717.5, 102727.7, 102728.3, 102708.4, 102684.2, 102655.6, 102618.3, 
    102577.4,
  102215.9, 102336.8, 102440.9, 102527.2, 102605.4, 102668.9, 102719.8, 
    102756.2, 102774, 102773.3, 102758.5, 102731.8, 102699.6, 102660.1, 
    102613.3,
  102212.4, 102339.9, 102450.7, 102540.1, 102620.2, 102689.3, 102744.6, 
    102784.7, 102803.2, 102807.1, 102799.5, 102778.6, 102746.9, 102709, 
    102657.9,
  102200.8, 102336.5, 102454.9, 102549.5, 102634, 102704, 102761.5, 102805.1, 
    102829.3, 102837.1, 102833.6, 102816.8, 102788.3, 102750, 102703.5,
  102181.7, 102327.7, 102455.8, 102555.1, 102642.5, 102715.6, 102779.3, 
    102828.7, 102854.4, 102866.4, 102864.4, 102849.3, 102826.4, 102793.5, 
    102745.8,
  102152.4, 102311.9, 102449, 102558.2, 102646.6, 102723.2, 102789.8, 
    102837.7, 102868.1, 102887.5, 102885.8, 102874.1, 102854.9, 102826.4, 
    102785.5,
  102117.3, 102287.6, 102434.1, 102550.3, 102645.6, 102726.2, 102796.9, 
    102848.6, 102883.9, 102903.6, 102905.5, 102899.7, 102880.4, 102853.4, 
    102820.3,
  102076.5, 102257.8, 102410.3, 102538.7, 102637.2, 102723.9, 102799.2, 
    102853, 102894.7, 102917.5, 102926.5, 102920.6, 102902.4, 102877.6, 102844,
  102281.2, 102363, 102437.6, 102493.9, 102534.5, 102563.3, 102577, 102583.5, 
    102575.6, 102562.1, 102541.8, 102509.5, 102467.9, 102422.5, 102373.5,
  102287.4, 102371.3, 102455.4, 102522.9, 102572.5, 102602, 102621.4, 
    102631.5, 102627.5, 102615.7, 102591.9, 102560.6, 102520.3, 102473, 
    102423.2,
  102297.8, 102393, 102483.8, 102555.1, 102608.6, 102644.2, 102669.3, 
    102680.5, 102683.8, 102667.9, 102646.1, 102615.2, 102574.4, 102526.3, 
    102474.4,
  102301.2, 102401.9, 102497, 102575.8, 102637.3, 102680.4, 102708.4, 
    102728.8, 102733.1, 102721.4, 102697.4, 102667.6, 102627.4, 102579.3, 
    102522.9,
  102305, 102408.9, 102511.3, 102594.9, 102662.5, 102717.1, 102755.4, 
    102775.4, 102787.1, 102771.4, 102749.5, 102718.8, 102677.2, 102631.7, 
    102573.1,
  102302, 102410.6, 102516.3, 102608.2, 102683.8, 102746.6, 102789.7, 
    102818.3, 102829.3, 102819.1, 102798.5, 102767.2, 102725.8, 102682, 
    102625.6,
  102294.9, 102409.2, 102518.7, 102616.4, 102701, 102768.2, 102818.5, 
    102852.7, 102867.3, 102866.1, 102844.3, 102809.3, 102774.5, 102730.5, 
    102678.9,
  102286.1, 102401.7, 102515.2, 102618.8, 102709.5, 102785.1, 102843.7, 
    102882.7, 102897.7, 102901.3, 102883.8, 102853, 102815.7, 102777.3, 
    102730.6,
  102273.4, 102391, 102507.8, 102616.5, 102713.6, 102793.9, 102858.3, 
    102903.2, 102930.6, 102936.3, 102919.6, 102892.5, 102859.2, 102818.3, 
    102772,
  102254.2, 102374, 102494.6, 102608.2, 102709.5, 102795.2, 102870.9, 
    102922.8, 102952.6, 102959.7, 102949.7, 102924.1, 102893.8, 102860.9, 
    102813.8,
  102261.7, 102317.9, 102366.3, 102405, 102435.7, 102456, 102462.1, 102459.2, 
    102445.8, 102426.6, 102404.3, 102376.8, 102344.7, 102308.4, 102266.1,
  102338.2, 102395.1, 102442.7, 102482.5, 102513.4, 102531.7, 102537.3, 
    102531.8, 102517.6, 102497.2, 102471.3, 102439.3, 102401.9, 102362.8, 
    102318.2,
  102417.8, 102474.7, 102521.6, 102560.4, 102591, 102607, 102609.1, 102602.9, 
    102588.6, 102569.5, 102541.9, 102505.8, 102465.2, 102420.4, 102373.8,
  102490.3, 102546, 102594.4, 102630.4, 102661.9, 102676.7, 102681.2, 
    102675.4, 102662.3, 102642.6, 102613.1, 102574.9, 102528.6, 102477.3, 
    102427.8,
  102561.5, 102614.8, 102666.1, 102699.9, 102728.1, 102746.6, 102752.6, 
    102749.6, 102735.1, 102710.9, 102679.9, 102641.7, 102594.4, 102538.7, 
    102483.3,
  102622.5, 102676.8, 102730, 102767.4, 102796.6, 102810.9, 102820.8, 
    102819.9, 102805.4, 102771.9, 102740.1, 102703, 102655.8, 102601.2, 
    102543.2,
  102676.4, 102737.9, 102792.7, 102830.4, 102859.9, 102878.7, 102892.6, 
    102892.5, 102877.1, 102842.5, 102804.9, 102766.3, 102717.8, 102662.8, 
    102603.8,
  102722.5, 102788.2, 102846.7, 102888.8, 102924.1, 102944.8, 102957.5, 
    102962.1, 102946.1, 102916.5, 102871.1, 102830.3, 102777.9, 102722.8, 
    102665.1,
  102767.7, 102832.6, 102894.6, 102939.5, 102974.9, 102999.9, 103016, 
    103019.7, 103008.4, 102982.7, 102936.9, 102890.4, 102838.1, 102779.3, 
    102722.9,
  102803.1, 102865.7, 102929.2, 102977, 103020.2, 103051.1, 103065.7, 
    103068.5, 103058.6, 103034, 102996.7, 102944.2, 102888.8, 102832.1, 
    102773.4,
  101583.6, 101686.2, 101791.8, 101879.6, 101950.4, 102025, 102090.6, 
    102134.9, 102173.2, 102198.3, 102213.1, 102214.3, 102207.9, 102194.1, 
    102170.4,
  101594.1, 101718.8, 101826.9, 101921.4, 101993.5, 102070.4, 102131.8, 
    102179.2, 102216.5, 102240.4, 102254, 102255.2, 102250.2, 102230.9, 
    102206.6,
  101647.9, 101773, 101879.4, 101978.4, 102046.4, 102122.9, 102182.7, 102232, 
    102266.5, 102287.6, 102298.6, 102297.7, 102289.1, 102270.2, 102247.6,
  101703.1, 101827, 101943, 102037.5, 102108.2, 102187.3, 102243, 102290.8, 
    102321.7, 102341.1, 102348.4, 102349.3, 102337.2, 102315.9, 102285.7,
  101769.9, 101892.2, 102009.9, 102094.6, 102174.8, 102249.1, 102304, 102351, 
    102381.4, 102399.8, 102406.4, 102403.5, 102388.7, 102366.6, 102336,
  101836.8, 101966.2, 102076, 102161.9, 102247.3, 102316.8, 102373.9, 
    102418.5, 102446.2, 102462.9, 102467.4, 102461.4, 102443, 102419.4, 
    102384.9,
  101915.2, 102047, 102149, 102243.9, 102323.1, 102392.4, 102446.8, 102486, 
    102509.7, 102522.5, 102523.5, 102515.7, 102496, 102466.9, 102435.4,
  102008.1, 102136.1, 102235.8, 102333.5, 102408.7, 102474.4, 102523.7, 
    102557.5, 102575.9, 102583.6, 102579.1, 102569.4, 102547.1, 102514.5, 
    102478,
  102108.2, 102229.4, 102327.9, 102418.4, 102489.1, 102550.5, 102595.3, 
    102629.8, 102647.6, 102650.3, 102639.8, 102621.9, 102594.2, 102561.2, 
    102520.3,
  102211.4, 102327.5, 102417.4, 102502.4, 102567.6, 102624.7, 102662.8, 
    102691.2, 102701.3, 102705.1, 102695.4, 102676.1, 102643.6, 102607.6, 
    102564.4,
  101842.8, 101832.9, 101845.7, 101875.8, 101880.7, 101932.2, 102010.8, 
    102079.3, 102118.4, 102157.3, 102178.3, 102181.1, 102173.5, 102158.4, 
    102135.6,
  101837, 101862.4, 101870.7, 101894.6, 101905.4, 101949.3, 102027.8, 
    102080.7, 102139, 102183.1, 102199.8, 102205.9, 102200.3, 102184.1, 
    102162.4,
  101883.8, 101898.8, 101888.1, 101916.6, 101927.3, 101945.4, 102050.9, 
    102098.4, 102164.2, 102201.4, 102226.4, 102236.2, 102231.2, 102214.7, 
    102196,
  101909, 101929.8, 101909, 101936.7, 101948, 101962.6, 102077.4, 102119.2, 
    102189.4, 102225.5, 102255.3, 102263.4, 102260.1, 102245.4, 102222.3,
  101943, 101959.5, 101930.9, 101947.8, 101967.7, 101996.8, 102105.9, 
    102142.8, 102217.6, 102250.9, 102284.6, 102294.8, 102293.7, 102276.4, 
    102253.1,
  101983.5, 101976.3, 101964.4, 101977.8, 102008.5, 102035, 102135.2, 
    102176.6, 102249.6, 102280.9, 102314.9, 102323.5, 102328.2, 102315.2, 
    102287.4,
  102012.1, 101999.6, 102012.7, 102014.1, 102057.1, 102084.8, 102176.4, 
    102217, 102282, 102313.1, 102345.9, 102359.5, 102363.4, 102345.4, 102320.5,
  102031.7, 102037.9, 102046, 102053.1, 102106, 102128.5, 102220, 102257.9, 
    102319.4, 102348.2, 102378.2, 102389.7, 102394.6, 102375.3, 102345.2,
  102054.8, 102081.3, 102076.7, 102108.2, 102150.6, 102184.6, 102275.6, 
    102311.8, 102366.1, 102393.2, 102416, 102423.6, 102421.6, 102399.6, 
    102372.7,
  102090.9, 102125.7, 102130.8, 102163.3, 102207.2, 102252.7, 102328.8, 
    102357.7, 102409.2, 102431.8, 102454.1, 102451, 102443.7, 102423.2, 
    102391.9,
  100691.3, 100763.6, 100911.4, 101052.6, 101213.6, 101367.1, 101501.9, 
    101607.4, 101690.9, 101749.7, 101795.7, 101827.9, 101852.4, 101871.5, 
    101875.4,
  100679.1, 100773, 100904.1, 101047.9, 101208.9, 101371.2, 101514.3, 
    101623.5, 101706.3, 101768.4, 101813.1, 101849.2, 101875.7, 101893.7, 
    101903.1,
  100699.4, 100798.3, 100929.1, 101069.9, 101227.5, 101388.7, 101526.8, 
    101639.6, 101728.9, 101793.4, 101842.1, 101875.1, 101901, 101917.3, 
    101927.5,
  100707.2, 100825.2, 100953.1, 101091.5, 101248.5, 101406.4, 101542.6, 
    101663.3, 101751.8, 101820.6, 101867.2, 101899.4, 101926.6, 101944.8, 
    101957.2,
  100727.9, 100862.5, 100977.8, 101126.3, 101268.7, 101424.7, 101560.4, 
    101684.2, 101771.8, 101846.2, 101889.8, 101929.9, 101953.9, 101973.1, 
    101981.4,
  100757.4, 100890.1, 101003.7, 101155.4, 101293.9, 101450.2, 101588.2, 
    101712.4, 101804.9, 101878.7, 101929, 101969.1, 101987.4, 101996.8, 
    101998.4,
  100802, 100921, 101044.3, 101189.5, 101331.8, 101486.4, 101622, 101740.6, 
    101835.4, 101908, 101957.3, 101991.9, 102013.8, 102028.8, 102022.8,
  100851.1, 100952.4, 101101.1, 101235.1, 101383.7, 101531.5, 101662.3, 
    101776.7, 101872.8, 101939.4, 101989.5, 102027.3, 102047, 102062, 102063.4,
  100908.9, 101006.7, 101166.8, 101292.2, 101443.8, 101585.4, 101709, 
    101818.1, 101907.7, 101971.2, 102016.3, 102050.1, 102076.6, 102088.9, 
    102093.2,
  100976.5, 101073.9, 101239, 101358.1, 101509.2, 101646.2, 101763.5, 101867, 
    101948.2, 102005.1, 102053.2, 102087.7, 102105.7, 102120.1, 102124.2,
  99911.81, 100035.6, 100194.2, 100378.9, 100570.7, 100744.4, 100910.6, 
    101062.3, 101197.4, 101313.1, 101408.8, 101488.3, 101557.3, 101622.9, 
    101672.3,
  99845.77, 99973.11, 100107.7, 100290.7, 100475, 100663.2, 100837.1, 
    100996.7, 101148.4, 101277.8, 101385.9, 101474, 101550.8, 101616.4, 
    101672.8,
  99805.54, 99910.85, 100051.8, 100223.8, 100412.3, 100605.1, 100786.7, 
    100956.2, 101113.7, 101251.6, 101368.1, 101466.5, 101551.1, 101623.7, 
    101684.6,
  99770.18, 99855.58, 100001.1, 100167, 100357.4, 100544.6, 100735.3, 100913, 
    101081.6, 101231.4, 101358.3, 101462.6, 101552.6, 101629.7, 101691.5,
  99752.31, 99809.85, 99974.76, 100133.5, 100327.2, 100505, 100699, 100880.7, 
    101057.9, 101213.8, 101348.1, 101458, 101554.7, 101634.9, 101700.5,
  99738.05, 99787.72, 99960.49, 100122.8, 100314.8, 100480.2, 100670.3, 
    100855.3, 101038.4, 101200, 101342.2, 101458.1, 101563, 101647, 101716.6,
  99733.47, 99798.04, 99964.48, 100133.3, 100323.6, 100483.8, 100664.7, 
    100847.8, 101030, 101197.2, 101341.5, 101464.8, 101571.6, 101658.9, 
    101731.5,
  99747.66, 99825.28, 99983.64, 100160.7, 100345.7, 100504.9, 100673.9, 
    100852.7, 101031, 101200.5, 101347.8, 101475.1, 101586, 101676.4, 101751.2,
  99781.02, 99880.09, 100022.8, 100205.2, 100378.9, 100541.5, 100703.6, 
    100877.8, 101050.6, 101217.9, 101366.1, 101500.2, 101612.7, 101703.2, 
    101775.7,
  99833.41, 99945.55, 100079.8, 100260.5, 100424.2, 100587.9, 100746.5, 
    100916.4, 101082.2, 101247.9, 101397.4, 101529.6, 101639.6, 101730.3, 
    101803.5,
  101241.1, 101307.8, 101412.7, 101495.3, 101563.9, 101623.6, 101665.5, 
    101699.8, 101721.5, 101735.7, 101742, 101740.2, 101736.5, 101732.1, 
    101749.2,
  101168.4, 101282.4, 101389.8, 101484.4, 101559.3, 101621.6, 101670.3, 
    101708.8, 101735.7, 101753.5, 101759.7, 101760.3, 101759, 101759.6, 
    101769.7,
  101106.5, 101221.8, 101341, 101444.5, 101533.5, 101606.1, 101664.9, 101709, 
    101740.9, 101763.3, 101773.7, 101771.7, 101768.9, 101775.9, 101776.6,
  101013.5, 101143.2, 101287.2, 101405.6, 101508.9, 101593, 101658.9, 
    101710.6, 101749.1, 101774.6, 101791.9, 101791.3, 101785.1, 101795.1, 
    101793.3,
  100885.5, 101039.8, 101201.6, 101339.2, 101458.1, 101556.2, 101633.5, 
    101695, 101745.1, 101774.7, 101799.5, 101804.5, 101798.2, 101799.9, 
    101808.8,
  100733.8, 100906.2, 101089.5, 101254.2, 101391.8, 101508.5, 101604.1, 
    101677.1, 101734.9, 101774.5, 101804.7, 101815, 101813.3, 101816.5, 
    101820.2,
  100567.4, 100758.1, 100962.9, 101146.8, 101312.7, 101449.7, 101561.9, 
    101648.5, 101718, 101767.8, 101805.9, 101821.1, 101823.2, 101828.4, 
    101831.4,
  100388.8, 100604.8, 100830.8, 101032.9, 101218.9, 101378.4, 101512.1, 
    101614.5, 101697.1, 101758.4, 101801.5, 101825.9, 101832.5, 101841.4, 
    101849,
  100225.8, 100459.9, 100695.6, 100915, 101121.2, 101301.4, 101452.8, 101574, 
    101669.4, 101741.3, 101791.9, 101824.6, 101836.4, 101855.6, 101863.5,
  100095.4, 100325.5, 100563.7, 100801.9, 101021, 101219.2, 101386.7, 101526, 
    101635.1, 101720.2, 101779, 101819, 101839.7, 101860.2, 101877.2,
  100126.2, 100314.8, 100487.9, 100646, 100802.9, 100941.4, 101069, 101177.7, 
    101270.1, 101348.8, 101421.1, 101489.8, 101553, 101601.8, 101641.9,
  100107.6, 100275.4, 100458.3, 100622.6, 100778.7, 100918.1, 101046.8, 
    101159.8, 101253.2, 101334.5, 101404.5, 101477, 101542.2, 101597.8, 
    101647.8,
  100128.4, 100304.6, 100487.3, 100638.2, 100796, 100927.6, 101047.7, 
    101150.3, 101249.8, 101336.8, 101413.3, 101485.8, 101548, 101603, 101653.6,
  100156.1, 100328.1, 100497.4, 100649.1, 100801.5, 100923.6, 101041.6, 
    101144.2, 101246.5, 101332.1, 101409.1, 101480.8, 101543.5, 101604.7, 
    101659.6,
  100211.3, 100374.1, 100534.7, 100683.7, 100821.8, 100944, 101056.7, 
    101159.2, 101260.8, 101348.8, 101427, 101495.7, 101556.3, 101616.2, 
    101673.9,
  100273.4, 100429.6, 100583.3, 100722.3, 100853.6, 100969.5, 101077.7, 
    101182.5, 101280, 101368.6, 101444.9, 101509.9, 101568.5, 101629.9, 101696,
  100346.5, 100495.9, 100641.5, 100774.1, 100898.9, 101008.2, 101117.4, 
    101218.6, 101314.3, 101401.6, 101473.5, 101537.7, 101593.4, 101661, 101726,
  100428, 100565.4, 100701.6, 100828.1, 100945.3, 101051.5, 101160.1, 
    101258.2, 101354.8, 101435.9, 101502.2, 101563.5, 101625, 101690.2, 
    101752.8,
  100512.4, 100637, 100766.6, 100883.4, 100995.4, 101103.5, 101208.3, 
    101308.5, 101402, 101474.8, 101538.9, 101602.2, 101666, 101729.1, 101788,
  100598.9, 100711.4, 100835.3, 100941.2, 101052.7, 101156.8, 101260.8, 
    101363.8, 101452.9, 101519.1, 101582.5, 101650.1, 101712, 101770.6, 
    101827.7,
  100631.7, 100743.1, 100855.3, 100976.2, 101094.7, 101213.4, 101337.1, 
    101450, 101545.3, 101629.7, 101696.3, 101754, 101797.7, 101831.9, 101854.5,
  100534.2, 100655.6, 100774.4, 100900.3, 101020.3, 101144.5, 101259.5, 
    101374.9, 101474.9, 101571, 101643.7, 101703.5, 101753.6, 101793.1, 
    101819.4,
  100445.7, 100568.8, 100682.9, 100809.6, 100938.1, 101061.8, 101188.2, 
    101309, 101418.3, 101516.2, 101598, 101663.5, 101719.5, 101763.5, 101795.7,
  100371.5, 100491.3, 100609.4, 100741.9, 100870.6, 100995.2, 101122.5, 
    101241.9, 101357, 101458.5, 101546.4, 101617.3, 101677.8, 101725.9, 
    101762.4,
  100298.2, 100418.5, 100535.8, 100667.7, 100801.2, 100928.9, 101058.6, 
    101177.5, 101298, 101406.9, 101498.8, 101577.8, 101643.2, 101695.9, 
    101735.1,
  100235.3, 100350.9, 100473.9, 100607.3, 100737.8, 100871.4, 100996.4, 
    101121.1, 101241.4, 101349.7, 101451.8, 101536.5, 101610.7, 101661.9, 
    101705.2,
  100178, 100289.4, 100414.6, 100549.8, 100682.5, 100813.6, 100941, 101068.6, 
    101188, 101303.5, 101409.7, 101506.3, 101578.8, 101628.3, 101676.2,
  100119.4, 100236.6, 100363.4, 100496, 100630.8, 100764.4, 100888.6, 101018, 
    101136.5, 101256.1, 101369.7, 101471.5, 101538.4, 101591, 101648.9,
  100061.4, 100190.8, 100315.1, 100450, 100582.8, 100714.6, 100843.5, 
    100972.6, 101090.5, 101217.9, 101340.7, 101432.3, 101498.8, 101559.5, 
    101624.8,
  100009.8, 100150.7, 100272.2, 100407.7, 100538.8, 100672.8, 100804.9, 
    100933.7, 101054.1, 101194.4, 101302.3, 101388.5, 101459.8, 101532.7, 
    101603.2,
  100348.3, 100564.3, 100793, 101003.2, 101190.1, 101351.6, 101494.3, 
    101611.7, 101708.5, 101786.8, 101851.1, 101888.7, 101917.5, 101929.3, 
    101929,
  100258.2, 100502.6, 100733.5, 100941.5, 101139, 101315.2, 101460.3, 
    101587.1, 101696, 101778.6, 101847.3, 101886.3, 101911.2, 101926.3, 
    101934.4,
  100228.8, 100464.6, 100683.2, 100896.8, 101095.8, 101271.4, 101425.5, 
    101558.8, 101669.7, 101763.5, 101840.9, 101880.8, 101913.2, 101928.7, 
    101935.9,
  100194, 100431.5, 100656.3, 100868.1, 101068.1, 101252, 101412.8, 101550.8, 
    101666.2, 101763.7, 101839.5, 101880.1, 101911.2, 101930, 101935.9,
  100167.4, 100411.3, 100638.7, 100848.4, 101045.8, 101228.8, 101389, 
    101528.7, 101647.1, 101746.5, 101822.9, 101874.1, 101907.3, 101927.8, 
    101936.8,
  100151.4, 100398.8, 100627.2, 100836.9, 101035.1, 101217.4, 101378.2, 
    101518.6, 101637.4, 101742.8, 101820.9, 101876.1, 101907.7, 101930.2, 
    101940.8,
  100148.7, 100396, 100622.9, 100832.9, 101031.2, 101212, 101371.1, 101510.4, 
    101629.2, 101734.6, 101813.9, 101870.1, 101904.2, 101930.7, 101942,
  100160.2, 100405, 100626.3, 100836.5, 101032.4, 101214.3, 101372.6, 
    101509.6, 101629, 101730.5, 101811.1, 101871.4, 101907.3, 101930.6, 
    101947.9,
  100183.5, 100422, 100635.6, 100842.5, 101039.2, 101218.7, 101375.1, 
    101511.5, 101628.8, 101730.3, 101811.3, 101871.5, 101911.6, 101935.8, 
    101950.9,
  100213.9, 100451.6, 100656.2, 100858.3, 101048.2, 101226.1, 101380.3, 
    101516.6, 101633.8, 101734.5, 101815, 101875.9, 101915.4, 101939.4, 
    101955.5,
  99812.53, 99981.09, 100167.6, 100342.6, 100531, 100709.9, 100878.5, 
    101030.6, 101172.5, 101291.3, 101396.5, 101482.2, 101554.1, 101605.8, 
    101644.5,
  99801.02, 99984.23, 100173.5, 100346.6, 100526.1, 100714.5, 100885.7, 
    101042.9, 101185.9, 101305.5, 101415.8, 101505.5, 101573.8, 101625.4, 
    101668.6,
  99850.79, 100023.5, 100209.7, 100370.2, 100560.4, 100747.5, 100918.1, 
    101077.4, 101219.4, 101341.8, 101449.2, 101532.4, 101597.6, 101652.6, 
    101696.4,
  99891.62, 100063.9, 100247.6, 100413.6, 100599.6, 100785.2, 100956.2, 
    101114.2, 101252.1, 101372.9, 101478.2, 101557.5, 101623.3, 101677, 101720,
  99932.3, 100113.2, 100302.1, 100471.3, 100656.2, 100837.4, 101001.6, 
    101152.6, 101288.2, 101403.9, 101504.4, 101586.5, 101652, 101705.3, 
    101748.7,
  99970.23, 100163.2, 100358.3, 100537.6, 100718.8, 100894.4, 101053.3, 
    101196.3, 101328.9, 101441.9, 101543.1, 101624.9, 101688.5, 101737.6, 
    101781.3,
  100016.8, 100223.6, 100424.9, 100615.1, 100788.9, 100959.7, 101111.1, 
    101250.1, 101377.9, 101489.6, 101583.8, 101661, 101720.7, 101774, 101811.5,
  100075.8, 100295.7, 100496.9, 100690.4, 100859.1, 101024.1, 101171.6, 
    101306.4, 101431.2, 101538.6, 101627.4, 101699.3, 101760.5, 101811.6, 
    101843.1,
  100151.6, 100374, 100574.1, 100768.1, 100930.5, 101088.2, 101232.1, 
    101367.1, 101489, 101590.8, 101672.5, 101744.3, 101806, 101848.1, 101879.2,
  100237.5, 100452.4, 100651.8, 100838.5, 100999, 101150.9, 101296.3, 
    101429.3, 101547.7, 101643.7, 101727.1, 101797, 101852.7, 101893.2, 
    101923.3,
  99451.16, 99587.04, 99731.44, 99816.57, 99925.51, 100024.2, 100149.9, 
    100270.2, 100413.4, 100556.5, 100682.2, 100807.2, 100933, 101045.4, 
    101147.6,
  99414.78, 99561.61, 99682.12, 99782.02, 99871.15, 99970.26, 100109.3, 
    100248.5, 100403.2, 100544.1, 100681.4, 100813.1, 100937.8, 101053.4, 
    101163.4,
  99393.43, 99585, 99686.92, 99815.88, 99840.89, 99976.52, 100115.6, 
    100259.6, 100419.4, 100565.2, 100712.9, 100844.4, 100975.2, 101094, 
    101200.2,
  99398.16, 99594.47, 99672.08, 99802.12, 99796.5, 99957.99, 100095.3, 
    100261.5, 100421.5, 100578.2, 100733.1, 100870.5, 101004.3, 101126.3, 
    101230.3,
  99437.96, 99607.51, 99687.24, 99789.78, 99805.78, 99958.08, 100105.4, 
    100282.7, 100444.3, 100611.1, 100769.1, 100915.9, 101048.5, 101170.9, 
    101269.7,
  99485.67, 99623.7, 99700.15, 99769.53, 99806.97, 99966.52, 100126, 
    100307.8, 100470.9, 100646.8, 100808, 100960.2, 101097.5, 101214.8, 
    101307.2,
  99543.4, 99633.2, 99727.12, 99759.49, 99844.35, 99995.37, 100174.1, 
    100345.7, 100516, 100696.7, 100865.5, 101021.3, 101154, 101265, 101353,
  99607.49, 99652.11, 99762.06, 99756.03, 99893.59, 100035.1, 100224.8, 
    100389.7, 100569.8, 100755.7, 100929.1, 101084, 101213, 101318.8, 101403.6,
  99657.51, 99672.87, 99794.28, 99797.09, 99949.73, 100090.8, 100279.5, 
    100447.3, 100643.2, 100830.2, 101006.6, 101156.8, 101280.8, 101380.1, 
    101460.6,
  99676.26, 99699.23, 99801.99, 99856.85, 100009.5, 100158.6, 100347.2, 
    100526.3, 100728.1, 100912.7, 101089, 101232.2, 101351.4, 101444.5, 
    101521.8,
  100242.1, 100329.1, 100422.7, 100505.8, 100591.1, 100676.1, 100752.3, 
    100831.9, 100900.5, 100978.6, 101056.4, 101123.3, 101176.8, 101222.2, 
    101264.3,
  100157.4, 100249.9, 100349.6, 100438.1, 100522.1, 100602.6, 100676.5, 
    100746, 100817.2, 100906.1, 100982.5, 101052.2, 101113.3, 101165.7, 
    101213.4,
  100089.2, 100188.9, 100283.8, 100368.9, 100446.8, 100532.2, 100607.8, 
    100680.5, 100758, 100847, 100928.8, 101006.1, 101066.2, 101120.1, 101174.7,
  100030.8, 100134.7, 100226.7, 100313.3, 100390.1, 100469.1, 100537.9, 
    100617.7, 100696.6, 100789.2, 100870.9, 100951.3, 101014.8, 101072.1, 
    101133.7,
  99985.75, 100090.4, 100181.7, 100262.2, 100338.2, 100410.6, 100475.7, 
    100564.9, 100653.2, 100739, 100823.5, 100900.8, 100969.2, 101025.6, 
    101095.4,
  99954.57, 100059.6, 100151.9, 100226.7, 100296.8, 100359.9, 100426.5, 
    100515.8, 100608.1, 100691.3, 100768, 100850.2, 100920.7, 100981.5, 
    101059.6,
  99937.37, 100040.6, 100134, 100203.6, 100261.9, 100324.4, 100390.1, 
    100480.8, 100568.3, 100642.6, 100723.4, 100805.8, 100878.6, 100947.3, 
    101032.1,
  99929.84, 100031.6, 100121.2, 100192.5, 100246.7, 100303.5, 100365.9, 
    100446.4, 100521.7, 100597.8, 100678.7, 100759.9, 100840.4, 100918.5, 
    101008.8,
  99927.54, 100030.3, 100110, 100192.3, 100245.2, 100291.3, 100346, 100413.9, 
    100484.2, 100551.6, 100636.1, 100720.9, 100814.1, 100899.4, 100998.4,
  99944.16, 100035.1, 100116.3, 100202.8, 100237.3, 100286.5, 100322.6, 
    100382, 100444.8, 100518.1, 100600.7, 100692.7, 100795.9, 100890.4, 
    100997.6,
  101570.8, 101626.4, 101694, 101765.4, 101817.6, 101868.8, 101906.5, 
    101938.8, 101959.8, 101973.4, 101977.6, 101976.9, 101965, 101953, 101931.1,
  101541, 101608.3, 101684.1, 101746, 101801.4, 101852.1, 101890.8, 101926.3, 
    101951.8, 101969.3, 101976.8, 101982.8, 101975.7, 101964.9, 101948.9,
  101522.2, 101580.1, 101650.6, 101719.1, 101777.3, 101829.8, 101872, 
    101909.9, 101934.4, 101957.4, 101969.4, 101977.4, 101972.8, 101962.6, 
    101949.5,
  101477.9, 101542.6, 101621.2, 101688.4, 101749.2, 101803.1, 101849.5, 
    101888.9, 101921.9, 101946.3, 101964.9, 101972.7, 101974.5, 101966, 
    101955.4,
  101416.8, 101490, 101567.5, 101637.6, 101703.8, 101761.7, 101813.8, 
    101857.6, 101894.9, 101924.2, 101946.5, 101959.2, 101963.6, 101959.7, 
    101952.4,
  101344.7, 101420.8, 101499.2, 101576.8, 101646.6, 101713.4, 101769.3, 
    101822.9, 101863.2, 101898.7, 101925.2, 101942.1, 101953.2, 101952.8, 
    101948,
  101259.9, 101339.2, 101419.1, 101501.9, 101578.8, 101649.8, 101714.7, 
    101772.1, 101823.2, 101862.2, 101896.8, 101918.9, 101935.7, 101940.5, 
    101939.4,
  101167.9, 101252.1, 101328.9, 101416.6, 101498.8, 101578.6, 101649.4, 
    101713.4, 101772.2, 101820.8, 101862.3, 101890.5, 101913.8, 101925.4, 
    101928.7,
  101072.5, 101160.1, 101239.1, 101325, 101409.1, 101497.5, 101575.7, 
    101645.9, 101714.1, 101771.4, 101821.1, 101857.4, 101885.2, 101906, 
    101913.2,
  100973.3, 101060.1, 101141, 101228.3, 101315.2, 101407.2, 101494.6, 
    101573.2, 101648.2, 101713.5, 101771.8, 101816.9, 101852.2, 101879.8, 
    101892.5,
  101029.6, 101052.8, 101149.1, 101227.9, 101332, 101427.9, 101517.3, 
    101592.8, 101656.2, 101709.4, 101751.2, 101788.4, 101820.4, 101840.9, 
    101853.9,
  100981.4, 101025.4, 101133.1, 101221.8, 101326.6, 101425.1, 101514.4, 
    101591.7, 101664.2, 101716.5, 101763.1, 101798.4, 101827.9, 101849.8, 
    101865.9,
  100953.2, 101032.4, 101132.1, 101230.4, 101341.8, 101444.4, 101537.3, 
    101615.6, 101683.4, 101739.6, 101784.9, 101824.6, 101855.1, 101880.3, 
    101896.9,
  100942.6, 101044.1, 101138.5, 101249.7, 101359.6, 101463, 101554, 101634.1, 
    101699.5, 101760.1, 101807.9, 101848.7, 101877.9, 101902.3, 101915.1,
  100940.8, 101072.3, 101162.3, 101285.5, 101390.5, 101492.6, 101583, 
    101666.8, 101732.9, 101793.6, 101841.1, 101880.3, 101909.5, 101933.1, 
    101945,
  100957.4, 101117.1, 101202.5, 101334.8, 101430.2, 101534.4, 101620.6, 
    101705, 101769.2, 101829.3, 101875.1, 101913.6, 101943.4, 101963.8, 
    101974.7,
  101011.1, 101180.6, 101259.3, 101393.6, 101485.9, 101587.2, 101672.3, 
    101754, 101818.1, 101875.4, 101921.7, 101960.3, 101986.5, 102001.3, 
    102009.3,
  101101.2, 101257.5, 101338.7, 101466.4, 101550.8, 101652.7, 101732.1, 
    101809.7, 101871.8, 101925, 101970.6, 102006.3, 102029.7, 102042.3, 
    102044.6,
  101228.1, 101352.1, 101437.2, 101550.8, 101631.4, 101725.9, 101795.1, 
    101868.3, 101927.4, 101978.2, 102023.6, 102055.5, 102075, 102084.2, 
    102080.9,
  101357.3, 101452.9, 101537.5, 101635.5, 101713, 101796.6, 101861.2, 
    101927.5, 101983.6, 102033.3, 102074, 102102.3, 102119.3, 102122.3, 
    102116.7,
  101511.1, 101637.7, 101749.4, 101844, 101921.4, 101982, 102031.8, 102066.5, 
    102090.9, 102097.1, 102093.8, 102083.4, 102067.2, 102044.3, 102020.7,
  101494.6, 101623.1, 101731.1, 101826.7, 101906.2, 101970.6, 102021.6, 
    102056.7, 102078.1, 102091, 102091.8, 102085.5, 102074.1, 102054.9, 
    102032.5,
  101490, 101608.4, 101712.8, 101806, 101887.5, 101950.3, 102002.4, 102039.8, 
    102065.5, 102076.9, 102078.3, 102075.1, 102060.3, 102043.8, 102023.2,
  101468.3, 101586.7, 101696.9, 101792.5, 101873.9, 101937.8, 101990.7, 
    102028, 102050, 102062, 102066.6, 102063, 102053.2, 102038.3, 102020.2,
  101447.2, 101558.8, 101670.5, 101763.1, 101844.3, 101911.2, 101961.6, 
    101997.7, 102023.1, 102037.9, 102043.8, 102041.6, 102037.2, 102021.7, 
    102009.3,
  101419.7, 101529.1, 101642.7, 101734.7, 101816.6, 101882.7, 101935.8, 
    101972.2, 101996.8, 102010.9, 102016.4, 102017.8, 102014.3, 102005.2, 
    101997,
  101389.6, 101501.8, 101612.5, 101703.8, 101785.1, 101850.1, 101903.4, 
    101938.7, 101960.3, 101976.7, 101983.9, 101987.6, 101986.8, 101984.6, 
    101979.4,
  101351.2, 101462.6, 101576.1, 101666.8, 101749, 101813, 101864.5, 101904.5, 
    101927.9, 101944.3, 101954.1, 101957.6, 101959.7, 101961.7, 101963.6,
  101302.3, 101420.2, 101531.7, 101622.8, 101705.9, 101772.9, 101827.2, 
    101867.7, 101895.5, 101915.2, 101922.4, 101927.9, 101932.2, 101937.1, 
    101941.2,
  101256.8, 101381.9, 101490.6, 101584.1, 101667.5, 101736.3, 101793.7, 
    101834.9, 101866.7, 101883.9, 101900.4, 101902.6, 101909.4, 101916.3, 
    101926.2,
  101067.4, 101241.9, 101401.3, 101539.8, 101660.8, 101759.3, 101845, 101911, 
    101964.4, 102003.1, 102029.2, 102041.8, 102043.9, 102038.4, 102031.2,
  101051.4, 101248.9, 101418.6, 101555.5, 101678.2, 101780.8, 101869.2, 
    101940.6, 101996.1, 102033.6, 102059.6, 102070.8, 102070, 102063.2, 
    102052.2,
  101119.9, 101291.2, 101445.4, 101586.3, 101710.8, 101810.2, 101898.6, 
    101965.3, 102019.2, 102055.3, 102079.3, 102089, 102089, 102081.2, 102068.5,
  101167.4, 101331.1, 101488.9, 101625.3, 101739.7, 101840.5, 101925, 
    101994.6, 102047.9, 102083.8, 102105.1, 102113.3, 102111.2, 102101.2, 
    102086.9,
  101225.4, 101384.7, 101536.3, 101661.8, 101773.1, 101868.2, 101952, 
    102020.1, 102073, 102109.8, 102127.2, 102133.9, 102130.3, 102119.1, 
    102103.5,
  101284.2, 101435.9, 101581.2, 101702.7, 101810.7, 101903.8, 101984.5, 
    102051.6, 102102.6, 102135.6, 102152.7, 102156, 102150.3, 102136.7, 
    102119.7,
  101345, 101489.2, 101630.3, 101746.8, 101852.4, 101939.6, 102015.9, 
    102077.9, 102127.2, 102158.5, 102174.1, 102176.4, 102168.5, 102151.8, 
    102132,
  101409.8, 101544.5, 101680.4, 101792, 101892.2, 101975.4, 102048.7, 
    102108.9, 102153.4, 102181.9, 102192.5, 102194, 102182.5, 102163.8, 102141,
  101474.3, 101601, 101729.4, 101835.8, 101932, 102012.8, 102081, 102135.7, 
    102176.3, 102200.2, 102208.7, 102206.5, 102192.2, 102172.2, 102146.2,
  101538, 101656.4, 101777.9, 101878.4, 101968.8, 102044.8, 102109.2, 
    102161.2, 102197.3, 102214.7, 102221.2, 102213.3, 102196.3, 102174.1, 
    102146.8,
  100493.9, 100577.6, 100721.3, 100816.2, 100930, 101042.9, 101152, 101261.9, 
    101357.5, 101441.1, 101513.1, 101580.3, 101634.2, 101680.9, 101726.6,
  100415.8, 100516.2, 100662.1, 100761.5, 100875.9, 100988.3, 101102, 
    101216.8, 101319.3, 101412.3, 101489.7, 101561.5, 101622, 101676.9, 
    101722.4,
  100361.4, 100484.2, 100620.1, 100727.5, 100844.8, 100961.7, 101081.2, 
    101191.9, 101299.8, 101395.6, 101478.6, 101552.1, 101618.7, 101674, 
    101721.1,
  100328.3, 100450.7, 100585, 100697.5, 100816.7, 100936.6, 101058.2, 
    101180.1, 101291.9, 101389.5, 101475.1, 101551.6, 101618.9, 101678.7, 
    101732,
  100318.4, 100435.2, 100567.9, 100682.9, 100807.4, 100928.9, 101051.7, 
    101175.3, 101288.9, 101386.5, 101477.7, 101553.3, 101621.7, 101685.5, 
    101739.2,
  100321.2, 100433.3, 100570.3, 100686.8, 100811.8, 100929.7, 101051.1, 
    101179.6, 101296.1, 101396.5, 101484.7, 101564.5, 101632.6, 101697.2, 
    101753.9,
  100337, 100451.6, 100587.8, 100706.1, 100832.3, 100947.5, 101073.2, 
    101201.2, 101316, 101416.7, 101502.1, 101580.2, 101650.8, 101715.7, 
    101772.8,
  100364.8, 100481, 100623.3, 100744.9, 100867.3, 100984.5, 101109.7, 
    101235.2, 101346.6, 101444, 101526.6, 101606.9, 101675.2, 101737.6, 
    101790.1,
  100417.2, 100532.2, 100675.5, 100791.3, 100915, 101036.2, 101162.2, 
    101282.6, 101380.1, 101477.8, 101562.8, 101639.2, 101704.3, 101762.3, 
    101812.3,
  100482.2, 100600.7, 100740.5, 100856.4, 100981.6, 101101.1, 101218.8, 
    101324.6, 101427.9, 101522.9, 101603.1, 101675.4, 101738.5, 101793.2, 
    101836.1,
  101651.2, 101707.4, 101774, 101838.9, 101892.4, 101939.1, 101975.1, 
    102003.1, 102014.7, 102021.2, 102015.3, 102004.2, 101986.9, 101968.1, 
    101934.3,
  101613.1, 101678.9, 101746.5, 101805.2, 101859.9, 101907.1, 101945.5, 
    101978.1, 102001.3, 102010.8, 102010.6, 102006, 101997.8, 101969.7, 
    101944.2,
  101575.6, 101637.1, 101695.8, 101753.4, 101809.5, 101859.7, 101900.4, 
    101932.9, 101956.7, 101972.4, 101981.3, 101981.4, 101975.8, 101963.4, 
    101942.7,
  101537.5, 101592.6, 101658, 101721.9, 101774, 101826.4, 101866.2, 101901.7, 
    101929.1, 101952.5, 101965.6, 101969.4, 101970.5, 101961.3, 101943.4,
  101490.3, 101543.8, 101606.2, 101668, 101724.4, 101772.3, 101813.3, 101848, 
    101881.7, 101907.7, 101930.4, 101937.2, 101944.8, 101945.5, 101934.3,
  101443.3, 101494, 101551.9, 101610.3, 101672.7, 101720.4, 101761.8, 
    101796.9, 101832.8, 101862.5, 101892.2, 101907.4, 101925.2, 101930, 
    101923.8,
  101395.8, 101440.8, 101492.3, 101545.4, 101607.9, 101658.1, 101696, 
    101731.9, 101769.3, 101805.1, 101844.8, 101867.3, 101893.9, 101907.8, 
    101907.7,
  101346.9, 101387.9, 101431.8, 101480.6, 101536.8, 101589.7, 101625, 
    101660.2, 101704, 101747.9, 101793.5, 101824.8, 101855.1, 101881.1, 
    101887.2,
  101302.6, 101330, 101368.3, 101413.2, 101466.3, 101514.1, 101546.3, 
    101582.4, 101634.2, 101682.1, 101731.7, 101773.8, 101810.7, 101847, 
    101863.1,
  101261, 101273.2, 101308.6, 101343.1, 101385.2, 101427.6, 101466.2, 
    101511.8, 101560.5, 101608, 101666.3, 101718.6, 101766.7, 101808.1, 
    101836.5,
  100587.7, 100774.1, 100914.6, 101049.2, 101157.2, 101248.8, 101331.1, 
    101407.9, 101474.5, 101537.7, 101582.9, 101625.5, 101653.9, 101675, 
    101687.4,
  100710.9, 100894.9, 101019.8, 101139, 101240.2, 101330.6, 101411.6, 
    101486.4, 101549.8, 101604.8, 101650, 101684, 101711.8, 101725.1, 101732.6,
  100870.6, 101020.1, 101134.2, 101243.9, 101339.8, 101423.4, 101501.7, 
    101568.9, 101625.3, 101673.7, 101714.7, 101745, 101769.5, 101775.6, 
    101780.8,
  101022.7, 101149.9, 101259.8, 101358.7, 101442.8, 101522.9, 101596.2, 
    101655.6, 101708.3, 101751.4, 101786.4, 101813.5, 101827.5, 101833.1, 
    101833.7,
  101168.3, 101282.1, 101384, 101472.9, 101554.2, 101629.7, 101694.6, 
    101749.3, 101795.4, 101831.2, 101860.7, 101879, 101889.2, 101888.2, 
    101884.6,
  101305.7, 101406.9, 101500.8, 101584, 101664.1, 101730.6, 101790, 101837.4, 
    101879.4, 101909.7, 101936.6, 101951.2, 101956.4, 101951.4, 101941.4,
  101440.4, 101527.4, 101619.2, 101697, 101769.7, 101828.9, 101882.9, 
    101925.4, 101961, 101986.7, 102006.6, 102017.4, 102018, 102012, 101995.2,
  101566.7, 101643.5, 101730.1, 101799.9, 101865.4, 101920.9, 101968.5, 
    102007.3, 102038.8, 102061.6, 102077.5, 102085.3, 102081.2, 102074.1, 
    102053.3,
  101683.1, 101753.8, 101831.7, 101896.4, 101957.3, 102007.1, 102050.2, 
    102083.8, 102111, 102130.1, 102143.2, 102146.6, 102140.4, 102130, 102107.9,
  101789.3, 101852.1, 101922.7, 101981.5, 102035.5, 102081.5, 102120.9, 
    102151.6, 102175.1, 102190.3, 102200.1, 102203, 102195.4, 102184.5, 
    102160.4,
  100149.8, 100286.9, 100443, 100569.1, 100680.1, 100787.2, 100869.7, 100935, 
    100995.5, 101057.6, 101114.9, 101186.2, 101255.8, 101320.9, 101369.2,
  100080.1, 100226.2, 100383.5, 100517.5, 100642, 100751, 100838.8, 100912, 
    100980.8, 101052.1, 101120.2, 101200.6, 101269.4, 101337.4, 101392.5,
  100047, 100216.2, 100368.2, 100501.1, 100624.5, 100741.5, 100829.3, 100907, 
    100987, 101068.8, 101131.6, 101220.2, 101297.6, 101376.4, 101428.7,
  100033.8, 100197.7, 100332.8, 100471.8, 100600.3, 100717.7, 100812.2, 
    100903.8, 100988.9, 101084.1, 101154.6, 101247.1, 101330.4, 101409.9, 
    101468.2,
  100036.2, 100188.2, 100319, 100462, 100583.9, 100704.3, 100810.1, 100909, 
    101003.3, 101106.6, 101179.3, 101275.5, 101362.2, 101446.2, 101510,
  100059.5, 100195.9, 100328.9, 100457.7, 100578.7, 100700.8, 100810.4, 
    100921.2, 101028.2, 101136.4, 101209.6, 101307.5, 101402.9, 101488.6, 
    101554.5,
  100102.8, 100217.5, 100353.7, 100473, 100592.9, 100709.2, 100828.9, 
    100942.1, 101063.7, 101171.5, 101245.5, 101348.3, 101442.8, 101533.3, 
    101596.7,
  100160.2, 100262, 100399.7, 100513.5, 100626.6, 100734.6, 100854.9, 
    100973.6, 101112.6, 101211.4, 101288.8, 101392.4, 101488.2, 101580.3, 
    101645.9,
  100238, 100334.1, 100462.6, 100580.7, 100679.7, 100780.4, 100891.3, 
    101016.5, 101167.3, 101253.7, 101340.4, 101442.9, 101543.5, 101633.4, 
    101695.2,
  100339.3, 100431.5, 100550.3, 100667.3, 100758.3, 100847.4, 100946, 
    101073.2, 101224.7, 101305.1, 101404.1, 101501.5, 101606.6, 101687.7, 
    101751.4,
  99348.19, 99474.01, 99590.03, 99711.38, 99831.59, 99950.94, 100071.1, 
    100186.9, 100306, 100426, 100536.4, 100650, 100758, 100866.1, 100959.7,
  99529.9, 99638.59, 99726.8, 99832.66, 99935.5, 100044.3, 100151.5, 100262, 
    100370.2, 100480.4, 100591.7, 100708.1, 100816.1, 100924.2, 101019.6,
  99698.59, 99789.36, 99876.68, 99972.92, 100067.2, 100163.4, 100261.3, 
    100356.2, 100454.6, 100559.2, 100666.9, 100781.8, 100894.5, 101000.7, 
    101088.4,
  99863.36, 99951.1, 100030.5, 100110.8, 100191.7, 100278.6, 100361.6, 
    100449.9, 100543, 100645.4, 100746.6, 100863.9, 100973.4, 101069.6, 
    101150.6,
  100029.4, 100110.8, 100178.8, 100255.1, 100327.4, 100401, 100477.6, 100563, 
    100650.8, 100754.3, 100850, 100955.8, 101055.2, 101144.9, 101221.1,
  100188.1, 100264.2, 100332.9, 100404, 100468.5, 100536.5, 100606.5, 
    100685.6, 100768.7, 100867.3, 100950.6, 101042.8, 101136.4, 101219.2, 
    101290.6,
  100350, 100426.6, 100490.2, 100557.3, 100619.4, 100681.1, 100745.3, 
    100818.5, 100895.5, 100984.4, 101056.1, 101132.7, 101217.5, 101295.9, 
    101363.3,
  100525.9, 100593.5, 100652.9, 100714.1, 100767.5, 100820.9, 100879, 
    100948.9, 101020.8, 101099, 101158.1, 101221.3, 101299.4, 101372.2, 
    101437.1,
  100698.6, 100757.3, 100810.9, 100863.7, 100911.4, 100958.6, 101012.7, 
    101071.3, 101144.4, 101209.5, 101256.9, 101310.2, 101380.6, 101449.7, 
    101509.8,
  100859.7, 100909.3, 100957, 101000.9, 101045.3, 101086.1, 101130.5, 
    101180.9, 101257.1, 101305.8, 101344.7, 101397.4, 101459.8, 101526.5, 
    101581.1,
  99723.67, 99903.55, 100095.5, 100255.6, 100416.1, 100558.7, 100688.3, 
    100802, 100901, 100993, 101083.4, 101164.2, 101222.4, 101271.2, 101316.8,
  99704.91, 99879.6, 100063, 100224, 100378.3, 100515.2, 100643.9, 100758.3, 
    100866.3, 100963.7, 101051.6, 101130.8, 101194.9, 101246.2, 101294.8,
  99714.91, 99893.8, 100068, 100227.7, 100377.7, 100511.2, 100643.9, 
    100758.4, 100872.8, 100971.6, 101056.5, 101129.6, 101182.4, 101232.8, 
    101290,
  99729.48, 99899.66, 100060.9, 100217.6, 100355.4, 100494.1, 100620.9, 
    100738.7, 100848.8, 100947.5, 101033.5, 101095.8, 101156.9, 101216.9, 
    101284.6,
  99757.62, 99926.09, 100070.7, 100223, 100360.9, 100494.9, 100618.2, 
    100735.9, 100841.9, 100934.9, 101014.2, 101082.9, 101148, 101216.5, 
    101294.4,
  99814.21, 99964.21, 100095, 100235.3, 100363.1, 100490.8, 100610, 100726.1, 
    100825.1, 100919.1, 101001.7, 101077.2, 101147.5, 101226, 101308.9,
  99878.91, 100001.5, 100123.6, 100248.2, 100376.8, 100497.5, 100616.3, 
    100727, 100824.9, 100921.8, 101007, 101088.5, 101165.3, 101251.7, 101335.9,
  99945.71, 100044.9, 100156.7, 100279.1, 100396.4, 100518.8, 100632.9, 
    100739.2, 100839.2, 100934.3, 101027.6, 101112, 101196, 101283, 101377.1,
  100014.1, 100101.3, 100213.6, 100331.3, 100452.6, 100564.9, 100667, 
    100773.1, 100869.5, 100973.3, 101067.1, 101154.4, 101242.4, 101330.7, 
    101429.3,
  100095.3, 100193.5, 100304.1, 100419.6, 100520.7, 100623.2, 100723.8, 
    100829.2, 100930.6, 101029.8, 101124.6, 101213.8, 101300, 101395.2, 
    101484.6,
  101281.3, 101362.4, 101438.5, 101501.4, 101569.4, 101632.1, 101690.3, 
    101741.5, 101783, 101810.5, 101840.2, 101859.5, 101880.9, 101891.5, 
    101895.1,
  101322.2, 101404.6, 101481, 101544.7, 101610.1, 101663.8, 101717, 101762.8, 
    101808.4, 101838.6, 101859.1, 101881.8, 101895.2, 101907.9, 101906,
  101363.2, 101445.6, 101523.3, 101589.8, 101650, 101702.9, 101756.4, 
    101795.6, 101834.7, 101863.8, 101882.8, 101903.9, 101912.2, 101927.6, 
    101925.6,
  101407.5, 101490.8, 101574, 101636.1, 101694.8, 101749, 101795.6, 101836.3, 
    101871.9, 101902.3, 101918.6, 101932.7, 101938.9, 101948.4, 101945.4,
  101449.3, 101530, 101612.5, 101677.4, 101740.7, 101789.8, 101836.5, 
    101872.5, 101904.8, 101933.1, 101944.5, 101961.1, 101961.2, 101966, 101963,
  101490.8, 101571.5, 101656.6, 101720.4, 101781.8, 101829.4, 101876.1, 
    101911.2, 101940.5, 101969.4, 101976.8, 101987.3, 101988.4, 101988.7, 
    101987.1,
  101528.6, 101612.8, 101698.1, 101764.1, 101822.8, 101870.5, 101912.5, 
    101946.4, 101972.5, 101998.9, 102008.9, 102015.6, 102011.3, 102006.3, 
    102003.1,
  101560.8, 101648.8, 101734.3, 101802.8, 101861.3, 101909.4, 101946.5, 
    101978.6, 102004.3, 102025.8, 102032.7, 102039.2, 102034.7, 102028.9, 
    102015.4,
  101589.1, 101682.5, 101768.5, 101837, 101896.8, 101942.5, 101978.3, 
    102008.8, 102028.8, 102048.8, 102052.6, 102057.7, 102056.3, 102042.1, 
    102030,
  101613.8, 101710, 101793.1, 101865.8, 101924.8, 101975, 102006.8, 102033.3, 
    102052.2, 102069.2, 102068.8, 102069.3, 102072.7, 102044.2, 102053.6,
  101419.5, 101506.1, 101603.6, 101679.7, 101747.7, 101802, 101848.1, 
    101885.1, 101911.2, 101929.8, 101943, 101965.7, 101975.3, 101976.6, 101979,
  101378.4, 101478, 101579.6, 101658.9, 101737.4, 101798.8, 101844.8, 
    101887.7, 101922, 101941.2, 101959.4, 101968.5, 101977.5, 101982.3, 
    101986.6,
  101363, 101450.6, 101544.4, 101630.7, 101715.3, 101781.2, 101834.5, 101878, 
    101912.4, 101936.4, 101953.3, 101967.5, 101979.8, 101979.4, 101981.4,
  101345.3, 101428.1, 101527.1, 101616.1, 101702.6, 101772.1, 101833.4, 
    101878.6, 101917.9, 101942.6, 101962.2, 101973, 101984.2, 101981.7, 
    101985.3,
  101329.1, 101409.4, 101504.9, 101590.7, 101676.4, 101748.1, 101812, 
    101860.7, 101901.9, 101929.8, 101950, 101963.2, 101974.8, 101980.6, 
    101982.1,
  101319.5, 101395.7, 101485.4, 101571.4, 101656.5, 101731.4, 101797.7, 
    101850.3, 101892.9, 101924.8, 101947.5, 101963.6, 101974, 101980.1, 
    101982.1,
  101316.8, 101389.5, 101476.9, 101557.8, 101640, 101713.3, 101782.5, 
    101836.8, 101880.3, 101909.6, 101939.2, 101953.9, 101968.7, 101976.8, 
    101980.3,
  101329, 101394.8, 101478.8, 101556.1, 101634.1, 101705, 101774.4, 101827.6, 
    101868.4, 101903.4, 101933.8, 101950.7, 101962, 101975.7, 101975.7,
  101352.9, 101412.7, 101491.2, 101560.5, 101637.2, 101705.2, 101768.6, 
    101822.3, 101860, 101891.1, 101918.5, 101939.7, 101952.4, 101960.3, 
    101965.4,
  101388.9, 101443.6, 101512.3, 101578.2, 101649.5, 101715.4, 101776.3, 
    101820.4, 101850.4, 101883.1, 101906.9, 101930, 101939.8, 101941.9, 
    101956.9,
  100669.8, 100771.6, 100889.4, 100994.6, 101107.2, 101200.8, 101298.2, 
    101387.4, 101476, 101546.8, 101613.1, 101668.4, 101718.5, 101755.4, 
    101778.2,
  100642.1, 100764, 100896.2, 101000.8, 101111.2, 101203.9, 101287.8, 
    101375.6, 101455.7, 101530.6, 101593.6, 101653.7, 101704.2, 101746.1, 
    101770.7,
  100658.1, 100767.4, 100874.8, 100975.3, 101083.4, 101185.4, 101281.4, 
    101370.4, 101452.1, 101522.7, 101589.6, 101644.9, 101694.1, 101737.2, 
    101765.4,
  100668.7, 100789, 100899.4, 101000.7, 101103.5, 101201.9, 101296.5, 
    101384.7, 101468.5, 101537.7, 101599.2, 101651.8, 101698.2, 101739.8, 
    101762.1,
  100691.2, 100809, 100907.6, 101013.1, 101106.5, 101209.4, 101299.2, 
    101390.9, 101472.8, 101543.4, 101603.5, 101653, 101695.6, 101736.6, 
    101756.9,
  100726.2, 100839, 100935.5, 101033.1, 101124.9, 101221.4, 101315.5, 
    101399.9, 101484.8, 101557.3, 101619.2, 101665.8, 101706, 101738.5, 
    101759.9,
  100772.7, 100878, 100967.5, 101059.7, 101144.5, 101237.3, 101325.8, 
    101413.1, 101492.8, 101567.9, 101632.9, 101676.9, 101714.4, 101741.3, 
    101762.2,
  100827.3, 100923.9, 101010.5, 101095.1, 101176, 101259.5, 101346.6, 
    101427.7, 101506.9, 101580.9, 101643.6, 101690.7, 101727.5, 101748.4, 
    101764.4,
  100885.5, 100972.8, 101054.2, 101133.3, 101210.5, 101287.3, 101362.2, 
    101444.6, 101517.3, 101588, 101650.1, 101696.1, 101733.5, 101754.8, 
    101764.6,
  100949.4, 101027, 101107.4, 101180.2, 101252.4, 101320.7, 101387.4, 
    101458.9, 101528.2, 101596.6, 101652.1, 101697.6, 101732.8, 101758.1, 
    101765.6,
  99720.2, 99878.04, 100070.6, 100245.7, 100410.1, 100552.3, 100667.2, 
    100797.3, 100905.8, 101026.5, 101136.3, 101234.6, 101319.3, 101390.8, 
    101448.8,
  99595.58, 99794.96, 99990.4, 100165.5, 100337.3, 100488.2, 100611.8, 
    100750.2, 100877.7, 100986.3, 101103.5, 101208, 101297.5, 101372.3, 
    101433.9,
  99567.84, 99762.32, 99931.78, 100109.5, 100275.3, 100436.4, 100561.6, 
    100693.6, 100829.4, 100949.7, 101071.7, 101181.5, 101275.5, 101354.6, 
    101420.3,
  99512.12, 99701.61, 99881.38, 100055.7, 100221.3, 100387.2, 100521.9, 
    100650.5, 100788.6, 100924.4, 101045.8, 101161.1, 101258.7, 101340.4, 
    101408,
  99468.49, 99663.29, 99834.84, 100014.3, 100174.5, 100341.7, 100483.6, 
    100609.7, 100744.2, 100888.5, 101014.1, 101135, 101235.5, 101318.7, 
    101391.1,
  99429.54, 99622.05, 99786.43, 99968.8, 100128.5, 100300.1, 100448.4, 
    100576.5, 100708, 100851.5, 100985.1, 101108.1, 101213.5, 101301.5, 
    101377.3,
  99407.27, 99586.8, 99750.49, 99931.54, 100093.4, 100261.7, 100416.3, 
    100544, 100678.6, 100818.3, 100961.4, 101084.2, 101190.4, 101283.8, 
    101362.9,
  99386.69, 99558.97, 99720.04, 99897.42, 100057.2, 100227.7, 100385.7, 
    100517.2, 100653.8, 100791.2, 100935, 101057.7, 101170.3, 101268.4, 
    101348.9,
  99371.99, 99534.48, 99695.25, 99867.96, 100031.1, 100198.7, 100358.8, 
    100491.4, 100630.1, 100767.6, 100910.8, 101035.1, 101150.6, 101252.9, 
    101338,
  99360.3, 99514.96, 99673.24, 99845.48, 100003.9, 100173, 100334.6, 
    100467.4, 100609.8, 100747.1, 100889.9, 101015.7, 101135.9, 101238.9, 
    101327.1,
  99157.64, 99302.55, 99491.04, 99674.84, 99857.27, 100040, 100205, 100362.2, 
    100498.5, 100644.7, 100772.3, 100896.3, 101004.7, 101109.4, 101200.1,
  99068.55, 99227.91, 99399.66, 99581.02, 99766.19, 99946.55, 100117.3, 
    100277.8, 100413.1, 100562.6, 100699.3, 100828.3, 100945.6, 101056.5, 
    101156.8,
  98994.73, 99146.67, 99314.23, 99498.06, 99681.65, 99865.96, 100033.6, 
    100202.6, 100353.7, 100496.7, 100640.8, 100775.2, 100899.8, 101016.5, 
    101124,
  98918.03, 99072.23, 99246.08, 99428.04, 99612.58, 99791.22, 99957.05, 
    100130.4, 100291.5, 100434.9, 100587.8, 100728.5, 100857, 100982.8, 101096,
  98835.09, 99000.25, 99177.92, 99360.8, 99550.29, 99723.91, 99887.51, 
    100065.1, 100236.8, 100390.7, 100541.5, 100685, 100818.9, 100949.7, 
    101068.7,
  98751.01, 98928.8, 99115.3, 99304.73, 99495.55, 99659.5, 99826.51, 
    100001.1, 100178.3, 100346.5, 100491.1, 100649.1, 100784, 100919.2, 
    101043.5,
  98675.91, 98864.7, 99058.29, 99257.69, 99447.95, 99611.53, 99776.65, 
    99950.99, 100132.8, 100309.8, 100457.7, 100617.3, 100753.6, 100895.2, 
    101023,
  98629.6, 98812.79, 99022.92, 99222.36, 99412.88, 99571.96, 99732.76, 
    99906.75, 100094, 100268.7, 100428.7, 100588.4, 100730.4, 100877.1, 
    101006.3,
  98600.49, 98787.94, 99006.16, 99201.2, 99390.39, 99546.84, 99697.51, 
    99873.03, 100061.8, 100239.5, 100408.8, 100566.7, 100712, 100863.1, 
    100995.3,
  98602.49, 98804.69, 99003.57, 99198.33, 99382.91, 99529.38, 99674.26, 
    99846.55, 100038.5, 100217.2, 100391.6, 100551.6, 100703.6, 100858.1, 
    100991.7,
  99504.46, 99686.88, 99895.42, 100092.4, 100274.6, 100456, 100622, 100774.4, 
    100916, 101038.7, 101156.9, 101256.4, 101346.3, 101414.2, 101463.2,
  99396.12, 99618.77, 99833.45, 100026.5, 100216.7, 100395.4, 100562, 
    100718.2, 100867.5, 101005.1, 101130.7, 101230.4, 101322.1, 101395.1, 
    101450.2,
  99371.22, 99560.91, 99752.99, 99941.59, 100133.1, 100315.5, 100494.5, 
    100663.4, 100810.8, 100954, 101076.7, 101187.7, 101283.9, 101366.1, 
    101429.8,
  99325.53, 99509.35, 99696.16, 99886.33, 100074.7, 100257.3, 100439.8, 
    100612.7, 100778.5, 100928.3, 101062.5, 101174.9, 101273.6, 101356.8, 
    101422.9,
  99286.47, 99468.77, 99647.79, 99834.27, 100014, 100202.6, 100383.2, 
    100563.1, 100730.9, 100888.5, 101027, 101145.8, 101247.3, 101331.8, 
    101402.1,
  99248.13, 99424.27, 99599.42, 99787, 99968.46, 100156.3, 100332.9, 
    100517.4, 100690.3, 100855.2, 100999.1, 101123, 101227.4, 101312.9, 
    101388.7,
  99207.88, 99381.16, 99558.65, 99745.02, 99924.94, 100110.9, 100288.5, 
    100471.4, 100649.9, 100817.2, 100965.9, 101094.8, 101204.5, 101293.4, 
    101371.5,
  99156.5, 99331.64, 99511.44, 99700.46, 99887.53, 100068, 100246.1, 
    100433.1, 100612, 100782.3, 100935.5, 101067.3, 101183.2, 101273.6, 
    101356.2,
  99090.98, 99273.6, 99464.58, 99655.84, 99843.91, 100024.7, 100207.9, 
    100395.1, 100576.4, 100746.4, 100903.6, 101039.3, 101158.2, 101254.2, 
    101338.4,
  99011.07, 99211.27, 99413.15, 99607.11, 99796.43, 99982.77, 100170, 
    100357.9, 100541.5, 100713.2, 100873, 101011.7, 101132.2, 101233.8, 
    101321.2,
  99044.85, 99232.66, 99473.56, 99679.65, 99879.65, 100063.4, 100216.8, 
    100367.2, 100506.4, 100636.8, 100764, 100890.6, 101006.1, 101114.7, 
    101213.8,
  98854.25, 99096.27, 99348.71, 99574.07, 99781.55, 99968.76, 100129.5, 
    100286, 100429.5, 100568.1, 100694.2, 100828.3, 100954.7, 101071.5, 
    101175.1,
  98736.77, 98981.76, 99228.26, 99465.85, 99677.44, 99881.41, 100055.6, 
    100210.6, 100360.8, 100506.8, 100634.2, 100774, 100907.2, 101029.2, 
    101138.8,
  98596.54, 98853.67, 99110.43, 99354.03, 99584.82, 99791.88, 99977.14, 
    100138.1, 100298, 100452.7, 100590.8, 100733.2, 100868.7, 100996.1, 
    101112.6,
  98475.23, 98744.35, 99000.2, 99258.77, 99490.95, 99708.84, 99903.83, 
    100076, 100235.3, 100400.4, 100543.6, 100690.4, 100830.8, 100962, 101080.9,
  98372.62, 98638.98, 98899.41, 99160.14, 99397.98, 99627.63, 99834.09, 
    100014.1, 100178.6, 100347.8, 100503, 100651.9, 100794.9, 100931.2, 
    101055.4,
  98284.68, 98550.59, 98814.66, 99073.6, 99320.93, 99559.13, 99770.27, 
    99961.95, 100131.2, 100302.7, 100467.9, 100617.8, 100766.1, 100904.5, 
    101033.8,
  98201.29, 98472.71, 98741.74, 99001.99, 99253.07, 99499.46, 99715.49, 
    99910.8, 100090.6, 100268, 100436.5, 100591.3, 100742.5, 100883.9, 
    101016.7,
  98134.1, 98405.7, 98681.34, 98941.22, 99201.66, 99447.23, 99668.5, 
    99871.47, 100059.2, 100238.5, 100415.6, 100570.2, 100724.7, 100868, 
    101000.9,
  98084.22, 98351.98, 98631.82, 98895.62, 99161.78, 99406.73, 99625.38, 
    99839.8, 100032.5, 100217, 100398.4, 100556.9, 100711.7, 100856.8, 
    100993.1,
  100423.6, 100446.2, 100550.4, 100653.2, 100769, 100901.8, 101035.7, 
    101164.9, 101276.7, 101377.6, 101457.4, 101524.9, 101576.2, 101618.1, 
    101648.7,
  100311.7, 100376.7, 100466.4, 100556, 100667.1, 100796.6, 100914.4, 
    101050.4, 101166.7, 101281.1, 101375.9, 101457.4, 101517.6, 101568.9, 
    101608.5,
  100233.6, 100275, 100349.9, 100443, 100543.2, 100657.8, 100791.9, 100922.7, 
    101049.9, 101170.4, 101276.2, 101372, 101447.3, 101511.5, 101558.2,
  100148.6, 100195.9, 100256.6, 100347.3, 100441.9, 100553.3, 100678.5, 
    100808.8, 100945.8, 101070.5, 101190.2, 101294.6, 101382.1, 101453.4, 
    101512.5,
  100050.2, 100105.7, 100155.9, 100242.8, 100331.4, 100442.6, 100560.4, 
    100694.4, 100826.7, 100961.3, 101084.4, 101200.4, 101301, 101381.7, 101452,
  99950.01, 100005.2, 100048.8, 100139.6, 100223.2, 100333.5, 100449.1, 
    100578.2, 100712, 100849.2, 100981.1, 101106, 101216.9, 101309, 101390.6,
  99849.37, 99890.54, 99929.38, 100026.7, 100112.6, 100219.2, 100334.1, 
    100462, 100595, 100733.8, 100868, 101001, 101125.6, 101230.8, 101323,
  99737.8, 99773.45, 99807.43, 99903.38, 99996.66, 100108.3, 100225.1, 
    100354.2, 100480, 100619.5, 100762.7, 100901.1, 101034.1, 101150.3, 
    101254.1,
  99605.41, 99644.23, 99678.16, 99772.87, 99871.62, 99993.22, 100108.1, 
    100238.4, 100365.7, 100508.5, 100649.3, 100796.6, 100936.9, 101064.8, 
    101180.4,
  99456.15, 99508.41, 99540.05, 99633.3, 99743.78, 99872.84, 99992.37, 
    100124.5, 100252, 100394.3, 100547.5, 100695.9, 100845.2, 100982.3, 
    101106.3,
  101226.5, 101338.3, 101472.9, 101592.6, 101692.4, 101783.5, 101859.1, 
    101927.5, 101983.9, 102035.3, 102087.2, 102133.8, 102166.7, 102180.7, 
    102183.1,
  101118.4, 101268.2, 101408.6, 101529.9, 101636.5, 101730.4, 101811.6, 
    101879.1, 101946.7, 102003.2, 102057.1, 102109.3, 102151.4, 102174.9, 
    102185.5,
  101062.9, 101214.9, 101347.8, 101471.8, 101586.3, 101686.9, 101779.3, 
    101854.6, 101924.3, 101985.6, 102040.8, 102096.3, 102141.3, 102169.7, 
    102183.6,
  101007.6, 101151.4, 101288.1, 101418.7, 101536.2, 101639, 101737.6, 
    101820.9, 101892.9, 101958.9, 102015.7, 102075.2, 102127, 102161.9, 
    102179.6,
  100951.3, 101098.1, 101233.5, 101369.8, 101482.8, 101597.9, 101697.1, 
    101787.5, 101867.2, 101934.6, 101996.7, 102057.8, 102111.5, 102151.3, 
    102173.4,
  100894.2, 101041.1, 101185.9, 101317.4, 101436.8, 101554.1, 101657.6, 
    101752.6, 101834.6, 101908.5, 101973.8, 102033.7, 102093.6, 102140, 
    102165.8,
  100840.6, 100990.5, 101133.4, 101269.9, 101389.7, 101507.9, 101618.9, 
    101718.2, 101803.7, 101883.2, 101950.4, 102013.8, 102074.4, 102124.8, 
    102155.1,
  100796.5, 100938.9, 101084.2, 101221.1, 101341.6, 101464.9, 101577.3, 
    101678.5, 101771.6, 101853.8, 101923, 101991.2, 102051.6, 102105.7, 
    102141.2,
  100753.9, 100890.9, 101035.8, 101170.6, 101298.7, 101420.4, 101532.7, 
    101638.9, 101735, 101822.1, 101896.1, 101964.3, 102028.8, 102082.7, 
    102123.3,
  100718.4, 100849.8, 100986.8, 101121.6, 101253.3, 101373.3, 101488.1, 
    101596.2, 101694.4, 101788, 101865.4, 101936.1, 102003, 102058.3, 102101.9,
  101732.6, 101863.7, 101994.5, 102106.5, 102207.4, 102292.4, 102360.8, 
    102407.8, 102438.2, 102449.8, 102452.9, 102468.1, 102485.7, 102503.6, 
    102492.9,
  101656.4, 101798.8, 101935.8, 102052.4, 102156.5, 102243.3, 102319.1, 
    102376.9, 102415.2, 102437.7, 102444, 102455.8, 102477.9, 102504.1, 
    102500.6,
  101583.4, 101731.6, 101868.8, 101993.8, 102106, 102203.8, 102285.3, 
    102349.3, 102396.5, 102425.5, 102437.7, 102451, 102471.1, 102502.4, 
    102506.1,
  101515.7, 101664.9, 101809.2, 101940.8, 102057.3, 102157.3, 102245.7, 
    102318.8, 102373.8, 102410.9, 102430, 102439.5, 102458.7, 102494, 102507.8,
  101442.4, 101596.9, 101745, 101881.9, 102003.2, 102109.6, 102202.8, 
    102282.6, 102343.9, 102390.5, 102416.3, 102431.2, 102450.6, 102482.4, 
    102505.6,
  101367.2, 101525.4, 101679.4, 101821.5, 101948.5, 102059.7, 102158.2, 
    102244.2, 102311.9, 102364.9, 102399.7, 102418.4, 102436.7, 102468.3, 
    102496.7,
  101296.4, 101452.2, 101611.1, 101758.7, 101891.2, 102009.3, 102112, 
    102202.4, 102278.2, 102337, 102379.2, 102405.9, 102423.3, 102456.1, 
    102488.4,
  101224.1, 101377.1, 101542.8, 101693.2, 101831.9, 101954.9, 102065.4, 
    102160.1, 102241.6, 102305.6, 102355.4, 102386, 102407.2, 102437.1, 
    102475.8,
  101148.1, 101308.2, 101469.9, 101623.6, 101769.1, 101899, 102015.5, 
    102115.6, 102202.5, 102273.1, 102327.6, 102365.9, 102390.7, 102418.7, 
    102456.7,
  101073.6, 101233.9, 101398.2, 101553.7, 101703.8, 101838.2, 101962.1, 
    102069.3, 102161.4, 102237.2, 102298, 102342.2, 102368.6, 102400, 102434.2,
  101966.8, 102052.4, 102130.6, 102196.7, 102247, 102294.3, 102326.6, 
    102345.4, 102361.4, 102365.3, 102359.3, 102364.2, 102362.8, 102356.5, 
    102325,
  101998.7, 102082.3, 102155.4, 102220.2, 102276.9, 102324.2, 102352.7, 
    102376.7, 102391.5, 102400.8, 102397.9, 102391.2, 102384, 102384.1, 
    102360.5,
  102038.9, 102113.2, 102184.4, 102246.6, 102305.3, 102350.9, 102382.7, 
    102405.2, 102425.3, 102432.1, 102429.8, 102418.6, 102409.1, 102401.8, 
    102394.3,
  102071.7, 102139.6, 102211.3, 102272.3, 102327.9, 102372.3, 102410.6, 
    102430.7, 102451.4, 102464.3, 102463, 102454.1, 102432.5, 102418.6, 
    102414.3,
  102103.5, 102167.3, 102235.9, 102290.3, 102343.9, 102385.1, 102426.8, 
    102454.8, 102470.3, 102486.1, 102485.8, 102484.9, 102462.8, 102438.5, 
    102426.5,
  102125.1, 102185, 102252, 102306.9, 102352.9, 102397.2, 102433.8, 102466.5, 
    102489.9, 102506.8, 102502.4, 102505.4, 102493.4, 102467.7, 102442.6,
  102139, 102196.2, 102260.7, 102313.6, 102355.7, 102403.1, 102437.5, 
    102464.6, 102488.4, 102511.9, 102524.4, 102521.6, 102507.2, 102493.2, 
    102460.8,
  102141.5, 102198.6, 102257.1, 102307, 102349.4, 102398.6, 102434.7, 
    102458.3, 102473.7, 102492.8, 102516.4, 102523.8, 102522, 102508.5, 
    102481.4,
  102142, 102187.1, 102241.2, 102294.7, 102338.2, 102382.4, 102418.4, 
    102446.3, 102467.6, 102485.9, 102492.1, 102511.9, 102516.5, 102506.9, 
    102494.5,
  102128, 102172.4, 102221.8, 102272.8, 102318.8, 102356.2, 102392.4, 
    102422.9, 102443.6, 102469.4, 102476, 102492.9, 102500.7, 102506.7, 
    102493.6,
  100965.3, 101059.2, 101163.3, 101269.4, 101366.6, 101459, 101553.4, 
    101647.7, 101719.7, 101779.5, 101827.4, 101873.8, 101913.4, 101940.5, 
    101962.5,
  101021.8, 101124.2, 101227.1, 101328.8, 101412, 101500, 101587.5, 101678.4, 
    101756.6, 101814.6, 101862.9, 101903, 101940.5, 101970.6, 101994.1,
  101084.9, 101188.8, 101280.4, 101380.1, 101463.6, 101549.2, 101636.1, 
    101720.1, 101794.3, 101853.8, 101907, 101948.7, 101986.8, 102013.5, 
    102034.9,
  101183.5, 101276.8, 101366.1, 101455.5, 101534, 101611.7, 101688.6, 
    101767.6, 101844.3, 101903.4, 101948.9, 101985.1, 102020.9, 102049.4, 
    102070.9,
  101295.9, 101384.2, 101468.8, 101550.8, 101618.9, 101690.3, 101765.3, 
    101837.8, 101907.9, 101964.3, 102010.9, 102044.4, 102072.7, 102096.3, 
    102109.5,
  101455.7, 101529.5, 101600.2, 101663.9, 101726, 101793.4, 101860.4, 
    101926.4, 101993.3, 102044.6, 102083.2, 102114, 102133.5, 102141.9, 
    102150.1,
  101621.9, 101672.7, 101729.2, 101777.6, 101832.8, 101887.8, 101947.2, 
    102006.4, 102068.8, 102118.2, 102160.1, 102185.1, 102205.7, 102208, 102201,
  101775.6, 101811.6, 101856.5, 101894.6, 101942.4, 101988.7, 102034.3, 
    102085.4, 102135.1, 102182.6, 102218, 102244.4, 102259.7, 102266.8, 102261,
  101907.9, 101938.3, 101977, 102014.2, 102051.2, 102088.6, 102125.1, 
    102165.3, 102204.2, 102242.8, 102265.3, 102290.9, 102302.3, 102307.7, 
    102299.5,
  102027.1, 102054.4, 102083.2, 102114.3, 102142.3, 102172.9, 102199.9, 
    102227.6, 102256.7, 102288.4, 102311.9, 102325.7, 102335.2, 102342.9, 
    102329.3,
  101541, 101608.2, 101687, 101749.9, 101810, 101859, 101901.7, 101934.2, 
    101957.1, 101970.2, 101974.6, 101974, 101952, 101928.1, 101910.9,
  101508.1, 101583.9, 101664.5, 101729.5, 101791, 101841.1, 101885.5, 
    101921.5, 101947, 101963.3, 101972, 101975, 101962.5, 101944.6, 101933,
  101481, 101552.1, 101633.4, 101699.4, 101763.6, 101815.7, 101864.8, 
    101903.4, 101935.8, 101957, 101969.1, 101977.4, 101968.4, 101945, 101940.5,
  101451.1, 101522, 101602.6, 101671.6, 101739.6, 101793.5, 101847.7, 101892, 
    101926.5, 101951, 101965, 101975.5, 101966.4, 101948.2, 101946.4,
  101410.1, 101481.4, 101564.9, 101637.2, 101707, 101767.8, 101822.6, 
    101868.7, 101905.9, 101934.5, 101952, 101961, 101958, 101945.4, 101942.2,
  101356.2, 101432.6, 101521.1, 101599.5, 101671.8, 101733.5, 101790.9, 
    101843.6, 101883.8, 101916.2, 101936, 101946.9, 101951.1, 101944.3, 
    101953.9,
  101303.2, 101396.8, 101479.9, 101560.3, 101635.9, 101702.4, 101764.8, 
    101816.6, 101860.8, 101893.4, 101919.1, 101933.4, 101944.1, 101944, 
    101960.8,
  101271, 101369.1, 101449, 101536.6, 101610.8, 101678.6, 101744.1, 101796.1, 
    101840.2, 101874.4, 101904.9, 101923.4, 101940.9, 101954.6, 101974.4,
  101263.5, 101354.1, 101430, 101518.8, 101592.1, 101665.4, 101732.8, 
    101785.7, 101830.4, 101868.1, 101898.4, 101919.7, 101944.3, 101969.5, 
    101983.4,
  101280.4, 101361.3, 101437.1, 101519.7, 101592.2, 101669.1, 101732.1, 
    101788.6, 101831.6, 101866, 101901.3, 101927.9, 101955.6, 101985, 101998,
  100935, 101016.3, 101114.5, 101204.6, 101293.2, 101382.2, 101459.5, 
    101532.4, 101598.1, 101654.7, 101701.1, 101741.4, 101767.4, 101792.4, 
    101811.8,
  101040.4, 101120.4, 101212.5, 101295.9, 101379.8, 101455.1, 101527.2, 
    101598, 101654.8, 101709.9, 101750.5, 101787.8, 101813.3, 101836, 101850.9,
  101167.1, 101237, 101316.8, 101394.4, 101472.2, 101545.2, 101612.3, 
    101672.6, 101724.9, 101767.7, 101803.4, 101832.2, 101853, 101871.1, 
    101883.9,
  101299.2, 101365.2, 101436.3, 101502.5, 101571.9, 101636, 101698.7, 101752, 
    101794.8, 101831.2, 101859.4, 101883.2, 101899.1, 101912.5, 101922.7,
  101441.3, 101494.8, 101554.2, 101610.8, 101672.6, 101729.7, 101785.6, 
    101831.2, 101867, 101893.8, 101915.8, 101934, 101945.2, 101953.7, 101962.5,
  101569.9, 101612.2, 101668.1, 101717.2, 101772.9, 101823.1, 101874.9, 
    101909, 101938.7, 101959.6, 101975.3, 101986, 101994.9, 102001.4, 102010.8,
  101686.5, 101723.8, 101774.2, 101817.9, 101866.7, 101911.9, 101955.8, 
    101984.3, 102010.8, 102023.8, 102035.9, 102039.6, 102043.6, 102045.2, 
    102049.8,
  101791.2, 101825.6, 101870.1, 101909.8, 101953.7, 101993.7, 102031.4, 
    102055.9, 102076.8, 102084.3, 102089.8, 102088.7, 102090.9, 102088.2, 
    102093.5,
  101882.5, 101916.6, 101958.2, 101994.8, 102035, 102069.6, 102099.5, 
    102122.1, 102135.7, 102139.5, 102141.2, 102132.6, 102131.1, 102123.9, 
    102132.3,
  101958.9, 101993.6, 102032.9, 102069.7, 102106.2, 102136.8, 102162.8, 
    102180, 102190.9, 102188.9, 102187.4, 102178.2, 102169.3, 102166.6, 
    102167.8,
  101256.9, 101319.5, 101418.7, 101488.5, 101559, 101611.7, 101650, 101687.2, 
    101711.2, 101738.4, 101775.1, 101810, 101851.1, 101897.4, 101927.5,
  101212.3, 101282.4, 101379.7, 101446.4, 101515.7, 101581, 101627.8, 
    101665.6, 101698.3, 101732.7, 101774.6, 101818.1, 101856.5, 101909.6, 
    101945,
  101184, 101242.7, 101335.2, 101408.5, 101484.8, 101546.4, 101599.5, 101649, 
    101694.1, 101736, 101781.4, 101837.7, 101870.5, 101936.6, 101971.1,
  101143.9, 101214.5, 101301.7, 101379, 101460.9, 101530.5, 101586.2, 
    101641.2, 101693.3, 101741.5, 101789.6, 101853.1, 101891.6, 101958.5, 
    101996.4,
  101098.3, 101179.6, 101269, 101360, 101440.3, 101509.2, 101570.2, 101628.4, 
    101689.5, 101746.1, 101797.5, 101864.1, 101911.4, 101978.6, 102021.2,
  101079.5, 101166.3, 101254.5, 101342.9, 101424, 101499, 101562.3, 101625, 
    101690.1, 101753.8, 101811.3, 101879.2, 101933.2, 102004, 102050.6,
  101072.3, 101160.3, 101249, 101335.9, 101418.9, 101494.2, 101559.9, 
    101623.5, 101693.5, 101765.1, 101833.4, 101903.3, 101958.2, 102030.4, 
    102081.2,
  101098.6, 101179.5, 101263.5, 101346.9, 101427.2, 101501.2, 101568.8, 
    101636, 101705.8, 101779.8, 101858.7, 101930.5, 101985.9, 102058.6, 
    102108.5,
  101168.9, 101228.9, 101303.9, 101373.2, 101448.9, 101522, 101588.2, 
    101660.1, 101728.4, 101804.5, 101885.7, 101960.8, 102018.5, 102090.7, 
    102143.4,
  101251.8, 101298.3, 101366.1, 101427.2, 101494.1, 101561.7, 101625.1, 
    101695.9, 101762.9, 101837.9, 101913.8, 101991.2, 102054, 102126, 102179.9,
  101614.2, 101682.6, 101765.2, 101831.3, 101895.2, 101951.2, 101997.3, 
    102038.5, 102066.2, 102091.9, 102119.4, 102140.1, 102166.2, 102189.8, 
    102202.2,
  101630.3, 101717.1, 101799.8, 101867.5, 101929.4, 101979.8, 102021.9, 
    102064.1, 102090.4, 102114.7, 102135.6, 102158.9, 102178.6, 102205.5, 
    102219.6,
  101689.8, 101768.3, 101841.9, 101906.1, 101965.2, 102015.4, 102057.5, 
    102096.2, 102117.6, 102137.4, 102156.6, 102179.8, 102191.9, 102221.9, 
    102241.3,
  101730.4, 101809.1, 101886.5, 101944.8, 102002, 102048.7, 102089.3, 
    102123.9, 102146.6, 102161.7, 102177.8, 102196.5, 102205.8, 102242.5, 
    102258.9,
  101777.4, 101851.7, 101923.4, 101978.1, 102031.9, 102077.1, 102118.4, 
    102151.2, 102176.2, 102186.5, 102196.9, 102215.1, 102223, 102252.6, 
    102276.2,
  101812, 101884.3, 101956, 102009.6, 102064.6, 102109.4, 102149.6, 102180, 
    102205, 102214.3, 102221.2, 102234.1, 102235.7, 102266, 102289.8,
  101845.5, 101910.6, 101981.7, 102039, 102091.6, 102135.1, 102173.1, 
    102204.7, 102228.3, 102240.6, 102240.2, 102251.4, 102246.7, 102277.1, 
    102307.2,
  101862.1, 101925.4, 102000.4, 102057.3, 102108.9, 102155.7, 102192.5, 
    102224.4, 102249.7, 102264, 102259.3, 102268.9, 102262.5, 102283.7, 
    102318.9,
  101870.7, 101937.4, 102007.3, 102066.2, 102119.9, 102164.9, 102203.9, 
    102237.4, 102264.4, 102285, 102273.7, 102280.1, 102282.3, 102284, 102326.5,
  101866.8, 101936.3, 102008, 102069.3, 102118.4, 102166, 102206.9, 102244.7, 
    102270, 102296.4, 102287.3, 102290.1, 102299.5, 102286.3, 102333.1,
  101839.2, 101857.7, 101902.8, 101944.4, 101991.4, 101997.2, 102012.1, 
    102036, 102082.7, 102141.4, 102197.5, 102246, 102279.3, 102300, 102306.8,
  101775.5, 101817.1, 101880.6, 101922.6, 101978.3, 101996.5, 102020.5, 
    102034.9, 102066.6, 102133.1, 102198.5, 102253.3, 102290.4, 102312.9, 
    102322.6,
  101743.5, 101785.9, 101845.5, 101899.7, 101961.4, 101988.4, 102025, 
    102045.7, 102069.3, 102137.2, 102209.3, 102259.7, 102297.8, 102325.7, 
    102339.1,
  101690.3, 101741.6, 101816.5, 101878.6, 101944.5, 101980.1, 102018.7, 
    102048.2, 102071.2, 102138.8, 102212.9, 102264.4, 102304.8, 102338.4, 
    102356.1,
  101640.6, 101704.8, 101785, 101848.7, 101917.4, 101965.3, 102003.7, 102047, 
    102077.2, 102140.1, 102212.6, 102266, 102312.8, 102349, 102368.4,
  101592.7, 101668.3, 101752.4, 101825.4, 101894.9, 101955.5, 102001.8, 
    102048.6, 102080.2, 102136.9, 102210.1, 102266.8, 102323.2, 102359.9, 
    102386.8,
  101553.7, 101637, 101725, 101802.8, 101874, 101940, 101996.9, 102051.2, 
    102086.3, 102134, 102205.4, 102264.8, 102327.5, 102366.9, 102400.2,
  101520.6, 101610.6, 101702.9, 101784.7, 101858.2, 101930.6, 101992.4, 
    102054.1, 102093.9, 102135.6, 102201.4, 102262.7, 102328, 102373, 102413.8,
  101499.5, 101589.9, 101685.6, 101771.8, 101849.5, 101922.5, 101986.8, 
    102055.3, 102101.1, 102139.8, 102200.2, 102262.1, 102327.2, 102374.3, 
    102412.4,
  101487.4, 101578.5, 101679.7, 101763.8, 101844.5, 101918.7, 101984, 
    102053.9, 102105.3, 102146.5, 102202.8, 102264.4, 102327, 102372.9, 
    102410.5,
  102159.9, 102191.8, 102228.6, 102259.5, 102284.9, 102283.6, 102260.3, 
    102229.3, 102231.7, 102233, 102265.8, 102292.8, 102310.5, 102317, 102320.7,
  102142.8, 102184.5, 102220.1, 102257.3, 102287.9, 102306.6, 102309.2, 
    102265.7, 102252.3, 102242.9, 102269, 102304.1, 102322.4, 102331.9, 
    102337.9,
  102136, 102182.2, 102217.6, 102254.1, 102295.8, 102309.2, 102325.3, 
    102302.5, 102272.5, 102264.8, 102276.4, 102306.3, 102328.5, 102347.7, 
    102354.9,
  102118.7, 102173.6, 102217.2, 102255.4, 102292.3, 102320.6, 102334.1, 
    102336.5, 102300, 102277.7, 102281.2, 102308.4, 102342.3, 102363.8, 
    102371.1,
  102086.1, 102156.8, 102204.9, 102249.4, 102282.6, 102318.8, 102335.2, 
    102333.7, 102314.4, 102287, 102283.7, 102312.3, 102350.6, 102373.3, 
    102388.6,
  102043.6, 102124.3, 102189.6, 102236.3, 102275.7, 102313, 102334.9, 
    102351.5, 102336.8, 102292.5, 102284.6, 102314.1, 102356.8, 102397.5, 
    102420.2,
  101991.6, 102081.3, 102161.8, 102218.8, 102263, 102300.8, 102329.1, 102348, 
    102342.1, 102296.8, 102295.1, 102308.3, 102360.9, 102397, 102425.8,
  101928.3, 102032.8, 102124.7, 102191.4, 102242.9, 102287.6, 102317.1, 
    102345.2, 102348, 102303.1, 102302.9, 102298.4, 102356, 102399.8, 102438.7,
  101856.5, 101977.8, 102078, 102156.7, 102213.8, 102267.3, 102301.3, 
    102329.8, 102351.5, 102317.1, 102300.4, 102291.5, 102346.5, 102392.5, 
    102430.2,
  101777.9, 101914.9, 102024.2, 102112.2, 102181.9, 102239.6, 102282.7, 
    102315.7, 102334.8, 102321.4, 102296.2, 102286.6, 102334.6, 102390, 
    102425.2,
  101886.8, 101939.4, 102004.1, 102049.4, 102083.7, 102087.2, 102099.7, 
    102134, 102176.5, 102223, 102263.6, 102296.3, 102301.1, 102300.9, 102295.3,
  101856.3, 101919.8, 101987.8, 102040.7, 102088.6, 102092.5, 102083.1, 
    102126.9, 102172.8, 102216.8, 102256.1, 102297.1, 102312.3, 102321, 
    102314.8,
  101859, 101926.1, 101986.8, 102035.1, 102082.9, 102106.4, 102090.3, 
    102117.6, 102169, 102216.2, 102263.3, 102306.3, 102328.9, 102338.4, 102328,
  101863.1, 101933.5, 101995, 102039, 102083, 102112.2, 102098.8, 102120, 
    102170.2, 102215.6, 102269.3, 102315.2, 102341.9, 102357.7, 102347.5,
  101875.2, 101948.5, 102005.6, 102047.9, 102084.1, 102109.1, 102104.7, 
    102131.2, 102175.4, 102220.2, 102272.6, 102320.2, 102353.6, 102373.8, 
    102374.4,
  101892, 101967.2, 102023.2, 102065.6, 102097.4, 102121.1, 102114.8, 
    102138.7, 102176.5, 102222, 102279.2, 102329.7, 102378.6, 102394.1, 
    102394.1,
  101914.9, 101987.8, 102046.2, 102087.7, 102117.5, 102130.4, 102120.6, 
    102146.1, 102184.5, 102231.9, 102284.6, 102337.9, 102389.7, 102409.2, 
    102412.5,
  101938.6, 102009.9, 102070.3, 102113.8, 102145, 102151.1, 102136.1, 
    102156.8, 102205.1, 102248.9, 102301, 102345.4, 102393.7, 102412.2, 
    102417.4,
  101963.5, 102031.9, 102094.6, 102138.7, 102173.8, 102179.5, 102160.5, 
    102172.1, 102223.1, 102264.3, 102314.6, 102341.5, 102396.3, 102413.2, 
    102426.3,
  101983.7, 102054.9, 102117.9, 102166.2, 102204, 102209.1, 102198.4, 
    102194.5, 102243.5, 102285.9, 102323.3, 102353.7, 102395.6, 102424.7, 
    102437.9,
  102077.4, 102112.6, 102143.8, 102150.8, 102159.1, 102159.2, 102204.9, 
    102252.7, 102295.6, 102331.8, 102360.3, 102379.8, 102378.2, 102363.5, 
    102347.7,
  102048, 102094.1, 102131.1, 102148.8, 102160, 102157.3, 102199.5, 102251.4, 
    102297.6, 102340.8, 102375.8, 102400.2, 102400.2, 102389.3, 102375.8,
  102024.5, 102075.7, 102116.7, 102141.2, 102160.7, 102166.3, 102206.9, 
    102266.3, 102309.1, 102354.1, 102389.7, 102416.6, 102430, 102412.8, 
    102398.7,
  102006.2, 102064.1, 102111, 102136.6, 102157.2, 102171.8, 102209.4, 
    102270.1, 102320.6, 102362.1, 102399.7, 102427.9, 102435.4, 102435.8, 
    102422.4,
  101982.3, 102042.4, 102099.2, 102128.7, 102147.4, 102177.4, 102221.6, 
    102280, 102333.5, 102370.6, 102411.2, 102438.6, 102453.7, 102462, 102449.7,
  101957.7, 102022.7, 102089.5, 102130.1, 102150.6, 102185, 102234, 102287.1, 
    102341.9, 102378, 102419.5, 102455.8, 102474.1, 102482.1, 102469.9,
  101933.3, 102001.5, 102075.1, 102124.2, 102151.9, 102196, 102246.7, 
    102298.5, 102351.2, 102386.5, 102430.8, 102470.8, 102499.7, 102498, 
    102486.8,
  101907.5, 101978.2, 102059.7, 102114.8, 102154.4, 102204.5, 102253.7, 
    102305.5, 102353.7, 102394.8, 102437, 102489.2, 102529.1, 102514.8, 
    102506.9,
  101880.4, 101955.9, 102042.4, 102103.3, 102151.1, 102208.2, 102257.3, 
    102308.7, 102358.8, 102397.7, 102448.6, 102505.8, 102541.5, 102530.3, 
    102527.5,
  101850.8, 101932.6, 102022.6, 102089.4, 102147, 102204.2, 102250.7, 
    102304.6, 102357.8, 102402.6, 102459.3, 102516.4, 102545.3, 102544.5, 
    102541.2,
  101951.3, 102065.9, 102156.7, 102226.2, 102281.9, 102345.1, 102390.9, 
    102434.9, 102463.9, 102478.4, 102467.6, 102455, 102431.5, 102408.3, 
    102377.9,
  101928.8, 102042.6, 102137.6, 102214.3, 102275.2, 102342.8, 102398.8, 
    102449.1, 102484, 102499.1, 102501.3, 102484.9, 102460, 102438.6, 102408.4,
  101907.9, 102028.8, 102127.8, 102212.1, 102279.7, 102348.2, 102410.2, 
    102461.6, 102500.4, 102519.2, 102527.2, 102510.4, 102493.4, 102470.6, 
    102440.7,
  101883.7, 102010.3, 102111.2, 102200.2, 102273.5, 102347, 102415.8, 
    102472.1, 102519.1, 102551, 102544.4, 102539.9, 102521.5, 102500.7, 
    102472.3,
  101862.3, 101992.7, 102097, 102188.9, 102266.8, 102347.2, 102420.9, 
    102483.2, 102536, 102564, 102567.7, 102567.5, 102553.4, 102532.6, 102506.7,
  101840.5, 101974.7, 102082, 102175.3, 102253.9, 102342.2, 102419.5, 
    102493.3, 102551.9, 102579.5, 102593.2, 102593.4, 102581.2, 102561.6, 
    102537.3,
  101820.9, 101957.7, 102068.7, 102164, 102242.9, 102336.3, 102420.4, 
    102499.7, 102562.6, 102595.1, 102613.5, 102616.1, 102606.9, 102590.5, 
    102567.6,
  101803.2, 101943, 102057.2, 102153.8, 102234.4, 102330.8, 102420.8, 
    102505.8, 102573.1, 102615.4, 102644.8, 102649.3, 102643.3, 102616.2, 
    102594.2,
  101788.3, 101931.1, 102049, 102147.8, 102231.1, 102328.4, 102421.5, 
    102510.7, 102586.2, 102636.7, 102671.4, 102682, 102667.2, 102647.3, 
    102624.1,
  101778.2, 101922.2, 102042.2, 102142.4, 102234, 102332.4, 102426.5, 
    102518.1, 102597, 102653.5, 102688.9, 102708.4, 102693.9, 102679.1, 
    102653.9,
  102281.2, 102380.1, 102447.2, 102483.3, 102521.7, 102552.2, 102575.3, 
    102581, 102572.9, 102555.9, 102540.9, 102509.4, 102471.8, 102431.7, 
    102385.6,
  102271.4, 102368.2, 102438.5, 102484.7, 102530.3, 102566.3, 102596.5, 
    102600.2, 102602.8, 102586, 102569.1, 102543.6, 102506.7, 102465.6, 
    102417.6,
  102255.5, 102362.1, 102441.4, 102490.9, 102539, 102583.8, 102616.5, 
    102633.6, 102626.4, 102623, 102602.1, 102577.9, 102541.4, 102499.2, 
    102451.2,
  102240.3, 102354.1, 102439.7, 102494.5, 102544.8, 102600.2, 102633.9, 
    102656.6, 102657.6, 102658, 102635.4, 102612.9, 102575.6, 102534.5, 
    102485.2,
  102223.5, 102341.7, 102434.7, 102499.1, 102551.1, 102613.2, 102652.8, 
    102678.1, 102694, 102682.7, 102669.9, 102650.1, 102612.8, 102569.7, 
    102519.8,
  102205.1, 102328.7, 102427.8, 102497.6, 102553.6, 102622, 102670.4, 
    102701.3, 102729.2, 102721.2, 102703.3, 102688.5, 102653.1, 102608.9, 
    102554.7,
  102188, 102313.2, 102418.4, 102495.8, 102555.5, 102626.7, 102681.7, 
    102726.7, 102744, 102737.1, 102735.2, 102722.2, 102691.7, 102647.4, 
    102589.8,
  102169.9, 102300, 102406.8, 102491.5, 102555.7, 102629.6, 102692.7, 
    102745.9, 102765.6, 102776.5, 102773.7, 102754.3, 102728.8, 102687.5, 
    102628,
  102153.6, 102288.8, 102395.3, 102485.7, 102553.4, 102631.1, 102699.7, 
    102762.1, 102786.8, 102804.3, 102803.4, 102791.3, 102764.3, 102721.9, 
    102664.1,
  102138.1, 102277.3, 102384.6, 102478.2, 102551, 102628.6, 102702.4, 
    102769.9, 102802.5, 102826.7, 102831.5, 102825.5, 102799, 102754.5, 
    102698.1,
  102569.4, 102655.5, 102700.1, 102724.3, 102751.1, 102771.3, 102764.5, 
    102740.7, 102720.6, 102691.6, 102652.4, 102605, 102555.2, 102498.8, 
    102442.3,
  102557.7, 102645.7, 102690.8, 102728.7, 102764.4, 102784.9, 102789.2, 
    102784.3, 102751.5, 102728, 102691.5, 102644.3, 102595.6, 102535.9, 
    102478.9,
  102536.7, 102635.7, 102688, 102734.7, 102775.7, 102799.7, 102811.4, 
    102808.3, 102791.8, 102761.5, 102730.3, 102683.3, 102634.2, 102577.9, 
    102516.2,
  102517.1, 102626.5, 102682.5, 102735.6, 102783.6, 102808.2, 102828, 
    102828.7, 102822.1, 102803.3, 102769.8, 102726.3, 102674.2, 102617.3, 
    102554.5,
  102496.6, 102614.3, 102675.9, 102735, 102788.9, 102824.6, 102850.4, 102856, 
    102859.6, 102839.7, 102809.8, 102764.7, 102715.6, 102655.6, 102592.8,
  102477.5, 102602.4, 102669.7, 102732.8, 102793.8, 102834.5, 102867.4, 
    102887.1, 102891.3, 102878.3, 102850.7, 102803.2, 102755.1, 102694.8, 
    102629.6,
  102458.4, 102588.4, 102662.4, 102728.4, 102796.4, 102843.1, 102886.7, 
    102910.8, 102915.1, 102913.8, 102890.3, 102839.9, 102789.3, 102731.7, 
    102663.6,
  102440.5, 102574.5, 102655.1, 102721.8, 102795.8, 102850.6, 102899.6, 
    102919.7, 102934.4, 102935, 102915.9, 102877, 102818.8, 102763.2, 102695.2,
  102422.9, 102557.9, 102647.1, 102714.8, 102791.9, 102852, 102905.5, 
    102931.5, 102951.2, 102952.2, 102936.2, 102903.8, 102849.8, 102794, 
    102722.3,
  102402.9, 102541.2, 102637.8, 102706.6, 102786.6, 102850.6, 102907.6, 
    102939.5, 102955.8, 102966.8, 102958.3, 102919.9, 102869.1, 102820.2, 
    102750.7,
  102706.8, 102767.9, 102801, 102821.6, 102838.9, 102838.5, 102831.5, 
    102804.3, 102780, 102740.5, 102693.7, 102643.1, 102583.8, 102521.6, 
    102460.3,
  102707.7, 102773.1, 102810, 102839.5, 102863.2, 102867.9, 102861.4, 
    102843.2, 102813.4, 102780.4, 102733.7, 102684, 102626.9, 102564, 102501.3,
  102704.8, 102775.2, 102817.9, 102851.4, 102881.7, 102885.4, 102893.6, 
    102882.9, 102853.8, 102819.5, 102773.5, 102723.2, 102664.8, 102602.6, 
    102538,
  102701.5, 102775.9, 102828.5, 102860.5, 102899.7, 102909.8, 102923.3, 
    102911, 102892.1, 102859.8, 102811, 102762.2, 102703.7, 102640.8, 102576.9,
  102693.6, 102773.4, 102831.1, 102867.4, 102908.8, 102929, 102945.4, 102945, 
    102924.2, 102895.9, 102846.2, 102796.3, 102739.9, 102676.5, 102611.8,
  102685, 102770, 102834, 102875, 102915.1, 102942.3, 102964.1, 102971, 
    102956.7, 102924.8, 102880.5, 102827.2, 102773, 102709.1, 102644,
  102673.3, 102761.8, 102830.6, 102877.6, 102915.4, 102954.1, 102973.5, 
    102990.8, 102979.4, 102948.1, 102911.3, 102856.4, 102800.7, 102739.3, 
    102671.6,
  102658, 102749.5, 102821.4, 102879.5, 102915.6, 102951, 102977.6, 102996.6, 
    102996.9, 102965.9, 102935.4, 102882.6, 102825.3, 102764.3, 102696,
  102639.6, 102733.1, 102809.3, 102870.6, 102917.3, 102948.1, 102975.6, 
    102994.6, 103001.1, 102984.1, 102952.1, 102904.7, 102847.7, 102786.9, 
    102719.6,
  102617.5, 102712.1, 102795, 102860.1, 102908.3, 102943.2, 102971.3, 
    102991.9, 102998.8, 102991.7, 102963.9, 102920.5, 102864.5, 102804.1, 
    102738.9,
  102256.4, 102350.2, 102429.5, 102487.4, 102529.5, 102558.5, 102563.7, 
    102562.9, 102551.5, 102533.5, 102507.1, 102472.6, 102430.7, 102384.2, 
    102336.7,
  102274.4, 102367.8, 102445, 102505.9, 102550.2, 102576.4, 102590.2, 
    102594.5, 102585.6, 102565.7, 102534.6, 102498.7, 102457.8, 102408.9, 
    102360.8,
  102297.5, 102394, 102475, 102541.7, 102589.8, 102614.4, 102622, 102625.2, 
    102616.1, 102594.3, 102563.7, 102525.3, 102484.5, 102434.8, 102384.4,
  102321.7, 102417.7, 102501.9, 102565.2, 102608.5, 102635.1, 102651.9, 
    102654, 102645.6, 102625.4, 102590.8, 102552.9, 102510, 102460.1, 102407,
  102350.5, 102443.1, 102525.4, 102591.1, 102637.7, 102671.9, 102682.8, 
    102681.6, 102670.9, 102650.4, 102618, 102579.4, 102534.6, 102484.6, 
    102428.8,
  102377.8, 102467, 102548.2, 102614.2, 102665, 102698.6, 102715.5, 102714.8, 
    102700.1, 102677.3, 102645.5, 102606.6, 102558.7, 102508.7, 102451,
  102405, 102492.8, 102572.4, 102636.8, 102688.2, 102719.1, 102735.1, 
    102737.7, 102723.5, 102699.7, 102666, 102627.7, 102579.3, 102529.1, 
    102471.2,
  102428.2, 102515.3, 102591.5, 102653, 102705.8, 102734.2, 102753.6, 
    102753.5, 102741.3, 102719, 102683.7, 102645.8, 102596.4, 102544, 102486.3,
  102450.9, 102537, 102612.1, 102669.1, 102721.9, 102752.9, 102756, 102764.1, 
    102750.4, 102728, 102694.4, 102657.3, 102608.8, 102558.5, 102499,
  102468.5, 102555.5, 102626.2, 102682.6, 102729.9, 102758, 102760.1, 
    102768.2, 102752.5, 102731.1, 102699.9, 102663.8, 102616.7, 102566.1, 
    102508,
  102140.9, 102124.8, 102153.3, 102162.6, 102170.7, 102180.4, 102184.8, 
    102190.6, 102203.6, 102219.7, 102231, 102225.6, 102215.3, 102187.9, 
    102162.9,
  102068, 102068.2, 102112.1, 102124.3, 102146.2, 102160.6, 102171.2, 
    102186.1, 102199.6, 102214.8, 102226, 102228.6, 102222.2, 102196.2, 
    102169.4,
  102007.7, 102024, 102073.6, 102092.5, 102128.6, 102150, 102169.5, 102184.9, 
    102197.5, 102216, 102227.5, 102230.5, 102224.1, 102200, 102174.6,
  101954.1, 101979.3, 102030.4, 102061, 102105.2, 102133.4, 102158.6, 
    102177.9, 102193.5, 102214.8, 102227.4, 102235.6, 102224.6, 102206.9, 
    102181.4,
  101898.6, 101933.9, 101988.9, 102032.4, 102080, 102117.6, 102147.5, 
    102170.4, 102194.4, 102216.5, 102232.9, 102238.1, 102227.6, 102210.7, 
    102185.8,
  101846.1, 101889.2, 101950.4, 102002.4, 102054.9, 102101.1, 102140.3, 
    102170.8, 102196, 102219.6, 102236.7, 102238.7, 102227.6, 102214.7, 
    102189.1,
  101800.6, 101847.6, 101919.5, 101977.9, 102037.8, 102093.7, 102133.6, 
    102170.5, 102197, 102223.3, 102233, 102240.3, 102232.1, 102214.7, 102190.6,
  101759.6, 101814.4, 101894.2, 101958.5, 102026.6, 102084.9, 102130, 
    102167.3, 102197.9, 102223.2, 102238.1, 102242.9, 102228.4, 102215.9, 
    102188.2,
  101724.4, 101789.7, 101877.4, 101946.7, 102020.4, 102081.5, 102130.8, 
    102173.8, 102202.3, 102223.1, 102235.1, 102239.1, 102223.1, 102212.1, 
    102176.9,
  101703, 101775.3, 101866.9, 101941.6, 102017.4, 102078.1, 102128, 102172.4, 
    102203.8, 102221.5, 102234.1, 102230.6, 102211.1, 102191.2, 102157.4,
  102148.3, 102165.9, 102178.5, 102190.1, 102185.6, 102178.3, 102165, 102140, 
    102109.9, 102067.2, 102031.4, 102011.9, 102020.2, 102028.3, 102027.4,
  102139.8, 102161.7, 102184.4, 102188.3, 102181.8, 102167.9, 102149.6, 
    102120.5, 102094, 102060.8, 102031.1, 102005.1, 102008.3, 102016.6, 
    102021.2,
  102134.2, 102148.4, 102169.5, 102173.1, 102166.3, 102152.2, 102141.2, 
    102108.2, 102083.1, 102043.7, 102016.2, 101991.2, 101993, 102002.8, 
    102012.5,
  102118.8, 102136.5, 102157.2, 102158.1, 102152.5, 102138.6, 102126.9, 
    102093.4, 102066.3, 102027.2, 102001, 101977.2, 101974.9, 101988.7, 102003,
  102101.7, 102114.1, 102133.7, 102136.3, 102133.8, 102124.8, 102109, 
    102083.8, 102044, 102015.3, 101983.3, 101962.5, 101956.7, 101975, 101992.7,
  102090.5, 102096, 102111.8, 102115.1, 102114.6, 102103.5, 102088.7, 
    102062.6, 102029.2, 101993.7, 101964.7, 101943.6, 101940.5, 101960.9, 
    101980.7,
  102081, 102076.1, 102087.1, 102086, 102087.7, 102079.8, 102065.3, 102036.3, 
    102009.9, 101968.3, 101943.4, 101926.6, 101924.5, 101948.4, 101971.6,
  102067.8, 102050.5, 102058.8, 102057.6, 102054.1, 102050.9, 102034.2, 
    102011.4, 101981.5, 101944.2, 101919.5, 101902.5, 101907.5, 101936.6, 
    101958.2,
  102027.2, 102017.2, 102022.9, 102023.9, 102020.6, 102016.7, 102002.9, 
    101983.8, 101954.4, 101925.3, 101899.1, 101889.7, 101891.8, 101922.8, 
    101951.8,
  101974.1, 101969.3, 101984.7, 101980.3, 101982.1, 101981, 101973.8, 
    101954.3, 101928.4, 101900.6, 101878.9, 101866.2, 101882.2, 101913.6, 
    101937.2,
  100941.6, 101067, 101207.7, 101321.5, 101429.8, 101524.6, 101605.8, 
    101670.8, 101718.9, 101759.2, 101790.6, 101812.3, 101835.2, 101860.7, 
    101880.5,
  100849.1, 100987.2, 101133.3, 101254.8, 101362.5, 101461.4, 101548, 
    101618.3, 101676.3, 101722.6, 101764.8, 101790.1, 101807.1, 101828, 
    101851.8,
  100786.3, 100927.3, 101064.5, 101182.6, 101300.8, 101404.9, 101499, 
    101578.3, 101641, 101688.8, 101731.9, 101767.1, 101789.8, 101805.6, 
    101828.9,
  100751.1, 100890.2, 101024.4, 101146.6, 101265.6, 101369.2, 101467.3, 
    101542.4, 101606.5, 101660.7, 101706.7, 101743.1, 101774.3, 101787.1, 
    101804.2,
  100722.7, 100858.1, 100988.9, 101111.4, 101225.2, 101329.5, 101427.8, 
    101504.8, 101571, 101631.6, 101679.6, 101721, 101748.9, 101767.2, 101785.7,
  100720.4, 100844, 100969.2, 101084.4, 101196.1, 101300.4, 101400.3, 101477, 
    101541.8, 101603.5, 101652, 101698.2, 101730.3, 101750.2, 101766.4,
  100733.1, 100847.5, 100962.1, 101070.3, 101179.3, 101278.7, 101376.7, 
    101448.9, 101519.7, 101579.8, 101629.6, 101675.8, 101708.2, 101731.6, 
    101752.1,
  100766.6, 100866.9, 100975.1, 101073.7, 101174.3, 101269.6, 101356, 
    101433.2, 101501.7, 101559.6, 101607.3, 101651.9, 101685, 101709.2, 
    101736.5,
  100816, 100902.9, 100997.1, 101086.7, 101175.6, 101266.3, 101343.8, 101426, 
    101486.5, 101545, 101590.8, 101634.4, 101666.5, 101689.9, 101723.6,
  100880.9, 100953.3, 101038.3, 101116.6, 101195.3, 101271.6, 101348.1, 
    101419.8, 101482.2, 101533.5, 101581.8, 101618.6, 101644, 101668.6, 
    101711.1,
  101467.4, 101540, 101623.7, 101691.3, 101745.4, 101793.3, 101833.1, 101869, 
    101892.9, 101909.8, 101911.8, 101899.5, 101894.9, 101885.9, 101883.3,
  101355.5, 101445.5, 101540.4, 101610.9, 101676.8, 101733.3, 101779.4, 
    101817.6, 101848.1, 101865.9, 101873.9, 101867.5, 101861.3, 101855.5, 
    101855.7,
  101247.2, 101346.3, 101431.7, 101517.2, 101591.9, 101659, 101714, 101760.1, 
    101792.7, 101817.5, 101830, 101834.9, 101833.6, 101831.7, 101834.8,
  101133.3, 101245.3, 101340.4, 101441.1, 101517.9, 101589.8, 101650.2, 
    101703, 101740, 101766.9, 101782.4, 101794.5, 101799.5, 101803.7, 101806.1,
  101014.5, 101137.3, 101234.1, 101343, 101423, 101499.5, 101570.1, 101630.3, 
    101677.2, 101712.2, 101736.6, 101755.2, 101761.4, 101770.5, 101776.5,
  100901.7, 101028, 101135.6, 101249.4, 101337.3, 101423, 101493.5, 101562.1, 
    101614.9, 101659.6, 101687.4, 101712.2, 101723.7, 101735.2, 101745.2,
  100792.1, 100919.2, 101036.6, 101153.9, 101247.8, 101338.7, 101417.8, 
    101487.7, 101546.7, 101599.3, 101634.8, 101664.3, 101681.8, 101698.7, 
    101713.7,
  100684.9, 100817.8, 100940.3, 101058.5, 101163.7, 101257.2, 101341.7, 
    101417.6, 101480.3, 101538.4, 101579.8, 101613.1, 101638.4, 101661.1, 
    101679.3,
  100583, 100720.5, 100846.2, 100968.8, 101075.1, 101178.4, 101264.7, 
    101344.6, 101413.5, 101475.4, 101524.8, 101564.4, 101596.3, 101625, 
    101646.8,
  100488.9, 100630.1, 100757.6, 100883.7, 100994.1, 101098.8, 101191.4, 
    101275.5, 101349.8, 101414, 101469.3, 101515.1, 101552.3, 101586.8, 
    101614.5,
  101902.9, 101994.3, 102084.8, 102163.1, 102235.6, 102295, 102345.5, 
    102374.7, 102384, 102379.4, 102361.9, 102333.7, 102306.7, 102269.8, 102226,
  101867.8, 101962.5, 102054.1, 102134.2, 102210.4, 102274, 102326.4, 
    102366.8, 102382.3, 102371.7, 102367.7, 102349.5, 102322.4, 102282.3, 
    102242.9,
  101849.9, 101943.5, 102032.8, 102116.8, 102192.7, 102259.8, 102313.6, 
    102351.3, 102376.1, 102380.3, 102371.7, 102349.3, 102321.9, 102286.8, 
    102254.5,
  101832, 101923.2, 102014.7, 102098.6, 102173, 102242.1, 102303.2, 102340.6, 
    102361.6, 102372.2, 102369.5, 102352.7, 102322.2, 102285.3, 102263.2,
  101813.8, 101905.1, 101994.8, 102079.4, 102154, 102224.4, 102284.9, 
    102328.5, 102352.8, 102365.7, 102364.4, 102350.7, 102319.1, 102291.9, 
    102269.3,
  101792.2, 101885.1, 101975.7, 102059.9, 102138.4, 102211.2, 102272.3, 
    102314.6, 102344.6, 102354.1, 102353.7, 102341.8, 102317.2, 102292.5, 
    102272.5,
  101771.8, 101865, 101956.9, 102042, 102122.7, 102193.7, 102251.9, 102296.9, 
    102324.6, 102337.1, 102338, 102332.3, 102309.3, 102293, 102273.3,
  101750.7, 101841.1, 101937.1, 102020.1, 102101.4, 102174.4, 102233.7, 
    102276.9, 102304.6, 102321.6, 102322.4, 102317.1, 102303.7, 102289, 
    102271.4,
  101724.1, 101817.9, 101916.5, 102001.2, 102078.3, 102151.7, 102206.3, 
    102251.5, 102282.5, 102300.1, 102309.4, 102304.3, 102295, 102284.3, 
    102263.2,
  101695.1, 101791.2, 101890.8, 101976.9, 102052.7, 102122.5, 102178, 
    102223.9, 102259.7, 102278.4, 102288.7, 102286.9, 102284.9, 102275.1, 
    102256.3,
  102230.6, 102309, 102414.3, 102480.5, 102548.6, 102593.2, 102631, 102641.5, 
    102637.7, 102608, 102573.7, 102533.5, 102488.6, 102441.5, 102396.2,
  102216.6, 102290.3, 102397.7, 102478.6, 102553.1, 102603.5, 102642.4, 
    102663.1, 102666.3, 102642.4, 102608, 102564.2, 102523.3, 102472, 102422,
  102205.8, 102299.8, 102409.6, 102493.9, 102566.5, 102620.3, 102659, 
    102684.5, 102685.7, 102673.7, 102638.1, 102595.1, 102550, 102502.1, 
    102450.7,
  102191.6, 102301.9, 102406.8, 102496.3, 102570.1, 102635.1, 102678.1, 
    102707.4, 102713.3, 102704.4, 102672.6, 102628.5, 102579.2, 102533.5, 
    102478.4,
  102189, 102311.5, 102412.3, 102507.1, 102584.7, 102650.6, 102699.1, 
    102727.9, 102739.6, 102728.2, 102699.2, 102659.5, 102612.1, 102563.1, 
    102509.2,
  102190.5, 102316.6, 102415.5, 102514.4, 102592.3, 102663.8, 102720.8, 
    102754.3, 102767.4, 102754, 102724.1, 102685.7, 102641.9, 102593.4, 
    102541.2,
  102197.2, 102325.6, 102424.7, 102522.3, 102606.6, 102681.6, 102739.2, 
    102777.5, 102793.3, 102779, 102748, 102714.7, 102668.3, 102620.9, 102567.5,
  102206, 102335.5, 102433.6, 102530.3, 102618.7, 102696, 102752.8, 102797.3, 
    102812.4, 102801.7, 102777.7, 102742.1, 102695.7, 102646.4, 102592.9,
  102217.3, 102347.1, 102444.7, 102541.1, 102630.5, 102713.9, 102774.3, 
    102822.3, 102832.6, 102822.3, 102800.8, 102765.1, 102720.3, 102674.6, 
    102616.2,
  102229.5, 102358.1, 102455.8, 102553.3, 102644.6, 102729.2, 102787.9, 
    102837.7, 102845.3, 102844.3, 102817.1, 102788.1, 102743.5, 102699.5, 
    102642.6,
  102707, 102719.6, 102727.6, 102730.6, 102726.8, 102718.5, 102725.5, 
    102719.9, 102707.6, 102663.7, 102624.1, 102578.7, 102540.3, 102493.2, 
    102448.3,
  102684.4, 102700, 102716, 102719.5, 102725.7, 102726.9, 102737.1, 102738.7, 
    102733.9, 102692.6, 102657.7, 102610.9, 102571.4, 102525.5, 102477.7,
  102667.3, 102693.8, 102715.6, 102716.8, 102731.2, 102737.6, 102751.3, 
    102762.1, 102756.3, 102721.4, 102683.4, 102639.3, 102601, 102558, 102510.5,
  102647.1, 102673.7, 102706.6, 102707.5, 102725.4, 102741.6, 102757.4, 
    102780.9, 102773.3, 102745.4, 102711.1, 102670.2, 102627, 102586.4, 
    102540.1,
  102613.7, 102647.3, 102691, 102702.9, 102722.2, 102743.3, 102767.3, 
    102787.6, 102788.6, 102768.4, 102733.4, 102696.4, 102655.6, 102613.4, 
    102564.6,
  102574.6, 102612.7, 102670.1, 102692, 102718.1, 102742.8, 102773.7, 
    102797.6, 102802.6, 102789.6, 102760.4, 102723.9, 102684, 102639.5, 102591,
  102528.8, 102577.4, 102643.9, 102681.6, 102716.2, 102746.8, 102780.8, 
    102806.7, 102816.6, 102808.2, 102782.3, 102750.4, 102706.9, 102665.4, 
    102617.5,
  102479.9, 102539.2, 102613.9, 102668.1, 102709.1, 102748.4, 102786.3, 
    102820.7, 102834.3, 102834, 102806.6, 102774.3, 102733.3, 102687.7, 
    102640.7,
  102432.4, 102497.7, 102585.1, 102652.2, 102704.3, 102751.4, 102791.3, 
    102832.9, 102848.5, 102848.5, 102825.6, 102794.9, 102757.9, 102712.1, 
    102664,
  102383.2, 102459.3, 102560.5, 102637.6, 102700.5, 102752.9, 102800.2, 
    102842.6, 102865.9, 102864.1, 102850.3, 102811.7, 102784.3, 102734.4, 
    102690.8,
  102891.6, 102891.1, 102889.8, 102875.1, 102859.4, 102831.5, 102814.8, 
    102782.3, 102743.9, 102697.2, 102659, 102617.3, 102573.8, 102526.7, 
    102475.5,
  102959.1, 102952.1, 102952.1, 102937.1, 102923.2, 102889.8, 102864.1, 
    102836.3, 102802.6, 102754, 102706.7, 102660, 102614.2, 102564, 102511.8,
  103016.6, 103010.2, 103005.6, 102986, 102971, 102942.5, 102910.5, 102882, 
    102847.4, 102799.4, 102751, 102702.7, 102655.6, 102608, 102548.5,
  103069.8, 103066, 103059.5, 103038.5, 103020.3, 102992, 102954.1, 102927, 
    102894.2, 102849.4, 102798.3, 102747.2, 102696.3, 102646.5, 102589.4,
  103114, 103113.3, 103104.4, 103086.3, 103061.7, 103029.7, 102987.3, 
    102962.9, 102932.8, 102892.5, 102840.7, 102790.7, 102739, 102689.1, 
    102630.5,
  103157.9, 103152.6, 103147.6, 103125.1, 103104.5, 103066, 103030, 102996.8, 
    102970, 102935, 102881, 102833, 102780.3, 102729.4, 102674.4,
  103191, 103183.4, 103183.3, 103158.5, 103140.8, 103101, 103068.6, 103019.9, 
    102999.6, 102971.6, 102918.3, 102870.9, 102819.7, 102765.9, 102713.7,
  103214.3, 103207.9, 103213.3, 103186.3, 103171.7, 103133.7, 103104, 
    103049.4, 103026, 103003, 102953.2, 102904, 102855.2, 102798, 102746.1,
  103226.6, 103226, 103230.9, 103212.3, 103194.5, 103162.7, 103124.7, 
    103079.4, 103045.6, 103026.6, 102984.6, 102936, 102890.7, 102831.3, 
    102778.1,
  103230.5, 103237.4, 103240.8, 103228, 103212, 103185.4, 103141.3, 103097.2, 
    103063.3, 103043.9, 103008.8, 102961.8, 102919.3, 102859.5, 102803.4,
  102332.9, 102368.7, 102402.4, 102419.9, 102433.2, 102436.3, 102434.9, 
    102428.8, 102420.4, 102405, 102389.2, 102365.2, 102339.5, 102312.2, 
    102281.7,
  102446.1, 102477.2, 102506, 102517, 102525.5, 102523.3, 102518.6, 102506.6, 
    102491.7, 102471, 102451, 102427.2, 102394.8, 102355.8, 102321.3,
  102563.9, 102581.8, 102601.5, 102610.6, 102614.7, 102609.1, 102599.2, 
    102583.5, 102563, 102539.5, 102512.8, 102482.5, 102449.4, 102407.2, 
    102364.8,
  102676.5, 102688.2, 102703.8, 102704.5, 102702.2, 102692.9, 102679.6, 
    102659.4, 102635.8, 102603.8, 102572.9, 102537.5, 102501.3, 102457, 
    102410.1,
  102778.5, 102788, 102797.7, 102794.3, 102788.1, 102773.2, 102757, 102730.1, 
    102704.7, 102667.4, 102633.1, 102592.6, 102552.3, 102508.2, 102457.2,
  102879.6, 102888.2, 102896, 102890.3, 102881.1, 102856.2, 102834.1, 
    102801.3, 102770, 102729.2, 102688, 102645, 102601.7, 102556.5, 102505.7,
  102983, 102988.6, 102994.8, 102986.4, 102975.2, 102946.5, 102912.1, 
    102870.6, 102832.5, 102789.1, 102742, 102695.8, 102650.3, 102602.4, 
    102553.1,
  103082.1, 103083.5, 103086.6, 103075.5, 103060.8, 103032.7, 102999, 
    102948.4, 102899, 102847.1, 102796.7, 102742.7, 102693.9, 102643.5, 
    102595.7,
  103174.8, 103171.5, 103171.4, 103155.7, 103134.9, 103104.5, 103070.7, 
    103024.8, 102967.7, 102909.5, 102853.6, 102793, 102737.2, 102681.5, 102632,
  103260.9, 103252.9, 103247.6, 103228.7, 103205.4, 103169.3, 103128.9, 
    103089.2, 103035.2, 102972.2, 102911.9, 102845.6, 102782.6, 102719.3, 
    102664.7,
  101624.4, 101627.3, 101670.2, 101710.3, 101757.5, 101802.1, 101852.9, 
    101896.6, 101940.4, 101964.6, 101994.7, 102020.4, 102044, 102053.1, 
    102058.2,
  101714.6, 101741.6, 101776.1, 101811.9, 101852.6, 101888.5, 101928, 
    101960.5, 101995.4, 102023.1, 102049.1, 102065.5, 102078.7, 102085.1, 
    102090.1,
  101886.2, 101903, 101908.2, 101929.5, 101957.2, 101985.2, 102017, 102043.8, 
    102069.3, 102088.9, 102105.2, 102117, 102126.3, 102128.5, 102126.5,
  102078.1, 102077.5, 102079.4, 102086.1, 102095.3, 102109.6, 102124.9, 
    102139, 102152.5, 102162.4, 102169.8, 102173.8, 102174.2, 102169.8, 
    102162.2,
  102281.9, 102263.7, 102254, 102245.3, 102244.6, 102242.1, 102240.6, 
    102238.8, 102241, 102240, 102239.7, 102236.9, 102231.5, 102220.1, 102202.6,
  102460.9, 102436.7, 102419.6, 102403.1, 102390.5, 102375.8, 102363.7, 
    102348.1, 102334.8, 102320.3, 102309.5, 102297.7, 102284.7, 102268.3, 
    102245.5,
  102611.4, 102585.3, 102568.1, 102545.6, 102528.1, 102504.6, 102484.3, 
    102458.3, 102432.5, 102405.9, 102381.1, 102358.8, 102339.4, 102316.7, 
    102288.7,
  102736.8, 102708.2, 102686.7, 102660.1, 102637.6, 102612.6, 102590.9, 
    102562.7, 102531, 102495.7, 102459, 102426.6, 102391.4, 102363.8, 102331.7,
  102851.7, 102818.2, 102792, 102762.3, 102734.1, 102705.7, 102676.3, 
    102646.2, 102612.3, 102574.9, 102535.6, 102495.3, 102450.2, 102412.4, 
    102373.9,
  102954.6, 102916.3, 102884.8, 102849.4, 102816.7, 102780.1, 102746.6, 
    102715.5, 102679.9, 102639.7, 102597.9, 102556, 102507, 102456.8, 102419.6,
  102242.7, 102250.7, 102287, 102302.4, 102318.6, 102324.7, 102325.4, 
    102317.6, 102303.9, 102275.6, 102256.9, 102219.3, 102185.7, 102146.7, 
    102088.4,
  102190.5, 102221.3, 102258.7, 102275.5, 102293.1, 102302.1, 102303.9, 
    102294.7, 102281.2, 102259.6, 102229.5, 102190.2, 102170.5, 102134.1, 
    102103.3,
  102160.2, 102190.6, 102223.8, 102252.1, 102271.4, 102278.4, 102279.8, 
    102272.6, 102259.1, 102238.1, 102207.2, 102181.6, 102157, 102115.4, 
    102096.7,
  102137.3, 102172.2, 102192.8, 102223, 102240.5, 102248.2, 102250.6, 
    102244.9, 102236.2, 102212.3, 102191.5, 102166.4, 102137.8, 102114.7, 
    102111.1,
  102133.9, 102167.5, 102183.9, 102207.1, 102220.8, 102232.8, 102234.9, 
    102229.8, 102213.1, 102197.4, 102177, 102157.5, 102134.6, 102128.9, 
    102136.4,
  102168.7, 102186, 102196.9, 102211.4, 102218.1, 102220.6, 102220.1, 
    102211.2, 102203.8, 102192.7, 102175.7, 102152.1, 102151.3, 102155.9, 
    102153,
  102216.2, 102224.2, 102225.9, 102227.6, 102232.6, 102231.1, 102226.5, 
    102217.9, 102209, 102185.5, 102161.8, 102165.9, 102176.9, 102180.9, 
    102176.6,
  102273.9, 102267.8, 102264.8, 102259.3, 102255.4, 102246.1, 102232.8, 
    102216.5, 102203.7, 102203.9, 102207.8, 102207.6, 102206.1, 102201.9, 
    102194,
  102336, 102317.8, 102307.8, 102294.1, 102286, 102275.4, 102268.5, 102260.9, 
    102254.1, 102246.7, 102242.5, 102240.6, 102233.8, 102235, 102218.1,
  102398, 102376, 102362, 102351.2, 102337.1, 102326.6, 102310.6, 102303.1, 
    102294.4, 102296.4, 102290.1, 102269.4, 102251.3, 102240.5, 102222.6,
  102881.7, 102846, 102807.7, 102766.5, 102722.3, 102666.8, 102611.5, 
    102552.3, 102498.2, 102435.7, 102376.2, 102329.6, 102290, 102210.9, 102142,
  102890.7, 102865.7, 102825.4, 102780.2, 102729.9, 102681.5, 102626.6, 
    102568.9, 102509.9, 102447.5, 102387.3, 102327.2, 102278.6, 102218.7, 
    102174.8,
  102899.6, 102866.8, 102830.2, 102788.1, 102739.2, 102687.5, 102629, 102567, 
    102507.7, 102450.7, 102391.6, 102333.8, 102288.3, 102221.3, 102175.8,
  102899.8, 102866.4, 102831.1, 102789.7, 102744.7, 102690.1, 102630.5, 
    102569.6, 102505.3, 102449.8, 102389.9, 102343, 102286, 102225, 102200.4,
  102891.9, 102857.9, 102823.1, 102783.5, 102737.3, 102680.8, 102622, 
    102562.9, 102495.6, 102438.3, 102384.9, 102346.9, 102277.6, 102238.2, 
    102229.5,
  102872.5, 102838.5, 102807.5, 102765.7, 102719.7, 102667.6, 102614.9, 
    102552, 102484.3, 102427.6, 102382.4, 102322.8, 102271.3, 102264.3, 
    102239.6,
  102843.9, 102811.1, 102780, 102739, 102698.4, 102645.3, 102598, 102538.4, 
    102477.7, 102422.6, 102353.2, 102305.7, 102288.7, 102277.9, 102253.2,
  102802.2, 102769.8, 102742.3, 102705.4, 102669.8, 102626.9, 102579.7, 
    102520.3, 102449.5, 102386.4, 102340.3, 102323.7, 102308.7, 102285.7, 
    102263.4,
  102749.7, 102717.2, 102689.8, 102656.2, 102624.4, 102581.5, 102534.9, 
    102482.4, 102432.8, 102385.5, 102366.6, 102348.8, 102320.6, 102294.1, 
    102268.1,
  102683.2, 102650.2, 102629.3, 102598.6, 102566.1, 102533.5, 102497.6, 
    102461.3, 102429.4, 102402.8, 102376.6, 102351.3, 102324.5, 102292.4, 
    102262.2,
  102706.2, 102646.1, 102588.9, 102518.6, 102444.6, 102379.5, 102321.1, 
    102274.7, 102231.7, 102175.4, 102133.7, 102089.3, 102052.2, 102028.2, 
    102005,
  102764.3, 102704, 102641.6, 102583.9, 102518.3, 102452, 102385.3, 102317.4, 
    102267.5, 102217.1, 102179.5, 102131, 102090.2, 102057.3, 102030.7,
  102804.9, 102744.5, 102680.1, 102623.5, 102558.9, 102499.6, 102434.5, 
    102364.4, 102308.2, 102256.8, 102205.7, 102161.8, 102119.6, 102085.9, 
    102067,
  102839.7, 102777.2, 102713.8, 102660.2, 102598.6, 102543.3, 102488.9, 
    102411.3, 102345.1, 102287.1, 102236, 102189.2, 102151.2, 102118.1, 
    102091.7,
  102861.6, 102798.5, 102732.3, 102678.6, 102623.2, 102567.5, 102513.8, 
    102456.1, 102382.3, 102328.2, 102257.7, 102209.7, 102177.6, 102150.5, 
    102116.5,
  102871.4, 102809, 102742.3, 102690.7, 102636.5, 102582.8, 102531.1, 
    102481.4, 102419.2, 102363.9, 102293.9, 102236, 102209.4, 102176.8, 
    102140.7,
  102869.3, 102805.8, 102744.1, 102686.8, 102635, 102582.9, 102534.5, 
    102486.8, 102439, 102382.6, 102321.3, 102267.6, 102242.2, 102199.7, 
    102162.8,
  102853.4, 102791.3, 102731, 102678.1, 102624.7, 102573.7, 102526.6, 
    102482.4, 102443.9, 102394, 102344.3, 102294.6, 102265.2, 102221.6, 
    102179.5,
  102831.4, 102772.8, 102713, 102655.7, 102605.1, 102553.7, 102507.8, 
    102471.6, 102433.4, 102390.9, 102346, 102302.6, 102270.3, 102225.8, 
    102186.5,
  102801, 102739.4, 102686.2, 102629.8, 102581, 102528.4, 102483.4, 102443, 
    102408.1, 102369.4, 102331.9, 102297.9, 102258.8, 102225.3, 102185.8,
  101962.5, 101932.5, 101911.4, 101901.4, 101896, 101882.9, 101873.2, 101869, 
    101868.6, 101859.1, 101850.7, 101834.4, 101818.9, 101796, 101772.9,
  102070.3, 102044.3, 102025.7, 102011.9, 102003.9, 101993, 101969.7, 
    101950.1, 101935.9, 101918.6, 101911.1, 101889.1, 101869.6, 101838.9, 
    101815.1,
  102180, 102142.8, 102118, 102101.4, 102087, 102073.4, 102056.2, 102028.1, 
    102007.5, 101975.7, 101958.2, 101939.5, 101913.4, 101879.6, 101852.1,
  102274.4, 102226.5, 102192.3, 102166.2, 102151.9, 102138.8, 102126.7, 
    102091, 102078.4, 102051.4, 102015.6, 101988.9, 101967.1, 101928, 101891,
  102354.8, 102305.5, 102264.4, 102230.3, 102202.3, 102179.4, 102164.6, 
    102143.5, 102114.8, 102096.2, 102068.8, 102029.3, 102008.1, 101973.1, 
    101927.1,
  102421.3, 102365.1, 102319.8, 102281.9, 102249.9, 102221.2, 102195.1, 
    102177.4, 102146.6, 102121.9, 102104.1, 102063.7, 102042.6, 102009.4, 
    101963.9,
  102478, 102421.2, 102367.8, 102325.3, 102287.1, 102250.1, 102221.4, 
    102193.8, 102167.2, 102139, 102110.5, 102082, 102058.7, 102029.4, 101996.3,
  102526.5, 102463.9, 102410.2, 102363.5, 102322, 102280.1, 102245.2, 
    102214.7, 102186.8, 102160.4, 102130.2, 102099.9, 102074.8, 102050.6, 
    102023.1,
  102564.2, 102499.8, 102443.6, 102390.5, 102347.5, 102303.8, 102266, 
    102230.1, 102199.3, 102172.9, 102149.7, 102117.2, 102086.9, 102067.6, 
    102042.1,
  102594.6, 102527.9, 102471.2, 102416, 102369.3, 102322, 102281.4, 102247.2, 
    102210.6, 102182.1, 102159, 102137, 102111.5, 102083.7, 102055.2,
  101772.4, 101783.3, 101822.1, 101843.4, 101809.7, 101760.2, 101767.3, 
    101788.1, 101779.9, 101765.6, 101756.2, 101752.1, 101747.6, 101740.4, 
    101729.1,
  101771.7, 101792, 101815.6, 101801.4, 101805.3, 101826.9, 101826.8, 
    101812.4, 101807.6, 101808, 101804.4, 101798, 101784.1, 101769.9, 101758.6,
  101797.5, 101824.6, 101818.2, 101824.9, 101857.2, 101867.3, 101866.9, 
    101871.7, 101873.7, 101862.6, 101847.4, 101834.3, 101826.9, 101813.2, 
    101797.4,
  101843.2, 101850.4, 101876.4, 101896.7, 101902.6, 101914.7, 101922, 
    101927.4, 101922.2, 101906.8, 101894, 101880.3, 101867.3, 101852, 101832.2,
  101907.6, 101922.8, 101942.2, 101954.5, 101967.5, 101980.7, 101983.1, 
    101979.5, 101970.2, 101948.3, 101935.5, 101921.3, 101908.5, 101888.5, 
    101866.1,
  101981.5, 101992.8, 101996, 102002.1, 102010.7, 102017.3, 102013.6, 
    102013.9, 102000.6, 101985, 101972.3, 101963.9, 101948.3, 101929, 101896.2,
  102065.8, 102066.1, 102061.8, 102063, 102061.6, 102058.2, 102048.4, 
    102044.4, 102028.4, 102018.8, 102005.6, 101997.7, 101980.7, 101960.3, 
    101932.7,
  102142.1, 102124.3, 102117.6, 102109.4, 102101.4, 102094.1, 102089.9, 
    102086, 102068, 102057, 102037, 102026.3, 102008.2, 101984, 101958,
  102206.7, 102181.6, 102175, 102157.5, 102147, 102128.7, 102119.3, 102118.6, 
    102110.5, 102093.8, 102070.5, 102052.1, 102033.7, 102011.5, 101987.2,
  102271.3, 102240.9, 102225.8, 102201.2, 102182, 102164.5, 102151, 102145.6, 
    102134, 102119.4, 102105.7, 102084.9, 102061.7, 102032.7, 102010.9,
  101593.2, 101575.7, 101605.1, 101656.1, 101620.4, 101531.5, 101506.6, 
    101520.9, 101525.5, 101543, 101562.8, 101584.2, 101598.5, 101608, 101616,
  101667.3, 101701.1, 101649.1, 101587.8, 101518.2, 101523.7, 101536.9, 
    101550, 101557, 101575.3, 101586.6, 101604.1, 101618.9, 101632.9, 101643.5,
  101647.8, 101627.1, 101532.6, 101516.4, 101547.4, 101561.9, 101570.4, 
    101595.2, 101613.2, 101631.6, 101639.4, 101654.5, 101665.4, 101670.1, 
    101673.3,
  101679.4, 101613.2, 101645.4, 101618.8, 101587.8, 101611.4, 101625.8, 
    101644, 101655.4, 101667.6, 101676.5, 101689.3, 101695.3, 101698.6, 
    101702.2,
  101710.8, 101693.3, 101674, 101659.9, 101676.5, 101685.6, 101695.8, 
    101701.7, 101716.2, 101724.9, 101731.7, 101734.3, 101735.9, 101735.6, 
    101735.4,
  101774.9, 101774.9, 101750.2, 101750.7, 101746, 101746.8, 101756.7, 
    101762.9, 101774.2, 101777.7, 101775.4, 101776.8, 101772.3, 101770.6, 
    101767.4,
  101868.6, 101868.8, 101844.1, 101838.2, 101827.1, 101823.5, 101825.1, 
    101825.6, 101824.6, 101825, 101821.3, 101817.9, 101812.4, 101807.5, 
    101800.2,
  101966.7, 101949.2, 101932.7, 101916.8, 101909.7, 101902.2, 101896.8, 
    101892, 101885.2, 101874.4, 101866.8, 101859.9, 101848.1, 101842.8, 
    101833.5,
  102054.5, 102014.5, 102009.9, 101987.9, 101980.5, 101971, 101973.3, 
    101965.9, 101956.6, 101933.6, 101918.2, 101903.7, 101888.6, 101880.1, 
    101867.7,
  102137.5, 102090.2, 102084.3, 102055.5, 102046.9, 102028.4, 102027.7, 
    102013.2, 102007.5, 101979.2, 101969.1, 101947.9, 101930.2, 101914.7, 
    101902.6,
  100906.6, 100998.7, 101071.1, 101152.1, 101228.9, 101282.3, 101328.3, 
    101364.3, 101386.2, 101403.5, 101417.3, 101433.4, 101446, 101460.4, 101471,
  100889.7, 100973.1, 101034.8, 101117.9, 101180.8, 101243.5, 101283.7, 
    101316.7, 101339.4, 101364.6, 101381.4, 101404.7, 101419.2, 101441.4, 
    101459.4,
  100942.5, 101006.1, 101058.1, 101128.6, 101177.5, 101226.8, 101255.7, 
    101283.9, 101307.3, 101333, 101355.6, 101391.3, 101414.3, 101443.3, 
    101466.3,
  100941.9, 101018.8, 101061, 101109.8, 101149, 101191.3, 101216.9, 101251.8, 
    101281.4, 101313, 101342.5, 101374.4, 101404, 101435.8, 101467.5,
  101030.6, 101057.6, 101075.1, 101111, 101132.9, 101164.8, 101189.3, 
    101227.5, 101260.4, 101300.1, 101335.3, 101372.6, 101410.7, 101446.2, 
    101478.3,
  101077.5, 101072.7, 101076.7, 101097.6, 101119.9, 101151.1, 101182.4, 
    101219.1, 101262.1, 101306.8, 101340.4, 101386.3, 101424.6, 101462.6, 
    101500.3,
  101204.4, 101178.9, 101161.7, 101162, 101173.4, 101193.9, 101222.9, 
    101258.5, 101293.8, 101333.1, 101375.3, 101415.3, 101451.5, 101495.7, 
    101533,
  101375, 101318.5, 101283.4, 101267.4, 101264.4, 101279.3, 101300.6, 
    101323.7, 101355.2, 101390.1, 101418.5, 101455.8, 101496.4, 101537.8, 
    101575.1,
  101540.9, 101478.3, 101435.4, 101407.6, 101392.4, 101394, 101401.6, 
    101417.5, 101434.1, 101454.2, 101480.5, 101516, 101551.2, 101588.1, 
    101623.3,
  101705.8, 101639, 101590.6, 101555.2, 101537.6, 101527.8, 101527.2, 
    101527.9, 101534.3, 101545.5, 101562.3, 101587.4, 101614, 101646.6, 101675,
  100509.4, 100613.5, 100731.4, 100870.6, 100976.5, 101069.9, 101143.9, 
    101205.8, 101257.7, 101306.9, 101353.1, 101391.7, 101418.8, 101436.3, 
    101437.7,
  100523.7, 100619.4, 100709.9, 100826.5, 100924.8, 101020.7, 101092.2, 
    101162.1, 101216.8, 101274.8, 101315.3, 101353.7, 101382.4, 101407.4, 
    101411.5,
  100598, 100661, 100716.6, 100816.2, 100901.9, 100992.6, 101065.4, 101136.4, 
    101189.5, 101244, 101286.1, 101326.8, 101357.4, 101382, 101388.9,
  100672.5, 100723.1, 100759.1, 100834, 100904.4, 100986.4, 101053.3, 
    101118.7, 101171.9, 101225, 101261.7, 101298.3, 101329.3, 101350.4, 
    101368.2,
  100741, 100776.5, 100807.9, 100861.6, 100919.2, 100987, 101046.8, 101105.1, 
    101153.7, 101197.7, 101235.1, 101274.6, 101301, 101325.5, 101355.9,
  100790.1, 100821.6, 100849.6, 100895.9, 100939.5, 100993.4, 101042.8, 
    101093.9, 101135.9, 101179.7, 101216.1, 101246.4, 101274.3, 101315.1, 
    101335.9,
  100829.1, 100852.8, 100886.2, 100919.4, 100957, 100997.2, 101044.2, 
    101087.3, 101125.2, 101165.7, 101190.2, 101224.3, 101262.5, 101301.8, 
    101315.9,
  100865.3, 100875.6, 100903.7, 100933.5, 100969.9, 101005, 101047.2, 
    101081.1, 101110.4, 101147.4, 101175.1, 101210.2, 101250.2, 101280.5, 
    101304.3,
  100879.2, 100898, 100913.4, 100940.5, 100975.7, 101004.2, 101041.9, 
    101073.1, 101104.4, 101135.3, 101161.9, 101196.8, 101229.1, 101263.8, 
    101307.7,
  100940.4, 100906.1, 100910.7, 100935.4, 100961.1, 100995, 101028.1, 
    101062.4, 101093.7, 101120.9, 101155.1, 101183.2, 101228.1, 101275.6, 
    101327.2,
  100965.6, 101016.8, 101106.7, 101184.9, 101258.4, 101328.9, 101396.6, 
    101458.6, 101505.6, 101546.7, 101577.7, 101604.3, 101621.6, 101633.7, 
    101641.7,
  100865, 100918, 101005.8, 101108, 101196.1, 101274.9, 101340.9, 101407.6, 
    101461.7, 101511.8, 101547.4, 101577.5, 101598.7, 101614.5, 101629.9,
  100810.4, 100862.9, 100918.2, 101012.3, 101112.2, 101207, 101286.8, 
    101360.4, 101425.4, 101479.6, 101521.8, 101556.5, 101583.2, 101603, 
    101619.3,
  100773.4, 100805.2, 100841.6, 100940.3, 101047.8, 101152.4, 101241.3, 
    101319.2, 101386.8, 101447.2, 101494, 101531.8, 101560.9, 101586.6, 
    101606.7,
  100754.6, 100779.6, 100791.3, 100874, 100972.8, 101085, 101186.6, 101271.6, 
    101344.8, 101413.2, 101465.1, 101509.1, 101541.4, 101573.3, 101593.2,
  100739.5, 100760.5, 100769.2, 100824.3, 100915.4, 101028, 101135.6, 
    101230.2, 101307.9, 101379.9, 101438.3, 101486.9, 101522.8, 101561.6, 
    101581,
  100727.4, 100738, 100752.3, 100792.7, 100871.5, 100978.9, 101087, 101186.2, 
    101269.9, 101348.6, 101413.4, 101465, 101508.8, 101548.1, 101573.9,
  100711.9, 100722.3, 100738.4, 100774.8, 100842.5, 100942.3, 101048, 
    101151.7, 101240.7, 101321.7, 101390.4, 101446.8, 101496, 101535.2, 101569,
  100714.6, 100716.5, 100727.7, 100761.1, 100827, 100915.2, 101020.2, 
    101123.4, 101214.7, 101300.5, 101370.1, 101432.9, 101483.4, 101524.5, 
    101558.6,
  100703.8, 100714.2, 100726.3, 100759.1, 100824.5, 100906.4, 101005.3, 
    101106.1, 101201.3, 101285.6, 101356.9, 101422.9, 101472.7, 101515, 
    101550.4,
  101320.5, 101357, 101392, 101423.3, 101458.5, 101490.9, 101522.8, 101553.5, 
    101579.6, 101601.6, 101624.3, 101639.3, 101660.6, 101675.4, 101690,
  101378.2, 101408.8, 101446.7, 101478.6, 101510.3, 101539.1, 101567.7, 
    101595.5, 101619.2, 101640.8, 101662.4, 101676.4, 101693.6, 101703.7, 
    101713.3,
  101430.5, 101461, 101498.1, 101525.2, 101553.8, 101581.2, 101607.1, 
    101633.5, 101650.7, 101670.8, 101693, 101710.3, 101721.7, 101730.6, 
    101738.5,
  101464.3, 101498.5, 101534.7, 101562.4, 101592, 101615, 101639.2, 101662.4, 
    101682.9, 101702.6, 101722.5, 101741.2, 101748.9, 101755.7, 101758.5,
  101489.1, 101528.8, 101566.2, 101596.1, 101626, 101651.5, 101670.8, 
    101692.3, 101710.3, 101731.7, 101748.2, 101763.5, 101775.8, 101781.2, 
    101779,
  101503.7, 101546.8, 101588.1, 101620, 101653.4, 101677.9, 101702.7, 
    101722.7, 101741.1, 101761.9, 101779.1, 101791.1, 101798.1, 101804.2, 
    101798.6,
  101515.5, 101561.9, 101608, 101644.2, 101678.3, 101704.4, 101730.6, 101752, 
    101771.8, 101788.3, 101803.6, 101819, 101826.8, 101821.2, 101822.7,
  101518, 101571.5, 101622.2, 101661.5, 101700, 101725.5, 101754.6, 101781.2, 
    101800.1, 101816.4, 101826.5, 101839.2, 101844.9, 101846.9, 101845.4,
  101518.8, 101577.9, 101632.6, 101676.2, 101715.6, 101745.3, 101774.4, 
    101802.7, 101823.8, 101840.2, 101850, 101860, 101866.1, 101869.3, 101865.6,
  101514.1, 101580.5, 101636.1, 101684, 101726.1, 101758.1, 101790, 101819.3, 
    101844.3, 101859.7, 101871.2, 101881.6, 101886.6, 101890.8, 101887.2,
  101078.9, 101161.2, 101250.1, 101325.4, 101391.8, 101440.4, 101483.1, 
    101506.8, 101531.4, 101543.7, 101548.2, 101551.3, 101562.3, 101566.3, 
    101578.3,
  101078.6, 101158.1, 101236.4, 101299.5, 101357.3, 101401.6, 101444.4, 
    101467.4, 101495.9, 101509.7, 101522.9, 101529.1, 101540.2, 101552.4, 
    101582.4,
  101088.2, 101150.3, 101220.2, 101282.5, 101338.4, 101380.3, 101422.6, 
    101449.9, 101475.7, 101497.1, 101511.8, 101530, 101545, 101567.6, 101596,
  101102.8, 101160.1, 101225.2, 101276, 101326.6, 101364.9, 101403.2, 
    101429.9, 101458.5, 101485, 101509, 101530.6, 101549.1, 101579.9, 101607.4,
  101147.7, 101190.7, 101244.8, 101287.5, 101334.6, 101366.9, 101404.2, 
    101432.1, 101461.4, 101488.5, 101515.7, 101542.2, 101567.3, 101602, 
    101623.7,
  101202.7, 101233, 101278.4, 101310.7, 101350.9, 101377.2, 101410.5, 
    101433.9, 101467.2, 101492.6, 101529.6, 101562.9, 101588.4, 101622.2, 
    101650.3,
  101262.8, 101283.3, 101316.6, 101345.1, 101379.9, 101403.2, 101432.9, 
    101457.5, 101490.5, 101524.9, 101558.9, 101583.8, 101623.2, 101653.4, 
    101683.4,
  101319.1, 101339.1, 101363.9, 101385.9, 101412.9, 101432.5, 101460.6, 
    101490.2, 101528.1, 101553.9, 101581, 101613.4, 101652.7, 101684.9, 
    101719.2,
  101396.6, 101413.2, 101430, 101448.6, 101469.7, 101489.5, 101519.4, 
    101545.7, 101569.7, 101589.2, 101621, 101657.1, 101691.2, 101726.3, 
    101757.8,
  101485.6, 101498.8, 101511.8, 101525.3, 101541.7, 101555.3, 101573.8, 
    101594.8, 101618.2, 101646.4, 101677.3, 101707.7, 101737.1, 101769.4, 
    101797.5,
  101795.2, 101875.7, 101948.8, 102006.8, 102054.9, 102094.4, 102119.2, 
    102135.6, 102133.1, 102125, 102105.3, 102072.8, 102034.4, 101988.1, 101939,
  101769.9, 101849.8, 101925.1, 101986.7, 102035.1, 102075.9, 102105.7, 
    102119.6, 102124, 102115.7, 102096, 102065.6, 102024.3, 101982.1, 101930,
  101762.4, 101841.4, 101912.2, 101970.5, 102022.2, 102061.4, 102089.8, 
    102108.8, 102107.6, 102101.6, 102078.6, 102041.9, 102000.9, 101959.1, 
    101913,
  101755.2, 101829.2, 101898.2, 101959.6, 102008.3, 102047.4, 102074.2, 
    102086.8, 102090.4, 102076.3, 102053.8, 102018.8, 101978.9, 101932.1, 
    101890.5,
  101748, 101818.2, 101883.8, 101941.5, 101988.7, 102022.6, 102048.2, 
    102057.6, 102057.6, 102041.3, 102016.5, 101984, 101939.9, 101900, 101864.5,
  101740.3, 101804.4, 101867.7, 101919.6, 101963.4, 101996.4, 102018.6, 
    102028.8, 102024.9, 102014.2, 101986.3, 101949.9, 101911.6, 101876.1, 
    101833.5,
  101729.7, 101785.5, 101846.1, 101891.4, 101930.9, 101960.7, 101982, 
    101991.2, 101987.7, 101966.4, 101940, 101912.2, 101881.1, 101839.8, 
    101808.3,
  101717.1, 101755.7, 101812.7, 101855.2, 101897.9, 101923.3, 101943.4, 
    101941.4, 101936.9, 101926, 101911.5, 101888.9, 101849.2, 101807.4, 
    101770.8,
  101684.1, 101723.2, 101777.2, 101811.2, 101846.1, 101864.6, 101883.6, 
    101892.7, 101895.9, 101892.4, 101872.1, 101830.6, 101804.1, 101787.4, 
    101773.9,
  101651.1, 101682.7, 101723.7, 101757.7, 101796.8, 101825.1, 101843.8, 
    101853.1, 101843.4, 101839.8, 101817.2, 101802.4, 101799.8, 101791.9, 
    101771.3,
  102073.7, 102167.8, 102246.9, 102317.1, 102370.9, 102413.3, 102433.3, 
    102448.6, 102445.7, 102431, 102405.3, 102368, 102329.1, 102287.3, 102241.1,
  102089.2, 102189.3, 102265.5, 102333.9, 102388.5, 102427.7, 102451.3, 
    102465.9, 102467.6, 102451.5, 102428.2, 102392, 102351.4, 102312, 102267.8,
  102103.2, 102199.7, 102276.8, 102348.1, 102406.2, 102446.6, 102469.7, 
    102489.2, 102488.9, 102472.6, 102448.4, 102410.5, 102359.3, 102321.2, 
    102278.8,
  102114.2, 102211.1, 102292.4, 102362.1, 102419.8, 102459.2, 102489.8, 
    102507.2, 102499.9, 102485.9, 102460.6, 102420.8, 102373.8, 102332.6, 
    102285.6,
  102127.5, 102221, 102299.8, 102368.6, 102426.9, 102462.4, 102491.3, 
    102510.3, 102508.7, 102494.6, 102472, 102426, 102377.5, 102331.1, 102280.3,
  102139, 102230.3, 102310, 102375.6, 102429.4, 102465.8, 102492.7, 102507.8, 
    102509, 102505, 102476.1, 102424.4, 102378.9, 102325.2, 102269.3,
  102148.1, 102237.2, 102315.3, 102376.5, 102427.6, 102465.7, 102487, 
    102504.6, 102509.1, 102503.8, 102471.7, 102421.1, 102371, 102303.2, 
    102242.4,
  102155.1, 102240.7, 102315.9, 102375.2, 102428.2, 102464, 102485.1, 
    102502.8, 102506.5, 102497.1, 102461.8, 102412.7, 102353, 102283, 102218.8,
  102156.2, 102239.4, 102313.2, 102371, 102422.4, 102457.9, 102480.6, 
    102500.4, 102500.1, 102483, 102448.1, 102395.4, 102329.1, 102255.9, 102197,
  102157.6, 102239.1, 102309.2, 102363.7, 102414, 102451, 102473.1, 102489.3, 
    102490.8, 102470.1, 102430.3, 102372.8, 102310.1, 102242.7, 102158.6,
  101902.6, 102025.1, 102118.2, 102204.3, 102270, 102325.1, 102359.4, 
    102378.8, 102383.5, 102376.7, 102364.2, 102344, 102319, 102289.9, 102256.9,
  101927.4, 102053.3, 102150.3, 102240, 102308, 102361.1, 102396.9, 102415.9, 
    102419.3, 102410.6, 102392, 102372.1, 102343.3, 102315.2, 102279.2,
  101965.7, 102094.7, 102195.3, 102284.3, 102351.9, 102402.8, 102438.4, 
    102452.3, 102450.7, 102440.1, 102419, 102396.6, 102365.4, 102332.8, 
    102294.2,
  101993.6, 102125.7, 102230.2, 102319.8, 102387.1, 102439.1, 102469.5, 
    102483.6, 102482.9, 102472.5, 102447.6, 102418.4, 102386.6, 102350.4, 
    102304.9,
  102024.2, 102156, 102264, 102352.1, 102421.8, 102470.9, 102499.1, 102512.5, 
    102511.8, 102497.5, 102471.6, 102439.5, 102401.8, 102361.5, 102315.1,
  102049.6, 102184.7, 102292.7, 102384, 102452.3, 102501.1, 102532.1, 
    102543.2, 102540.6, 102525.2, 102494, 102460.7, 102416.6, 102373, 102322.8,
  102076.2, 102212.3, 102320.1, 102409.3, 102476.9, 102528, 102557.8, 
    102571.1, 102569.6, 102550.8, 102517.5, 102479.9, 102431.4, 102382.6, 
    102331.5,
  102103.3, 102235.9, 102341.2, 102430.9, 102502.5, 102550, 102584.1, 
    102600.7, 102598.7, 102578.8, 102537.2, 102500.7, 102446.6, 102391.1, 
    102337.1,
  102129, 102258.4, 102361, 102451.8, 102521.3, 102572.1, 102609.7, 102627.1, 
    102624.3, 102607.8, 102563.6, 102523.6, 102464.4, 102409.6, 102346.2,
  102154.3, 102279.9, 102381, 102470, 102539.9, 102591, 102629, 102649.1, 
    102649.1, 102626.8, 102590, 102546.1, 102482.3, 102430, 102354.7,
  101671.6, 101714.7, 101775.8, 101823.6, 101868, 101915.6, 101962.7, 
    102016.2, 102070.5, 102117.7, 102148.2, 102171.1, 102179, 102163.4, 
    102144.9,
  101636.3, 101691.6, 101762.9, 101814.9, 101868.1, 101920.1, 101972.6, 
    102027.8, 102080.7, 102124.2, 102159.1, 102182.3, 102177.7, 102169, 
    102156.1,
  101625.6, 101679.1, 101758.8, 101821.7, 101887.2, 101944.3, 102000.1, 
    102053.2, 102103.1, 102142.2, 102172, 102190.2, 102192.9, 102177.6, 102164,
  101609.9, 101673.4, 101767.4, 101836.4, 101912.3, 101971, 102028.7, 
    102080.2, 102125.9, 102162, 102189.1, 102199.6, 102196.8, 102188.9, 
    102181.4,
  101602.1, 101679.8, 101776.4, 101853.3, 101933.2, 101998.6, 102062.5, 
    102110.8, 102151.4, 102182.9, 102199.3, 102200.2, 102199.8, 102198.1, 
    102195.4,
  101605.7, 101690.3, 101787.7, 101875.2, 101961.7, 102031, 102097.6, 
    102142.9, 102181.3, 102204.7, 102212.6, 102207.6, 102207.4, 102209.4, 
    102210.4,
  101615.5, 101709, 101814.5, 101910.1, 101995.5, 102069.8, 102133, 102178.1, 
    102210.7, 102228.6, 102233.8, 102226.6, 102222.1, 102224.3, 102228,
  101637.2, 101742.5, 101847.5, 101947.9, 102034.9, 102111.7, 102170, 
    102212.6, 102240.2, 102251.3, 102251, 102249.2, 102245.5, 102247.1, 102242,
  101670.5, 101782.4, 101889.7, 101994.6, 102080.5, 102152.5, 102206, 
    102250.5, 102271.6, 102286.5, 102287.2, 102286.4, 102278.9, 102269.3, 
    102265.6,
  101710.1, 101831.1, 101935.2, 102040.9, 102123.4, 102195.4, 102248.2, 
    102290.4, 102315.7, 102333, 102338.3, 102330.9, 102321.6, 102300.7, 
    102278.1,
  102209.5, 102221.6, 102244.5, 102256.5, 102261.6, 102255.2, 102240.5, 
    102209.6, 102180.8, 102152.1, 102146.9, 102170.2, 102178.9, 102171.4, 
    102165,
  102163.7, 102187.2, 102222.3, 102234, 102244.3, 102241.7, 102228.4, 
    102205.5, 102183.7, 102162.4, 102143.5, 102165.4, 102180.5, 102171.3, 
    102173,
  102143.1, 102168.4, 102199, 102214.1, 102233.1, 102229.2, 102222.3, 
    102204.7, 102179.2, 102167.4, 102147.4, 102166.2, 102181.4, 102177.5, 
    102183.6,
  102114.2, 102140.9, 102177.1, 102195, 102209.8, 102210.3, 102206.3, 
    102193.7, 102171, 102165.1, 102150.4, 102164.8, 102176.9, 102186.3, 
    102190.1,
  102081.4, 102111.3, 102148.7, 102168.6, 102182.5, 102189, 102184.3, 
    102176.4, 102162, 102160, 102151.6, 102166.3, 102176.3, 102192, 102204.3,
  102048, 102080.2, 102118, 102139.5, 102158.2, 102167.2, 102161, 102158.2, 
    102151.9, 102155.1, 102150, 102165.7, 102178.2, 102197.8, 102212.7,
  102010.9, 102045.4, 102084.9, 102109.1, 102130.2, 102139.4, 102137.9, 
    102140.2, 102141, 102146.2, 102149.2, 102160.8, 102180.5, 102201.6, 
    102218.2,
  101973.3, 102005.2, 102048.7, 102076.4, 102099.4, 102111.2, 102118, 
    102122.7, 102130.1, 102137.7, 102141.4, 102156.3, 102180.1, 102202.9, 
    102217.6,
  101931, 101967.1, 102011.2, 102039.7, 102065.9, 102086.4, 102095.9, 
    102107.8, 102117.5, 102131.1, 102135.1, 102157.9, 102180.3, 102205.4, 
    102226.9,
  101886.9, 101925.7, 101971.5, 102002.4, 102035.5, 102058.4, 102077.1, 
    102091.5, 102109.8, 102121.6, 102133.7, 102161.9, 102190.2, 102215.6, 
    102238.7,
  102359.6, 102372.3, 102396.5, 102405.7, 102412.1, 102406.4, 102405.3, 
    102384, 102366.4, 102340, 102320.3, 102329.8, 102331.1, 102319.5, 102303.5,
  102399.3, 102412.5, 102437.5, 102445.6, 102450.3, 102438.4, 102434.2, 
    102412.3, 102389.1, 102369.7, 102332.2, 102329.6, 102338.6, 102327.2, 
    102314.3,
  102445.1, 102450.9, 102468.8, 102472.3, 102481.2, 102462.2, 102452.8, 
    102436.5, 102401.2, 102392.9, 102353.8, 102322.4, 102334.4, 102342.5, 
    102332,
  102496.6, 102490.6, 102499.2, 102500.8, 102501.2, 102494.8, 102472.3, 
    102461.6, 102418.8, 102401.3, 102374.7, 102320.5, 102334.2, 102348.6, 
    102347.2,
  102546.1, 102529.7, 102528.9, 102528.4, 102523.6, 102513.6, 102492.3, 
    102476.3, 102444, 102413, 102377.2, 102329.8, 102342.2, 102342.7, 102355.9,
  102601.7, 102570.1, 102561.8, 102552.1, 102545.8, 102536.1, 102513.1, 
    102488.2, 102461.9, 102426.9, 102399.4, 102340.5, 102344.3, 102345.5, 
    102357.4,
  102646.8, 102609.9, 102587.3, 102574, 102563.1, 102548.6, 102534.7, 
    102498.6, 102476.8, 102433.8, 102408.6, 102344.6, 102343.3, 102343.9, 
    102360.7,
  102686.8, 102651.3, 102614.7, 102594.8, 102576.5, 102561.6, 102549.7, 
    102510.3, 102487.9, 102439.7, 102415.2, 102349.2, 102343, 102338.9, 
    102365.4,
  102706.6, 102685.8, 102642.8, 102615.1, 102592.4, 102574.1, 102558.2, 
    102522.1, 102492.6, 102445.3, 102418.2, 102353.7, 102338.7, 102340.9, 
    102362.2,
  102718.2, 102699, 102666.4, 102625, 102604.6, 102580, 102565.6, 102531.3, 
    102496.5, 102451.4, 102415.9, 102363.9, 102340, 102349.1, 102378.9,
  101666.5, 101724.7, 101797, 101865.7, 101934.2, 101999.4, 102060.6, 102113, 
    102164.3, 102213.9, 102259, 102292.6, 102310.4, 102317.8, 102295.9,
  101638.4, 101699.3, 101766.9, 101838.2, 101909.7, 101977.8, 102040.8, 
    102100, 102151.6, 102198.2, 102241.1, 102280, 102302.9, 102317.3, 102299.6,
  101626.9, 101684.1, 101747.1, 101818.5, 101892.9, 101964.3, 102029, 
    102090.6, 102143, 102188.6, 102231, 102259.8, 102299.8, 102320.7, 102308.8,
  101625.6, 101682, 101740.9, 101808, 101882.7, 101956.6, 102021.3, 102081.5, 
    102134.6, 102181.1, 102223.6, 102248.9, 102289.6, 102321, 102313.6,
  101634.3, 101687.3, 101737.2, 101801.6, 101875.8, 101949, 102015.3, 
    102077.7, 102128.8, 102172.2, 102210.8, 102234.2, 102273.5, 102301.6, 
    102306.7,
  101657.7, 101703.3, 101755.4, 101813.6, 101879.3, 101950.2, 102018.2, 
    102076.2, 102130, 102171.3, 102214.2, 102228.2, 102259.2, 102295.6, 
    102304.4,
  101694.1, 101735, 101781.6, 101832.6, 101895.8, 101958.7, 102025.4, 
    102079.2, 102135.4, 102172.2, 102212.9, 102222.8, 102247.2, 102277.3, 
    102303.5,
  101752.1, 101783.1, 101823.2, 101865.9, 101923.8, 101981.8, 102043.8, 
    102089.1, 102146.4, 102177.2, 102209.7, 102222.8, 102239.6, 102264.6, 
    102308.3,
  101826.6, 101851, 101884.7, 101922, 101972, 102021.1, 102072.8, 102108, 
    102162.4, 102184.9, 102212.6, 102215, 102217.6, 102252.3, 102298.4,
  101919.1, 101934.3, 101958.5, 101991.7, 102029.4, 102074.1, 102112.6, 
    102146.1, 102181.4, 102199.2, 102218.4, 102207.3, 102200.8, 102250.3, 
    102298.5,
  102123.3, 102185.4, 102235.1, 102272.9, 102289.1, 102300.2, 102304.5, 
    102291.2, 102276.2, 102261.2, 102247.1, 102246.7, 102250.7, 102259.8, 
    102274.7,
  102097.3, 102159.6, 102210.1, 102250, 102267.8, 102286.5, 102293.4, 
    102285.3, 102270.5, 102254.2, 102234.2, 102229.1, 102229.1, 102244.3, 
    102260.2,
  102075.5, 102132.4, 102182.6, 102221.3, 102241.7, 102258.9, 102271.4, 
    102268.5, 102258.6, 102242.7, 102227.3, 102219.8, 102224, 102237.5, 
    102262.1,
  102050.2, 102101.1, 102151.2, 102192.6, 102221, 102237, 102248.9, 102247.1, 
    102242.9, 102225.6, 102214.4, 102206.2, 102211.1, 102223.3, 102254.5,
  102016.7, 102065.4, 102117.1, 102151.1, 102183.8, 102206.8, 102214.7, 
    102221, 102220.4, 102205, 102202.8, 102195.1, 102198.8, 102217.9, 102240.7,
  101983.1, 102029.9, 102079, 102114.3, 102144.5, 102171.8, 102185.8, 
    102197.2, 102200.1, 102184.6, 102184.9, 102179.1, 102188.6, 102203.6, 
    102224.9,
  101942.9, 101984.7, 102033.8, 102071.3, 102100.5, 102128.8, 102147.7, 
    102162.1, 102173.2, 102162.9, 102164.5, 102161.9, 102171.9, 102192.5, 
    102216.5,
  101889.5, 101930.8, 101974.5, 102016, 102052.5, 102080.3, 102102.7, 
    102122.9, 102140.2, 102140.6, 102143.2, 102140.4, 102157.6, 102174.2, 
    102205.2,
  101827.5, 101866.7, 101910.1, 101950.8, 101992.6, 102025.8, 102055.1, 
    102077, 102098.2, 102109.8, 102118, 102122.6, 102137.7, 102155.3, 102187.8,
  101761.9, 101792.6, 101833.6, 101873.6, 101921.8, 101964.9, 102000, 
    102029.5, 102056.9, 102078.5, 102092.1, 102102.7, 102118.1, 102138.2, 
    102173,
  102111.1, 102181.2, 102253.6, 102322.4, 102380.3, 102426.3, 102456.2, 
    102475.5, 102478.4, 102469.7, 102449, 102419.5, 102383, 102328.6, 102286.9,
  102065.9, 102143.8, 102216.7, 102286.1, 102346.3, 102396.5, 102436.1, 
    102466, 102478.4, 102474.8, 102454.6, 102427, 102385.7, 102335.4, 102294.8,
  102030.6, 102106.4, 102183.7, 102254.3, 102317.1, 102369.9, 102413.1, 
    102445, 102469.1, 102470, 102447.3, 102426.1, 102385.4, 102333.9, 102294.1,
  101995.6, 102073.2, 102153.2, 102220.5, 102285.6, 102340.9, 102392.6, 
    102430.5, 102450.3, 102459.5, 102447.7, 102420.9, 102384.8, 102336.6, 
    102296.7,
  101962.7, 102038.5, 102116.7, 102187.4, 102253.5, 102309.9, 102363.9, 
    102408.6, 102435.9, 102448.8, 102444.6, 102415.8, 102384, 102335.3, 
    102297.8,
  101933.1, 102006.4, 102083.9, 102154.7, 102221.6, 102282.3, 102335.6, 
    102383.1, 102413.6, 102432.2, 102429.4, 102403.3, 102379.3, 102339.9, 
    102295.6,
  101909.3, 101980.8, 102055.1, 102123.7, 102191.2, 102253.7, 102306.6, 
    102361.1, 102396.2, 102418.8, 102415.9, 102402.7, 102373.1, 102336.8, 
    102289.7,
  101887.7, 101959.9, 102031.6, 102097.2, 102162.8, 102225.7, 102282.2, 
    102330, 102373.1, 102399, 102399.5, 102388.8, 102361.6, 102328, 102288.2,
  101865.5, 101941.3, 102007.7, 102073.5, 102136.7, 102196.9, 102254.9, 
    102302, 102341.1, 102372.8, 102385.7, 102377.7, 102351.4, 102323.7, 
    102283.1,
  101845.1, 101918.6, 101984.8, 102049.7, 102111.1, 102170.9, 102227.4, 
    102274.7, 102312.4, 102348.7, 102362.6, 102358.5, 102337.6, 102311.9, 
    102277.3,
  102314.5, 102398.7, 102472.6, 102529.8, 102577.3, 102610.7, 102634.5, 
    102642.2, 102629.5, 102612, 102583.3, 102550.7, 102510.3, 102455.8, 
    102406.8,
  102273.4, 102363.5, 102444.5, 102507.4, 102557.5, 102594.5, 102626.8, 
    102638.2, 102640.1, 102626.1, 102599.5, 102570.3, 102532.5, 102482.5, 
    102435.8,
  102241.2, 102336.6, 102419.8, 102489.2, 102542.3, 102580.9, 102612.9, 
    102629.7, 102636.4, 102631.4, 102610.4, 102585.1, 102550.4, 102499.9, 
    102451.6,
  102210.2, 102307.6, 102395, 102465.3, 102520.6, 102563.7, 102596.2, 
    102619.2, 102628.6, 102628.9, 102619, 102594.4, 102562.9, 102520.4, 
    102472.9,
  102182.7, 102280.2, 102368.4, 102440.7, 102500, 102547.3, 102578.7, 
    102603.2, 102620.5, 102624.8, 102619.8, 102598.6, 102568.4, 102533.9, 
    102485.6,
  102158.9, 102252.8, 102341.1, 102415.1, 102477.6, 102526.6, 102564.1, 
    102587.9, 102606.1, 102613.1, 102614.8, 102596.5, 102575.9, 102546, 
    102499.5,
  102141.8, 102229.2, 102316.1, 102388.1, 102451.4, 102505.1, 102541.7, 
    102572.3, 102590.1, 102600.3, 102600.8, 102588.6, 102577, 102548.6, 
    102505.8,
  102127.5, 102206.8, 102290.9, 102360.3, 102423.6, 102480.8, 102521.2, 
    102551.3, 102570.3, 102584.9, 102586.5, 102582.4, 102569.9, 102546.2, 
    102511.5,
  102113.7, 102186.4, 102268, 102335.6, 102396.3, 102450.9, 102494.4, 
    102527.7, 102549.4, 102566, 102568.3, 102567.2, 102557.1, 102541.8, 102512,
  102097.7, 102162.5, 102239.4, 102307.6, 102368.3, 102420.2, 102464.2, 
    102498.3, 102526.4, 102543.7, 102549.5, 102550.1, 102543.2, 102532.2, 
    102508.7,
  102028.6, 102097.9, 102161.6, 102220.1, 102274.6, 102316, 102339.8, 
    102352.8, 102355.8, 102349, 102338.5, 102316.6, 102288.9, 102258.5, 
    102226.6,
  102069.5, 102139.8, 102205.2, 102261, 102311.7, 102348.1, 102372.5, 
    102388.7, 102390.5, 102385.3, 102372, 102350.2, 102323.2, 102291.3, 
    102252.8,
  102113.4, 102181.7, 102249.2, 102299, 102346.6, 102380.4, 102404.2, 
    102414.7, 102419.3, 102416, 102401.7, 102380.3, 102351.5, 102321.6, 102287,
  102145.1, 102214.4, 102281.3, 102332.9, 102378.5, 102408.6, 102434.7, 
    102444.9, 102448.8, 102444.5, 102434.4, 102413.5, 102382.3, 102350.9, 
    102314.3,
  102170.6, 102237, 102306.8, 102357.3, 102402.8, 102430.9, 102457.6, 102466, 
    102475.2, 102476.9, 102460.7, 102441.7, 102410.9, 102377.8, 102340.3,
  102180, 102248.5, 102320.3, 102373.5, 102417.8, 102449.6, 102477.2, 
    102493.2, 102495.6, 102501.7, 102486.8, 102466.7, 102436, 102401.9, 
    102365.6,
  102187.7, 102254.3, 102326.9, 102381.9, 102431.1, 102464.4, 102494.9, 
    102510.6, 102517, 102522.8, 102503.8, 102488.5, 102457.6, 102423.9, 
    102388.4,
  102191.7, 102258.1, 102330.3, 102383.2, 102437.4, 102474.9, 102511, 
    102531.1, 102538.4, 102540.5, 102529.5, 102505.5, 102481.3, 102442.7, 
    102407.9,
  102204, 102261.3, 102331.3, 102385.5, 102439.8, 102479.4, 102515.6, 
    102539.4, 102550.7, 102552.5, 102544.8, 102525.1, 102497.1, 102459.1, 
    102423.1,
  102210.5, 102264.3, 102334.4, 102386.3, 102439.8, 102481.5, 102519.4, 
    102545.1, 102559.5, 102564.4, 102556.4, 102539.4, 102514.8, 102475.7, 
    102437.7,
  102186.2, 102208.7, 102238.4, 102248.1, 102252.2, 102244.6, 102233.6, 
    102217.4, 102199.8, 102204.1, 102202.6, 102189.9, 102175.6, 102160.8, 
    102140.9,
  102119.2, 102154.5, 102195.1, 102213.9, 102228.4, 102231.8, 102231.3, 
    102233.6, 102219.8, 102217.4, 102218.7, 102219.7, 102205, 102180.7, 
    102156.4,
  102058.8, 102110.7, 102161.5, 102191.9, 102219.2, 102232.1, 102245.8, 
    102254.2, 102246.2, 102243.7, 102246.5, 102237.5, 102224.9, 102208.4, 
    102183.3,
  102002.1, 102067.3, 102124.4, 102167.8, 102202.6, 102225.8, 102249.6, 
    102261.4, 102262.5, 102265.1, 102270.3, 102263.8, 102251.2, 102229, 
    102202.9,
  101953.5, 102028.6, 102095, 102150.6, 102193.7, 102229.1, 102258.9, 
    102273.4, 102281.9, 102288.9, 102292.7, 102289.8, 102275.4, 102253, 102228,
  101913.9, 101998.9, 102073.3, 102137.2, 102186, 102227.2, 102262.6, 
    102286.3, 102302.8, 102315.1, 102324, 102315.7, 102301.8, 102278.5, 
    102248.9,
  101883.3, 101976.7, 102058.6, 102129.5, 102185.1, 102234.9, 102275.4, 
    102305.9, 102326.6, 102344.8, 102350.1, 102346.1, 102324.7, 102305.2, 
    102274,
  101863.5, 101965.2, 102051.9, 102130.4, 102191.2, 102245, 102288, 102321.5, 
    102344.9, 102360.7, 102367.2, 102364.3, 102348.1, 102326.1, 102300.2,
  101853.1, 101960, 102051.3, 102133, 102199.3, 102252.6, 102299.9, 102336.4, 
    102365.8, 102385.6, 102393.8, 102391.2, 102379.7, 102351, 102319.6,
  101853, 101960.2, 102053.8, 102137.1, 102204.6, 102264.3, 102313.8, 
    102353.2, 102386.6, 102404.1, 102412.5, 102415.2, 102398.1, 102373.7, 
    102337.2,
  103113.2, 103048.3, 102967.4, 102881, 102794.6, 102717.5, 102620.3, 
    102537.9, 102467.2, 102416.3, 102387.4, 102339.1, 102303.1, 102260.9, 
    102215.3,
  103153.5, 103089.6, 103015.6, 102932.5, 102841.4, 102770.8, 102675, 
    102588.4, 102505, 102438.5, 102416.8, 102378.9, 102335, 102287.3, 102240,
  103173.2, 103114.3, 103041.8, 102970.7, 102879.8, 102802, 102707.8, 
    102626.3, 102544.9, 102475.3, 102446.2, 102403.5, 102362.8, 102318, 102270,
  103190.3, 103135.5, 103071.5, 103004.9, 102915, 102842.3, 102748.5, 
    102663.4, 102577.4, 102500.6, 102470.4, 102437.1, 102393.3, 102345.8, 
    102296.4,
  103203, 103148.7, 103090.4, 103024, 102943.1, 102869.1, 102778.5, 102698.2, 
    102607.8, 102531.6, 102494.1, 102464.1, 102419.1, 102373.2, 102325.1,
  103207.5, 103155, 103103.8, 103037.9, 102966, 102891, 102804.8, 102724.3, 
    102638.2, 102559.7, 102517, 102491.6, 102446.2, 102401.1, 102348.1,
  103199, 103154.3, 103104.9, 103045.7, 102976.5, 102904.8, 102826.4, 
    102744.6, 102664.8, 102583.7, 102539.9, 102514, 102469.9, 102426.3, 
    102372.1,
  103188.4, 103144.5, 103100, 103047.2, 102982.5, 102916.8, 102842.2, 
    102761.1, 102679.8, 102603.9, 102558.3, 102528.8, 102495.1, 102446.5, 
    102393.5,
  103165.2, 103129.9, 103087.2, 103041, 102982, 102920.7, 102842.9, 102771.5, 
    102691.8, 102622.8, 102578.3, 102547.9, 102513.9, 102466.1, 102413.5,
  103130.2, 103105, 103068.4, 103028.6, 102976.4, 102917.3, 102846.8, 
    102773.4, 102699.5, 102636.9, 102581.9, 102562.1, 102528, 102481, 102429.4,
  102818.1, 102772.9, 102734.2, 102695.7, 102656.8, 102616.4, 102573.2, 
    102530.5, 102492.4, 102456.2, 102414.9, 102367.5, 102317.9, 102267.9, 
    102215.8,
  102931.9, 102878.7, 102833.8, 102791.4, 102750, 102700.5, 102644.3, 
    102585.9, 102537.5, 102495.7, 102454.4, 102405.9, 102353.9, 102301.8, 
    102250.6,
  103041.1, 102978.8, 102930.3, 102868.4, 102818, 102762.7, 102710.9, 
    102649.2, 102590.2, 102536, 102492.6, 102441.6, 102388.1, 102332.6, 
    102278.8,
  103137.3, 103078.2, 103025.1, 102962.9, 102902.7, 102845.1, 102772.6, 
    102708.5, 102640.5, 102579.9, 102529.9, 102477.3, 102420.5, 102364, 
    102307.3,
  103222.9, 103163.9, 103106, 103047.2, 102976.3, 102913, 102845.4, 102768.5, 
    102701.4, 102627, 102566.7, 102509.9, 102451.3, 102389.9, 102332,
  103309, 103245.9, 103185, 103122.1, 103056.6, 102983.7, 102901.5, 102820.4, 
    102756.9, 102676.4, 102606.9, 102542.6, 102482, 102417.8, 102357.4,
  103381.2, 103318.4, 103255.6, 103187.1, 103120, 103048.7, 102972.1, 
    102885.5, 102809, 102725.5, 102646.8, 102576.6, 102509, 102441.7, 102379.5,
  103447.7, 103382.4, 103316.3, 103252, 103180.3, 103107.3, 103026, 102939, 
    102853.8, 102772.5, 102686.7, 102610.3, 102536, 102466.9, 102401.8,
  103499.9, 103439.2, 103370.8, 103302.9, 103233.1, 103159.2, 103080.8, 
    102997, 102903.9, 102813.7, 102727, 102641.8, 102562.4, 102489.3, 102420.7,
  103538.7, 103483.2, 103416.2, 103344.6, 103273.8, 103199.3, 103126.2, 
    103038, 102949.2, 102853.7, 102764.4, 102674.8, 102588.5, 102512, 102440.1,
  102008.6, 102079.8, 102120.1, 102166.4, 102198.7, 102206.9, 102209, 
    102197.5, 102181.5, 102155.2, 102126.5, 102093.1, 102057.4, 102021.6, 
    101981.9,
  102078, 102162, 102205.8, 102245.9, 102267.4, 102273.5, 102270.7, 102251.2, 
    102228.7, 102199.7, 102166.9, 102129.4, 102089.1, 102051, 102008.9,
  102188.4, 102251.8, 102290.1, 102319.7, 102337.8, 102340.8, 102335.7, 
    102313.1, 102283.1, 102245.3, 102207.3, 102168.2, 102125.6, 102084.4, 
    102041,
  102297.9, 102342.5, 102384.1, 102402.8, 102411.2, 102413.2, 102400.3, 
    102376.8, 102345.5, 102301.4, 102255.7, 102211.2, 102162.8, 102117.2, 
    102069.3,
  102416.9, 102446.4, 102484.1, 102492.8, 102496.1, 102483.6, 102460.9, 
    102432.3, 102400, 102359.6, 102307.8, 102258.2, 102204.5, 102155.3, 
    102102.3,
  102526.9, 102545.1, 102574.2, 102575.8, 102576.6, 102558.3, 102535.1, 
    102487.8, 102453.8, 102410.4, 102361.6, 102307.3, 102251.4, 102194.3, 
    102137.2,
  102636.8, 102645.6, 102666.2, 102659, 102652.3, 102628.6, 102599.1, 102555, 
    102504.3, 102460.7, 102410.6, 102356.6, 102297.4, 102236.7, 102177.2,
  102744.1, 102740.1, 102751.3, 102740.2, 102722.3, 102695.6, 102663.9, 
    102620.5, 102562.5, 102508.9, 102460.4, 102403.1, 102344.9, 102277.9, 
    102214.3,
  102843, 102834, 102834.6, 102816.8, 102794.5, 102761.4, 102726, 102678.1, 
    102627.1, 102559, 102510.7, 102449.3, 102387.4, 102321.1, 102249.8,
  102929.1, 102918.1, 102908.8, 102887.2, 102860.9, 102823.4, 102783.9, 
    102733.5, 102677.5, 102613, 102557.6, 102495.2, 102433.1, 102360.2, 
    102286.5,
  101428.2, 101536.1, 101578.5, 101655.7, 101714.3, 101763.1, 101797.2, 
    101822.8, 101835.1, 101841.7, 101839.5, 101830.2, 101816.3, 101797.6, 
    101770.6,
  101481.2, 101610, 101659.8, 101741.2, 101788.3, 101835.1, 101860.7, 
    101878.7, 101885.7, 101888.5, 101881.3, 101871, 101851, 101829.1, 101800.4,
  101586.8, 101703.9, 101751.3, 101819.6, 101860.7, 101905.2, 101925.8, 
    101940.6, 101942.8, 101939.5, 101928, 101913.2, 101890.6, 101866.4, 
    101834.9,
  101697.3, 101789.3, 101845.7, 101905, 101943.1, 101979.2, 101997.5, 
    102005.8, 102003.4, 101994.4, 101978.9, 101958.8, 101931.9, 101903.8, 
    101869.1,
  101817.2, 101888.3, 101947.2, 101994.1, 102028.9, 102055.4, 102065.9, 
    102068.7, 102063.6, 102050.4, 102032, 102009.8, 101979.2, 101946.5, 
    101909.2,
  101932.5, 101991.4, 102048.1, 102086.6, 102113.9, 102132, 102139.4, 102137, 
    102127, 102108, 102085.1, 102060.7, 102029.7, 101993.2, 101949.8,
  102041.3, 102098.4, 102143.8, 102174.9, 102196.5, 102208.7, 102209.9, 
    102204.4, 102191, 102173.1, 102145, 102113.1, 102081.7, 102042.8, 101993.8,
  102140.3, 102193.3, 102228.2, 102258.2, 102275.6, 102282.3, 102280.8, 
    102268.2, 102257.1, 102237.1, 102206.3, 102167.6, 102131.3, 102089.8, 
    102038.6,
  102240.8, 102292, 102326.6, 102348.9, 102359.7, 102358, 102351.3, 102334.6, 
    102315.9, 102293.4, 102263.2, 102219.9, 102177.2, 102134.9, 102079.8,
  102345.7, 102378.7, 102412, 102423.6, 102433.2, 102426.5, 102417, 102396.5, 
    102371.4, 102342, 102305.8, 102264.1, 102214.7, 102172.4, 102118.8,
  101321.1, 101330.2, 101336, 101338.6, 101356, 101402, 101463, 101507, 
    101552.4, 101590.1, 101619.6, 101640.9, 101650.4, 101650.5, 101641.5,
  101298.5, 101361.5, 101352.3, 101388.8, 101402.9, 101448.8, 101499.4, 
    101552.9, 101601.9, 101638.7, 101664.8, 101677.6, 101682.5, 101678.9, 
    101668.7,
  101448.5, 101320.9, 101371.5, 101398.9, 101460.2, 101511.7, 101574.3, 
    101622.7, 101661.4, 101690.4, 101711.4, 101723.1, 101724.5, 101716.4, 
    101703.2,
  101369.5, 101312.6, 101434.7, 101459.6, 101524.2, 101585.6, 101645, 
    101685.9, 101719.8, 101744.5, 101761.7, 101767.5, 101763.6, 101752.1, 
    101735.1,
  101394.8, 101426.3, 101494.1, 101538.5, 101615.3, 101672.4, 101723.9, 
    101759, 101790.7, 101809.6, 101817.9, 101817.4, 101807.5, 101791.2, 
    101769.9,
  101449.9, 101538.3, 101575.5, 101651.9, 101711.1, 101764.4, 101805.1, 
    101838.8, 101858.3, 101871.2, 101872.6, 101868, 101854.7, 101835.2, 
    101811.8,
  101541.4, 101666.8, 101691.9, 101768.7, 101808.9, 101861.1, 101892.5, 
    101917.9, 101932.5, 101937.4, 101929.9, 101916.9, 101900.4, 101877.8, 
    101848.3,
  101679.3, 101789.4, 101812.7, 101879, 101912.2, 101953.1, 101974.1, 
    101992.7, 101997.6, 101994.2, 101982.4, 101964.5, 101945.4, 101921.7, 
    101893.2,
  101831.5, 101900.5, 101937.3, 101984.7, 102013.4, 102042.9, 102058.4, 
    102068.2, 102063.9, 102051.7, 102034.7, 102010.2, 101987.1, 101964.1, 
    101936,
  101982.4, 102020.4, 102059.7, 102087.2, 102111.2, 102128.7, 102134.8, 
    102133.2, 102120.6, 102101.8, 102081.2, 102055.8, 102032.2, 102007.7, 
    101974.3,
  101446.6, 101437, 101483.5, 101525.2, 101543, 101540.5, 101561, 101571.6, 
    101579.2, 101587.2, 101599.7, 101609.2, 101623.7, 101649.4, 101666.8,
  101363.1, 101405.6, 101445.3, 101464.1, 101480.1, 101487.9, 101519.1, 
    101532.6, 101546, 101563.7, 101587.1, 101608.4, 101632.1, 101646.4, 
    101664.1,
  101372.1, 101395, 101421.9, 101451.1, 101442.3, 101466.4, 101488.1, 
    101509.6, 101536.4, 101568.8, 101595.4, 101617.1, 101646, 101666.1, 
    101687.1,
  101353.7, 101381.8, 101400.4, 101387.6, 101412.8, 101422.5, 101453.2, 
    101486.3, 101528.7, 101568.2, 101597.4, 101629.6, 101657.4, 101681.3, 
    101702.6,
  101359.7, 101328.5, 101335.9, 101348.7, 101379, 101402, 101451.4, 101494.4, 
    101536.2, 101573.4, 101614.4, 101652.1, 101684, 101708.9, 101722.9,
  101294.6, 101266.2, 101328.7, 101345.3, 101382.4, 101422.8, 101468.1, 
    101504.4, 101552.5, 101599.8, 101647.6, 101685.5, 101714.2, 101736.8, 
    101750.3,
  101295.1, 101324.7, 101344.7, 101375.3, 101417.5, 101455.1, 101501.7, 
    101552.1, 101605.8, 101652.9, 101693.4, 101727.8, 101753.1, 101769.8, 
    101780.7,
  101299.2, 101379.7, 101390.5, 101442.3, 101476, 101525.7, 101576.7, 
    101627.4, 101673.1, 101714, 101749.2, 101776.6, 101795.7, 101809.4, 
    101815.2,
  101411.3, 101486.6, 101496.8, 101548.3, 101573.3, 101627.7, 101664.7, 
    101710.2, 101743.5, 101777.6, 101803.6, 101826.8, 101840.3, 101847.3, 
    101841.3,
  101569.6, 101608.9, 101624, 101663.6, 101689.8, 101728.3, 101759.6, 
    101794.3, 101819.5, 101843.6, 101860.1, 101873.3, 101879.2, 101879.7, 
    101876.1,
  102103.3, 102092.2, 102087.5, 102088.6, 102087.8, 102085.5, 102081.9, 
    102069.7, 102055.7, 102035.4, 102009.1, 101982.2, 101944.5, 101899.9, 
    101856.2,
  101995.9, 101994.7, 101999.2, 102001.2, 102010.8, 102011.9, 102012.2, 
    102009.2, 101999.7, 101986.6, 101962.9, 101936.3, 101905.5, 101876.4, 
    101835.4,
  101913.7, 101913.4, 101917, 101921.6, 101933.9, 101942, 101950.5, 101953.9, 
    101948.7, 101937.3, 101920.9, 101900.3, 101874.8, 101847.5, 101813.7,
  101830.1, 101833, 101840.6, 101849.1, 101862.2, 101874.3, 101883.8, 
    101892.1, 101891.4, 101883.7, 101873.5, 101853.4, 101834.7, 101810.8, 
    101784.5,
  101766.3, 101758.8, 101769.5, 101782.2, 101794.1, 101807.9, 101819.3, 
    101829, 101831.9, 101832.1, 101824.9, 101811.1, 101796, 101779.4, 101763.6,
  101719.2, 101710.7, 101714.5, 101725.3, 101736.5, 101749.3, 101763.3, 
    101776.6, 101783.2, 101783.3, 101777.5, 101768.4, 101758.8, 101749.2, 
    101738.9,
  101655.6, 101652.9, 101656.2, 101667.7, 101680.1, 101695.1, 101713, 
    101724.1, 101729.7, 101732.2, 101730.8, 101726.3, 101721.2, 101719.4, 
    101722.4,
  101597.8, 101602.2, 101615.3, 101623, 101644.5, 101653, 101667.3, 101671.5, 
    101677.6, 101684.4, 101684.5, 101686, 101688.7, 101696.1, 101710.3,
  101542.3, 101557.8, 101574, 101584.1, 101597.5, 101601.6, 101615.9, 
    101621.7, 101629.9, 101636.6, 101645.3, 101653.8, 101666.3, 101685.2, 
    101712.1,
  101490.3, 101519.3, 101528.7, 101542.4, 101548.8, 101558.9, 101569.9, 
    101582.9, 101594.4, 101610.7, 101625.5, 101645, 101663.3, 101687.7, 
    101717.4,
  102361.7, 102402, 102412.1, 102407.4, 102396.8, 102381.2, 102359.4, 
    102333.5, 102303.1, 102270.5, 102234.9, 102196.8, 102156.9, 102114.5, 
    102065,
  102296, 102325.4, 102332.7, 102328.1, 102319.3, 102306.3, 102289.2, 102267, 
    102240.6, 102212.3, 102182.2, 102150.5, 102118.7, 102079.7, 102038.6,
  102228.8, 102246.6, 102256.4, 102249.1, 102239.1, 102227.6, 102211, 
    102192.2, 102171.1, 102148.3, 102124.9, 102099.6, 102070.5, 102038.2, 
    102003.8,
  102159.2, 102164.8, 102175.7, 102165.1, 102162.4, 102147.1, 102132.5, 
    102114.5, 102096.1, 102080.5, 102060, 102042.7, 102020, 101994, 101963.9,
  102087.9, 102087.2, 102098.1, 102087.7, 102083, 102068, 102051.8, 102038.2, 
    102020.8, 102009.4, 101994.7, 101982.9, 101961.2, 101946.9, 101919.3,
  102016.1, 102011.1, 102019.8, 102010.1, 102000.9, 101984.6, 101970.6, 
    101958.5, 101944.5, 101934.8, 101923.8, 101916, 101904.6, 101891.3, 
    101874.2,
  101936.5, 101945.8, 101949.1, 101946.5, 101932.6, 101918, 101899.3, 
    101885.1, 101869.2, 101864.9, 101855.5, 101848.8, 101841.3, 101836.1, 
    101821.7,
  101856.3, 101877, 101885, 101883.7, 101870.5, 101854.3, 101835.1, 101821.1, 
    101803.8, 101795.9, 101788.8, 101784.8, 101782.4, 101778.2, 101770.2,
  101806.9, 101821.8, 101826.6, 101825.2, 101821.9, 101805.8, 101787.1, 
    101765.5, 101750.9, 101738.4, 101728.2, 101722, 101718.9, 101717.9, 
    101710.7,
  101722.1, 101760.7, 101768.9, 101774, 101771.2, 101759.4, 101740.4, 
    101720.2, 101705.9, 101690.8, 101676.4, 101666.8, 101660.2, 101656.9, 
    101655.9,
  102197.2, 102191, 102186.1, 102174.8, 102166, 102152.8, 102140.3, 102125.8, 
    102109.4, 102091.2, 102074.6, 102055.1, 102032.2, 102000.8, 101963.8,
  102158.9, 102151.1, 102143.5, 102136.2, 102125, 102108.6, 102092.7, 
    102076.6, 102062.6, 102051.6, 102039.4, 102023.3, 102002.5, 101974, 
    101940.8,
  102109.4, 102113, 102100.4, 102085.6, 102067.6, 102055, 102045.9, 102037.5, 
    102029, 102017.5, 102003.5, 101986.3, 101965.4, 101943.1, 101914.8,
  102084.1, 102069.3, 102056.8, 102051, 102042.1, 102032.1, 102018.8, 
    102002.4, 101984.9, 101967, 101951.9, 101932.6, 101913.1, 101893.7, 
    101872.9,
  102040.5, 102045.3, 102050.8, 102050.4, 102034.6, 102016.4, 101990.6, 
    101969.8, 101945.7, 101926.3, 101906.7, 101890.5, 101871.3, 101853.8, 
    101832,
  102037, 102059.8, 102050.5, 102035, 102007.4, 101976.6, 101942.2, 101915.5, 
    101889.8, 101869.7, 101853.6, 101835.5, 101819.4, 101805, 101788.8,
  102041.5, 102058.1, 102035.7, 102001.8, 101962.3, 101921.4, 101876.7, 
    101840.5, 101809.7, 101792, 101777.5, 101768.6, 101760.5, 101749.6, 
    101740.5,
  102061.1, 102049.3, 102013.8, 101969.8, 101916, 101859.9, 101800.4, 
    101754.3, 101720.2, 101704.8, 101700.8, 101698.2, 101694.5, 101690, 
    101690.5,
  102047.7, 102020.2, 101983.1, 101924.2, 101847.1, 101774.3, 101701.1, 
    101642, 101599.2, 101582.9, 101591.8, 101609.7, 101623.4, 101625.3, 
    101629.4,
  102024.9, 102004.7, 101947.2, 101872.7, 101788.6, 101697.7, 101613.2, 
    101533.8, 101477.5, 101453.8, 101476.1, 101531.1, 101562.7, 101572.7, 
    101580.4,
  102103.1, 102131.8, 102136.6, 102130.8, 102112.4, 102093.6, 102064.3, 
    102026.8, 101990.5, 101952.5, 101914.6, 101876.6, 101853.1, 101829.4, 
    101808.8,
  102083.8, 102110.1, 102108, 102104.3, 102089.8, 102066.9, 102035.6, 
    101999.8, 101966.8, 101932, 101901.5, 101873.8, 101850.1, 101824.1, 
    101796.9,
  102073, 102094, 102097.4, 102088.3, 102047.8, 102019.1, 101989.9, 101958.3, 
    101933.9, 101909.7, 101882.1, 101857.5, 101831.9, 101812.6, 101788.5,
  102078.6, 102082.7, 102058.5, 102038.9, 102011.2, 101988.5, 101966, 
    101940.5, 101911.2, 101884, 101856.5, 101832.6, 101809.5, 101789.3, 
    101764.8,
  102057.4, 102058.4, 102039.8, 102027.3, 101998.2, 101962.2, 101926.4, 
    101892.6, 101857.4, 101829.3, 101809.1, 101790.5, 101775.3, 101759.6, 
    101749.9,
  102048.4, 102056.2, 102037.4, 102007.2, 101967, 101917.8, 101869.9, 
    101829.1, 101792.6, 101766.4, 101745.1, 101731.8, 101726.7, 101723.5, 
    101720.8,
  102059.8, 102051.1, 102023.8, 101973.2, 101919.8, 101859.9, 101803.5, 
    101753.6, 101705.8, 101674, 101657.4, 101651.8, 101655.4, 101666.8, 
    101676.6,
  102064.1, 102037.6, 101987.9, 101924.7, 101871.7, 101807.9, 101748.5, 
    101679.7, 101626.4, 101589.1, 101564.8, 101557.7, 101570.7, 101594.5, 
    101619.5,
  102055.9, 102019.2, 101966.7, 101904.3, 101842.5, 101774.5, 101695.7, 
    101614.7, 101564.3, 101516.5, 101476.8, 101458.9, 101474.4, 101518, 
    101558.9,
  102063.1, 102018.3, 101957.2, 101888.8, 101826.9, 101746.2, 101664.3, 
    101587.7, 101527.7, 101462.6, 101393.5, 101348, 101361.8, 101426.6, 
    101491.9,
  101915.7, 101919.3, 101947.5, 101960.9, 101977.3, 101995.7, 102010.5, 
    102016.3, 102021, 102011.6, 102005.7, 101990, 101967.5, 101944.4, 101910.5,
  101849.4, 101866.8, 101898.7, 101917.4, 101935.8, 101952.5, 101973.1, 
    101987.5, 101998.5, 101995.9, 101997.9, 101987.8, 101969.1, 101944.8, 
    101913.8,
  101805, 101834.4, 101865.3, 101890.2, 101915.1, 101934.1, 101952.1, 
    101969.5, 101978.8, 101981.5, 101985.1, 101974.2, 101957.2, 101938, 
    101912.8,
  101758.3, 101795, 101826.4, 101854.4, 101879.2, 101901.4, 101922.9, 
    101944.3, 101962.3, 101961, 101967.4, 101958.7, 101946.4, 101928.1, 
    101907.6,
  101722.9, 101762.4, 101793.4, 101828.2, 101855.7, 101879.2, 101900.9, 
    101918.6, 101929.2, 101936.4, 101932.6, 101928.4, 101912.5, 101899.6, 
    101885.1,
  101696, 101738.9, 101769.4, 101808.7, 101837.1, 101857.9, 101871.9, 
    101888.5, 101893, 101896.8, 101894.1, 101888.9, 101882.2, 101874.2, 
    101867.2,
  101686.9, 101726.7, 101755.7, 101786.5, 101799.5, 101818.2, 101831.5, 
    101845.7, 101848.3, 101853.4, 101849.3, 101844.7, 101842.9, 101842.3, 
    101841.7,
  101685.5, 101720, 101734.4, 101748.3, 101773.1, 101788.8, 101798.8, 101804, 
    101808.5, 101813.5, 101822.7, 101830.8, 101835.5, 101831, 101823.6,
  101679.4, 101703.6, 101711.1, 101721.8, 101740.2, 101741.3, 101756.6, 
    101764.8, 101779.6, 101790.3, 101795.5, 101806.7, 101811.8, 101812.5, 
    101816.1,
  101689.2, 101699.3, 101703.1, 101706, 101721.8, 101718.8, 101736, 101749.9, 
    101762.7, 101766.4, 101772, 101774.3, 101779.6, 101786.3, 101798.1,
  102060.6, 102087.8, 102136.2, 102172.9, 102208.5, 102228.8, 102233.7, 
    102225.9, 102220.2, 102208, 102196.4, 102178, 102165.5, 102146.1, 102121.7,
  101954, 102002.1, 102075.8, 102111.9, 102143.3, 102166.1, 102176.6, 
    102177.9, 102177.2, 102169.6, 102168, 102158.3, 102155.4, 102149.3, 
    102127.1,
  101873.1, 101932.2, 101990.8, 102034.5, 102077.7, 102107.4, 102130, 
    102137.6, 102147.7, 102148.2, 102153.5, 102150.7, 102151.7, 102144.6, 
    102127.9,
  101802.7, 101863.2, 101921.4, 101973.9, 102020.8, 102050.5, 102077.3, 
    102090, 102106.1, 102116.9, 102128.3, 102138, 102146.7, 102153.7, 102131.1,
  101730.4, 101785.5, 101848.8, 101906.5, 101952.4, 101985.3, 102020.3, 
    102044.6, 102066.7, 102092.3, 102107.8, 102120.8, 102128.4, 102134.5, 
    102119,
  101658.8, 101717.7, 101782, 101837.9, 101886.9, 101928.8, 101963.3, 
    102002.4, 102029, 102060.8, 102079, 102099.8, 102113.6, 102116.7, 102110.4,
  101594.4, 101657.7, 101719, 101777, 101830.5, 101875.6, 101912.5, 101961, 
    101995, 102033.1, 102057, 102077, 102088.2, 102096.4, 102099.9,
  101534.7, 101597.1, 101657.6, 101719, 101772.8, 101823.4, 101868.8, 
    101921.9, 101962.3, 102005.7, 102031.1, 102050.9, 102077.9, 102101.3, 
    102094.6,
  101483.5, 101547.1, 101602.5, 101669.6, 101726.9, 101777.9, 101829.3, 
    101886.3, 101932, 101978.4, 102005.8, 102041, 102074.4, 102096.1, 102103.9,
  101435.9, 101498.2, 101560.8, 101626.9, 101688, 101740.8, 101800.5, 101854, 
    101905.7, 101956, 101988.2, 102029, 102068.8, 102090.8, 102110.6,
  102405.3, 102437.1, 102482.1, 102509, 102525.7, 102531.8, 102535.5, 
    102511.7, 102489.5, 102458.9, 102410.5, 102366.7, 102293.3, 102225.9, 
    102167.7,
  102329.3, 102372.1, 102424, 102457.4, 102483.2, 102497.4, 102503.5, 
    102493.3, 102478.3, 102453.5, 102410.3, 102355.9, 102301, 102242.2, 
    102180.4,
  102259, 102315, 102369.9, 102411, 102446.3, 102466.9, 102480.7, 102476.5, 
    102470.3, 102448.6, 102412.1, 102361, 102309.5, 102247.7, 102188.4,
  102182.2, 102248.5, 102312.2, 102361.3, 102403.5, 102426, 102448.4, 
    102453.7, 102448.9, 102437.6, 102407.3, 102357.4, 102312.2, 102252.8, 
    102196.7,
  102104.9, 102178, 102249.5, 102307.5, 102354.9, 102385.4, 102416.4, 
    102428.4, 102429.4, 102421.2, 102396.1, 102364.6, 102312, 102250.4, 
    102199.1,
  102024.9, 102108.3, 102186.1, 102251.5, 102306.1, 102346.5, 102381, 
    102399.2, 102408, 102402.4, 102382.3, 102352.4, 102302.3, 102253.5, 
    102203.3,
  101950.8, 102040.9, 102122.6, 102194.6, 102253.5, 102304.5, 102340.5, 
    102369.4, 102381.4, 102385.4, 102371, 102341.2, 102300.3, 102249.9, 
    102199.9,
  101878.3, 101975.6, 102060.2, 102139.8, 102202.6, 102260.9, 102303.4, 
    102333.7, 102354.7, 102363, 102353.3, 102329.9, 102288.2, 102247.4, 
    102196.2,
  101812.1, 101914.1, 102001.5, 102083.9, 102152.5, 102217.1, 102264.2, 
    102299.5, 102323.1, 102338.2, 102331.1, 102317.1, 102277, 102236.8, 
    102193.4,
  101749.2, 101853.1, 101945.7, 102031.1, 102105.1, 102171.8, 102224.4, 
    102264.4, 102293.7, 102312, 102309.3, 102298, 102262.6, 102229.1, 102186.2,
  102588.3, 102608.5, 102612, 102614.4, 102597.5, 102573.7, 102553.1, 102491, 
    102445.3, 102406, 102346.6, 102284.7, 102221.1, 102147.3, 102066.5,
  102562.1, 102582.9, 102597.7, 102605.2, 102591.2, 102568.9, 102553.3, 
    102513, 102464.6, 102421.7, 102367, 102303.2, 102241, 102180.2, 102095.7,
  102544.6, 102567.9, 102586.9, 102594.3, 102591.8, 102584.6, 102558.7, 
    102523.4, 102479.3, 102438.9, 102390, 102326.5, 102252.8, 102194.3, 
    102112.5,
  102525.8, 102548.3, 102572.4, 102590.8, 102596, 102575.9, 102569.5, 
    102528.1, 102496.4, 102454.2, 102403.7, 102341.1, 102272.5, 102210.5, 
    102134.6,
  102498, 102530.4, 102552.6, 102582.1, 102595.7, 102581.4, 102571.3, 
    102540.3, 102512.8, 102466.7, 102417.1, 102360.4, 102294.3, 102220.7, 
    102147.4,
  102465.5, 102508.5, 102533.9, 102565, 102587.2, 102579.4, 102577.2, 
    102549.4, 102524.6, 102484.2, 102433.8, 102379.6, 102309.1, 102239.2, 
    102172.1,
  102433.6, 102483.4, 102514.5, 102541.3, 102570, 102574.3, 102574, 102552.5, 
    102519.1, 102495.2, 102445.5, 102402, 102319.5, 102262.2, 102186.5,
  102404.9, 102458.3, 102493.6, 102524.5, 102551.4, 102574.6, 102568.5, 
    102552, 102531.1, 102504, 102456.2, 102424, 102339.2, 102279.6, 102207.4,
  102378.6, 102433.1, 102472.7, 102507.1, 102537.3, 102564.7, 102567.5, 
    102556.6, 102528, 102515.3, 102466.1, 102435.5, 102356.3, 102297.9, 
    102222.3,
  102351.4, 102408.2, 102453.6, 102491.4, 102524.3, 102550.2, 102562.7, 
    102559.2, 102536.5, 102521.8, 102479, 102448.1, 102368.6, 102316.6, 
    102232.7,
  102746.1, 102729.1, 102700.1, 102669.4, 102621.4, 102581.7, 102529.9, 
    102461.4, 102399.2, 102334.5, 102269, 102205.8, 102131.8, 102039.4, 
    101972.5,
  102734.2, 102726, 102713.4, 102692.8, 102647.2, 102597.8, 102549.3, 
    102487.3, 102428.2, 102362.1, 102287.6, 102209.4, 102155.1, 102070.2, 
    101994.5,
  102733.2, 102736.1, 102722.6, 102708.9, 102669.5, 102620.8, 102573.8, 
    102505.7, 102449.4, 102384.6, 102315.5, 102243.9, 102180, 102080.8, 
    102003.9,
  102734.3, 102734.2, 102728.9, 102720.7, 102691.4, 102644.7, 102602.1, 
    102532.9, 102477.1, 102406.4, 102341.2, 102268.1, 102195, 102103.6, 
    102028.6,
  102741.9, 102740.3, 102736.9, 102727.5, 102711.7, 102664.3, 102625.5, 
    102558.2, 102498.2, 102429.4, 102373, 102301.1, 102213.3, 102128.1, 
    102054.3,
  102744.3, 102745, 102740.1, 102733.7, 102724.7, 102683.5, 102648.4, 
    102585.4, 102524.1, 102458.6, 102396.4, 102332.7, 102236.5, 102162, 
    102084.5,
  102742.5, 102749.7, 102744.4, 102740, 102738.2, 102705.1, 102665.5, 
    102607.4, 102549, 102485.4, 102422.8, 102357, 102266.9, 102196.7, 102116.2,
  102743.3, 102750.7, 102751.3, 102741.6, 102740.4, 102720.7, 102690.3, 
    102634.6, 102580.5, 102516.1, 102451.4, 102391.6, 102296.9, 102235.4, 
    102151.8,
  102746.8, 102752.9, 102765, 102742.3, 102749.5, 102735.3, 102715.8, 102665, 
    102612.5, 102548, 102486.9, 102423.2, 102332.4, 102276.6, 102191.8,
  102745.6, 102751.3, 102766.9, 102749.6, 102751.6, 102750.6, 102739.6, 
    102699, 102648.6, 102583.4, 102521.2, 102461.8, 102371.6, 102316.5, 
    102233.9,
  102921.4, 102851.8, 102798.5, 102737, 102664.2, 102594.6, 102521.9, 102448, 
    102385.2, 102333.1, 102252.2, 102173.6, 102108.4, 102074.2, 102037.1,
  102926.2, 102880.7, 102838, 102776.7, 102696, 102622, 102546.2, 102467.6, 
    102386.6, 102308.6, 102239.5, 102195, 102142.8, 102085.5, 102045.6,
  102937.6, 102905, 102861.4, 102805.1, 102730.7, 102644.4, 102567.6, 
    102483.3, 102403, 102316.7, 102262.5, 102198.3, 102142.6, 102109.8, 
    102083.1,
  102945.7, 102922.4, 102887.5, 102833.5, 102767.9, 102681.7, 102603.6, 
    102513.5, 102424.8, 102318.2, 102253.8, 102200.3, 102162.1, 102139.1, 
    102110.2,
  102962.9, 102941.2, 102906.6, 102861.5, 102797.2, 102719.9, 102644.3, 
    102561.3, 102471, 102361, 102288, 102227.9, 102195.5, 102171.9, 102144.8,
  102980.8, 102960.8, 102924.9, 102891.5, 102831.9, 102768.1, 102692.6, 
    102622.3, 102533.7, 102419.4, 102321.4, 102259, 102234.5, 102208.3, 
    102183.8,
  103001.7, 102982.7, 102940.9, 102915.6, 102869.6, 102808.8, 102743.4, 
    102678, 102623.4, 102548.5, 102428.5, 102326.2, 102279.1, 102257.1, 
    102228.1,
  103023.7, 103001.1, 102960.7, 102935.2, 102904.5, 102853.3, 102803.7, 
    102726.2, 102673.1, 102601, 102481.8, 102399.4, 102333.6, 102302.9, 
    102276.5,
  103041.6, 103017, 102990.1, 102954, 102930.3, 102889, 102844.7, 102787.8, 
    102722.5, 102656.4, 102548.3, 102473.6, 102394.4, 102367.3, 102327.9,
  103056.2, 103030.9, 103009.8, 102972.2, 102946, 102921.5, 102876.5, 
    102823.1, 102768.1, 102697.7, 102599, 102536, 102464.7, 102421, 102375.5,
  102964.7, 102883.2, 102810.8, 102729.3, 102643.2, 102566, 102487.7, 
    102404.7, 102325.7, 102266.5, 102225, 102197.4, 102157.2, 102103, 102086,
  102957.5, 102898.9, 102849.5, 102772, 102683.5, 102595.4, 102504.1, 102406, 
    102316.1, 102262.3, 102235.7, 102203.4, 102169.2, 102129.9, 102106.7,
  102973.5, 102915.8, 102860, 102789.9, 102721.5, 102632.9, 102543.1, 102439, 
    102315.9, 102224.1, 102214.8, 102196.6, 102176.6, 102152.1, 102141.9,
  102979.1, 102932, 102892.3, 102821.7, 102758.2, 102668.9, 102576.1, 
    102462.7, 102316.3, 102190.5, 102200, 102204.7, 102188.1, 102194.9, 
    102173.7,
  103014, 102953.7, 102911.9, 102854.9, 102787.2, 102713.1, 102628.4, 
    102526.6, 102351.2, 102205.3, 102195, 102208.7, 102214.1, 102220, 102204.4,
  103034, 102986.8, 102937.8, 102884.7, 102819, 102751.9, 102674, 102604.8, 
    102451.3, 102286.4, 102218.8, 102249.4, 102255.3, 102255.4, 102234.8,
  103069.9, 103017.5, 102958.8, 102916.1, 102860.3, 102797, 102717.2, 
    102661.3, 102592.4, 102458.8, 102349.3, 102306.7, 102297.8, 102289, 
    102270.9,
  103112.7, 103051.4, 102993.8, 102936.4, 102887.5, 102821.3, 102769.2, 
    102681.9, 102657.7, 102536.8, 102448.7, 102364.1, 102343.4, 102330.6, 
    102307.3,
  103133, 103069.1, 103020.6, 102963.4, 102914, 102846.7, 102799, 102720.6, 
    102697.4, 102624.9, 102518.7, 102429.6, 102386.4, 102367.3, 102341.1,
  103149, 103090.4, 103043.2, 102983.6, 102930.7, 102871.8, 102821.5, 
    102749.7, 102705.9, 102674.8, 102587.2, 102499.9, 102432.8, 102401.7, 
    102371.6,
  102927.9, 102863.4, 102802, 102737.4, 102651.8, 102568, 102477.5, 102379.1, 
    102280.5, 102177.6, 102100.7, 102064.9, 102031.9, 101993.1, 101989.1,
  102964.5, 102902, 102836.6, 102774.4, 102690.3, 102600.8, 102507.4, 
    102401.5, 102292.8, 102174.6, 102100.9, 102057.2, 102040, 102004.2, 
    102001.9,
  103007.7, 102941.5, 102871.2, 102801.1, 102720.8, 102630.4, 102533.6, 
    102421.3, 102310.5, 102179.5, 102077.5, 102039.9, 102021.6, 102009.6, 
    102032.4,
  103044.5, 102978.8, 102906.2, 102834.6, 102756.7, 102666.2, 102570.7, 
    102454.8, 102335, 102190, 102070.3, 102024.2, 102026.2, 102022.6, 102037.1,
  103082.3, 103009.9, 102935.7, 102861.3, 102783.4, 102698.3, 102604.9, 
    102495.9, 102379.1, 102232.2, 102094.3, 102025, 102019.2, 102041.2, 
    102041.9,
  103107.6, 103033.6, 102962.9, 102887.7, 102813.2, 102730, 102640.5, 
    102542.8, 102439.5, 102293.6, 102152.4, 102068.6, 102052, 102062.6, 102058,
  103120.8, 103053.1, 102979.2, 102905.3, 102834.1, 102752.4, 102673.6, 
    102576.6, 102492.7, 102394.7, 102271.6, 102168.8, 102111.9, 102094.2, 
    102078.8,
  103119.5, 103054.2, 102986.6, 102914.6, 102848.9, 102771.8, 102697, 
    102609.4, 102535.3, 102444.7, 102355.1, 102274.6, 102194.5, 102139.3, 
    102107,
  103110.8, 103044.2, 102976.1, 102912, 102847.9, 102778.8, 102709.6, 
    102632.5, 102555.4, 102495.4, 102410.5, 102340.1, 102260.5, 102183.9, 
    102135.8,
  103089.5, 103020.2, 102955.6, 102893.5, 102833.1, 102772.4, 102707.7, 
    102642.6, 102570.1, 102506, 102445.7, 102377.4, 102310.4, 102227.9, 
    102167.1,
  102845.4, 102786.8, 102736.2, 102668.9, 102601.9, 102529, 102450.6, 
    102361.3, 102262.7, 102145.7, 102036.2, 101960.5, 101926.4, 101900.9, 
    101883,
  102894.1, 102836.6, 102782, 102719.3, 102652.3, 102580.6, 102504.7, 
    102422.6, 102335, 102234.6, 102120.9, 101999.9, 101923, 101908.5, 101892.3,
  102929.7, 102869.9, 102811, 102749.1, 102682.8, 102614.2, 102542.5, 
    102462.4, 102373.6, 102275.1, 102166, 102069.7, 101973.3, 101928.2, 
    101914.4,
  102955.4, 102903.4, 102842.3, 102784.1, 102718.1, 102650.1, 102581.4, 
    102507.4, 102426.3, 102340.1, 102231.5, 102133.7, 102028.5, 101955.4, 
    101934,
  102975.7, 102917.6, 102861, 102796.4, 102736.7, 102671.1, 102605.7, 
    102534.4, 102457.4, 102378.7, 102284.9, 102188.1, 102093.8, 102006.7, 
    101966,
  102982.1, 102922.5, 102866.8, 102804.5, 102749.5, 102688.6, 102624.5, 
    102559.9, 102489.9, 102417, 102331.2, 102242.4, 102157.5, 102064.9, 
    102009.9,
  102973.5, 102917.7, 102859.5, 102797.1, 102742, 102687.7, 102626.7, 
    102564.4, 102499.2, 102439.5, 102358.6, 102285, 102209.1, 102121.9, 
    102051.3,
  102960.8, 102903.6, 102842.2, 102779.8, 102726.7, 102673.2, 102617.7, 
    102563.2, 102503.1, 102445.7, 102376.8, 102309.7, 102242.9, 102172.3, 
    102100.9,
  102933, 102874, 102812.8, 102755.4, 102698.2, 102642.8, 102590.4, 102537.6, 
    102487.1, 102434.1, 102379.3, 102317, 102256.7, 102201.7, 102135,
  102893.8, 102832.5, 102774.4, 102715.3, 102658.9, 102602, 102549, 102498.3, 
    102455.6, 102408.1, 102357.7, 102311, 102254.6, 102208.9, 102155.2,
  102675.6, 102644.5, 102624.7, 102596.1, 102551, 102506.6, 102458.4, 
    102407.5, 102339.7, 102254.4, 102166.2, 102084, 102022.5, 101968.2, 
    101929.9,
  102708.4, 102687.1, 102655.3, 102631.6, 102596.6, 102548.5, 102504, 
    102449.2, 102390.3, 102325.2, 102244, 102175.9, 102092.8, 102003.8, 
    101950.6,
  102726.2, 102705.5, 102674.8, 102646.1, 102617.7, 102571.9, 102530.2, 
    102478.1, 102423.5, 102362.6, 102285.7, 102205.9, 102148.9, 102090.8, 
    102002.8,
  102745.2, 102721.2, 102694.7, 102669.3, 102632.1, 102591.8, 102549.8, 
    102499.8, 102448.5, 102400.6, 102335.7, 102265.3, 102192.8, 102131.3, 
    102052.1,
  102755.1, 102729.5, 102700.6, 102674.1, 102638.1, 102599.5, 102563.9, 
    102516, 102461, 102416.4, 102363.9, 102304.3, 102239, 102163.5, 102102.1,
  102758.3, 102730, 102696.1, 102666, 102636.2, 102601.3, 102560.1, 102519.5, 
    102473.1, 102424.2, 102379.5, 102328.7, 102275, 102212.8, 102144.7,
  102747, 102710.7, 102688.6, 102651.8, 102619.7, 102580.3, 102544.8, 
    102508.7, 102469.7, 102423.3, 102378.8, 102338.8, 102291.8, 102235.8, 
    102178.4,
  102716.4, 102688, 102660.9, 102627.2, 102595.2, 102556.5, 102521.3, 
    102486.1, 102450.8, 102413.7, 102372.8, 102331.8, 102297.8, 102250.6, 
    102201.9,
  102670.9, 102639.9, 102615, 102584.4, 102551.5, 102515.2, 102485.6, 
    102449.8, 102419.2, 102387.4, 102349.2, 102318, 102286.5, 102246.6, 102207,
  102611.7, 102579.7, 102552, 102520.5, 102489.5, 102458.2, 102427.1, 
    102400.6, 102374.4, 102347.5, 102319.2, 102291.7, 102264.7, 102229.7, 
    102193.7,
  102722.3, 102731.9, 102748.2, 102750.1, 102741.3, 102723, 102687.2, 
    102650.1, 102610.5, 102553.5, 102495.2, 102423.7, 102357.3, 102288.7, 
    102222.9,
  102764.1, 102773.5, 102787.7, 102783.9, 102767.3, 102749.2, 102720.8, 
    102678.1, 102639.8, 102592.7, 102538.2, 102477.9, 102414.6, 102344.7, 
    102274.2,
  102783.6, 102789.6, 102805.8, 102799, 102793.1, 102773.4, 102745.8, 
    102709.9, 102671.6, 102623.6, 102575.2, 102522.5, 102450.5, 102400.9, 
    102321.2,
  102808.3, 102824.5, 102840.6, 102832.3, 102815.3, 102793.8, 102764.5, 
    102730.9, 102697.6, 102645.2, 102601.3, 102556.6, 102501.1, 102437.4, 
    102374.2,
  102829.8, 102836.1, 102837.3, 102835.5, 102821.3, 102800.8, 102778, 
    102740.8, 102709, 102664.4, 102617, 102572.2, 102527.5, 102476.3, 102410.9,
  102837.4, 102837.1, 102839.6, 102834.4, 102810, 102799.3, 102773.6, 
    102739.7, 102704.6, 102671.1, 102633.8, 102583.1, 102539.6, 102495.1, 
    102443.9,
  102825.7, 102823.4, 102824.3, 102819.6, 102805.9, 102791.1, 102757.5, 
    102734.6, 102689, 102660.4, 102623.4, 102581.5, 102538.8, 102503.2, 
    102455.3,
  102805.1, 102799.9, 102796.3, 102788.6, 102779.5, 102754.9, 102737.6, 
    102709.1, 102673.2, 102637, 102606.1, 102571.2, 102529.9, 102494.1, 
    102456.2,
  102770.2, 102759.6, 102762.7, 102752.7, 102736.9, 102713.9, 102693.3, 
    102668.8, 102644.4, 102612.6, 102582.1, 102551.4, 102516.7, 102478.3, 
    102444.6,
  102717, 102712.6, 102714.7, 102706.9, 102693.5, 102675.3, 102655.4, 
    102633.2, 102610.2, 102580.7, 102553.6, 102526.4, 102492.1, 102461.1, 
    102428.9,
  102866.9, 102921.5, 102940.9, 102964.7, 102976.6, 102976.2, 102947.2, 
    102913, 102867.2, 102805.8, 102754, 102695.3, 102644.2, 102571.2, 102515.8,
  102854.4, 102917.2, 102956.9, 102993.2, 103001.5, 102999.5, 102971.5, 
    102935.5, 102894.3, 102836.4, 102782, 102725.7, 102672.6, 102606.4, 
    102546.5,
  102847.2, 102912.7, 102956.3, 103000.4, 103003.4, 103017.2, 102989.4, 
    102954, 102913.2, 102857.2, 102802.9, 102744, 102688.1, 102629.8, 102568.9,
  102839.3, 102905.7, 102961.6, 103013.5, 103027.5, 103020.4, 103014.1, 
    102969.9, 102929.4, 102876.1, 102816.9, 102756, 102697.7, 102645.1, 
    102585.6,
  102833.2, 102904, 102959.6, 103006.9, 103028.3, 103019.2, 103020.3, 
    102977.6, 102941.4, 102880.8, 102825.2, 102760.9, 102703.4, 102648.2, 
    102594.4,
  102831, 102898.8, 102960.5, 103000.4, 103023, 103024.2, 103018, 102981.8, 
    102943.9, 102891.6, 102833.9, 102771, 102708, 102653.9, 102598,
  102839, 102897.6, 102957, 102992.7, 103013.5, 103014.1, 103003.5, 102979.6, 
    102942.3, 102888.4, 102832.5, 102772.9, 102713.5, 102656.7, 102603.5,
  102848, 102900.1, 102951.5, 102978.4, 103000.3, 102997.5, 102988, 102965.7, 
    102933.9, 102886.8, 102828.5, 102774.7, 102715.1, 102658.5, 102606,
  102862.9, 102910.7, 102946.4, 102961.8, 102980.2, 102979.5, 102966.1, 
    102954.2, 102920.2, 102879.5, 102827.6, 102773.4, 102715.4, 102662.4, 
    102609.2,
  102870.3, 102908.3, 102939.8, 102951.5, 102953.4, 102955, 102946.9, 
    102928.9, 102902.8, 102865.2, 102816.3, 102766.2, 102712.9, 102662.8, 
    102609.9,
  102752.6, 102775.3, 102808.4, 102826.2, 102850.9, 102851.7, 102829.5, 
    102780.9, 102738.1, 102678.5, 102616.5, 102554.9, 102490.4, 102430.1, 
    102370.9,
  102718.6, 102748.2, 102794.8, 102839.1, 102857.8, 102852, 102842.4, 
    102815.6, 102770.6, 102720.6, 102653.7, 102588.4, 102519.4, 102457.2, 
    102394.9,
  102700.8, 102725.7, 102775.1, 102818.5, 102854.1, 102848, 102848.4, 
    102831.9, 102786.9, 102742, 102678.3, 102613.4, 102538.7, 102475.6, 
    102414.4,
  102690, 102695.8, 102751.2, 102793, 102842.6, 102843.3, 102849.6, 102841.6, 
    102802.8, 102763.5, 102700.1, 102636.4, 102560.2, 102498.5, 102435.6,
  102667.5, 102672.8, 102723.8, 102766.6, 102818.9, 102833.5, 102843.7, 
    102844.4, 102808.5, 102775.1, 102714.8, 102654.2, 102578.7, 102513.6, 
    102453.6,
  102637, 102649.3, 102694.4, 102737.1, 102792.5, 102825.4, 102843.9, 
    102841.4, 102811, 102784.7, 102729, 102673.6, 102596.2, 102532.4, 102471.1,
  102603.4, 102619.9, 102661.9, 102705.4, 102764.2, 102805.7, 102839, 
    102832.6, 102812.1, 102784.8, 102738.4, 102680.4, 102608.1, 102545.1, 
    102484.8,
  102565.2, 102591.8, 102629, 102675.8, 102734.2, 102781.9, 102814, 102822.4, 
    102801.8, 102783.7, 102739.6, 102685.8, 102618.2, 102555.6, 102496,
  102525.4, 102560.5, 102604.2, 102646.5, 102704.7, 102758.7, 102793.2, 
    102807.7, 102804.2, 102781.2, 102738, 102689, 102624.4, 102562, 102506.1,
  102493.8, 102539.5, 102582.6, 102628.1, 102677.5, 102735.4, 102772.5, 
    102789.2, 102784.2, 102772.3, 102726.7, 102687.8, 102627.9, 102565.7, 
    102513.2,
  102483, 102534.3, 102574.4, 102610.7, 102634.6, 102657.5, 102642.2, 
    102610.5, 102583, 102541.6, 102489.4, 102407.8, 102347.4, 102295, 102237.4,
  102445.2, 102501.4, 102551, 102586.1, 102617.1, 102637.7, 102640.4, 
    102625.9, 102604.2, 102568.7, 102511.9, 102449.2, 102380.5, 102324.1, 
    102264.6,
  102408.7, 102472.2, 102524.8, 102561.8, 102598.3, 102622.4, 102639.1, 
    102630.7, 102612.1, 102583.2, 102527.4, 102467.3, 102400.6, 102343.7, 
    102287,
  102374.8, 102435.3, 102489.6, 102529.3, 102573.4, 102600.9, 102612.6, 
    102632.8, 102612.6, 102590.4, 102546, 102496.6, 102426.6, 102367.2, 
    102309.6,
  102346.5, 102405.1, 102454.2, 102498.9, 102539, 102579.2, 102605.1, 
    102625.4, 102612.5, 102590.1, 102558.6, 102513.2, 102446.2, 102383.5, 
    102330.2,
  102326.3, 102382.8, 102425.7, 102464.3, 102504.3, 102554, 102586.8, 
    102609.5, 102610.3, 102599.7, 102566, 102525.2, 102469.1, 102402.9, 
    102347.6,
  102308.8, 102360.4, 102409.5, 102435.1, 102469.9, 102515.6, 102564.6, 
    102599.9, 102605.1, 102603.4, 102568.8, 102534.7, 102482.1, 102417.2, 
    102362.6,
  102301.9, 102342.9, 102388.8, 102414.2, 102440.1, 102479.1, 102532.9, 
    102574.8, 102589.2, 102598.2, 102572.3, 102543.7, 102491.4, 102429.7, 
    102374.8,
  102295.6, 102328.3, 102373.2, 102403.2, 102419.7, 102439.9, 102490.2, 
    102542, 102570.7, 102588, 102573.3, 102544.2, 102499.6, 102440.9, 102384.7,
  102272.2, 102301.8, 102340.6, 102378.1, 102402.3, 102415.7, 102448.1, 
    102500.8, 102544.8, 102567.2, 102571.4, 102544.5, 102508.9, 102450.7, 
    102394.3,
  102366, 102385.7, 102404.6, 102418.3, 102460.8, 102498.9, 102519.7, 
    102511.9, 102500.7, 102469.7, 102424.1, 102363.2, 102307.5, 102263.6, 
    102213.9,
  102312.6, 102341.4, 102376.9, 102397.3, 102436.7, 102479.9, 102506.1, 
    102514.5, 102509, 102475.7, 102448.3, 102401.4, 102336.2, 102287.4, 
    102237.8,
  102256.6, 102290.7, 102339.8, 102369.4, 102403.3, 102449.2, 102488.9, 
    102506.1, 102507.7, 102486.4, 102458.3, 102419.7, 102352, 102303.7, 
    102255.5,
  102191, 102230.4, 102287.4, 102331.7, 102372.7, 102415.9, 102462, 102488.3, 
    102500, 102492.8, 102464.4, 102430.8, 102370.5, 102322.8, 102275.2,
  102116.3, 102167, 102230, 102288, 102336.5, 102379.2, 102434.2, 102468.1, 
    102491.9, 102491.8, 102476.8, 102440.5, 102381.8, 102336.3, 102292.8,
  102046.7, 102103.8, 102170.7, 102231.5, 102296.4, 102342, 102400.7, 
    102448.7, 102477.7, 102493.8, 102470.6, 102446.9, 102395.8, 102351.4, 
    102310,
  101992.5, 102048.2, 102111.4, 102179.4, 102248.9, 102303.9, 102363.5, 
    102418.3, 102459.9, 102491, 102472, 102455.7, 102406.4, 102364.2, 102324.5,
  101954.5, 102001.9, 102062.2, 102127.3, 102201.6, 102262.8, 102324.6, 
    102382.7, 102428.6, 102462.8, 102474, 102458.1, 102415.7, 102376.3, 
    102338.5,
  101923.2, 101971.9, 102023.5, 102084.5, 102157.4, 102222.2, 102281.7, 
    102346.4, 102396.1, 102445.1, 102458.5, 102466.8, 102429.4, 102387.1, 
    102352,
  101915.8, 101953.3, 101992.5, 102052.2, 102116.6, 102183.7, 102241.6, 
    102306.5, 102363.3, 102419.4, 102435.9, 102467.7, 102439.9, 102401.2, 
    102363.3,
  102230.4, 102272.8, 102302.6, 102322.4, 102373.7, 102419.5, 102432.8, 
    102455.6, 102465.4, 102440.9, 102409.6, 102362.2, 102318.9, 102286, 
    102246.4,
  102219.1, 102269.7, 102314.6, 102332.5, 102351.2, 102402.1, 102434.1, 
    102445.4, 102455.5, 102447.9, 102437.9, 102390.6, 102340.8, 102306.5, 
    102266.6,
  102210.1, 102261.3, 102303.3, 102344.3, 102351.8, 102376.1, 102413.2, 
    102443, 102456.6, 102449.8, 102442, 102403.7, 102357.2, 102318.6, 102283.4,
  102201.4, 102242.9, 102286.6, 102326.7, 102353.3, 102358.9, 102391.6, 
    102430.4, 102448.2, 102464.9, 102447, 102410.6, 102369.9, 102336.2, 
    102301.1,
  102182.9, 102225.8, 102260.5, 102302.8, 102335.3, 102354.3, 102366.1, 
    102406.8, 102436.3, 102454.9, 102461.8, 102426.3, 102378.3, 102347.4, 
    102315.4,
  102158.9, 102196.9, 102232.2, 102268.4, 102305.7, 102336.5, 102354.8, 
    102377.1, 102411.6, 102434.8, 102448.7, 102429.3, 102394, 102362, 102331,
  102125.4, 102160, 102195.2, 102226.8, 102265.8, 102302.6, 102330.1, 
    102354.8, 102379.9, 102415, 102436.3, 102432.7, 102406.7, 102374, 102343.8,
  102090.6, 102117, 102149.4, 102179.8, 102214.7, 102255.8, 102290.7, 
    102322.7, 102349.6, 102386.7, 102418.9, 102423.3, 102418.9, 102381.4, 
    102356.8,
  102060.1, 102080.2, 102100, 102129.3, 102165.3, 102202.5, 102245.6, 
    102282.8, 102315.8, 102352.7, 102392.9, 102411.5, 102411.8, 102386.6, 
    102367.3,
  102027.1, 102038.3, 102052.5, 102078.6, 102108.1, 102147.9, 102192.2, 
    102238.4, 102279, 102319.2, 102357.7, 102389.9, 102403, 102390.3, 102372.1,
  101755.9, 101860.1, 101974.7, 102077.5, 102167.7, 102236.3, 102289.8, 
    102330.7, 102350.4, 102343.8, 102319.2, 102290.8, 102270.6, 102239.2, 
    102210.5,
  101714.4, 101830.8, 101948.3, 102054.1, 102148.8, 102226.7, 102280.9, 
    102318.8, 102344.6, 102348, 102341.3, 102306.4, 102288, 102262.5, 102235.9,
  101692.9, 101813.9, 101930.1, 102039.2, 102129.8, 102211.3, 102267, 
    102315.4, 102340.4, 102356.5, 102346.2, 102321.2, 102300.3, 102278.7, 
    102252.3,
  101671.4, 101795.5, 101914.1, 102020.8, 102111.1, 102190.5, 102251.7, 
    102305, 102336.8, 102354.4, 102361, 102335.8, 102315.3, 102297.1, 102272.2,
  101653.7, 101778.5, 101900.5, 102003.3, 102092.3, 102167, 102234.1, 
    102289.4, 102335.6, 102354.5, 102369.5, 102359.8, 102330.4, 102313.7, 
    102291.3,
  101639, 101767.3, 101887.9, 101988.7, 102079.3, 102150.4, 102218.1, 
    102279.2, 102326.1, 102353.7, 102380.1, 102367.9, 102355.6, 102329.1, 
    102310.1,
  101631.8, 101760.5, 101878.3, 101977.8, 102068.1, 102140, 102206.9, 102265, 
    102313.5, 102348, 102379.7, 102379.3, 102383.8, 102344.9, 102326.4,
  101625.1, 101756.5, 101869.1, 101967.5, 102057.2, 102133.4, 102204.6, 
    102260.1, 102301, 102332.1, 102362.6, 102372.3, 102371.4, 102356.4, 
    102338.8,
  101624.6, 101754.5, 101860.5, 101956.9, 102045.8, 102122.3, 102187.8, 
    102247.1, 102291.7, 102319.2, 102343.4, 102359.8, 102371.3, 102370.1, 
    102347.3,
  101627.1, 101752.3, 101855.1, 101946.8, 102030.6, 102105, 102168.2, 
    102226.7, 102272.6, 102307.2, 102326.4, 102341, 102362.1, 102365.6, 
    102347.3,
  101624.3, 101655, 101723, 101824, 101921.6, 102006.6, 102081.6, 102141.7, 
    102180.8, 102203.7, 102206.1, 102202.9, 102191.5, 102168.5, 102141.7,
  101605.7, 101637.8, 101688.6, 101785.5, 101889.2, 101981, 102063, 102133.4, 
    102181.5, 102203, 102214.2, 102215.3, 102208.8, 102192.7, 102171.1,
  101594.3, 101631.6, 101667.7, 101753.8, 101864.5, 101960.6, 102048.4, 
    102127.4, 102179.2, 102204.2, 102220.4, 102225.9, 102222, 102211.9, 
    102193.4,
  101586.9, 101624.2, 101656, 101723.8, 101834.7, 101937.2, 102030.8, 
    102114.1, 102171.2, 102204.3, 102220.4, 102234.9, 102234.3, 102231.1, 
    102214.9,
  101567.4, 101614.8, 101648.9, 101698.5, 101805.3, 101911.6, 102010.4, 
    102098.3, 102161.1, 102206.2, 102222.7, 102236.6, 102245.4, 102245.1, 
    102234,
  101550.7, 101603, 101643.1, 101677.3, 101773.9, 101886, 101989, 102082.4, 
    102146.3, 102199, 102224.7, 102236.7, 102253.4, 102258.3, 102254.2,
  101534.5, 101588, 101633.7, 101667.2, 101746.1, 101860.2, 101965.3, 102063, 
    102131.1, 102190.5, 102227.2, 102243, 102270.7, 102269.3, 102269.2,
  101513.1, 101570.8, 101620.9, 101660.7, 101720.8, 101835.5, 101940.5, 
    102041.8, 102112.6, 102179.9, 102226.9, 102247.9, 102275.5, 102278.8, 
    102279.6,
  101491.8, 101550.6, 101606, 101648.1, 101703.7, 101811, 101917.5, 102022.5, 
    102097.1, 102166.9, 102220.1, 102249.7, 102277.7, 102299.1, 102292.5,
  101471.8, 101527.6, 101591, 101631.8, 101693.7, 101788, 101897.4, 102002.4, 
    102083.3, 102155.6, 102213.2, 102250.6, 102283.2, 102300.1, 102299.5,
  101571.4, 101691.3, 101808.9, 101916, 102014.9, 102097.6, 102154.9, 102207, 
    102242.8, 102261, 102266.4, 102264.1, 102250.1, 102228.8, 102194.2,
  101531.3, 101654.6, 101773.4, 101883.9, 101986, 102076.5, 102142.4, 
    102200.5, 102241.6, 102262.7, 102273.1, 102280, 102269.6, 102254.4, 
    102226.4,
  101497.9, 101625.3, 101744.4, 101861.4, 101964.1, 102059.2, 102130.6, 
    102191.2, 102239.6, 102266.7, 102281.4, 102291.4, 102286.7, 102275.7, 
    102251.3,
  101467.7, 101598, 101717.4, 101835.4, 101940.8, 102037.6, 102116.5, 
    102179.8, 102234.7, 102266.2, 102283.4, 102298.7, 102302.7, 102295, 
    102275.5,
  101442, 101572.9, 101690.4, 101810.5, 101919.9, 102015.3, 102101.5, 102168, 
    102225.1, 102266.1, 102288.9, 102303.2, 102313.4, 102308.7, 102294.4,
  101418.7, 101552.4, 101668, 101783.4, 101895.9, 101995.8, 102083.3, 
    102157.9, 102217, 102261.8, 102287.8, 102304.8, 102314.6, 102316.9, 
    102310.2,
  101402.2, 101532.5, 101651.3, 101758.3, 101871.3, 101972, 102064.1, 
    102144.1, 102204.8, 102254.7, 102287.7, 102303.7, 102316.3, 102324.9, 
    102322.8,
  101392.7, 101517.5, 101637.5, 101738.6, 101846.6, 101950.3, 102044, 
    102127.5, 102191, 102244.9, 102281.8, 102307.4, 102315.4, 102322.5, 
    102322.1,
  101388.5, 101506.6, 101626, 101728.1, 101821.3, 101925.9, 102021.2, 
    102107.7, 102176.2, 102233.4, 102274.3, 102302.9, 102313.3, 102321.8, 
    102329.2,
  101389.2, 101501.6, 101616.8, 101717.7, 101803.5, 101901, 101996.7, 
    102085.5, 102158.9, 102219.9, 102263.8, 102294, 102306.8, 102320, 102332.8,
  101967.2, 102051.9, 102129.8, 102208.2, 102280, 102343, 102377.8, 102406.2, 
    102429.5, 102429, 102420.3, 102402.1, 102374, 102337.4, 102294.4,
  101923.3, 102017.2, 102104.4, 102186.2, 102262, 102330, 102372.9, 102406.1, 
    102431.8, 102436.7, 102436.7, 102419.1, 102392.8, 102359.9, 102319.8,
  101893.2, 101997.1, 102088.2, 102173.3, 102252, 102322.8, 102371.2, 
    102406.6, 102437.3, 102445.6, 102448.1, 102437, 102411.6, 102380.1, 
    102341.2,
  101867.8, 101973.6, 102069.1, 102155.8, 102236.4, 102311.1, 102367.7, 
    102404.4, 102438, 102454.4, 102454.9, 102451.6, 102427.5, 102397.7, 
    102361.2,
  101844.3, 101950.7, 102050.1, 102139.8, 102224, 102300.4, 102364.4, 
    102401.4, 102435.4, 102457, 102460.5, 102456.4, 102437.6, 102410.2, 
    102377.4,
  101821.4, 101925.1, 102030.9, 102121.8, 102208.9, 102288.8, 102356, 
    102403.7, 102433.5, 102456.7, 102467.4, 102463.4, 102448, 102420.8, 
    102389.9,
  101797.5, 101902.5, 102010.9, 102104, 102194.2, 102274.7, 102346.4, 
    102401.5, 102431.1, 102454.7, 102466.1, 102468.3, 102453, 102426.9, 
    102396.3,
  101774.3, 101880.3, 101991.7, 102086.9, 102178.7, 102260.9, 102334.6, 
    102393.2, 102429.2, 102461, 102469.3, 102471.8, 102459.2, 102435.2, 
    102399.8,
  101752.7, 101861.6, 101973.9, 102069.2, 102164.6, 102247.2, 102322.9, 
    102384, 102425, 102452.1, 102470.9, 102470.3, 102466.2, 102437.9, 102403.7,
  101732.7, 101843.6, 101956.9, 102053.5, 102149.3, 102232.9, 102309.4, 
    102372.5, 102417.6, 102446.5, 102461.4, 102469.5, 102464.2, 102439.2, 
    102406,
  102562.3, 102550.3, 102549.4, 102541.7, 102547.8, 102566.2, 102581.2, 
    102575.2, 102566.1, 102537, 102499.5, 102454.1, 102401, 102343.1, 102283.5,
  102524.6, 102527.4, 102537.7, 102534.5, 102539.7, 102561.4, 102575.1, 
    102576.7, 102567.4, 102544.1, 102510.2, 102469.6, 102417.1, 102360.8, 
    102300.7,
  102495.2, 102514.8, 102533.3, 102532.8, 102538.6, 102556.8, 102573.3, 
    102583.2, 102574.7, 102556.4, 102522.5, 102483.5, 102429.1, 102374.2, 
    102311.6,
  102467.3, 102489.3, 102514.5, 102523.2, 102531.9, 102552.7, 102566.8, 
    102584.9, 102577, 102562.8, 102533.1, 102492.7, 102441.5, 102387.1, 
    102325.8,
  102436.5, 102461.6, 102493, 102515.8, 102527, 102547.9, 102567.5, 102577.9, 
    102576.4, 102566.9, 102545.9, 102502.1, 102453.2, 102396.7, 102336,
  102407.9, 102432, 102465, 102495.9, 102516.6, 102537, 102562.1, 102579.7, 
    102586.2, 102574.4, 102552.9, 102509.5, 102462.3, 102407, 102346.9,
  102376.8, 102404, 102438.6, 102472.1, 102502.4, 102525.3, 102553.3, 
    102575.4, 102580.8, 102572.1, 102546.2, 102513.4, 102469.5, 102413.9, 
    102355.2,
  102344, 102371.8, 102412.1, 102447.6, 102485, 102511.7, 102541.9, 102566.8, 
    102576.4, 102571, 102558.9, 102520.5, 102475.1, 102421.4, 102362.2,
  102307.6, 102341.9, 102385.1, 102424.2, 102466, 102497.5, 102529.8, 
    102556.5, 102569.9, 102566.1, 102548.1, 102515.7, 102473.8, 102424.4, 
    102367.1,
  102269.3, 102310.3, 102355.2, 102398.1, 102444.7, 102481.2, 102515.4, 
    102541.4, 102558.4, 102557.6, 102536.4, 102512.5, 102472.9, 102424, 
    102368.6,
  102811, 102799.4, 102760.3, 102709.9, 102678.5, 102626, 102586.2, 102556.5, 
    102521.7, 102472, 102421.4, 102357.3, 102294.3, 102223.1, 102149.6,
  102826.8, 102819.6, 102786.4, 102740.4, 102705.6, 102647.1, 102594, 
    102571.6, 102537.5, 102486, 102440.4, 102378.4, 102316, 102246.2, 102173.4,
  102839.1, 102830.3, 102803, 102760.6, 102714.1, 102665.2, 102602.1, 
    102571.3, 102544.5, 102501.9, 102454.9, 102392.9, 102330.3, 102262.6, 
    102189.7,
  102834.9, 102831, 102816.8, 102784.8, 102734.3, 102690.1, 102625.6, 
    102583.9, 102551.2, 102513.9, 102468.3, 102409.6, 102345.7, 102278.8, 
    102206.3,
  102852.6, 102842.6, 102823.1, 102804.6, 102752.1, 102707.6, 102650.4, 
    102601.8, 102561.2, 102526.8, 102478.1, 102420.6, 102355.6, 102289.7, 
    102218.3,
  102844.3, 102844.9, 102833.6, 102810.4, 102770.1, 102723.2, 102673.7, 
    102625.1, 102580.1, 102538.1, 102487.3, 102430, 102366.3, 102300, 102228.3,
  102835.9, 102844, 102836.6, 102814.2, 102780.3, 102734.1, 102689.4, 
    102635.4, 102587.6, 102543.9, 102493.1, 102436.6, 102372.7, 102305.3, 
    102234.9,
  102817.8, 102830.1, 102830, 102814.4, 102777, 102743, 102694.9, 102645.4, 
    102592.7, 102548.4, 102497.2, 102440.5, 102378.2, 102310.9, 102240.2,
  102801.8, 102817.6, 102820.7, 102806, 102775.5, 102739.9, 102697.4, 
    102646.8, 102597.8, 102549, 102497.4, 102440.4, 102381.1, 102314.2, 
    102242.8,
  102773, 102796.4, 102800.8, 102791.1, 102763.7, 102729.1, 102691.1, 102641, 
    102593.4, 102542, 102492.8, 102438.9, 102379.4, 102312.5, 102244.4,
  102484.2, 102510, 102511.7, 102495.1, 102473.4, 102441.3, 102413.7, 
    102383.5, 102347.4, 102295.5, 102239.8, 102177.4, 102112.1, 102042.2, 
    101973.6,
  102497.5, 102523.8, 102536.8, 102526.8, 102507, 102484.4, 102446.3, 
    102397.8, 102362.1, 102317.2, 102263, 102198.9, 102134.2, 102066.3, 
    101997.7,
  102510.9, 102542.7, 102555.6, 102553.9, 102530.4, 102509.2, 102484.6, 
    102437.7, 102390.8, 102339.8, 102279.8, 102216.8, 102153.4, 102083.4, 
    102016.2,
  102524.5, 102558, 102578.6, 102580.3, 102570.1, 102542.9, 102514.7, 102465, 
    102413.6, 102360.9, 102298, 102234.9, 102169.5, 102101.4, 102035.4,
  102539.2, 102573.3, 102594.7, 102602.6, 102586.4, 102568.6, 102532.1, 
    102487, 102436.8, 102378.8, 102312.9, 102246.4, 102180, 102113.6, 102048.7,
  102556.1, 102595.5, 102618.4, 102621.3, 102612.6, 102584.9, 102546.7, 
    102501.8, 102447.6, 102391.5, 102324.2, 102256.4, 102190.3, 102124.4, 
    102061.3,
  102570.6, 102611.9, 102629.6, 102633.1, 102626.1, 102601.5, 102564.8, 
    102519, 102458.5, 102399.6, 102330.9, 102263.6, 102195.7, 102130.9, 
    102067.2,
  102586.3, 102630.6, 102651, 102652.5, 102638.8, 102610.8, 102573.5, 
    102533.6, 102472.3, 102407.6, 102339.1, 102269.8, 102202.7, 102136.6, 
    102074.2,
  102603.4, 102647.6, 102669.3, 102665.6, 102651.1, 102623.5, 102588.4, 
    102541.6, 102486.7, 102419.1, 102346.6, 102275.2, 102209.5, 102141.1, 
    102077.8,
  102616, 102661.6, 102686.7, 102684, 102662.3, 102636.2, 102600.2, 102552.1, 
    102497.5, 102430.7, 102354.7, 102285.1, 102214.7, 102148.3, 102081.9,
  102187.1, 102242.9, 102271, 102292.6, 102316.9, 102323, 102306.2, 102276.8, 
    102242.8, 102196.4, 102140.6, 102089.4, 102033.7, 101975.9, 101919.8,
  102183.1, 102246.5, 102286.2, 102314.2, 102334.4, 102331.5, 102320.2, 
    102296.9, 102264.9, 102210.8, 102148.9, 102096.7, 102045.9, 101992.2, 
    101933.9,
  102192.3, 102260.2, 102300.8, 102340.9, 102360.3, 102362, 102344, 102306.6, 
    102263.9, 102217.8, 102163.6, 102112.5, 102060.3, 102003.1, 101945,
  102207.9, 102277.4, 102325.5, 102372, 102386.2, 102379.1, 102355.3, 102325, 
    102282.2, 102242, 102175.8, 102126.7, 102073.6, 102017.1, 101957.9,
  102225.7, 102298, 102356.4, 102395.5, 102399.1, 102394.1, 102377.3, 
    102338.8, 102299.6, 102254.2, 102194.1, 102142.9, 102086.1, 102030.9, 
    101970.1,
  102247.9, 102324.4, 102380.4, 102408.3, 102418.1, 102413.6, 102393.7, 
    102360.3, 102315.9, 102271.8, 102211.4, 102161.3, 102102.1, 102047.1, 
    101984.8,
  102276.4, 102349.4, 102397.5, 102427.2, 102440.1, 102437.5, 102415.6, 
    102381.9, 102335.3, 102289.7, 102233.5, 102179.6, 102116.5, 102060, 101996,
  102301.7, 102368.7, 102416.1, 102447.3, 102457.5, 102452.1, 102435, 
    102404.4, 102358.6, 102309.3, 102256.2, 102198.2, 102132.9, 102074.7, 
    102010,
  102328, 102388.2, 102435.4, 102462, 102473.5, 102475.4, 102454, 102423.8, 
    102381, 102329.6, 102274.4, 102212.9, 102147.7, 102088.2, 102022.9,
  102348.4, 102405.4, 102453.4, 102481.5, 102494.6, 102488.9, 102471.2, 
    102438.1, 102398.3, 102343.1, 102290.1, 102228.2, 102161.2, 102102.6, 
    102037.7,
  102457.1, 102430.2, 102426, 102388.9, 102377.3, 102404.2, 102394.2, 102352, 
    102318, 102277.5, 102227.1, 102184, 102130, 102080.2, 102028.4,
  102425.8, 102403.1, 102399.4, 102376.2, 102387.9, 102394.5, 102401, 102372, 
    102329, 102286.6, 102238.6, 102194.1, 102144.4, 102096.8, 102043.5,
  102390.5, 102385.3, 102390.2, 102376.7, 102410, 102420, 102424.9, 102372.7, 
    102338.5, 102297.5, 102251.2, 102204, 102153.1, 102105.4, 102055.9,
  102361.1, 102365.5, 102376.6, 102388, 102428.3, 102429.6, 102424, 102378.3, 
    102349.6, 102313.5, 102266.9, 102217.7, 102167, 102120.4, 102072.1,
  102331.8, 102346.9, 102371, 102404.4, 102429.9, 102448.1, 102428.3, 
    102401.7, 102367, 102325.2, 102277.8, 102232.2, 102179.9, 102133.8, 
    102089.3,
  102309.5, 102337, 102373.8, 102410.4, 102430.5, 102442.8, 102437.3, 
    102418.5, 102382, 102339.7, 102294.6, 102246.1, 102195, 102148, 102099.1,
  102294.8, 102335.6, 102377.4, 102416.8, 102443.7, 102455.6, 102449.8, 
    102432.1, 102396, 102355.2, 102309.2, 102262.1, 102207.5, 102160.1, 
    102109.8,
  102283.1, 102337.9, 102382, 102425.5, 102458.9, 102469.5, 102465, 102445.1, 
    102413.1, 102367.6, 102321.2, 102277, 102224.3, 102175.2, 102126.3,
  102280.4, 102346.3, 102393.9, 102444.8, 102467.3, 102481.7, 102469.3, 
    102458.3, 102422.8, 102375.1, 102328.1, 102283, 102230, 102183.1, 102135.9,
  102284.1, 102355.3, 102404.4, 102452.9, 102477.1, 102488.7, 102487, 
    102464.7, 102434.7, 102380.8, 102332, 102285.8, 102234.5, 102187.3, 
    102140.6,
  102852.9, 102802.8, 102743.5, 102693, 102609.3, 102536, 102516.3, 102472.9, 
    102421.8, 102378.9, 102333.5, 102279.6, 102232, 102185, 102145.5,
  102839, 102799.9, 102742.3, 102689.4, 102610.9, 102543.6, 102522, 102490.1, 
    102449, 102400.9, 102346.6, 102294, 102246.9, 102200.4, 102157.3,
  102825.7, 102791.5, 102732.3, 102685.3, 102618.2, 102557.7, 102540.7, 
    102498.8, 102460.2, 102415.2, 102361.2, 102307, 102262.6, 102215.1, 
    102171.5,
  102815, 102776.8, 102732.5, 102681.2, 102620, 102561.9, 102541.4, 102509.8, 
    102482.1, 102433.4, 102376, 102323.8, 102276.7, 102229.4, 102181.3,
  102795.5, 102759.2, 102727.8, 102675.3, 102622.9, 102570.7, 102542.6, 
    102523.2, 102489.5, 102449.1, 102386.2, 102337, 102285.1, 102237.7, 
    102190.1,
  102766.2, 102737.6, 102708.2, 102660, 102613.8, 102557.4, 102551.1, 
    102531.9, 102504.2, 102459.8, 102395.2, 102344.3, 102286.6, 102238.6, 
    102194.7,
  102738.4, 102712.3, 102687, 102644.5, 102602.7, 102556.5, 102557, 102534.7, 
    102507, 102458.9, 102395, 102343.1, 102291.9, 102241.8, 102197.1,
  102704, 102687.5, 102664.7, 102622.6, 102587.6, 102561.1, 102555.7, 
    102542.7, 102512.9, 102458.1, 102392.5, 102339.8, 102287.1, 102239.4, 
    102194.5,
  102661.4, 102658.1, 102634.8, 102609, 102574.7, 102554.3, 102544.8, 102546, 
    102503.7, 102449.3, 102387.8, 102329.3, 102278, 102231.3, 102189.1,
  102618.8, 102620.3, 102603.6, 102586.5, 102561.9, 102555, 102552.3, 
    102541.9, 102504.2, 102444.8, 102382.7, 102324.2, 102268.7, 102217.6, 
    102176.8,
  102764.2, 102714.6, 102657.6, 102602.1, 102535.6, 102448.5, 102412.2, 
    102388.4, 102359.6, 102310.9, 102268, 102228.7, 102187.7, 102148.5, 
    102115.8,
  102800.9, 102746.4, 102686.9, 102632.4, 102563.8, 102480.8, 102429.8, 
    102400.1, 102379.6, 102321.5, 102270.8, 102225.6, 102190.5, 102155.7, 
    102122.4,
  102828.5, 102768.2, 102714.8, 102655.2, 102582.9, 102505.3, 102445.9, 
    102416.8, 102388.2, 102328.7, 102279.4, 102230.4, 102190.8, 102152.6, 
    102122.7,
  102862.3, 102796.2, 102743.6, 102683.4, 102604.5, 102526.3, 102466.6, 
    102433.6, 102399.5, 102341.5, 102283.2, 102230.6, 102189, 102151, 102121,
  102888.3, 102825.1, 102766.5, 102707.2, 102634.4, 102545.8, 102486.7, 
    102452, 102413.6, 102353.4, 102292.4, 102235.3, 102191.4, 102148, 102112.7,
  102916.3, 102848, 102793.3, 102725.8, 102664.9, 102570.9, 102508.2, 
    102470.2, 102429.2, 102365.6, 102303.7, 102243.6, 102193.2, 102148.2, 
    102110.5,
  102936.1, 102868.1, 102817.1, 102746, 102689.8, 102599.7, 102528, 102487.1, 
    102443, 102381, 102317.3, 102256.7, 102201.2, 102150.9, 102108.4,
  102948.5, 102883.7, 102836, 102765.5, 102717.8, 102624.7, 102551, 102503.9, 
    102455.5, 102394.9, 102335.3, 102274.2, 102214.4, 102158.7, 102112.4,
  102951.6, 102894.8, 102847.6, 102782.9, 102731, 102644.5, 102571.7, 
    102519.6, 102474.6, 102413.4, 102352.4, 102292.4, 102229.1, 102167.7, 
    102118.2,
  102946.8, 102899.8, 102853.5, 102792.3, 102739.5, 102658.3, 102586.3, 
    102531.9, 102483.3, 102424.5, 102368.5, 102308.1, 102246.1, 102180.7, 
    102128.2,
  101650.9, 101661.9, 101711, 101750.1, 101795, 101845.5, 101882.1, 101910.2, 
    101931.8, 101928.8, 101922.4, 101924, 101925.7, 101919.5, 101905,
  101653.3, 101685.9, 101735.2, 101767.1, 101807.9, 101851.2, 101893.5, 
    101909.7, 101910, 101910.4, 101916.8, 101919.4, 101917, 101910.5, 101895.9,
  101703.1, 101746.4, 101775.6, 101806.8, 101838.8, 101870.3, 101891.7, 
    101905.9, 101910.6, 101914.1, 101915.9, 101915.8, 101913, 101902.4, 
    101889.1,
  101774.7, 101815.7, 101830, 101853.2, 101868.9, 101883, 101903.8, 101909.4, 
    101916.9, 101920.4, 101917.5, 101916.3, 101910.9, 101899.6, 101883.1,
  101877, 101891.6, 101896.7, 101904.7, 101908.3, 101920.9, 101933.7, 
    101940.9, 101941.1, 101939.5, 101931.4, 101922.1, 101911.4, 101899.2, 
    101883.3,
  101990.4, 101975.2, 101972.3, 101968.2, 101966.3, 101965.1, 101971.1, 
    101977.2, 101973.1, 101965.1, 101953.7, 101938.2, 101923.7, 101908.8, 
    101886.5,
  102101.8, 102073, 102053.7, 102036.5, 102026, 102019.1, 102015, 102009.4, 
    102003.8, 101997, 101979.2, 101963, 101941.4, 101918.1, 101896.9,
  102213.2, 102172.7, 102145.7, 102118.8, 102096.9, 102079.6, 102066.3, 
    102052.4, 102041.1, 102025.5, 102007.3, 101980.3, 101960.6, 101934.4, 
    101910.2,
  102317.7, 102271, 102234.5, 102198.6, 102169.2, 102143, 102125.1, 102103, 
    102082.4, 102061.3, 102040.9, 102012.1, 101980.6, 101949.9, 101917.9,
  102411.1, 102366.4, 102320.6, 102283.3, 102249.7, 102207, 102181.9, 
    102151.6, 102124.8, 102098.7, 102072.4, 102038.3, 102001.2, 101962, 
    101926.8,
  101326.8, 101368.8, 101441.2, 101499.8, 101551.3, 101580.8, 101601.9, 
    101624, 101656.7, 101693.2, 101742.3, 101790.9, 101822.2, 101836.1, 101844,
  101210.9, 101273.9, 101373.1, 101433.8, 101495.7, 101539.6, 101569.6, 
    101596.1, 101634.3, 101674.2, 101725.8, 101772.4, 101809.6, 101830.2, 
    101837.4,
  101143.9, 101214.9, 101303.2, 101365.6, 101448, 101504.3, 101547.6, 101584, 
    101626, 101663.7, 101715.8, 101762.9, 101799, 101819.3, 101826.7,
  101046, 101141.3, 101230.6, 101320.9, 101408.4, 101470.4, 101524.6, 
    101566.5, 101607.6, 101654, 101705.7, 101751.5, 101785.8, 101815.2, 
    101818.9,
  100946.4, 101062.7, 101167.9, 101276.5, 101364.5, 101437.5, 101504, 
    101552.7, 101597.3, 101651, 101702.9, 101744.5, 101776.1, 101806.3, 
    101808.6,
  100859.2, 100997.9, 101115.9, 101232.4, 101330.7, 101415.4, 101489.2, 
    101543.6, 101593.4, 101649, 101700, 101741.8, 101774.3, 101799.2, 101805.8,
  100808.2, 100948.8, 101076.3, 101205.9, 101309.8, 101403.8, 101481.2, 
    101541, 101598.6, 101657.5, 101704, 101745, 101776.4, 101796.5, 101807.8,
  100819.6, 100937, 101065.7, 101195.6, 101309.1, 101401.5, 101484, 101549.6, 
    101610.8, 101669.6, 101714.9, 101757.9, 101787.2, 101810.9, 101830.7,
  100870.7, 100965.6, 101089.9, 101213.3, 101325.5, 101419.1, 101502.3, 
    101570.4, 101635.6, 101690.1, 101736.4, 101774.8, 101803.3, 101828.1, 
    101832.5,
  100961.7, 101046, 101152.5, 101264.7, 101363.2, 101455.7, 101537.2, 
    101603.5, 101670.3, 101718.1, 101764, 101791.5, 101815.4, 101824.7, 
    101830.3,
  102567.7, 102545.8, 102532.2, 102499.1, 102458.9, 102426.5, 102385.7, 
    102336.8, 102284.9, 102218.8, 102159.5, 102099, 102041.5, 102042.3, 
    102046.2,
  102511.8, 102494.2, 102498.1, 102471, 102449.2, 102414.9, 102381.7, 
    102338.4, 102289.1, 102226.5, 102164.4, 102108.4, 102053.3, 102040.3, 
    102042,
  102427.6, 102422.7, 102443.2, 102431, 102418.7, 102390.5, 102364.4, 
    102326.1, 102282, 102232.3, 102169.8, 102119.2, 102063.8, 102054.6, 
    102059.4,
  102313.7, 102330.2, 102367.7, 102375.7, 102378.6, 102360.1, 102340.8, 
    102314.2, 102277.2, 102231.2, 102171.4, 102122.8, 102072.1, 102063.5, 
    102056,
  102177.9, 102215.6, 102270.4, 102301.4, 102319.6, 102315.6, 102305.9, 
    102289.9, 102262.4, 102223, 102170.3, 102128.4, 102082.4, 102074.1, 
    102062.1,
  102014.7, 102074, 102157.2, 102206.9, 102248, 102260.8, 102266.1, 102258.8, 
    102241.3, 102210.2, 102164.6, 102127.4, 102087, 102073.4, 102066.5,
  101829, 101915, 102021.4, 102099.2, 102159, 102191.9, 102213, 102218.6, 
    102212.7, 102188.5, 102153.1, 102125.4, 102093.4, 102078.3, 102068.3,
  101623.7, 101741.6, 101870.8, 101974.3, 102058, 102112.6, 102150.8, 
    102171.7, 102174.9, 102160.5, 102136.1, 102116, 102090.2, 102076.5, 
    102081.7,
  101430.1, 101565.3, 101715.2, 101841.9, 101947.5, 102026.3, 102082.4, 
    102118.7, 102134.3, 102130.8, 102115.3, 102108.8, 102085.6, 102093.4, 
    102086.2,
  101265.9, 101409.9, 101568.7, 101709.4, 101836.7, 101935.9, 102010.8, 
    102063, 102087.1, 102100.3, 102092.2, 102095.6, 102083.3, 102088.6, 
    102079.6,
  103253.5, 103205.2, 103153.5, 103096.9, 103036.3, 102968.8, 102899.4, 
    102833.8, 102751.6, 102687.8, 102604.5, 102523.4, 102412.2, 102328.9, 
    102261.1,
  103248.7, 103204, 103154.4, 103103.2, 103048.1, 102984.6, 102918.4, 
    102855.3, 102778.3, 102715.6, 102630.8, 102558.8, 102464.9, 102369.6, 
    102284.1,
  103221.5, 103180.1, 103134.4, 103087.8, 103035.9, 102978.5, 102915.6, 
    102855.7, 102780.7, 102726.4, 102648.7, 102576.2, 102485.7, 102395.7, 
    102309.2,
  103188.4, 103150, 103110.7, 103066.7, 103021.2, 102972, 102914.1, 102857.6, 
    102786.3, 102733.8, 102661.7, 102591.8, 102509.9, 102423.4, 102333.1,
  103144.1, 103107, 103070.2, 103028.7, 102989, 102948.3, 102895.6, 102844.5, 
    102780.5, 102726.7, 102663.8, 102598.6, 102519.6, 102441.5, 102352.5,
  103084.9, 103052.7, 103021.9, 102984.8, 102949.4, 102913.6, 102871.9, 
    102827.5, 102767, 102714.2, 102654.3, 102596.8, 102525.1, 102453.7, 
    102366.3,
  103017.5, 102983.3, 102959, 102924.1, 102894.5, 102863.2, 102831.9, 
    102794.2, 102743.1, 102692.9, 102637.8, 102588.4, 102521.9, 102456.8, 
    102376,
  102931.5, 102902.3, 102885.4, 102855.5, 102830.7, 102804.4, 102781.3, 
    102749, 102713.9, 102666, 102616.2, 102569.2, 102512.6, 102456.3, 102377.8,
  102832.4, 102809.3, 102798.9, 102771.9, 102754.5, 102731.8, 102716.9, 
    102693.1, 102669.1, 102629, 102586.6, 102545, 102499.9, 102445.6, 102372,
  102719.1, 102702.5, 102695.9, 102676.6, 102665.7, 102647.7, 102641.6, 
    102627.7, 102616.4, 102585.2, 102550.4, 102512.5, 102477.8, 102428.1, 
    102363.1,
  103240, 103203.9, 103148.8, 103097.7, 103036.1, 102969.6, 102902.8, 
    102835.7, 102761.6, 102688.2, 102606.3, 102525.6, 102452, 102375.5, 
    102305.7,
  103258.5, 103224.2, 103172.7, 103120.7, 103061.4, 102997, 102931.4, 
    102864.8, 102789.4, 102718.7, 102637.2, 102559.3, 102477.8, 102402.7, 
    102329.4,
  103257, 103226.8, 103179.5, 103130.4, 103071.7, 103010.8, 102946.4, 
    102881.3, 102808.9, 102738.1, 102657.5, 102581.4, 102498.9, 102422.1, 
    102346.4,
  103252.6, 103229.3, 103188.3, 103140.4, 103083.2, 103023.9, 102963.1, 
    102897.4, 102824.9, 102756.7, 102681.1, 102602.7, 102521.7, 102440.6, 
    102364.6,
  103236.2, 103219.5, 103182.1, 103140.3, 103082.4, 103027.4, 102969.2, 
    102907, 102835.9, 102769, 102692.3, 102615.4, 102536.7, 102458.5, 102381.8,
  103220, 103205, 103175.1, 103135, 103084.8, 103029.3, 102975.5, 102911, 
    102842.2, 102775.3, 102701.5, 102626.3, 102547.7, 102471.8, 102396.2,
  103190.1, 103179.3, 103157.4, 103119.8, 103070.4, 103021.6, 102970, 
    102908.3, 102843.2, 102776.7, 102702.9, 102633.2, 102555.8, 102482.3, 
    102407.5,
  103148.8, 103144.2, 103125.7, 103096, 103052.4, 103008.3, 102959.8, 
    102904.1, 102840.5, 102776.4, 102701.4, 102630.9, 102555.7, 102486.4, 
    102412.6,
  103100.1, 103097.3, 103085, 103059.9, 103026.8, 102983.6, 102940.8, 
    102890.2, 102833.4, 102769.7, 102696, 102625.2, 102553.7, 102483.3, 
    102411.7,
  103043.3, 103047.2, 103038.1, 103019.5, 102988.9, 102951.2, 102913.8, 
    102870.6, 102817.9, 102754.7, 102684.9, 102614.2, 102545.2, 102475, 
    102408.9,
  103059, 103058.5, 103020.2, 102979.1, 102932.2, 102875.5, 102817.2, 
    102754.4, 102689.9, 102622.6, 102545.5, 102471.4, 102401.8, 102329.7, 
    102261.8,
  103059.5, 103073.5, 103041.8, 103006.6, 102966.4, 102907.3, 102856, 
    102790.4, 102728.1, 102664.6, 102588, 102511.5, 102436.8, 102363, 102290,
  103061.5, 103057.5, 103046.6, 103019.5, 102988.5, 102934, 102883.8, 
    102821.8, 102755.3, 102692.3, 102614.7, 102540.2, 102464.2, 102389.9, 
    102315.2,
  103048.7, 103052.9, 103055.8, 103032.4, 103001.9, 102959.3, 102911.7, 
    102852.9, 102790, 102724.7, 102648.3, 102573.5, 102496.1, 102418.6, 
    102344.8,
  103022.6, 103039.1, 103052, 103037.3, 103005.1, 102974.4, 102929.8, 
    102873.8, 102813.7, 102750.5, 102672, 102597.9, 102525, 102444.1, 102368.4,
  102984.1, 103016, 103033.4, 103031.9, 103013.1, 102980.7, 102943.4, 
    102892.4, 102835.9, 102775.6, 102700.2, 102624, 102549.7, 102471.9, 102394,
  102943.7, 102983.8, 103007.6, 103015.6, 103004.8, 102975.6, 102945.2, 
    102899.9, 102850.2, 102791.6, 102721, 102642.5, 102571.6, 102494.4, 
    102416.5,
  102892.1, 102938.8, 102972, 102987.5, 102988.9, 102970.7, 102945.3, 
    102902.7, 102856.2, 102806.3, 102738, 102659.9, 102589.5, 102517.7, 
    102437.5,
  102833.6, 102888.5, 102930.8, 102953, 102965.6, 102955.1, 102930.4, 
    102894.8, 102861.3, 102805.6, 102749.9, 102670.4, 102600.4, 102532.1, 
    102454.9,
  102764.5, 102828.8, 102879.4, 102910.1, 102927.2, 102930.5, 102910.7, 
    102887.8, 102855.9, 102802.5, 102752.4, 102682.3, 102610.1, 102543.5, 
    102473.6,
  103049.6, 103034, 103020.2, 102995.4, 102943.9, 102904.1, 102852.8, 
    102797.9, 102737.7, 102665.9, 102592.7, 102521.5, 102448.5, 102375.4, 
    102306,
  103069.4, 103063.1, 103057.1, 103025.1, 102977.5, 102933, 102889.5, 
    102835.1, 102780, 102717.5, 102640.7, 102564.8, 102491.9, 102415.9, 
    102344.8,
  103076.7, 103074.8, 103085.9, 103048.8, 103012.9, 102962.9, 102920.9, 
    102868.5, 102811.9, 102751.3, 102681.2, 102604.7, 102529, 102455.4, 
    102378.3,
  103073.4, 103086.7, 103101.1, 103086.9, 103044.4, 102989.4, 102949.4, 
    102898.4, 102843.3, 102785.4, 102718.4, 102645.2, 102567.6, 102492.2, 
    102418.1,
  103062.4, 103078.8, 103096.8, 103093.7, 103071.7, 103016.4, 102974.4, 
    102924.1, 102870.3, 102815.4, 102747.1, 102681.1, 102604.9, 102524.6, 
    102449,
  103039.2, 103069.6, 103085.5, 103092.1, 103078.6, 103038.3, 102997.2, 
    102946.2, 102895.4, 102839.9, 102775, 102711.1, 102639.4, 102560.4, 
    102481.3,
  103010.8, 103050, 103066.9, 103079.4, 103071.2, 103043.4, 103007.4, 
    102963.4, 102914.9, 102858.2, 102798.8, 102737.3, 102665.8, 102589.6, 
    102509,
  102981.1, 103015.4, 103041.3, 103057.9, 103056, 103045.1, 103017.7, 
    102975.8, 102929.4, 102874.9, 102815.5, 102758, 102689.7, 102617.6, 
    102538.2,
  102940, 102980.1, 103007, 103024.8, 103031.8, 103031, 103008.5, 102975.2, 
    102937.6, 102883.4, 102825.8, 102772.1, 102709.5, 102637.2, 102561.2,
  102887.4, 102933.6, 102970.4, 102990.9, 103001.2, 103005.1, 102993.6, 
    102968, 102933, 102884.4, 102834, 102780.5, 102723.9, 102655.3, 102582.9,
  103267.1, 103255.9, 103243.1, 103209.6, 103165.5, 103118.1, 103069.6, 
    103005.9, 102944.5, 102874.3, 102798.9, 102724.1, 102642.1, 102564.2, 
    102487.2,
  103277.5, 103279.8, 103276.2, 103245, 103203.7, 103150.8, 103107.2, 
    103044.2, 102983.7, 102914.7, 102840.9, 102766.7, 102689.7, 102608.8, 
    102526.4,
  103283.1, 103291.6, 103295.4, 103279.2, 103236.3, 103188.2, 103138.7, 
    103081.1, 103018.6, 102947.7, 102871.6, 102799.5, 102723.2, 102646.7, 
    102562.5,
  103279.1, 103295.3, 103308.6, 103288.7, 103258.9, 103215.9, 103169.1, 
    103108.1, 103049.9, 102982.9, 102904.6, 102830.7, 102761.3, 102684.1, 
    102599.2,
  103271.7, 103289.6, 103299.3, 103291.5, 103261, 103229.5, 103183.1, 
    103131.3, 103068.2, 103010.8, 102931.7, 102854.2, 102789.1, 102713.6, 
    102630.7,
  103262.8, 103281.5, 103289.5, 103287.1, 103269, 103234.3, 103194.1, 
    103140.4, 103082.5, 103025.2, 102953.4, 102878.9, 102812.6, 102741.2, 
    102659.1,
  103243.3, 103263.7, 103273.2, 103271.1, 103252.2, 103223.6, 103190.6, 
    103138.6, 103089.4, 103039.4, 102971.4, 102894.6, 102828.5, 102760.8, 
    102681.4,
  103214.8, 103241.5, 103251.6, 103252.1, 103238.7, 103212.1, 103178.6, 
    103135.7, 103085.9, 103039, 102980.3, 102902.4, 102842.1, 102772.9, 
    102696.7,
  103182.6, 103210.6, 103223.2, 103225.5, 103213.4, 103190.7, 103163.7, 
    103120.2, 103082, 103034, 102978.3, 102905.8, 102844.6, 102778, 102708.7,
  103144.7, 103173.5, 103189.8, 103191.7, 103184, 103164.2, 103137.7, 
    103105.1, 103068.1, 103019, 102965, 102900.3, 102840.5, 102777.5, 102712.5,
  103473.6, 103433.7, 103385.6, 103328.1, 103259, 103189, 103115.2, 103039, 
    102950.6, 102865.9, 102781.9, 102704.8, 102626.6, 102538.8, 102451.7,
  103485.1, 103446.1, 103400.9, 103348.4, 103283.1, 103214.5, 103143.4, 
    103070, 102986.2, 102902.5, 102810.8, 102729.1, 102650.3, 102569.6, 
    102483.5,
  103485.2, 103453.3, 103410.1, 103361.9, 103297.2, 103229.3, 103160, 
    103088.3, 103009.2, 102925.6, 102835.2, 102751.6, 102669.4, 102587.6, 
    102504.7,
  103479.4, 103452, 103409.2, 103364.8, 103305.9, 103241.8, 103175.3, 
    103105.1, 103027.1, 102946.9, 102858.9, 102770.8, 102688, 102608.4, 
    102525.4,
  103463.8, 103440.9, 103409.1, 103363.8, 103308.7, 103244.2, 103180, 103112, 
    103036, 102961.3, 102876.6, 102787.4, 102702.9, 102621.9, 102538.3,
  103437.9, 103424.9, 103397.9, 103355.5, 103302.9, 103244.1, 103182.1, 
    103113.4, 103040.3, 102968.9, 102887.1, 102795.4, 102714.9, 102633.9, 
    102548.6,
  103411.4, 103402.1, 103378.3, 103341, 103292.9, 103236.8, 103176.4, 
    103108.5, 103041.3, 102969.6, 102891.2, 102801.1, 102720.3, 102637, 
    102554.2,
  103384.4, 103371.8, 103353.2, 103319.4, 103277.5, 103223.7, 103165.9, 
    103099.8, 103035.1, 102965.5, 102886.9, 102798.6, 102718.5, 102636.8, 
    102553.8,
  103352.3, 103338.4, 103321.6, 103291.4, 103252.8, 103203.1, 103148.7, 
    103085, 103023.8, 102954.7, 102877.1, 102791.1, 102710.8, 102629.9, 
    102546.1,
  103315, 103298.5, 103281.2, 103255.4, 103220.8, 103175.8, 103124.4, 
    103066.7, 103004.4, 102936.2, 102856.2, 102777, 102698.3, 102616.7, 
    102533.5,
  103423.6, 103361.3, 103286, 103206.4, 103118.8, 103028.7, 102948.2, 
    102862.8, 102776.4, 102686.9, 102601.4, 102513.9, 102425.7, 102334.7, 
    102249.9,
  103458.5, 103390.8, 103316.5, 103238.4, 103152.3, 103060.8, 102974.8, 
    102890, 102801.7, 102712.7, 102622.1, 102534.5, 102450.7, 102359.1, 
    102272.3,
  103472, 103405.8, 103335.3, 103260.8, 103175.3, 103084.3, 102995.9, 
    102908.6, 102818.4, 102729.3, 102638.3, 102547.1, 102462.1, 102373.9, 
    102286.1,
  103489.9, 103425.2, 103354.7, 103279, 103194.9, 103104.1, 103016.7, 
    102928.6, 102836.7, 102748.9, 102654.9, 102561.9, 102475.2, 102388, 
    102300.7,
  103508.8, 103435, 103366.5, 103288.9, 103208.7, 103117.6, 103030.5, 
    102940.7, 102850.5, 102761.3, 102668.5, 102574.2, 102485.2, 102398.2, 
    102310.3,
  103518.9, 103444.2, 103376.9, 103297.9, 103216.4, 103125.1, 103037.6, 
    102949.3, 102860.5, 102772.9, 102679.2, 102583.4, 102493.9, 102405.1, 
    102317.4,
  103528.5, 103451.1, 103381.8, 103299.4, 103216, 103129, 103042.1, 102951.5, 
    102863.1, 102775, 102682.7, 102588.6, 102497.3, 102407.2, 102320.1,
  103525.7, 103454.2, 103380.9, 103294.7, 103212, 103125.2, 103039.1, 
    102949.2, 102862.2, 102773.9, 102682.3, 102587.9, 102496.4, 102405.6, 
    102320.4,
  103517.1, 103451.8, 103370, 103282.3, 103199.3, 103115.6, 103030.4, 
    102938.7, 102854.1, 102764.4, 102674.1, 102581.4, 102489.8, 102397.8, 
    102312.5,
  103499.3, 103431, 103347.7, 103262.2, 103182.8, 103099.4, 103013.8, 
    102924.5, 102839.2, 102748.8, 102659.5, 102569.8, 102478.8, 102388.4, 
    102301.9,
  103386.4, 103317.2, 103241.1, 103156.6, 103060.6, 102961.9, 102872.4, 
    102780.8, 102690.1, 102604.3, 102504.1, 102413.1, 102323.5, 102230.4, 
    102142.7,
  103430.8, 103356.1, 103276.9, 103196.4, 103103.5, 103000.5, 102907, 
    102813.4, 102721.6, 102636.6, 102537.5, 102446.1, 102357.2, 102265.2, 
    102174.7,
  103457.5, 103385.5, 103308, 103225.8, 103132.8, 103030.5, 102934.9, 
    102839.5, 102745.5, 102660.4, 102561.3, 102469.2, 102378.3, 102286.2, 
    102195.7,
  103485.9, 103414.4, 103337, 103255.9, 103159.7, 103059.8, 102962.5, 
    102864.9, 102770.2, 102682.4, 102584.4, 102490, 102400.2, 102310.5, 
    102219.3,
  103503.1, 103434.3, 103358.2, 103273.7, 103180.1, 103080, 102982.8, 102885, 
    102786.8, 102698, 102601.3, 102507.8, 102417.7, 102328.3, 102237,
  103513.9, 103449.1, 103373.1, 103288.9, 103194.9, 103096.9, 103000.1, 
    102901.2, 102801.9, 102710.9, 102615.9, 102519.7, 102427.5, 102341.8, 
    102253.3,
  103519.6, 103454.6, 103379.8, 103293.8, 103201.5, 103105.4, 103008.7, 
    102911.6, 102812.7, 102719.3, 102622.5, 102527.9, 102436.1, 102346.2, 
    102260.1,
  103517, 103452.9, 103379.9, 103290.9, 103202.9, 103108.8, 103013.1, 
    102916.6, 102818.1, 102722.6, 102625.9, 102531.5, 102437.8, 102347.9, 
    102262.7,
  103508.5, 103436.5, 103366.8, 103280.8, 103195.9, 103104, 103010, 102914.1, 
    102818.7, 102720.3, 102622.3, 102528.5, 102436.6, 102345.5, 102258.4,
  103485, 103414.2, 103347.2, 103263.4, 103182.8, 103093.8, 103000.9, 
    102905.7, 102809.2, 102710.2, 102613.5, 102519.2, 102429.2, 102340.7, 
    102254.2,
  103293.7, 103237, 103158.3, 103074.1, 102987.3, 102905.7, 102820.6, 
    102730.5, 102640.1, 102554.7, 102461.2, 102384.2, 102301.7, 102216, 
    102139.7,
  103340.2, 103279.7, 103202.3, 103117.1, 103027.4, 102944.8, 102859.1, 
    102769.5, 102677.1, 102591.7, 102497.6, 102411.6, 102328.5, 102248.3, 
    102165.7,
  103370.8, 103306.3, 103231.8, 103147.8, 103056.5, 102971.6, 102886.9, 
    102798.9, 102706.4, 102621.8, 102524.6, 102433.2, 102346.3, 102264.4, 
    102186.2,
  103402, 103336.7, 103266.5, 103179.3, 103088.2, 103000.5, 102915.4, 102827, 
    102733.3, 102648, 102553.3, 102458.2, 102362.7, 102281.3, 102203.8,
  103422.2, 103357.5, 103288.3, 103199.8, 103112, 103021.3, 102934.8, 
    102846.9, 102754.9, 102667.8, 102575.2, 102476.7, 102382.4, 102289.9, 
    102214.8,
  103438.1, 103375.1, 103307, 103221.8, 103134.7, 103043.7, 102953.8, 
    102865.6, 102773.6, 102684.9, 102591.8, 102495.5, 102398.1, 102304.1, 
    102224.4,
  103440.2, 103380.3, 103314.9, 103232.8, 103148.2, 103057.9, 102966.5, 
    102877, 102786.8, 102697.4, 102602.1, 102508.4, 102411.7, 102317.1, 
    102229.5,
  103433.2, 103376.8, 103315.3, 103239.8, 103158.5, 103069.5, 102977.7, 
    102886.8, 102797.1, 102704.4, 102609.7, 102515.5, 102421.9, 102325.7, 
    102237,
  103410.2, 103362.1, 103304.3, 103234.9, 103157.3, 103070.4, 102980.5, 
    102891, 102800.1, 102705.6, 102611.4, 102518.2, 102425.7, 102330.6, 
    102241.5,
  103379.5, 103337.3, 103285.1, 103220.1, 103147.8, 103064.6, 102977.5, 
    102888.5, 102795.3, 102699.3, 102608, 102515.6, 102422.1, 102330.4, 
    102242.9,
  103203.6, 103151.6, 103085.5, 103004.2, 102926.9, 102852.4, 102778.5, 
    102699.3, 102622, 102532.1, 102450, 102368.2, 102286.7, 102207.6, 102134.1,
  103238.9, 103183.3, 103118.2, 103044.6, 102961.1, 102879.8, 102806.6, 
    102730.4, 102654, 102571.8, 102484.7, 102398, 102316.4, 102234.8, 102161.2,
  103269.1, 103213.6, 103148.9, 103080.4, 102999.9, 102915.4, 102835.5, 
    102756.7, 102677.6, 102597, 102508.9, 102423.4, 102337.8, 102254.8, 
    102177.2,
  103293.2, 103231.4, 103168.3, 103100.4, 103023.2, 102940.4, 102858.5, 
    102778.1, 102698, 102619.1, 102535.6, 102446.9, 102360.1, 102276, 102196.7,
  103304.3, 103244.9, 103183.1, 103117.8, 103047.5, 102966.5, 102882.6, 
    102798.9, 102715.9, 102632.4, 102548.8, 102463.3, 102378.3, 102292.3, 
    102212.4,
  103309, 103247.6, 103190.2, 103123.4, 103055.8, 102978.4, 102899.3, 102814, 
    102730.2, 102646.3, 102561.5, 102477.8, 102392.5, 102308, 102225.2,
  103295.8, 103239.2, 103183.8, 103116.8, 103055.3, 102984.1, 102907.6, 
    102826.1, 102740.6, 102652.2, 102566, 102483.7, 102401.4, 102318.2, 
    102236.7,
  103275.4, 103220.7, 103170.4, 103103.9, 103044.2, 102975.2, 102905.6, 
    102828.6, 102746.3, 102656.1, 102569.7, 102485.6, 102405.1, 102324, 
    102242.4,
  103242.4, 103192.6, 103142.4, 103079.7, 103021.2, 102953.3, 102890.8, 
    102819, 102742.7, 102653.7, 102567.1, 102481.7, 102400.8, 102321, 102243.4,
  103197.2, 103151.8, 103104.3, 103048.4, 102988, 102923.2, 102862.9, 
    102795.7, 102724.6, 102642.5, 102558.6, 102473.4, 102390.9, 102312.2, 
    102237.6,
  103210.4, 103152, 103083.8, 103019.9, 102943.8, 102872, 102799, 102720.4, 
    102638.7, 102559.5, 102473.2, 102392.4, 102310, 102229.9, 102158.1,
  103228.7, 103165.6, 103094.1, 103029.5, 102953, 102884.1, 102810.3, 
    102732.2, 102650.6, 102571.4, 102489.6, 102408.8, 102327.1, 102247.2, 
    102172,
  103233.4, 103172.4, 103100.8, 103030.8, 102957.1, 102888.6, 102815, 
    102738.1, 102656.4, 102576, 102494.9, 102417.5, 102335.8, 102254.8, 102180,
  103236.1, 103173.9, 103099, 103028.9, 102955.2, 102885.2, 102812.4, 
    102733.2, 102652.8, 102573.3, 102493.8, 102414.8, 102337, 102258.8, 
    102185.9,
  103228.2, 103167.4, 103091.9, 103018.2, 102948.7, 102877.3, 102802.9, 
    102724.9, 102645.2, 102567.7, 102489.1, 102409.5, 102335, 102259, 102186.1,
  103216.1, 103152.2, 103078, 103002.9, 102932, 102859.8, 102786.1, 102707.7, 
    102627.8, 102552.1, 102476.7, 102399.3, 102326.9, 102252.5, 102182.8,
  103192.8, 103125.4, 103053.4, 102981, 102911.4, 102839.1, 102767, 102685.1, 
    102606.5, 102533.9, 102459.4, 102384, 102314.4, 102241.9, 102172,
  103160.7, 103097, 103028.1, 102955.9, 102883.1, 102809.7, 102737.5, 102656, 
    102580.4, 102508.7, 102435.5, 102364.2, 102296.1, 102225.1, 102157.8,
  103124.2, 103062.8, 102992.2, 102919.8, 102848.5, 102775.3, 102702.8, 
    102620.8, 102550.4, 102476.6, 102409, 102337.4, 102271.4, 102203.9, 
    102138.8,
  103082.3, 103020.5, 102951, 102879.2, 102806.9, 102732.9, 102658.8, 
    102581.9, 102513.4, 102441.3, 102376.6, 102307.2, 102242.8, 102177.8, 
    102117.6,
  103248.6, 103176.5, 103097.3, 102998.8, 102912, 102817.7, 102729.2, 
    102633.5, 102546.6, 102459, 102375.2, 102299.5, 102223.6, 102146.6, 
    102074.6,
  103257.5, 103184.8, 103102.6, 103005, 102920.5, 102824.7, 102736, 102646.1, 
    102559.8, 102474.1, 102387.9, 102312, 102235.1, 102159.6, 102086.7,
  103251.6, 103179.7, 103100.1, 103008, 102920.1, 102823.1, 102731.7, 
    102642.6, 102555.4, 102472.7, 102386.7, 102312.1, 102237.8, 102161.7, 
    102088.9,
  103241, 103171.5, 103094.3, 103004.7, 102912.4, 102819.5, 102730, 102640.8, 
    102555.4, 102473, 102391.2, 102316, 102240, 102168.8, 102093.9,
  103221.1, 103156.2, 103080.8, 102993.5, 102901.7, 102808.9, 102717.2, 
    102626.9, 102542.4, 102463, 102384.9, 102309.6, 102236.4, 102166.3, 
    102093.6,
  103192.2, 103132.6, 103059.5, 102975.5, 102884.5, 102793.5, 102703.8, 
    102613, 102529.6, 102452, 102376.6, 102302.1, 102229.9, 102162.4, 102092.3,
  103159.1, 103101.2, 103031.5, 102951.1, 102861.4, 102773, 102681.1, 
    102589.5, 102507.6, 102431.9, 102358.5, 102285.4, 102215.6, 102150.7, 
    102085.3,
  103116, 103064.5, 102999, 102921.9, 102835, 102746.7, 102653.3, 102565.9, 
    102480.4, 102406.7, 102334.8, 102263.9, 102197.4, 102135.3, 102072.4,
  103073.9, 103025.5, 102961.1, 102885.4, 102800.6, 102711.1, 102620.6, 
    102531.8, 102448.8, 102374.4, 102299.6, 102236.5, 102171, 102114.2, 
    102054.2,
  103025.5, 102977.2, 102915, 102841.7, 102758.8, 102672.1, 102582.5, 
    102494.2, 102409.7, 102333.4, 102259.6, 102200, 102139.6, 102085.9, 
    102033.5,
  103171, 103092, 103006.1, 102912.7, 102818.8, 102725.7, 102637, 102545.4, 
    102453.9, 102364.2, 102279.1, 102197.2, 102123.1, 102051.3, 101982.8,
  103186.8, 103107.6, 103018.4, 102929.2, 102833.5, 102738, 102647.2, 102558, 
    102470.4, 102379.1, 102290.4, 102207.3, 102131.7, 102062.7, 101993.9,
  103195.7, 103114.6, 103027.7, 102936.9, 102841.3, 102743.9, 102652.6, 
    102561.1, 102472.6, 102382.2, 102295.6, 102211, 102132.7, 102060, 101993.9,
  103205.6, 103123.2, 103033.8, 102944.8, 102848, 102750.2, 102657.6, 
    102565.3, 102476.9, 102386.8, 102300.7, 102210.7, 102135, 102063.6, 
    101997.3,
  103210.6, 103126.9, 103039.3, 102948, 102851.1, 102753.5, 102658.9, 102564, 
    102473.9, 102384.1, 102297.6, 102207.7, 102132.5, 102058.4, 101993.2,
  103212.2, 103127.5, 103039.6, 102947.4, 102852.8, 102753.5, 102658.3, 
    102562.4, 102471.2, 102379.1, 102292.5, 102201.3, 102126.4, 102054.3, 
    101988,
  103209.6, 103122.2, 103035.8, 102944.2, 102850.4, 102752.4, 102655.3, 
    102558.3, 102464.3, 102370.8, 102283.6, 102192.7, 102116, 102044.2, 
    101976.3,
  103200.9, 103112.9, 103028, 102937, 102844.9, 102746.9, 102651.6, 102551.8, 
    102457.6, 102361, 102273, 102179.6, 102102.5, 102030.9, 101964.5,
  103186.2, 103100.2, 103014.5, 102924.3, 102833.8, 102737.8, 102641.7, 
    102541.2, 102447.2, 102348.3, 102257.5, 102165.9, 102086.4, 102013.9, 
    101947.2,
  103163.2, 103078, 102993.4, 102905.1, 102817.7, 102723.9, 102627.5, 
    102527.5, 102431.7, 102330.8, 102238.9, 102147.4, 102065.3, 101993.3, 
    101927.9,
  103223.3, 103135, 103036.3, 102936.5, 102835.6, 102736.6, 102641.8, 
    102542.9, 102455.5, 102365.9, 102290.6, 102210.9, 102136.5, 102065.1, 
    102003,
  103267.1, 103177.7, 103076.2, 102979.6, 102878.5, 102780.4, 102682.4, 
    102581.3, 102486.8, 102395.7, 102313.8, 102236.5, 102159.1, 102085, 
    102015.6,
  103296.6, 103207.5, 103105.6, 103008.4, 102908.7, 102811.6, 102713.7, 
    102613.5, 102515.6, 102422, 102331.1, 102251.4, 102170.4, 102096.6, 
    102026.3,
  103330.3, 103243, 103141.8, 103039.4, 102938.7, 102844.1, 102745.5, 
    102644.5, 102542.8, 102446, 102354, 102270.3, 102189.8, 102112.8, 102039.6,
  103352.6, 103268.1, 103166.1, 103065.2, 102965.9, 102870.2, 102772.2, 
    102671.5, 102572.3, 102470.8, 102373.6, 102283.9, 102201.9, 102122.7, 
    102048,
  103372.6, 103290, 103189.5, 103090.5, 102991, 102895.7, 102796.6, 102695.7, 
    102593.5, 102492.1, 102391.4, 102300.9, 102216.6, 102136.2, 102058.8,
  103382, 103303.1, 103204.2, 103108.2, 103010.6, 102915.8, 102817.2, 
    102716.7, 102615.8, 102511.5, 102408.2, 102313.9, 102226, 102142.9, 
    102065.4,
  103382, 103309.4, 103216, 103124.6, 103029, 102932.1, 102833.5, 102734.6, 
    102631.5, 102528.9, 102423, 102328.9, 102234.9, 102151.7, 102070.7,
  103375.5, 103305.1, 103220.6, 103132.6, 103039.1, 102946.3, 102844.8, 
    102748.9, 102645.3, 102543.2, 102436.7, 102340.2, 102240.9, 102157.7, 
    102072.4,
  103360.6, 103291.8, 103217.7, 103137.7, 103045.8, 102952.6, 102852.3, 
    102756.2, 102653.3, 102553, 102449.1, 102352.1, 102249.7, 102162.6, 
    102075.5,
  103123.2, 103047, 102959.4, 102868.5, 102776.4, 102691.2, 102600.7, 
    102510.2, 102425.7, 102334.5, 102256.2, 102180.9, 102106.4, 102038.3, 
    101975.6,
  103163.2, 103090.4, 102998.8, 102914.5, 102823.4, 102733.2, 102644.8, 
    102553.1, 102465, 102374.3, 102292.9, 102213.8, 102138.6, 102065.9, 
    101994.7,
  103188.7, 103119.2, 103034.7, 102948.4, 102858.2, 102768.4, 102679.4, 
    102585, 102497.5, 102404.3, 102317.2, 102237.2, 102157.9, 102085.9, 
    102012.7,
  103211, 103146, 103064.7, 102980.9, 102892.1, 102802.8, 102713.8, 102622.9, 
    102532.6, 102437, 102346.8, 102265.6, 102184.9, 102111.2, 102036.9,
  103226, 103165.7, 103088.5, 103004.7, 102921.3, 102833.4, 102743.5, 
    102651.7, 102560.4, 102465.7, 102372, 102288.4, 102205, 102130.7, 102054.9,
  103237.2, 103176.7, 103107.4, 103026.9, 102944.9, 102859.1, 102769.4, 
    102678.1, 102588.8, 102494.8, 102398.4, 102311.7, 102228.5, 102150.2, 
    102073.7,
  103236.9, 103181.8, 103119, 103043, 102964.1, 102879.1, 102792.1, 102701.7, 
    102611.8, 102518.7, 102422.5, 102331.1, 102245.3, 102165.7, 102087.7,
  103227.6, 103180.1, 103121.9, 103052, 102976.8, 102896.3, 102808, 102720.4, 
    102631.2, 102538, 102446.6, 102350.5, 102262.7, 102178.9, 102101.1,
  103210.9, 103169.9, 103119.7, 103053.5, 102982.4, 102904.8, 102820.3, 
    102732.4, 102644.6, 102552.1, 102461.3, 102366.5, 102278.7, 102191.2, 
    102110.9,
  103183.4, 103151.4, 103106.7, 103049.7, 102981.5, 102908.4, 102826.3, 
    102740.2, 102650.9, 102559.6, 102474.5, 102378.9, 102288.6, 102203.7, 
    102120.1,
  103069.4, 103009.2, 102944.7, 102867.5, 102793.2, 102715.3, 102633.8, 
    102554.8, 102472.2, 102389.4, 102312.1, 102239.9, 102166.2, 102095.2, 
    102033.1,
  103108.3, 103048.7, 102981.1, 102909.4, 102835.2, 102755.2, 102674.5, 
    102594.4, 102513.4, 102428.4, 102346.8, 102271, 102196, 102121.5, 102054.9,
  103134.5, 103075.1, 103011.5, 102941.1, 102867, 102787.5, 102708.1, 
    102625.2, 102542.6, 102458.9, 102373.4, 102295.5, 102217.9, 102141.6, 
    102073.8,
  103162.6, 103102.4, 103044.8, 102975.1, 102900.2, 102822.5, 102743.8, 
    102661.5, 102577.9, 102492.4, 102405.2, 102323.5, 102243.8, 102165.5, 
    102098.4,
  103181, 103123.9, 103069.6, 103001.4, 102930, 102852.1, 102772.3, 102688.5, 
    102606.7, 102520.7, 102432.3, 102348, 102265.2, 102185.9, 102116.2,
  103192.8, 103141, 103091.4, 103022.9, 102957, 102879.7, 102802, 102718.8, 
    102634.6, 102550, 102459.9, 102373.1, 102288.2, 102205.8, 102132.6,
  103195.1, 103149.5, 103104.3, 103040.7, 102978, 102904.7, 102825.1, 
    102744.6, 102657.8, 102571, 102484.8, 102395.2, 102309.4, 102223, 102145,
  103187.9, 103150.4, 103109.9, 103051.5, 102996, 102923.9, 102848.9, 
    102767.8, 102681.3, 102592.5, 102504.7, 102417.3, 102331.9, 102242.4, 
    102161.8,
  103173.1, 103144, 103107.8, 103059.3, 103003.4, 102937.9, 102863.2, 
    102784.5, 102700.9, 102610.7, 102523.6, 102433, 102348.1, 102262.5, 
    102175.9,
  103143.4, 103126.3, 103095.9, 103053.3, 103003.6, 102944.2, 102873.6, 
    102793.9, 102714.3, 102626.4, 102537.7, 102449, 102362.2, 102274, 102188.6,
  103088.9, 103042.6, 102990.3, 102922.7, 102854.5, 102777.3, 102700.6, 
    102611.6, 102525.7, 102438.6, 102358, 102275.3, 102196.7, 102120.4, 
    102046.4,
  103119.1, 103071.5, 103021.4, 102960.3, 102892.8, 102816.5, 102737.3, 
    102651.2, 102568.6, 102479.9, 102394.8, 102308.1, 102228.1, 102148.6, 
    102071.3,
  103136.6, 103091, 103040.6, 102986, 102922.1, 102849.9, 102774, 102688.2, 
    102602.2, 102512.8, 102427.9, 102340.1, 102255.8, 102175.6, 102096.1,
  103153.1, 103117.4, 103062.9, 103013.3, 102949.8, 102881.4, 102807, 102725, 
    102639.4, 102548.4, 102462.7, 102373, 102284.7, 102202, 102121.7,
  103162.3, 103134.4, 103082.3, 103032.4, 102973.8, 102907, 102834.8, 
    102755.6, 102671.3, 102580.5, 102492.5, 102402.6, 102314, 102227.5, 
    102148.8,
  103170.1, 103144.3, 103096.8, 103053.9, 102993.2, 102930.3, 102861.3, 
    102781.7, 102699.9, 102612.1, 102524, 102433.4, 102344.4, 102255.5, 
    102173.1,
  103172.2, 103146.3, 103108.5, 103065.2, 103008.2, 102948.8, 102882.1, 
    102803.4, 102727.1, 102638.5, 102553, 102463.4, 102371.9, 102283.1, 
    102196.1,
  103167.4, 103149.7, 103115.7, 103068.8, 103024, 102964.1, 102900.4, 102828, 
    102752.8, 102667.2, 102580.3, 102491.2, 102400.5, 102311.8, 102219.9,
  103159.6, 103148.5, 103123.1, 103083.1, 103033.4, 102978.5, 102915, 
    102845.3, 102771.4, 102688.7, 102604.2, 102517, 102425.3, 102333.7, 
    102244.2,
  103143.6, 103135.9, 103122.2, 103086.4, 103045, 102993.5, 102931.1, 
    102859.6, 102786.9, 102705.8, 102625.2, 102539.3, 102449.3, 102355.6, 
    102266.5 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
