netcdf atmos_static_scalar_2.ak {
dimensions:
        lat = 4 ;
        lon = 5 ;
variables:
        float ak(lat, lon) ;
                ak:long_name = "vertical coordinate sigma value" ;
                ak:units = "unit" ;
                ak:missing_value = 1.e+20f ;
                ak:_FillValue = 1.e+20f ;
                ak:cell_methods = "time: point" ;
        float lat(lat) ;
        float lon(lon) ;
data:
  lat = 0, 1, 2, 3 ;
  lon = 0, 1, 2, 3, 4 ;
  ak =
   1, 2, 3, 4, 5,
   6, 7, 8, 9, 10,
   11, 12, 13, 14, 15,
   16, 17, 18, 19, 20 ;

}
