netcdf \00010101.atmos_daily.tile1.pv350K {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pv350K(time, grid_yt, grid_xt) ;
		pv350K:_FillValue = -1.e+10f ;
		pv350K:missing_value = -1.e+10f ;
		pv350K:units = "(K m**2) / (kg s)" ;
		pv350K:long_name = "350-K potential vorticity; needs x350 scaling" ;
		pv350K:cell_methods = "time: mean" ;
		pv350K:time_avg_info = "average_T1,average_T2,average_DT" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:53:52 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile1.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile1.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.1986115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9611561, 0.1583273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7949425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7552791, 0.2484612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.9872221, 0.4156101, 0.04560489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.8345782, 0.2958934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.7792858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9990003, 0.3505592, 0.06537855, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.8140894, 0.2409153, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.9453563, 0.02902743, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pv350K =
  -6.345782e-09, -6.824058e-09, -7.157473e-09, -7.714317e-09, -8.259162e-09, 
    -8.899335e-09, -1.020669e-08, -1.187854e-08, -1.354385e-08, 
    -1.468332e-08, -1.539314e-08, -1.648653e-08, -1.7746e-08, -1.983302e-08, 
    -2.13391e-08,
  -5.751619e-09, -6.632147e-09, -7.041045e-09, -7.378787e-09, -7.99286e-09, 
    -8.604391e-09, -9.27736e-09, -1.096393e-08, -1.269173e-08, -1.429016e-08, 
    -1.529036e-08, -1.609618e-08, -1.721403e-08, -1.898138e-08, -2.063958e-08,
  -5.340269e-09, -6.124341e-09, -6.898285e-09, -7.204083e-09, -7.663374e-09, 
    -8.303989e-09, -8.883058e-09, -9.870698e-09, -1.174704e-08, 
    -1.349389e-08, -1.489214e-08, -1.578684e-08, -1.68605e-08, -1.826493e-08, 
    -1.977458e-08,
  -5.104273e-09, -5.624179e-09, -6.483545e-09, -7.078458e-09, -7.452819e-09, 
    -7.995606e-09, -8.597795e-09, -9.235281e-09, -1.068449e-08, 
    -1.258998e-08, -1.431905e-08, -1.543829e-08, -1.642919e-08, 
    -1.767978e-08, -1.909094e-08,
  -4.983757e-09, -5.253679e-09, -5.982201e-09, -6.816753e-09, -7.327861e-09, 
    -7.732511e-09, -8.2753e-09, -8.874557e-09, -9.713975e-09, -1.149491e-08, 
    -1.346395e-08, -1.517161e-08, -1.623236e-08, -1.721985e-08, -1.833636e-08,
  -4.841342e-09, -5.101296e-09, -5.504532e-09, -6.298507e-09, -7.082266e-09, 
    -7.580407e-09, -8.047398e-09, -8.57677e-09, -9.172604e-09, -1.0358e-08, 
    -1.225582e-08, -1.423418e-08, -1.598161e-08, -1.714121e-08, -1.796971e-08,
  -4.789169e-09, -4.954333e-09, -5.311746e-09, -5.868492e-09, -6.578404e-09, 
    -7.28893e-09, -7.839696e-09, -8.393926e-09, -8.875502e-09, -9.576901e-09, 
    -1.103033e-08, -1.306964e-08, -1.50192e-08, -1.68259e-08, -1.775487e-08,
  -4.707742e-09, -4.831061e-09, -5.14282e-09, -5.624799e-09, -6.183014e-09, 
    -6.865959e-09, -7.569045e-09, -8.166554e-09, -8.596387e-09, 
    -9.078513e-09, -9.908805e-09, -1.164328e-08, -1.369107e-08, 
    -1.582742e-08, -1.755846e-08,
  -4.655432e-09, -4.681917e-09, -4.970518e-09, -5.492916e-09, -5.959785e-09, 
    -6.34874e-09, -7.154489e-09, -7.957977e-09, -8.495327e-09, -8.866614e-09, 
    -9.367081e-09, -1.037971e-08, -1.216798e-08, -1.415569e-08, -1.612164e-08,
  -4.489276e-09, -4.569956e-09, -4.798855e-09, -5.244501e-09, -5.833527e-09, 
    -6.262477e-09, -6.64102e-09, -7.510938e-09, -8.307995e-09, -8.719199e-09, 
    -9.0509e-09, -9.638994e-09, -1.100389e-08, -1.270545e-08, -1.460554e-08,
  -3.01113e-09, -3.222485e-09, -3.864106e-09, -5.039569e-09, -5.801964e-09, 
    -6.337572e-09, -7.022841e-09, -7.921589e-09, -8.822564e-09, 
    -9.637915e-09, -1.064089e-08, -1.16841e-08, -1.262587e-08, -1.354776e-08, 
    -1.43053e-08,
  -2.702818e-09, -3.131114e-09, -3.52571e-09, -4.309948e-09, -5.299523e-09, 
    -6.077494e-09, -6.783319e-09, -7.555413e-09, -8.404291e-09, 
    -9.202457e-09, -1.007413e-08, -1.099778e-08, -1.1991e-08, -1.297498e-08, 
    -1.384074e-08,
  -2.476192e-09, -2.895126e-09, -3.337952e-09, -3.897114e-09, -4.679022e-09, 
    -5.529267e-09, -6.366129e-09, -7.179092e-09, -7.97772e-09, -8.809854e-09, 
    -9.616342e-09, -1.045255e-08, -1.135872e-08, -1.236226e-08, -1.335225e-08,
  -2.487192e-09, -2.679825e-09, -3.100116e-09, -3.592757e-09, -4.198401e-09, 
    -4.972625e-09, -5.868954e-09, -6.736262e-09, -7.563936e-09, 
    -8.399461e-09, -9.220741e-09, -9.994372e-09, -1.083364e-08, 
    -1.181392e-08, -1.289038e-08,
  -2.596205e-09, -2.618154e-09, -2.908821e-09, -3.33702e-09, -3.855183e-09, 
    -4.515592e-09, -5.378526e-09, -6.275982e-09, -7.135958e-09, 
    -7.993876e-09, -8.852368e-09, -9.666135e-09, -1.042435e-08, -1.13089e-08, 
    -1.246062e-08,
  -2.740707e-09, -2.689281e-09, -2.839499e-09, -3.130149e-09, -3.57771e-09, 
    -4.182247e-09, -4.977735e-09, -5.880926e-09, -6.778761e-09, 
    -7.638105e-09, -8.509498e-09, -9.330769e-09, -1.014364e-08, 
    -1.100275e-08, -1.212588e-08,
  -2.795966e-09, -2.811507e-09, -2.888794e-09, -3.009232e-09, -3.350985e-09, 
    -3.917945e-09, -4.662315e-09, -5.547188e-09, -6.507251e-09, 
    -7.430313e-09, -8.306988e-09, -9.14882e-09, -9.92054e-09, -1.076319e-08, 
    -1.186193e-08,
  -2.721901e-09, -2.88058e-09, -2.932127e-09, -3.013019e-09, -3.213458e-09, 
    -3.757751e-09, -4.452037e-09, -5.313557e-09, -6.285614e-09, 
    -7.250819e-09, -8.155022e-09, -9.022476e-09, -9.795722e-09, 
    -1.060393e-08, -1.156935e-08,
  -2.608892e-09, -2.857421e-09, -3.037957e-09, -3.081435e-09, -3.171751e-09, 
    -3.606665e-09, -4.300953e-09, -5.112669e-09, -6.086284e-09, 
    -7.083464e-09, -7.994063e-09, -8.865132e-09, -9.611611e-09, 
    -1.041572e-08, -1.130709e-08,
  -2.545095e-09, -2.868231e-09, -3.030967e-09, -3.13607e-09, -3.309025e-09, 
    -3.608919e-09, -4.118966e-09, -4.959329e-09, -5.871504e-09, 
    -6.855484e-09, -7.798996e-09, -8.697939e-09, -9.461026e-09, 
    -1.022612e-08, -1.106662e-08,
  -3.101458e-09, -3.758049e-09, -4.419856e-09, -5.024257e-09, -5.618399e-09, 
    -6.112923e-09, -6.226802e-09, -6.667536e-09, -7.162672e-09, 
    -7.486135e-09, -7.779005e-09, -8.262323e-09, -9.157303e-09, 
    -1.047446e-08, -1.199223e-08,
  -2.339775e-09, -2.931135e-09, -3.475594e-09, -4.14767e-09, -4.935642e-09, 
    -5.693913e-09, -6.00849e-09, -5.941839e-09, -6.156167e-09, -6.352686e-09, 
    -6.517828e-09, -6.826866e-09, -7.369482e-09, -8.112879e-09, -9.083573e-09,
  -1.852831e-09, -2.225171e-09, -2.672673e-09, -3.247132e-09, -3.94064e-09, 
    -4.652918e-09, -5.042963e-09, -4.90209e-09, -4.712078e-09, -4.746975e-09, 
    -4.916471e-09, -5.020734e-09, -5.362811e-09, -5.857553e-09, -6.627664e-09,
  -1.432862e-09, -1.550079e-09, -2.003421e-09, -2.418745e-09, -2.885487e-09, 
    -3.491277e-09, -3.98398e-09, -4.102132e-09, -3.755392e-09, -3.593501e-09, 
    -3.68073e-09, -3.82712e-09, -3.932263e-09, -4.336174e-09, -5.00481e-09,
  -1.497001e-09, -1.050893e-09, -1.144312e-09, -1.580424e-09, -2.116e-09, 
    -2.587627e-09, -2.939257e-09, -3.057006e-09, -3.022119e-09, 
    -3.079184e-09, -3.331375e-09, -3.580673e-09, -3.760971e-09, 
    -3.914471e-09, -4.321924e-09,
  -2.190504e-09, -1.292674e-09, -7.818418e-10, -8.542861e-10, -1.319301e-09, 
    -1.75471e-09, -2.009443e-09, -2.160474e-09, -2.395842e-09, -2.79188e-09, 
    -2.979299e-09, -3.078997e-09, -3.24344e-09, -3.416513e-09, -3.6579e-09,
  -3.214031e-09, -2.161635e-09, -1.357947e-09, -8.235002e-10, -8.502126e-10, 
    -1.114051e-09, -1.288006e-09, -1.493392e-09, -1.848983e-09, 
    -2.205401e-09, -2.448537e-09, -2.786846e-09, -3.20382e-09, -3.279476e-09, 
    -3.313213e-09,
  -3.540064e-09, -2.975663e-09, -2.263025e-09, -1.59211e-09, -1.262842e-09, 
    -1.414351e-09, -1.56592e-09, -1.646964e-09, -1.906546e-09, -2.224537e-09, 
    -2.374975e-09, -2.59614e-09, -3.000322e-09, -3.204049e-09, -3.154637e-09,
  -3.808307e-09, -3.13559e-09, -2.597689e-09, -2.066259e-09, -1.701299e-09, 
    -1.626871e-09, -1.96049e-09, -2.294127e-09, -2.515319e-09, -2.82333e-09, 
    -3.013833e-09, -3.143676e-09, -3.299776e-09, -3.402888e-09, -3.300852e-09,
  -3.440547e-09, -3.350983e-09, -2.628994e-09, -2.125434e-09, -1.897856e-09, 
    -1.971979e-09, -2.201672e-09, -2.700157e-09, -3.143903e-09, 
    -3.554583e-09, -3.713019e-09, -3.692796e-09, -3.6381e-09, -3.593042e-09, 
    -3.493926e-09,
  -7.99593e-09, -9.15216e-09, -1.026673e-08, -1.073831e-08, -1.073747e-08, 
    -1.076978e-08, -1.0818e-08, -1.092891e-08, -1.118427e-08, -1.183846e-08, 
    -1.321146e-08, -1.484275e-08, -1.646251e-08, -1.792893e-08, -1.926311e-08,
  -6.365544e-09, -7.652623e-09, -8.708104e-09, -9.772688e-09, -1.054723e-08, 
    -1.076463e-08, -1.073566e-08, -1.08157e-08, -1.099782e-08, -1.119981e-08, 
    -1.153006e-08, -1.220573e-08, -1.330902e-08, -1.451501e-08, -1.57344e-08,
  -4.264577e-09, -5.73796e-09, -7.126923e-09, -8.242237e-09, -9.287128e-09, 
    -1.012194e-08, -1.05717e-08, -1.06039e-08, -1.060692e-08, -1.074659e-08, 
    -1.093803e-08, -1.123448e-08, -1.159418e-08, -1.213423e-08, -1.277419e-08,
  -3.40008e-09, -3.986353e-09, -5.158097e-09, -6.449959e-09, -7.704164e-09, 
    -8.728857e-09, -9.60852e-09, -1.028195e-08, -1.057534e-08, -1.05807e-08, 
    -1.057514e-08, -1.065541e-08, -1.079626e-08, -1.068241e-08, -1.066568e-08,
  -3.271817e-09, -3.357403e-09, -3.747745e-09, -4.645766e-09, -5.849103e-09, 
    -7.135373e-09, -8.284299e-09, -9.154401e-09, -9.943522e-09, 
    -1.042182e-08, -1.056618e-08, -1.044604e-08, -1.027728e-08, 
    -1.016038e-08, -1.009193e-08,
  -3.133645e-09, -3.179103e-09, -3.266231e-09, -3.613693e-09, -4.356006e-09, 
    -5.346726e-09, -6.58568e-09, -7.729587e-09, -8.680167e-09, -9.333419e-09, 
    -9.811992e-09, -1.018875e-08, -1.015861e-08, -9.819894e-09, -9.806922e-09,
  -2.872456e-09, -2.925033e-09, -3.035114e-09, -3.16902e-09, -3.516639e-09, 
    -4.072433e-09, -4.855616e-09, -5.835259e-09, -6.969441e-09, -7.97464e-09, 
    -8.803306e-09, -9.26953e-09, -9.306555e-09, -9.51301e-09, -9.672625e-09,
  -2.749572e-09, -2.752698e-09, -2.841646e-09, -2.890876e-09, -2.945599e-09, 
    -3.210377e-09, -3.691824e-09, -4.329286e-09, -5.203001e-09, 
    -6.179678e-09, -7.200874e-09, -7.792487e-09, -8.322107e-09, 
    -8.881402e-09, -9.157743e-09,
  -2.794071e-09, -2.664533e-09, -2.603883e-09, -2.58651e-09, -2.5988e-09, 
    -2.578199e-09, -2.818073e-09, -3.284575e-09, -3.908008e-09, 
    -4.652433e-09, -5.509495e-09, -6.385357e-09, -7.052951e-09, 
    -7.791108e-09, -8.472387e-09,
  -2.759092e-09, -2.841291e-09, -2.685481e-09, -2.484461e-09, -2.349613e-09, 
    -2.367494e-09, -2.573338e-09, -2.849682e-09, -3.189176e-09, 
    -3.726741e-09, -4.415618e-09, -5.187841e-09, -5.942625e-09, 
    -6.643034e-09, -7.089957e-09,
  -5.105246e-09, -5.145785e-09, -5.127548e-09, -4.799462e-09, -4.716342e-09, 
    -4.960783e-09, -5.646629e-09, -6.643437e-09, -7.528008e-09, 
    -8.186941e-09, -8.868432e-09, -9.465077e-09, -9.836822e-09, 
    -9.742344e-09, -9.399512e-09,
  -4.965839e-09, -4.906445e-09, -4.824365e-09, -4.910637e-09, -4.869324e-09, 
    -4.903933e-09, -5.170347e-09, -5.61108e-09, -6.322243e-09, -7.174996e-09, 
    -7.964796e-09, -8.583932e-09, -9.18924e-09, -9.761534e-09, -1.000195e-08,
  -4.342528e-09, -4.26317e-09, -4.141507e-09, -4.157024e-09, -4.353042e-09, 
    -4.432162e-09, -4.422659e-09, -4.655081e-09, -5.076139e-09, 
    -5.844781e-09, -6.796375e-09, -7.649477e-09, -8.397505e-09, 
    -8.990511e-09, -9.457252e-09,
  -3.643158e-09, -3.834533e-09, -3.960223e-09, -4.021519e-09, -4.082137e-09, 
    -4.209262e-09, -4.262025e-09, -4.304418e-09, -4.549938e-09, 
    -5.038428e-09, -5.742187e-09, -6.609385e-09, -7.415861e-09, -8.07866e-09, 
    -8.667513e-09,
  -2.871793e-09, -3.159081e-09, -3.574433e-09, -3.875797e-09, -3.964749e-09, 
    -4.078893e-09, -4.159072e-09, -4.194632e-09, -4.300797e-09, 
    -4.579099e-09, -5.016114e-09, -5.663024e-09, -6.532671e-09, -7.23126e-09, 
    -7.795038e-09,
  -2.280629e-09, -2.618662e-09, -3.029523e-09, -3.474572e-09, -3.711706e-09, 
    -3.849659e-09, -3.995353e-09, -4.09814e-09, -4.131198e-09, -4.309805e-09, 
    -4.555468e-09, -4.989693e-09, -5.661133e-09, -6.40229e-09, -7.028535e-09,
  -1.837491e-09, -2.183467e-09, -2.555393e-09, -2.980001e-09, -3.3284e-09, 
    -3.541386e-09, -3.774934e-09, -3.943429e-09, -3.99754e-09, -4.065126e-09, 
    -4.226851e-09, -4.530901e-09, -4.98932e-09, -5.605824e-09, -6.178356e-09,
  -1.443894e-09, -1.782168e-09, -2.19262e-09, -2.557067e-09, -2.962724e-09, 
    -3.22457e-09, -3.448204e-09, -3.726582e-09, -3.884132e-09, -3.88242e-09, 
    -3.962347e-09, -4.215748e-09, -4.590748e-09, -4.978881e-09, -5.448126e-09,
  -1.093205e-09, -1.263476e-09, -1.680457e-09, -2.191925e-09, -2.609112e-09, 
    -2.944149e-09, -3.051337e-09, -3.261288e-09, -3.607745e-09, 
    -3.721256e-09, -3.801063e-09, -3.982756e-09, -4.249697e-09, -4.54841e-09, 
    -4.882379e-09,
  -7.96095e-10, -7.296955e-10, -9.318507e-10, -1.491573e-09, -1.898463e-09, 
    -2.443878e-09, -2.813014e-09, -2.876773e-09, -3.129339e-09, 
    -3.445838e-09, -3.602711e-09, -3.76602e-09, -3.952171e-09, -4.182745e-09, 
    -4.406675e-09,
  -5.051225e-09, -4.451228e-09, -3.970282e-09, -3.843553e-09, -4.012195e-09, 
    -4.314144e-09, -4.535738e-09, -4.459039e-09, -4.087357e-09, 
    -3.821949e-09, -3.826393e-09, -3.834551e-09, -3.663894e-09, 
    -3.286341e-09, -2.89236e-09,
  -2.640413e-09, -2.381055e-09, -2.348067e-09, -2.749369e-09, -3.211211e-09, 
    -3.376996e-09, -3.180457e-09, -2.862675e-09, -2.666847e-09, -2.58455e-09, 
    -2.516702e-09, -2.578936e-09, -2.653239e-09, -2.791296e-09, -3.119876e-09,
  -1.903809e-09, -1.966462e-09, -2.056031e-09, -2.423019e-09, -2.514551e-09, 
    -2.374811e-09, -2.163437e-09, -2.064333e-09, -2.019475e-09, 
    -1.944376e-09, -1.974215e-09, -2.163466e-09, -2.448714e-09, 
    -2.752364e-09, -3.214998e-09,
  -1.112362e-09, -1.37389e-09, -1.700873e-09, -1.811469e-09, -1.764265e-09, 
    -1.708755e-09, -1.637153e-09, -1.502189e-09, -1.551401e-09, 
    -1.654491e-09, -1.702372e-09, -1.831265e-09, -2.132985e-09, 
    -2.495405e-09, -2.811591e-09,
  -7.03701e-10, -9.951284e-10, -1.37097e-09, -1.584334e-09, -1.635361e-09, 
    -1.662554e-09, -1.47501e-09, -1.276908e-09, -1.239617e-09, -1.243152e-09, 
    -1.415725e-09, -1.73728e-09, -2.051867e-09, -2.473154e-09, -2.806825e-09,
  -5.016336e-10, -7.685338e-10, -9.940687e-10, -1.220669e-09, -1.407822e-09, 
    -1.524658e-09, -1.525176e-09, -1.556528e-09, -1.509529e-09, 
    -1.602978e-09, -1.637133e-09, -1.803224e-09, -2.045047e-09, 
    -2.397454e-09, -2.685729e-09,
  -6.863382e-10, -7.791288e-10, -8.483858e-10, -8.642052e-10, -1.071543e-09, 
    -1.309028e-09, -1.627166e-09, -1.910452e-09, -2.087318e-09, 
    -2.144367e-09, -2.150525e-09, -2.087737e-09, -2.109119e-09, 
    -2.275914e-09, -2.523823e-09,
  -9.81101e-10, -9.986374e-10, -1.029593e-09, -9.702671e-10, -1.065909e-09, 
    -1.287422e-09, -1.548982e-09, -1.798297e-09, -2.009023e-09, 
    -2.130633e-09, -2.206741e-09, -2.159206e-09, -2.246789e-09, 
    -2.413857e-09, -2.715462e-09,
  -1.337471e-09, -1.314735e-09, -1.32954e-09, -1.417981e-09, -1.519665e-09, 
    -1.613014e-09, -1.695615e-09, -1.769827e-09, -1.958432e-09, 
    -2.031665e-09, -1.955359e-09, -1.893944e-09, -2.186455e-09, 
    -2.580799e-09, -2.960391e-09,
  -1.814666e-09, -1.851233e-09, -1.802712e-09, -1.807594e-09, -1.723844e-09, 
    -1.601585e-09, -1.478196e-09, -1.466336e-09, -1.682757e-09, 
    -1.946636e-09, -1.979034e-09, -2.007119e-09, -2.285818e-09, 
    -2.385387e-09, -2.387124e-09,
  -1.52709e-08, -1.554971e-08, -1.572285e-08, -1.590981e-08, -1.622007e-08, 
    -1.664874e-08, -1.708236e-08, -1.741688e-08, -1.749236e-08, 
    -1.732584e-08, -1.665743e-08, -1.582202e-08, -1.453544e-08, 
    -1.358833e-08, -1.277925e-08,
  -1.282204e-08, -1.321906e-08, -1.354681e-08, -1.379647e-08, -1.40469e-08, 
    -1.431632e-08, -1.44553e-08, -1.450543e-08, -1.432284e-08, -1.395731e-08, 
    -1.362596e-08, -1.340481e-08, -1.331938e-08, -1.318325e-08, -1.279492e-08,
  -9.424884e-09, -1.0266e-08, -1.10289e-08, -1.165218e-08, -1.19719e-08, 
    -1.206949e-08, -1.192182e-08, -1.154131e-08, -1.104929e-08, 
    -1.024263e-08, -1.014578e-08, -9.977356e-09, -1.001835e-08, 
    -9.976729e-09, -9.526985e-09,
  -5.750501e-09, -6.583953e-09, -7.361181e-09, -8.186437e-09, -8.807512e-09, 
    -9.20186e-09, -9.228003e-09, -9.117247e-09, -8.927276e-09, -8.356319e-09, 
    -8.360402e-09, -8.364797e-09, -8.419533e-09, -8.066155e-09, -7.489097e-09,
  -2.949791e-09, -3.534772e-09, -4.336445e-09, -5.090532e-09, -5.762514e-09, 
    -6.106357e-09, -6.580384e-09, -7.002568e-09, -7.056427e-09, 
    -7.013419e-09, -6.905013e-09, -6.76695e-09, -6.569154e-09, -6.124964e-09, 
    -5.571099e-09,
  -1.117323e-09, -1.148439e-09, -1.445822e-09, -2.013734e-09, -2.732264e-09, 
    -3.733035e-09, -4.558679e-09, -4.864056e-09, -5.035816e-09, 
    -5.264336e-09, -5.199477e-09, -5.116187e-09, -4.747937e-09, 
    -4.239716e-09, -3.747604e-09,
  -6.025896e-10, -2.78454e-10, -1.553925e-10, -3.216036e-10, -9.494995e-10, 
    -1.910074e-09, -2.723848e-09, -3.494538e-09, -3.891573e-09, -3.97936e-09, 
    -3.891287e-09, -3.651368e-09, -3.438196e-09, -3.102058e-09, -2.896833e-09,
  -6.336947e-10, -4.971721e-10, -5.059273e-10, -6.770047e-10, -7.870586e-10, 
    -1.192665e-09, -1.481595e-09, -1.850132e-09, -2.233433e-09, 
    -2.406621e-09, -2.53713e-09, -2.509998e-09, -2.379918e-09, -2.318022e-09, 
    -2.332889e-09,
  -7.404287e-10, -6.469575e-10, -6.686609e-10, -8.02437e-10, -8.479493e-10, 
    -9.117961e-10, -1.075378e-09, -9.58558e-10, -1.079904e-09, -1.221012e-09, 
    -1.366166e-09, -1.41265e-09, -1.510637e-09, -1.669858e-09, -1.752457e-09,
  -6.185718e-10, -6.467897e-10, -4.719234e-10, -3.779086e-10, -4.672195e-10, 
    -6.646592e-10, -1.028505e-09, -1.010378e-09, -8.780374e-10, -9.65474e-10, 
    -1.35097e-09, -1.201912e-09, -1.006935e-09, -1.084786e-09, -1.181159e-09,
  -1.550212e-08, -1.672344e-08, -1.769918e-08, -1.735011e-08, -1.655171e-08, 
    -1.552644e-08, -1.468877e-08, -1.451503e-08, -1.464496e-08, 
    -1.479424e-08, -1.505634e-08, -1.525341e-08, -1.524104e-08, 
    -1.506317e-08, -1.483763e-08,
  -1.381694e-08, -1.498059e-08, -1.620235e-08, -1.74031e-08, -1.818604e-08, 
    -1.83119e-08, -1.776015e-08, -1.677801e-08, -1.570311e-08, -1.503372e-08, 
    -1.493092e-08, -1.504084e-08, -1.524545e-08, -1.529964e-08, -1.51794e-08,
  -1.069092e-08, -1.192081e-08, -1.32776e-08, -1.465986e-08, -1.614255e-08, 
    -1.748459e-08, -1.841205e-08, -1.873233e-08, -1.844312e-08, 
    -1.769902e-08, -1.663433e-08, -1.583305e-08, -1.534002e-08, 
    -1.537735e-08, -1.55976e-08,
  -7.883875e-09, -8.528207e-09, -9.284456e-09, -1.049323e-08, -1.214297e-08, 
    -1.409095e-08, -1.584798e-08, -1.737608e-08, -1.846044e-08, 
    -1.907126e-08, -1.906587e-08, -1.853023e-08, -1.780998e-08, 
    -1.689726e-08, -1.618364e-08,
  -5.617756e-09, -6.18502e-09, -6.769643e-09, -7.405654e-09, -8.125847e-09, 
    -9.359503e-09, -1.100723e-08, -1.296771e-08, -1.472883e-08, 
    -1.629558e-08, -1.762921e-08, -1.858945e-08, -1.90916e-08, -1.908873e-08, 
    -1.873098e-08,
  -4.174386e-09, -4.395186e-09, -4.683763e-09, -4.914759e-09, -5.304663e-09, 
    -5.944479e-09, -6.958548e-09, -8.363874e-09, -1.024627e-08, 
    -1.230565e-08, -1.436569e-08, -1.59736e-08, -1.728472e-08, -1.818424e-08, 
    -1.883706e-08,
  -2.519775e-09, -2.622322e-09, -2.782756e-09, -2.835703e-09, -2.862782e-09, 
    -2.911001e-09, -3.181398e-09, -4.090707e-09, -5.441048e-09, 
    -7.061295e-09, -8.963005e-09, -1.103863e-08, -1.302157e-08, 
    -1.477595e-08, -1.600473e-08,
  -1.537425e-09, -1.201961e-09, -1.046881e-09, -1.322047e-09, -1.464856e-09, 
    -1.65693e-09, -1.897589e-09, -2.122608e-09, -2.69498e-09, -3.428786e-09, 
    -4.516471e-09, -5.913806e-09, -7.625764e-09, -9.397726e-09, -1.111329e-08,
  -1.134378e-09, -1.024044e-09, -9.183478e-10, -9.365839e-10, -9.081786e-10, 
    -9.941714e-10, -1.18913e-09, -1.361378e-09, -1.568117e-09, -1.897247e-09, 
    -2.294761e-09, -2.84472e-09, -3.741257e-09, -5.067388e-09, -6.660624e-09,
  -1.14632e-09, -1.035557e-09, -8.338579e-10, -7.938324e-10, -8.758441e-10, 
    -1.07206e-09, -1.269061e-09, -1.09914e-09, -9.816941e-10, -1.243844e-09, 
    -1.333741e-09, -1.665101e-09, -1.995612e-09, -2.560012e-09, -3.537114e-09,
  -1.020913e-08, -1.053552e-08, -1.098447e-08, -1.148597e-08, -1.180852e-08, 
    -1.174964e-08, -1.132429e-08, -1.070651e-08, -1.002512e-08, 
    -9.538558e-09, -9.240127e-09, -9.205869e-09, -9.637918e-09, 
    -1.014365e-08, -1.075479e-08,
  -9.869759e-09, -1.0182e-08, -1.046594e-08, -1.090874e-08, -1.142178e-08, 
    -1.199989e-08, -1.241912e-08, -1.246818e-08, -1.199837e-08, 
    -1.151397e-08, -1.086516e-08, -1.022242e-08, -9.801857e-09, 
    -9.921879e-09, -1.048884e-08,
  -9.050274e-09, -9.293126e-09, -9.491378e-09, -9.822271e-09, -1.024878e-08, 
    -1.074031e-08, -1.123652e-08, -1.177365e-08, -1.219196e-08, 
    -1.246742e-08, -1.231746e-08, -1.190198e-08, -1.136909e-08, 
    -1.065366e-08, -1.032587e-08,
  -8.0387e-09, -8.176578e-09, -8.329843e-09, -8.63325e-09, -8.881036e-09, 
    -9.208419e-09, -9.593007e-09, -1.021802e-08, -1.081753e-08, 
    -1.125483e-08, -1.170627e-08, -1.214703e-08, -1.228632e-08, 
    -1.211107e-08, -1.168865e-08,
  -6.519942e-09, -6.993527e-09, -7.421428e-09, -7.865319e-09, -8.052211e-09, 
    -8.108081e-09, -7.937742e-09, -8.363117e-09, -9.041983e-09, 
    -9.897814e-09, -1.052179e-08, -1.094216e-08, -1.146443e-08, 
    -1.200104e-08, -1.227585e-08,
  -4.913281e-09, -5.394051e-09, -6.040142e-09, -6.545796e-09, -6.781903e-09, 
    -6.847088e-09, -6.678127e-09, -6.391726e-09, -6.715969e-09, -7.59433e-09, 
    -8.697152e-09, -9.638232e-09, -1.040177e-08, -1.102997e-08, -1.174394e-08,
  -3.99437e-09, -4.472851e-09, -5.13072e-09, -5.535723e-09, -5.548763e-09, 
    -5.471265e-09, -5.534564e-09, -5.503557e-09, -5.56906e-09, -5.691474e-09, 
    -6.265196e-09, -7.12219e-09, -8.198722e-09, -9.461732e-09, -1.061895e-08,
  -3.076428e-09, -3.650251e-09, -4.177859e-09, -4.400385e-09, -4.564581e-09, 
    -4.433585e-09, -4.673081e-09, -4.932041e-09, -5.325141e-09, 
    -5.429114e-09, -5.434596e-09, -5.617459e-09, -6.078419e-09, 
    -6.849967e-09, -8.058882e-09,
  -2.359456e-09, -2.836191e-09, -3.340025e-09, -3.624582e-09, -3.738205e-09, 
    -3.911599e-09, -4.572944e-09, -5.071649e-09, -5.31386e-09, -5.415912e-09, 
    -5.689319e-09, -5.827496e-09, -5.852122e-09, -5.961668e-09, -6.210653e-09,
  -1.872368e-09, -2.229207e-09, -2.633051e-09, -2.997698e-09, -3.100942e-09, 
    -3.460711e-09, -4.075279e-09, -4.812249e-09, -5.147575e-09, 
    -5.461863e-09, -5.677165e-09, -5.892839e-09, -5.766472e-09, -5.92724e-09, 
    -6.127362e-09,
  -5.733561e-09, -5.7797e-09, -5.878449e-09, -6.111276e-09, -6.425147e-09, 
    -6.717283e-09, -6.964214e-09, -7.133561e-09, -7.281346e-09, 
    -7.447622e-09, -7.595908e-09, -7.705188e-09, -7.833893e-09, 
    -7.942557e-09, -8.072251e-09,
  -6.078009e-09, -6.162008e-09, -6.20427e-09, -6.26241e-09, -6.409739e-09, 
    -6.633726e-09, -6.925135e-09, -7.221414e-09, -7.487395e-09, 
    -7.684124e-09, -7.842801e-09, -7.988084e-09, -8.115165e-09, 
    -8.251599e-09, -8.292856e-09,
  -6.304259e-09, -6.365508e-09, -6.410256e-09, -6.467304e-09, -6.56636e-09, 
    -6.728304e-09, -6.912555e-09, -7.160848e-09, -7.434721e-09, 
    -7.694855e-09, -8.022668e-09, -8.25616e-09, -8.455282e-09, -8.606285e-09, 
    -8.704625e-09,
  -6.36808e-09, -6.399114e-09, -6.460461e-09, -6.579405e-09, -6.726015e-09, 
    -6.900265e-09, -7.069477e-09, -7.275313e-09, -7.477888e-09, 
    -7.751866e-09, -8.031147e-09, -8.509021e-09, -8.901288e-09, 
    -9.239701e-09, -9.515734e-09,
  -6.201291e-09, -6.20173e-09, -6.247478e-09, -6.426191e-09, -6.579481e-09, 
    -6.734487e-09, -6.93989e-09, -7.200464e-09, -7.540703e-09, -7.895858e-09, 
    -8.50464e-09, -9.331802e-09, -9.893426e-09, -9.933069e-09, -9.742309e-09,
  -5.919154e-09, -5.99796e-09, -6.060042e-09, -6.211244e-09, -6.417335e-09, 
    -6.56015e-09, -6.811888e-09, -7.071606e-09, -7.433985e-09, -7.685259e-09, 
    -8.304482e-09, -8.936819e-09, -8.31171e-09, -7.792201e-09, -8.111062e-09,
  -5.757936e-09, -5.887351e-09, -6.096207e-09, -6.312419e-09, -6.489476e-09, 
    -6.658594e-09, -6.915168e-09, -7.153357e-09, -7.456318e-09, 
    -7.633602e-09, -8.053525e-09, -8.616323e-09, -7.818957e-09, 
    -7.248622e-09, -6.231605e-09,
  -5.248532e-09, -5.323986e-09, -5.571287e-09, -5.857829e-09, -6.034435e-09, 
    -6.249236e-09, -6.42969e-09, -6.810958e-09, -7.202892e-09, -7.461766e-09, 
    -7.502139e-09, -7.657549e-09, -6.939008e-09, -6.100797e-09, -5.784607e-09,
  -4.302146e-09, -4.281663e-09, -4.53055e-09, -4.740795e-09, -4.993077e-09, 
    -5.13902e-09, -5.419983e-09, -5.611255e-09, -5.933937e-09, -6.298894e-09, 
    -6.444599e-09, -6.625588e-09, -6.970035e-09, -6.026424e-09, -5.183352e-09,
  -3.202282e-09, -3.237593e-09, -3.42011e-09, -3.632789e-09, -3.732829e-09, 
    -4.185043e-09, -4.685392e-09, -5.114976e-09, -5.22819e-09, -5.35774e-09, 
    -5.339329e-09, -5.463449e-09, -5.988295e-09, -6.397393e-09, -6.117669e-09,
  -1.886643e-09, -2.040453e-09, -2.213387e-09, -2.317341e-09, -2.538664e-09, 
    -2.770201e-09, -3.044391e-09, -3.407564e-09, -3.908258e-09, 
    -4.550922e-09, -5.229115e-09, -5.966655e-09, -6.705583e-09, 
    -7.394514e-09, -8.131592e-09,
  -1.693215e-09, -1.829195e-09, -2.002635e-09, -2.128004e-09, -2.193369e-09, 
    -2.38187e-09, -2.655553e-09, -2.949156e-09, -3.27893e-09, -3.722311e-09, 
    -4.319569e-09, -4.95519e-09, -5.615556e-09, -6.270096e-09, -6.941809e-09,
  -1.601858e-09, -1.683875e-09, -1.818934e-09, -1.971809e-09, -2.092919e-09, 
    -2.178443e-09, -2.375175e-09, -2.634808e-09, -2.936002e-09, -3.24228e-09, 
    -3.586917e-09, -4.109941e-09, -4.664175e-09, -5.271191e-09, -5.870348e-09,
  -1.614005e-09, -1.630594e-09, -1.727433e-09, -1.834903e-09, -1.98346e-09, 
    -2.094228e-09, -2.204108e-09, -2.386215e-09, -2.630124e-09, 
    -2.945571e-09, -3.242516e-09, -3.568778e-09, -3.962074e-09, 
    -4.393858e-09, -4.942306e-09,
  -1.754057e-09, -1.671899e-09, -1.677451e-09, -1.779165e-09, -1.91331e-09, 
    -2.081388e-09, -2.256751e-09, -2.391828e-09, -2.540303e-09, 
    -2.723635e-09, -2.959631e-09, -3.189833e-09, -3.481123e-09, 
    -3.841261e-09, -4.280884e-09,
  -2.042303e-09, -1.880484e-09, -1.807078e-09, -1.800946e-09, -1.869092e-09, 
    -1.969637e-09, -2.123922e-09, -2.314813e-09, -2.467163e-09, 
    -2.602744e-09, -2.724605e-09, -2.887302e-09, -3.098641e-09, 
    -3.390462e-09, -3.761327e-09,
  -2.447358e-09, -2.266651e-09, -2.10048e-09, -2.043999e-09, -2.043548e-09, 
    -2.095704e-09, -2.139319e-09, -2.230635e-09, -2.369296e-09, 
    -2.506469e-09, -2.627044e-09, -2.747846e-09, -2.9247e-09, -3.191735e-09, 
    -3.479427e-09,
  -3.133565e-09, -2.988701e-09, -2.842878e-09, -2.723294e-09, -2.6422e-09, 
    -2.634492e-09, -2.644936e-09, -2.670101e-09, -2.72088e-09, -2.804742e-09, 
    -2.925501e-09, -3.058236e-09, -3.199749e-09, -3.417604e-09, -3.648998e-09,
  -4.017012e-09, -3.845575e-09, -3.707252e-09, -3.587196e-09, -3.507198e-09, 
    -3.361022e-09, -3.291523e-09, -3.284019e-09, -3.365348e-09, 
    -3.496921e-09, -3.612987e-09, -3.776199e-09, -3.936146e-09, 
    -4.106145e-09, -4.237985e-09,
  -5.116019e-09, -4.852811e-09, -4.470941e-09, -4.295602e-09, -4.081905e-09, 
    -3.992971e-09, -3.944231e-09, -3.878305e-09, -3.794152e-09, 
    -3.899244e-09, -4.014354e-09, -4.141015e-09, -4.256868e-09, 
    -4.431267e-09, -4.655628e-09,
  -2.954891e-09, -2.940949e-09, -2.921849e-09, -2.894701e-09, -2.869269e-09, 
    -2.866761e-09, -2.886765e-09, -2.897795e-09, -2.92223e-09, -2.96884e-09, 
    -3.071658e-09, -3.191986e-09, -3.320083e-09, -3.469764e-09, -3.660686e-09,
  -2.950863e-09, -2.868604e-09, -2.792458e-09, -2.739342e-09, -2.691565e-09, 
    -2.644361e-09, -2.606945e-09, -2.603255e-09, -2.616883e-09, 
    -2.639262e-09, -2.68127e-09, -2.767619e-09, -2.86795e-09, -2.995206e-09, 
    -3.140493e-09,
  -3.103126e-09, -2.994723e-09, -2.831482e-09, -2.711942e-09, -2.626181e-09, 
    -2.554827e-09, -2.498036e-09, -2.451252e-09, -2.399995e-09, 
    -2.382589e-09, -2.356254e-09, -2.370777e-09, -2.407396e-09, 
    -2.485013e-09, -2.594615e-09,
  -3.291845e-09, -3.217761e-09, -3.012268e-09, -2.838621e-09, -2.665519e-09, 
    -2.561884e-09, -2.486811e-09, -2.441844e-09, -2.378839e-09, 
    -2.317664e-09, -2.263699e-09, -2.229034e-09, -2.223741e-09, 
    -2.240105e-09, -2.311338e-09,
  -3.511148e-09, -3.32348e-09, -3.119404e-09, -2.927018e-09, -2.759132e-09, 
    -2.686906e-09, -2.64951e-09, -2.601964e-09, -2.555009e-09, -2.465232e-09, 
    -2.358587e-09, -2.26457e-09, -2.214006e-09, -2.20983e-09, -2.207067e-09,
  -3.53402e-09, -3.392351e-09, -3.184587e-09, -2.891776e-09, -2.742826e-09, 
    -2.755337e-09, -2.747886e-09, -2.71534e-09, -2.711684e-09, -2.623325e-09, 
    -2.486432e-09, -2.36923e-09, -2.282368e-09, -2.244205e-09, -2.213608e-09,
  -3.613915e-09, -3.452199e-09, -3.162429e-09, -3.012645e-09, -3.104802e-09, 
    -3.071931e-09, -2.774565e-09, -2.569909e-09, -2.493376e-09, 
    -2.392827e-09, -2.294552e-09, -2.207567e-09, -2.162719e-09, 
    -2.145714e-09, -2.156533e-09,
  -3.983313e-09, -3.89735e-09, -3.657391e-09, -3.726662e-09, -3.744769e-09, 
    -3.128976e-09, -2.698903e-09, -2.483498e-09, -2.384094e-09, 
    -2.295228e-09, -2.184011e-09, -2.084536e-09, -1.995996e-09, 
    -1.979453e-09, -1.951913e-09,
  -4.61133e-09, -4.739479e-09, -4.315996e-09, -4.391627e-09, -4.309636e-09, 
    -3.521446e-09, -3.055701e-09, -2.678649e-09, -2.361655e-09, 
    -2.127399e-09, -1.939334e-09, -1.854638e-09, -1.793961e-09, -1.78774e-09, 
    -1.778321e-09,
  -5.691651e-09, -5.562049e-09, -5.237578e-09, -5.063903e-09, -4.633097e-09, 
    -3.771341e-09, -3.196157e-09, -2.693645e-09, -2.175682e-09, -1.88079e-09, 
    -1.716162e-09, -1.638482e-09, -1.59557e-09, -1.576156e-09, -1.579627e-09,
  -3.016034e-09, -3.161479e-09, -3.243857e-09, -3.305971e-09, -3.353313e-09, 
    -3.394517e-09, -3.438414e-09, -3.49367e-09, -3.543005e-09, -3.595555e-09, 
    -3.635405e-09, -3.649801e-09, -3.656526e-09, -3.628291e-09, -3.594393e-09,
  -2.609511e-09, -2.773197e-09, -2.925925e-09, -3.069835e-09, -3.180763e-09, 
    -3.261301e-09, -3.364538e-09, -3.464655e-09, -3.552847e-09, 
    -3.633626e-09, -3.689845e-09, -3.705181e-09, -3.696552e-09, -3.66598e-09, 
    -3.629999e-09,
  -2.385594e-09, -2.533595e-09, -2.631084e-09, -2.794766e-09, -2.928821e-09, 
    -3.055868e-09, -3.21233e-09, -3.381436e-09, -3.559826e-09, -3.674425e-09, 
    -3.781172e-09, -3.844081e-09, -3.871533e-09, -3.852538e-09, -3.82074e-09,
  -2.27506e-09, -2.368539e-09, -2.467447e-09, -2.662679e-09, -2.732005e-09, 
    -2.876299e-09, -3.00194e-09, -3.150969e-09, -3.305532e-09, -3.470674e-09, 
    -3.625206e-09, -3.747837e-09, -3.857926e-09, -3.92085e-09, -3.965761e-09,
  -2.186748e-09, -2.385402e-09, -2.570924e-09, -2.622191e-09, -2.754255e-09, 
    -2.927023e-09, -3.06753e-09, -3.159209e-09, -3.293315e-09, -3.420443e-09, 
    -3.595541e-09, -3.733911e-09, -3.851575e-09, -3.915659e-09, -3.993236e-09,
  -2.236304e-09, -2.39412e-09, -2.703276e-09, -2.804875e-09, -2.942314e-09, 
    -3.08367e-09, -3.172135e-09, -3.296262e-09, -3.386224e-09, -3.547344e-09, 
    -3.739461e-09, -3.857877e-09, -3.901829e-09, -3.935241e-09, -4.01382e-09,
  -2.345164e-09, -2.635604e-09, -2.837671e-09, -3.010244e-09, -3.239783e-09, 
    -3.555615e-09, -3.880376e-09, -3.987799e-09, -4.017121e-09, 
    -4.038519e-09, -3.97927e-09, -3.983699e-09, -3.928486e-09, -3.914479e-09, 
    -3.954454e-09,
  -2.978181e-09, -3.165616e-09, -3.25288e-09, -3.359889e-09, -3.764397e-09, 
    -4.315913e-09, -4.475548e-09, -4.466963e-09, -4.357026e-09, 
    -4.321959e-09, -4.231512e-09, -4.041447e-09, -3.88318e-09, -3.7789e-09, 
    -3.777964e-09,
  -3.721628e-09, -4.004878e-09, -4.255086e-09, -4.046065e-09, -4.498262e-09, 
    -4.824073e-09, -4.846346e-09, -4.748666e-09, -4.618213e-09, 
    -4.532833e-09, -4.427764e-09, -4.1837e-09, -4.006803e-09, -3.886337e-09, 
    -3.769366e-09,
  -5.259188e-09, -5.426754e-09, -5.675668e-09, -5.708565e-09, -5.46917e-09, 
    -5.705424e-09, -5.714087e-09, -5.297326e-09, -4.865874e-09, 
    -4.612994e-09, -4.476006e-09, -4.444025e-09, -4.399965e-09, 
    -3.874249e-09, -3.470902e-09,
  -3.155538e-09, -3.261269e-09, -3.299931e-09, -3.399931e-09, -3.56993e-09, 
    -3.691038e-09, -3.76237e-09, -3.763835e-09, -3.779188e-09, -3.782465e-09, 
    -3.802418e-09, -3.924499e-09, -4.089154e-09, -4.272478e-09, -4.492976e-09,
  -2.653279e-09, -2.668407e-09, -2.633767e-09, -2.745603e-09, -2.924256e-09, 
    -3.093225e-09, -3.218702e-09, -3.33324e-09, -3.390959e-09, -3.471677e-09, 
    -3.566297e-09, -3.649897e-09, -3.749674e-09, -3.843614e-09, -3.962393e-09,
  -2.242024e-09, -2.367571e-09, -2.344042e-09, -2.458177e-09, -2.468884e-09, 
    -2.491506e-09, -2.597065e-09, -2.760723e-09, -2.993922e-09, 
    -3.121084e-09, -3.312294e-09, -3.460189e-09, -3.570598e-09, 
    -3.661686e-09, -3.744426e-09,
  -2.122986e-09, -2.116425e-09, -2.225757e-09, -2.364768e-09, -2.385613e-09, 
    -2.354584e-09, -2.391044e-09, -2.49914e-09, -2.63347e-09, -2.766533e-09, 
    -2.927222e-09, -3.074443e-09, -3.173117e-09, -3.265497e-09, -3.372688e-09,
  -2.143158e-09, -2.097676e-09, -2.342308e-09, -2.378961e-09, -2.392126e-09, 
    -2.396757e-09, -2.481172e-09, -2.586905e-09, -2.616799e-09, 
    -2.655554e-09, -2.693357e-09, -2.727653e-09, -2.758246e-09, 
    -2.804468e-09, -2.89593e-09,
  -2.070054e-09, -2.071728e-09, -2.282758e-09, -2.527633e-09, -2.375899e-09, 
    -2.370307e-09, -2.47079e-09, -2.567897e-09, -2.541395e-09, -2.465225e-09, 
    -2.447469e-09, -2.416055e-09, -2.422499e-09, -2.47182e-09, -2.585288e-09,
  -1.96348e-09, -2.111958e-09, -2.125358e-09, -2.774299e-09, -2.748734e-09, 
    -2.524485e-09, -2.675466e-09, -2.665021e-09, -2.568046e-09, 
    -2.427916e-09, -2.324523e-09, -2.250246e-09, -2.206244e-09, 
    -2.311583e-09, -2.44113e-09,
  -1.580874e-09, -2.076543e-09, -2.302539e-09, -2.917296e-09, -2.991724e-09, 
    -2.769502e-09, -2.745921e-09, -2.729217e-09, -2.771085e-09, 
    -2.581698e-09, -2.373378e-09, -2.2862e-09, -2.257539e-09, -2.332575e-09, 
    -2.444908e-09,
  -1.216646e-09, -1.778196e-09, -2.442901e-09, -2.870945e-09, -3.262181e-09, 
    -2.662582e-09, -2.415549e-09, -2.5527e-09, -2.873828e-09, -2.837957e-09, 
    -2.666354e-09, -2.561916e-09, -2.4455e-09, -2.435341e-09, -2.548327e-09,
  -1.951385e-09, -2.25726e-09, -2.484988e-09, -2.788953e-09, -2.763113e-09, 
    -2.152204e-09, -2.246598e-09, -2.545892e-09, -3.077879e-09, 
    -3.156756e-09, -3.028151e-09, -2.789335e-09, -2.635641e-09, 
    -2.619869e-09, -2.79929e-09,
  -3.306555e-09, -3.292259e-09, -3.232535e-09, -3.124929e-09, -3.011076e-09, 
    -2.980696e-09, -3.11647e-09, -3.389801e-09, -3.670386e-09, -3.757218e-09, 
    -4.781026e-09, -5.30809e-09, -5.532786e-09, -5.395335e-09, -5.106909e-09,
  -3.429183e-09, -3.479369e-09, -3.365156e-09, -3.24241e-09, -3.156609e-09, 
    -3.071963e-09, -3.021265e-09, -3.066092e-09, -3.337151e-09, 
    -3.589484e-09, -3.873091e-09, -4.525659e-09, -5.043137e-09, 
    -5.175263e-09, -5.107345e-09,
  -3.63895e-09, -3.523503e-09, -3.417619e-09, -3.391493e-09, -3.346283e-09, 
    -3.264189e-09, -3.200054e-09, -3.092383e-09, -3.136363e-09, 
    -3.297059e-09, -3.543803e-09, -3.872131e-09, -4.488012e-09, 
    -4.938045e-09, -5.099539e-09,
  -3.540807e-09, -3.467413e-09, -3.426174e-09, -3.46542e-09, -3.506245e-09, 
    -3.485696e-09, -3.475054e-09, -3.413184e-09, -3.339035e-09, 
    -3.360969e-09, -3.446235e-09, -3.630308e-09, -3.988098e-09, 
    -4.476929e-09, -4.743738e-09,
  -3.372916e-09, -3.465827e-09, -3.75374e-09, -3.565416e-09, -3.516983e-09, 
    -3.56669e-09, -3.60196e-09, -3.651442e-09, -3.712449e-09, -3.695773e-09, 
    -3.618352e-09, -3.597862e-09, -3.749905e-09, -4.163003e-09, -4.448525e-09,
  -3.349242e-09, -3.45158e-09, -3.786461e-09, -3.999369e-09, -3.607246e-09, 
    -3.325524e-09, -3.342904e-09, -3.618566e-09, -3.788011e-09, 
    -3.907339e-09, -3.90327e-09, -3.779309e-09, -3.703124e-09, -3.82295e-09, 
    -4.119398e-09,
  -3.082628e-09, -3.194661e-09, -3.435283e-09, -3.576042e-09, -3.641279e-09, 
    -3.26715e-09, -2.971053e-09, -3.020476e-09, -3.36026e-09, -3.61059e-09, 
    -3.860606e-09, -3.930131e-09, -3.747291e-09, -3.661855e-09, -3.830126e-09,
  -2.80092e-09, -2.870225e-09, -3.197316e-09, -3.696865e-09, -3.418515e-09, 
    -3.004564e-09, -2.827565e-09, -2.795325e-09, -2.861694e-09, 
    -3.082385e-09, -3.29869e-09, -3.484583e-09, -3.522172e-09, -3.472241e-09, 
    -3.548896e-09,
  -2.620933e-09, -2.569655e-09, -2.991566e-09, -3.487849e-09, -3.540147e-09, 
    -3.540491e-09, -3.07318e-09, -2.603807e-09, -2.46994e-09, -2.650877e-09, 
    -2.909502e-09, -3.114668e-09, -3.388439e-09, -3.415395e-09, -3.484135e-09,
  -2.945344e-09, -2.578703e-09, -2.88615e-09, -3.07742e-09, -4.167118e-09, 
    -3.327002e-09, -2.743159e-09, -2.32983e-09, -2.216185e-09, -2.458701e-09, 
    -2.815578e-09, -3.069585e-09, -3.465699e-09, -3.48893e-09, -3.398771e-09,
  -2.039725e-09, -1.998261e-09, -2.038673e-09, -1.995121e-09, -1.947829e-09, 
    -1.957674e-09, -1.944516e-09, -1.918418e-09, -1.9611e-09, -2.041824e-09, 
    -2.062245e-09, -2.075675e-09, -2.072982e-09, -1.966784e-09, -1.79587e-09,
  -2.283202e-09, -2.159731e-09, -2.115366e-09, -2.062093e-09, -1.986506e-09, 
    -1.984615e-09, -1.939446e-09, -1.801446e-09, -1.75917e-09, -1.890854e-09, 
    -1.961485e-09, -1.969688e-09, -1.95424e-09, -1.856735e-09, -1.613238e-09,
  -2.285304e-09, -2.312305e-09, -2.435091e-09, -2.391582e-09, -2.32689e-09, 
    -2.181128e-09, -1.988117e-09, -1.815569e-09, -1.687385e-09, 
    -1.680705e-09, -1.769154e-09, -1.755408e-09, -1.703968e-09, -1.6442e-09, 
    -1.513393e-09,
  -2.123562e-09, -2.443729e-09, -2.435676e-09, -2.306198e-09, -2.488959e-09, 
    -2.540977e-09, -2.238167e-09, -2.088616e-09, -1.916839e-09, 
    -1.753062e-09, -1.666789e-09, -1.679106e-09, -1.65375e-09, -1.731338e-09, 
    -1.860363e-09,
  -2.361683e-09, -2.39802e-09, -2.435391e-09, -2.580916e-09, -2.580083e-09, 
    -2.808348e-09, -2.686732e-09, -2.309279e-09, -2.044564e-09, 
    -1.768984e-09, -1.612295e-09, -1.61327e-09, -1.632041e-09, -1.707164e-09, 
    -1.944102e-09,
  -2.671593e-09, -2.246518e-09, -2.58473e-09, -3.080577e-09, -2.472482e-09, 
    -2.515628e-09, -2.487012e-09, -2.163208e-09, -1.998875e-09, 
    -1.751693e-09, -1.66459e-09, -1.660118e-09, -1.625274e-09, -1.62696e-09, 
    -1.886568e-09,
  -2.686873e-09, -3.284095e-09, -3.972533e-09, -2.939414e-09, -2.295206e-09, 
    -1.522424e-09, -1.285374e-09, -1.756642e-09, -1.977182e-09, 
    -1.549973e-09, -1.435107e-09, -1.44894e-09, -1.546943e-09, -1.641893e-09, 
    -1.914493e-09,
  -4.22461e-09, -5.946557e-09, -3.380583e-09, -2.439527e-09, -8.522046e-10, 
    6.56255e-11, -1.272375e-09, -1.997765e-09, -1.988511e-09, -1.598589e-09, 
    -1.407052e-09, -1.506554e-09, -1.588791e-09, -1.585029e-09, -1.793741e-09,
  -5.3878e-09, -4.313411e-09, -1.857019e-09, -1.158102e-09, -6.288794e-10, 
    -1.350959e-09, -1.684841e-09, -1.951445e-09, -1.999427e-09, 
    -1.752937e-09, -1.556003e-09, -1.503079e-09, -1.572358e-09, 
    -1.651841e-09, -1.99656e-09,
  -4.053195e-09, -2.991349e-09, -2.220438e-09, -1.962383e-09, -1.880241e-09, 
    -1.574505e-09, -1.576196e-09, -1.692828e-09, -1.765676e-09, 
    -1.844704e-09, -1.615529e-09, -1.673932e-09, -1.948297e-09, -2.14147e-09, 
    -2.716215e-09,
  -2.555096e-09, -2.589148e-09, -2.606908e-09, -2.611684e-09, -2.587206e-09, 
    -2.562085e-09, -2.45698e-09, -2.34365e-09, -2.199797e-09, -1.981456e-09, 
    -1.860697e-09, -1.810035e-09, -1.683593e-09, -1.532175e-09, -1.571102e-09,
  -2.37543e-09, -2.451033e-09, -2.513099e-09, -2.547234e-09, -2.504485e-09, 
    -2.467566e-09, -2.236345e-09, -2.209729e-09, -2.25e-09, -2.238158e-09, 
    -2.168164e-09, -2.152614e-09, -2.237235e-09, -2.246977e-09, -2.18781e-09,
  -2.230901e-09, -2.208039e-09, -2.176022e-09, -2.187805e-09, -2.066485e-09, 
    -1.858434e-09, -2.04331e-09, -2.290471e-09, -2.399276e-09, -2.375179e-09, 
    -2.334932e-09, -2.255149e-09, -2.329039e-09, -2.47281e-09, -2.62225e-09,
  -1.89977e-09, -1.797064e-09, -1.750083e-09, -1.938054e-09, -1.904655e-09, 
    -1.753745e-09, -1.923273e-09, -2.155369e-09, -2.094615e-09, 
    -2.130006e-09, -2.14118e-09, -2.097591e-09, -2.068999e-09, -2.082475e-09, 
    -2.086151e-09,
  -1.75253e-09, -1.579559e-09, -1.725483e-09, -1.814323e-09, -2.02381e-09, 
    -2.251266e-09, -1.856707e-09, -1.659055e-09, -1.83889e-09, -2.085257e-09, 
    -2.153767e-09, -2.034148e-09, -1.943225e-09, -1.85041e-09, -1.603386e-09,
  -1.902769e-09, -1.882511e-09, -2.35297e-09, -2.809152e-09, -2.304468e-09, 
    -1.668779e-09, -1.56514e-09, -1.910041e-09, -1.876761e-09, -1.679192e-09, 
    -1.696904e-09, -1.763317e-09, -1.763301e-09, -1.649516e-09, -1.541952e-09,
  -2.554771e-09, -2.511118e-09, -1.869082e-09, -1.592746e-09, -1.262341e-09, 
    -1.281691e-09, -1.723706e-09, -1.559784e-09, -1.270474e-09, 
    -1.257832e-09, -1.465693e-09, -1.659565e-09, -1.485068e-09, 
    -1.548708e-09, -1.684178e-09,
  -1.621094e-09, -1.477792e-09, -1.204811e-09, -1.08138e-09, -1.492614e-09, 
    -1.479641e-09, -1.074082e-09, -8.764498e-10, -9.135354e-10, 
    -1.140981e-09, -1.261127e-09, -1.237929e-09, -2.064892e-09, 
    -1.708113e-09, -9.306119e-10,
  -5.363697e-10, -7.049131e-10, -1.156518e-09, -1.362205e-09, -1.178824e-09, 
    -7.245658e-10, -6.076452e-10, -7.132817e-10, -8.606493e-10, 
    -8.797332e-10, -1.461423e-09, -2.099575e-09, -1.131496e-09, 
    -8.702417e-10, -1.011683e-09,
  -4.325692e-10, -8.1725e-10, -1.111379e-09, -9.390672e-10, -8.280803e-10, 
    -6.724044e-10, -6.9359e-10, -7.303028e-10, -9.914616e-10, -1.504693e-09, 
    -1.739954e-09, -1.093189e-09, -9.908864e-10, -1.346412e-09, -1.63288e-09,
  -2.222755e-09, -2.274487e-09, -2.335517e-09, -2.401862e-09, -2.536918e-09, 
    -2.782205e-09, -3.15885e-09, -3.632773e-09, -4.149361e-09, -4.664565e-09, 
    -5.181763e-09, -5.6123e-09, -6.03733e-09, -6.335912e-09, -6.662908e-09,
  -2.176274e-09, -2.258468e-09, -2.319705e-09, -2.361009e-09, -2.409532e-09, 
    -2.490488e-09, -2.630207e-09, -2.837864e-09, -3.112045e-09, 
    -3.405332e-09, -3.719066e-09, -4.028483e-09, -4.328375e-09, 
    -4.628866e-09, -4.892773e-09,
  -2.114237e-09, -2.166877e-09, -2.213885e-09, -2.273157e-09, -2.297481e-09, 
    -2.289055e-09, -2.321879e-09, -2.378833e-09, -2.454038e-09, 
    -2.574952e-09, -2.738141e-09, -2.905262e-09, -3.083189e-09, 
    -3.285557e-09, -3.543519e-09,
  -2.023377e-09, -2.055899e-09, -2.089863e-09, -2.124556e-09, -2.137294e-09, 
    -2.146622e-09, -2.135457e-09, -2.117497e-09, -2.0656e-09, -2.046451e-09, 
    -2.098636e-09, -2.172802e-09, -2.268089e-09, -2.392914e-09, -2.62134e-09,
  -1.908237e-09, -1.948429e-09, -1.968281e-09, -1.999778e-09, -2.019071e-09, 
    -2.007901e-09, -1.988557e-09, -1.973945e-09, -1.968118e-09, 
    -1.947356e-09, -1.945116e-09, -2.023925e-09, -2.162539e-09, 
    -2.309331e-09, -2.411899e-09,
  -1.828552e-09, -1.891897e-09, -1.8814e-09, -1.89677e-09, -1.936588e-09, 
    -2.020855e-09, -2.043351e-09, -2.073689e-09, -2.152311e-09, 
    -2.220813e-09, -2.24188e-09, -2.243388e-09, -2.254444e-09, -2.251862e-09, 
    -2.243074e-09,
  -1.597353e-09, -1.822399e-09, -1.820934e-09, -1.817172e-09, -1.882417e-09, 
    -1.966241e-09, -2.063619e-09, -2.1097e-09, -2.108463e-09, -2.123844e-09, 
    -2.147351e-09, -2.172639e-09, -2.163033e-09, -2.158106e-09, -2.146608e-09,
  -1.295734e-09, -1.602509e-09, -1.75945e-09, -1.727752e-09, -1.789508e-09, 
    -1.861273e-09, -1.959834e-09, -2.054191e-09, -2.067748e-09, 
    -2.036925e-09, -2.026758e-09, -2.048591e-09, -2.101232e-09, 
    -2.134552e-09, -2.100674e-09,
  -1.152302e-09, -1.2393e-09, -1.484013e-09, -1.590765e-09, -1.695758e-09, 
    -1.834033e-09, -1.909008e-09, -1.997768e-09, -2.048618e-09, 
    -2.010308e-09, -1.976795e-09, -2.024132e-09, -1.991501e-09, 
    -1.920543e-09, -1.846077e-09,
  -1.014046e-09, -8.864668e-10, -9.707468e-10, -1.096862e-09, -1.322697e-09, 
    -1.682733e-09, -1.869052e-09, -1.895157e-09, -1.96161e-09, -1.984523e-09, 
    -1.977861e-09, -1.920304e-09, -1.810909e-09, -1.794417e-09, -1.751496e-09,
  -1.106868e-08, -1.143916e-08, -1.179993e-08, -1.200983e-08, -1.21454e-08, 
    -1.219509e-08, -1.198922e-08, -1.163846e-08, -1.118325e-08, 
    -1.070058e-08, -1.048104e-08, -1.05702e-08, -1.061973e-08, -1.046248e-08, 
    -1.011149e-08,
  -9.381151e-09, -9.742989e-09, -1.006262e-08, -1.033682e-08, -1.042822e-08, 
    -1.031985e-08, -1.00522e-08, -9.720798e-09, -9.286033e-09, -8.732184e-09, 
    -8.314907e-09, -8.004077e-09, -7.772527e-09, -7.393611e-09, -7.056633e-09,
  -7.639171e-09, -8.03846e-09, -8.28938e-09, -8.367515e-09, -8.335937e-09, 
    -8.267391e-09, -8.029858e-09, -7.744128e-09, -7.474632e-09, -6.91472e-09, 
    -6.4536e-09, -6.018749e-09, -5.661638e-09, -5.58558e-09, -5.67924e-09,
  -5.927781e-09, -6.3549e-09, -6.574364e-09, -6.696884e-09, -6.768308e-09, 
    -6.77454e-09, -6.699771e-09, -6.5324e-09, -6.273361e-09, -5.951911e-09, 
    -5.618057e-09, -5.289202e-09, -5.254234e-09, -5.47793e-09, -5.760196e-09,
  -4.18726e-09, -4.508204e-09, -4.83289e-09, -4.995239e-09, -5.182141e-09, 
    -5.292947e-09, -5.318822e-09, -5.204376e-09, -5.015852e-09, -4.70715e-09, 
    -4.478292e-09, -4.231009e-09, -4.213172e-09, -4.376774e-09, -4.56386e-09,
  -2.775967e-09, -3.102771e-09, -3.370113e-09, -3.626087e-09, -3.791688e-09, 
    -3.911488e-09, -3.857002e-09, -3.862862e-09, -3.745811e-09, 
    -3.573329e-09, -3.381352e-09, -3.190863e-09, -3.158199e-09, 
    -3.202225e-09, -3.273728e-09,
  -1.77296e-09, -2.00844e-09, -2.261348e-09, -2.468413e-09, -2.65733e-09, 
    -2.751601e-09, -2.807184e-09, -2.834249e-09, -2.839108e-09, 
    -2.725558e-09, -2.508544e-09, -2.305931e-09, -2.11894e-09, -2.01797e-09, 
    -1.910514e-09,
  -1.025773e-09, -1.203003e-09, -1.430049e-09, -1.56121e-09, -1.697248e-09, 
    -1.772524e-09, -1.778792e-09, -1.783609e-09, -1.850104e-09, 
    -1.831329e-09, -1.722755e-09, -1.628763e-09, -1.546866e-09, 
    -1.413928e-09, -1.272418e-09,
  -2.678949e-10, -4.815426e-10, -7.213425e-10, -9.383385e-10, -1.113843e-09, 
    -1.215771e-09, -1.248468e-09, -1.279537e-09, -1.340078e-09, 
    -1.346243e-09, -1.283384e-09, -1.240059e-09, -1.25374e-09, -1.251819e-09, 
    -1.241783e-09,
  1.371838e-10, -2.001673e-11, -1.911638e-10, -4.57793e-10, -6.034637e-10, 
    -7.217499e-10, -8.441111e-10, -9.80269e-10, -1.067311e-09, -1.224326e-09, 
    -1.296699e-09, -1.376957e-09, -1.48936e-09, -1.583639e-09, -1.658324e-09,
  -8.744129e-09, -9.434501e-09, -1.025197e-08, -1.116324e-08, -1.198188e-08, 
    -1.293902e-08, -1.352227e-08, -1.411864e-08, -1.468765e-08, 
    -1.529631e-08, -1.598183e-08, -1.677494e-08, -1.758032e-08, -1.83667e-08, 
    -1.908472e-08,
  -8.228923e-09, -9.201488e-09, -1.000644e-08, -1.093716e-08, -1.171427e-08, 
    -1.259397e-08, -1.347759e-08, -1.414434e-08, -1.481013e-08, 
    -1.536304e-08, -1.59893e-08, -1.661693e-08, -1.735854e-08, -1.81233e-08, 
    -1.873645e-08,
  -7.880043e-09, -8.807635e-09, -9.684801e-09, -1.054719e-08, -1.135596e-08, 
    -1.207135e-08, -1.302671e-08, -1.389153e-08, -1.447731e-08, 
    -1.516609e-08, -1.581839e-08, -1.645532e-08, -1.713491e-08, 
    -1.770463e-08, -1.820128e-08,
  -7.764823e-09, -8.500386e-09, -9.345624e-09, -1.021219e-08, -1.106961e-08, 
    -1.183418e-08, -1.261584e-08, -1.345722e-08, -1.410556e-08, 
    -1.471331e-08, -1.54639e-08, -1.61428e-08, -1.681958e-08, -1.739556e-08, 
    -1.78124e-08,
  -7.413255e-09, -8.170671e-09, -8.916439e-09, -9.728217e-09, -1.053806e-08, 
    -1.145034e-08, -1.231424e-08, -1.305892e-08, -1.365965e-08, 
    -1.421682e-08, -1.48997e-08, -1.557064e-08, -1.62283e-08, -1.686359e-08, 
    -1.738238e-08,
  -7.233186e-09, -7.805622e-09, -8.523875e-09, -9.250883e-09, -9.959434e-09, 
    -1.074865e-08, -1.153827e-08, -1.2389e-08, -1.291042e-08, -1.351304e-08, 
    -1.420667e-08, -1.480377e-08, -1.531043e-08, -1.583022e-08, -1.63056e-08,
  -6.885642e-09, -7.475679e-09, -8.151507e-09, -8.808247e-09, -9.389215e-09, 
    -1.004962e-08, -1.073477e-08, -1.155543e-08, -1.218958e-08, 
    -1.281179e-08, -1.351368e-08, -1.411993e-08, -1.449806e-08, 
    -1.484904e-08, -1.497923e-08,
  -6.549756e-09, -7.117165e-09, -7.740804e-09, -8.405256e-09, -8.877549e-09, 
    -9.364084e-09, -9.81689e-09, -1.056785e-08, -1.10269e-08, -1.158709e-08, 
    -1.215622e-08, -1.275637e-08, -1.313376e-08, -1.349239e-08, -1.375383e-08,
  -6.119833e-09, -6.665098e-09, -7.366682e-09, -8.108078e-09, -8.676238e-09, 
    -9.065485e-09, -9.335353e-09, -9.802525e-09, -1.004814e-08, -1.02807e-08, 
    -1.05534e-08, -1.102662e-08, -1.1417e-08, -1.170889e-08, -1.201553e-08,
  -5.301657e-09, -5.815664e-09, -6.426338e-09, -7.310535e-09, -7.920582e-09, 
    -8.427503e-09, -8.536963e-09, -8.831952e-09, -8.89201e-09, -8.842673e-09, 
    -8.951307e-09, -9.11587e-09, -9.288788e-09, -9.526016e-09, -9.713454e-09,
  -1.11465e-09, -1.17347e-09, -1.348765e-09, -1.505552e-09, -1.68157e-09, 
    -1.858276e-09, -2.122651e-09, -2.339664e-09, -2.591924e-09, 
    -2.886427e-09, -3.201635e-09, -3.533521e-09, -3.905944e-09, 
    -4.384628e-09, -4.880629e-09,
  -1.164447e-09, -1.194488e-09, -1.287971e-09, -1.398058e-09, -1.545218e-09, 
    -1.67933e-09, -1.89109e-09, -2.126468e-09, -2.411304e-09, -2.740092e-09, 
    -3.037588e-09, -3.345499e-09, -3.706026e-09, -4.107676e-09, -4.566905e-09,
  -1.260514e-09, -1.325827e-09, -1.35476e-09, -1.398035e-09, -1.464932e-09, 
    -1.577799e-09, -1.746312e-09, -1.986403e-09, -2.257843e-09, 
    -2.557212e-09, -2.853004e-09, -3.143785e-09, -3.482177e-09, 
    -3.873624e-09, -4.324726e-09,
  -1.417853e-09, -1.495419e-09, -1.544125e-09, -1.572732e-09, -1.544008e-09, 
    -1.59336e-09, -1.714595e-09, -1.901109e-09, -2.161128e-09, -2.42975e-09, 
    -2.677811e-09, -2.950739e-09, -3.304455e-09, -3.702313e-09, -4.1565e-09,
  -1.560085e-09, -1.625806e-09, -1.691541e-09, -1.767023e-09, -1.754229e-09, 
    -1.754954e-09, -1.80787e-09, -1.937176e-09, -2.133888e-09, -2.346484e-09, 
    -2.591963e-09, -2.843173e-09, -3.170895e-09, -3.60683e-09, -4.061067e-09,
  -1.662653e-09, -1.758743e-09, -1.803901e-09, -1.85478e-09, -1.907732e-09, 
    -1.952618e-09, -2.02205e-09, -2.083747e-09, -2.198323e-09, -2.354118e-09, 
    -2.569975e-09, -2.85517e-09, -3.200155e-09, -3.585179e-09, -4.040738e-09,
  -1.775889e-09, -1.858165e-09, -1.955067e-09, -2.017472e-09, -2.068972e-09, 
    -2.139258e-09, -2.242951e-09, -2.303656e-09, -2.405817e-09, 
    -2.508928e-09, -2.70343e-09, -2.983388e-09, -3.304935e-09, -3.696667e-09, 
    -4.127886e-09,
  -2.052774e-09, -2.09269e-09, -2.116962e-09, -2.201648e-09, -2.317022e-09, 
    -2.398075e-09, -2.496493e-09, -2.518203e-09, -2.612625e-09, 
    -2.765903e-09, -2.977731e-09, -3.212721e-09, -3.493358e-09, 
    -3.855521e-09, -4.267451e-09,
  -2.423783e-09, -2.497151e-09, -2.513099e-09, -2.576855e-09, -2.666716e-09, 
    -2.713471e-09, -2.859748e-09, -2.840947e-09, -2.968239e-09, 
    -3.135489e-09, -3.371555e-09, -3.547797e-09, -3.765916e-09, -4.11486e-09, 
    -4.559644e-09,
  -3.179063e-09, -3.12928e-09, -3.185228e-09, -3.18395e-09, -3.237868e-09, 
    -3.287947e-09, -3.224189e-09, -3.239641e-09, -3.348505e-09, 
    -3.487394e-09, -3.724191e-09, -3.977793e-09, -4.249599e-09, 
    -4.550919e-09, -4.944307e-09,
  -1.491467e-09, -1.423364e-09, -1.329277e-09, -1.23785e-09, -1.191517e-09, 
    -1.180943e-09, -1.218759e-09, -1.274837e-09, -1.394667e-09, 
    -1.555649e-09, -1.762253e-09, -1.986359e-09, -2.205697e-09, 
    -2.416345e-09, -2.65285e-09,
  -1.73715e-09, -1.677129e-09, -1.563274e-09, -1.468263e-09, -1.382941e-09, 
    -1.316615e-09, -1.286056e-09, -1.285788e-09, -1.30458e-09, -1.365903e-09, 
    -1.464785e-09, -1.593672e-09, -1.748869e-09, -1.916598e-09, -2.128185e-09,
  -1.982118e-09, -1.827596e-09, -1.627132e-09, -1.489617e-09, -1.443368e-09, 
    -1.426902e-09, -1.402519e-09, -1.381597e-09, -1.372118e-09, 
    -1.370932e-09, -1.40327e-09, -1.434909e-09, -1.502472e-09, -1.585344e-09, 
    -1.693997e-09,
  -2.043846e-09, -1.828141e-09, -1.573006e-09, -1.459211e-09, -1.388928e-09, 
    -1.372362e-09, -1.395414e-09, -1.421609e-09, -1.443314e-09, 
    -1.440566e-09, -1.454706e-09, -1.471692e-09, -1.48682e-09, -1.494973e-09, 
    -1.530015e-09,
  -1.978962e-09, -1.715734e-09, -1.60003e-09, -1.530464e-09, -1.442398e-09, 
    -1.390194e-09, -1.37262e-09, -1.39446e-09, -1.430366e-09, -1.482587e-09, 
    -1.488361e-09, -1.483165e-09, -1.481692e-09, -1.49915e-09, -1.480216e-09,
  -1.946354e-09, -1.760641e-09, -1.720201e-09, -1.665469e-09, -1.600813e-09, 
    -1.531252e-09, -1.448337e-09, -1.401312e-09, -1.391505e-09, 
    -1.420864e-09, -1.483899e-09, -1.53248e-09, -1.495018e-09, -1.46836e-09, 
    -1.458469e-09,
  -2.061849e-09, -1.951554e-09, -1.885494e-09, -1.823068e-09, -1.750725e-09, 
    -1.648407e-09, -1.549686e-09, -1.459052e-09, -1.415423e-09, 
    -1.404117e-09, -1.416891e-09, -1.483786e-09, -1.55165e-09, -1.53689e-09, 
    -1.48189e-09,
  -2.233616e-09, -2.145286e-09, -2.081869e-09, -1.903217e-09, -1.745575e-09, 
    -1.618034e-09, -1.497972e-09, -1.414623e-09, -1.369536e-09, 
    -1.374019e-09, -1.399934e-09, -1.42699e-09, -1.472451e-09, -1.525896e-09, 
    -1.559602e-09,
  -2.158134e-09, -2.057439e-09, -1.93557e-09, -1.810281e-09, -1.736774e-09, 
    -1.57706e-09, -1.425064e-09, -1.312136e-09, -1.263014e-09, -1.264972e-09, 
    -1.324252e-09, -1.416457e-09, -1.496473e-09, -1.549257e-09, -1.612454e-09,
  -2.315578e-09, -2.0837e-09, -1.90033e-09, -1.686461e-09, -1.664235e-09, 
    -1.649538e-09, -1.47533e-09, -1.329799e-09, -1.212664e-09, -1.173608e-09, 
    -1.202306e-09, -1.298185e-09, -1.428039e-09, -1.543448e-09, -1.617176e-09,
  -2.269967e-09, -2.396084e-09, -2.47126e-09, -2.543932e-09, -2.59953e-09, 
    -2.601684e-09, -2.56444e-09, -2.530852e-09, -2.504492e-09, -2.525367e-09, 
    -2.57561e-09, -2.61637e-09, -2.668155e-09, -2.724093e-09, -2.753375e-09,
  -1.650025e-09, -1.788869e-09, -1.824452e-09, -1.899948e-09, -1.990595e-09, 
    -2.078642e-09, -2.109541e-09, -2.214032e-09, -2.298717e-09, 
    -2.368041e-09, -2.427731e-09, -2.444604e-09, -2.469979e-09, 
    -2.494212e-09, -2.521716e-09,
  -1.028327e-09, -1.123324e-09, -1.144501e-09, -1.203518e-09, -1.237838e-09, 
    -1.325176e-09, -1.441397e-09, -1.634381e-09, -1.842471e-09, 
    -2.056823e-09, -2.199861e-09, -2.325886e-09, -2.410692e-09, 
    -2.470888e-09, -2.505849e-09,
  -6.075835e-10, -6.597185e-10, -6.656306e-10, -6.591284e-10, -7.166843e-10, 
    -8.168456e-10, -9.568063e-10, -1.135828e-09, -1.361674e-09, 
    -1.601942e-09, -1.835117e-09, -2.060473e-09, -2.237624e-09, 
    -2.351825e-09, -2.416111e-09,
  -4.440723e-10, -5.17678e-10, -6.288979e-10, -7.265889e-10, -7.747561e-10, 
    -7.411658e-10, -7.954126e-10, -9.073871e-10, -1.062556e-09, 
    -1.237145e-09, -1.412877e-09, -1.601722e-09, -1.784534e-09, 
    -1.972807e-09, -2.138614e-09,
  -4.612622e-10, -4.632212e-10, -5.993601e-10, -8.335813e-10, -1.018723e-09, 
    -1.203343e-09, -1.282443e-09, -1.244489e-09, -1.259607e-09, 
    -1.311867e-09, -1.369705e-09, -1.431166e-09, -1.526715e-09, 
    -1.652556e-09, -1.784384e-09,
  -6.496384e-10, -6.201064e-10, -7.602853e-10, -9.456094e-10, -1.050949e-09, 
    -1.1644e-09, -1.287921e-09, -1.371225e-09, -1.407815e-09, -1.45844e-09, 
    -1.499595e-09, -1.52008e-09, -1.528863e-09, -1.554264e-09, -1.586893e-09,
  -4.506292e-10, -4.63082e-10, -7.035515e-10, -1.04867e-09, -1.167113e-09, 
    -1.348657e-09, -1.427653e-09, -1.451016e-09, -1.466717e-09, 
    -1.547586e-09, -1.628819e-09, -1.682957e-09, -1.657092e-09, 
    -1.589531e-09, -1.533684e-09,
  -6.330184e-10, -7.005035e-10, -9.111387e-10, -1.116434e-09, -1.29384e-09, 
    -1.379973e-09, -1.38467e-09, -1.435519e-09, -1.51147e-09, -1.528002e-09, 
    -1.588323e-09, -1.613146e-09, -1.608904e-09, -1.557618e-09, -1.503082e-09,
  -8.830852e-10, -8.086389e-10, -1.037173e-09, -1.015313e-09, -1.024105e-09, 
    -1.058209e-09, -1.173944e-09, -1.238068e-09, -1.368139e-09, 
    -1.460089e-09, -1.50855e-09, -1.525449e-09, -1.476051e-09, -1.43764e-09, 
    -1.415678e-09,
  -4.46526e-09, -4.97096e-09, -5.495478e-09, -6.034491e-09, -6.50091e-09, 
    -6.801701e-09, -6.946362e-09, -6.949346e-09, -6.918773e-09, 
    -6.946534e-09, -6.985087e-09, -7.156838e-09, -7.502917e-09, -8.05863e-09, 
    -8.763252e-09,
  -2.68258e-09, -3.041821e-09, -3.425658e-09, -3.817352e-09, -4.14211e-09, 
    -4.409411e-09, -4.570742e-09, -4.640915e-09, -4.607595e-09, 
    -4.534919e-09, -4.537438e-09, -4.545967e-09, -4.627041e-09, 
    -4.709087e-09, -4.930385e-09,
  -1.458801e-09, -1.70586e-09, -1.950742e-09, -2.227786e-09, -2.485823e-09, 
    -2.739201e-09, -2.951359e-09, -3.10607e-09, -3.160987e-09, -3.166502e-09, 
    -3.141981e-09, -3.105927e-09, -3.059073e-09, -3.039419e-09, -3.070616e-09,
  -8.481388e-10, -9.459692e-10, -1.075019e-09, -1.213855e-09, -1.372284e-09, 
    -1.512279e-09, -1.669694e-09, -1.846272e-09, -2.008312e-09, 
    -2.125399e-09, -2.158322e-09, -2.062243e-09, -1.950095e-09, 
    -1.854151e-09, -1.919241e-09,
  -6.399226e-10, -6.922589e-10, -7.127013e-10, -7.49163e-10, -7.888798e-10, 
    -9.171713e-10, -1.032298e-09, -1.163042e-09, -1.239269e-09, 
    -1.265965e-09, -1.31579e-09, -1.371676e-09, -1.430008e-09, -1.515087e-09, 
    -1.629566e-09,
  -5.790295e-10, -5.663784e-10, -5.675382e-10, -4.308562e-10, -4.360505e-10, 
    -4.123605e-10, -4.38331e-10, -3.416866e-10, -4.742582e-10, -5.592284e-10, 
    -7.093408e-10, -6.941325e-10, -7.493238e-10, -8.896372e-10, -1.064548e-09,
  -5.722031e-10, -5.553778e-10, -4.881198e-10, -5.057865e-10, -4.834233e-10, 
    -2.535708e-10, -3.239568e-13, 2.384325e-10, 2.819483e-10, -1.346262e-12, 
    -2.123627e-10, -3.587256e-10, -5.11892e-10, -5.846199e-10, -6.11617e-10,
  -5.656129e-10, -6.114975e-10, -6.128967e-10, -6.586091e-10, -4.639477e-10, 
    -8.713901e-10, -7.613372e-10, -4.950702e-10, -2.302001e-10, 
    -3.192934e-10, -3.943098e-10, -4.050838e-10, -4.23308e-10, -4.957634e-10, 
    -4.755478e-10,
  -3.749456e-10, -4.710682e-10, -4.180454e-10, -4.533456e-10, -4.966783e-10, 
    -7.89941e-10, -7.004404e-10, -5.539087e-10, -5.004144e-10, -4.299543e-10, 
    -4.484476e-10, -3.818376e-10, -3.14214e-10, -2.334013e-10, -3.354121e-10,
  -2.227475e-10, -2.635347e-10, -3.515367e-10, -4.528094e-10, -4.545966e-10, 
    -4.506231e-10, -5.543744e-10, -5.655651e-10, -5.985316e-10, 
    -6.638791e-10, -4.799613e-10, -3.627758e-10, -3.144899e-10, 
    -3.201716e-10, -3.003337e-10,
  -9.736566e-09, -1.12937e-08, -1.251612e-08, -1.295291e-08, -1.400067e-08, 
    -1.556434e-08, -1.704017e-08, -1.786094e-08, -1.840601e-08, -1.83298e-08, 
    -1.867472e-08, -1.865918e-08, -1.940845e-08, -1.923718e-08, -1.606188e-08,
  -8.419026e-09, -9.310272e-09, -1.075566e-08, -1.186733e-08, -1.262258e-08, 
    -1.359989e-08, -1.497313e-08, -1.635155e-08, -1.737552e-08, 
    -1.829251e-08, -1.804978e-08, -1.87903e-08, -1.829143e-08, -1.596387e-08, 
    -1.204818e-08,
  -6.906658e-09, -8.070866e-09, -9.007429e-09, -1.020593e-08, -1.118274e-08, 
    -1.205548e-08, -1.30441e-08, -1.427161e-08, -1.50962e-08, -1.633992e-08, 
    -1.618812e-08, -1.641522e-08, -1.540819e-08, -1.293769e-08, -9.638477e-09,
  -5.162565e-09, -6.491826e-09, -7.734761e-09, -8.774458e-09, -9.836271e-09, 
    -1.055653e-08, -1.127491e-08, -1.236422e-08, -1.292154e-08, 
    -1.394476e-08, -1.414949e-08, -1.41715e-08, -1.349169e-08, -1.131389e-08, 
    -8.841996e-09,
  -3.360253e-09, -4.401467e-09, -5.708318e-09, -6.991869e-09, -8.22519e-09, 
    -9.316596e-09, -9.846029e-09, -1.05545e-08, -1.127786e-08, -1.177981e-08, 
    -1.227655e-08, -1.263969e-08, -1.187012e-08, -1.022345e-08, -8.406645e-09,
  -2.48311e-09, -3.006166e-09, -3.821718e-09, -4.883856e-09, -6.020448e-09, 
    -7.229118e-09, -8.246783e-09, -8.852023e-09, -9.393611e-09, 
    -9.962484e-09, -1.033494e-08, -1.067797e-08, -1.056443e-08, 
    -9.404521e-09, -8.983838e-09,
  -1.809932e-09, -2.207763e-09, -2.626672e-09, -3.350754e-09, -4.168764e-09, 
    -5.135093e-09, -6.152353e-09, -7.00815e-09, -7.682899e-09, -8.099443e-09, 
    -8.60549e-09, -8.449385e-09, -9.167488e-09, -9.921415e-09, -9.854606e-09,
  -1.244188e-09, -1.61624e-09, -1.902365e-09, -2.305737e-09, -2.862434e-09, 
    -3.496812e-09, -4.307789e-09, -5.166005e-09, -5.789509e-09, 
    -6.400048e-09, -6.789533e-09, -6.996839e-09, -6.924832e-09, 
    -7.067764e-09, -6.938448e-09,
  -8.96504e-10, -9.977333e-10, -1.303259e-09, -1.582661e-09, -1.967879e-09, 
    -2.366994e-09, -2.799551e-09, -3.414484e-09, -4.018216e-09, 
    -4.572479e-09, -5.012219e-09, -5.316014e-09, -5.402148e-09, 
    -5.316177e-09, -5.202257e-09,
  -8.622841e-10, -8.055488e-10, -8.501815e-10, -1.030863e-09, -1.249811e-09, 
    -1.630338e-09, -1.894692e-09, -2.250565e-09, -2.6507e-09, -3.026239e-09, 
    -3.360461e-09, -3.630807e-09, -3.822686e-09, -3.819644e-09, -3.733603e-09,
  -7.978847e-09, -8.408821e-09, -8.993651e-09, -9.60984e-09, -1.007844e-08, 
    -1.04325e-08, -1.090587e-08, -1.212862e-08, -1.414892e-08, -1.65153e-08, 
    -1.864777e-08, -2.0124e-08, -2.111634e-08, -2.160923e-08, -2.369554e-08,
  -7.465455e-09, -7.96765e-09, -8.432562e-09, -9.006958e-09, -9.682782e-09, 
    -9.993186e-09, -1.039201e-08, -1.084183e-08, -1.188102e-08, 
    -1.363466e-08, -1.598764e-08, -1.78338e-08, -2.009971e-08, -2.082476e-08, 
    -2.284333e-08,
  -6.949513e-09, -7.547533e-09, -7.993298e-09, -8.393534e-09, -9.087158e-09, 
    -9.601181e-09, -9.947367e-09, -1.028524e-08, -1.077553e-08, 
    -1.161389e-08, -1.326015e-08, -1.502623e-08, -1.75621e-08, -1.911319e-08, 
    -2.127169e-08,
  -6.265503e-09, -7.004754e-09, -7.612194e-09, -7.970858e-09, -8.478262e-09, 
    -9.073544e-09, -9.540345e-09, -9.851372e-09, -1.026323e-08, 
    -1.077176e-08, -1.153807e-08, -1.266079e-08, -1.433497e-08, 
    -1.597505e-08, -1.843495e-08,
  -5.583325e-09, -6.382751e-09, -7.140029e-09, -7.542257e-09, -8.004768e-09, 
    -8.50128e-09, -9.048891e-09, -9.439777e-09, -9.71577e-09, -1.016464e-08, 
    -1.070682e-08, -1.151083e-08, -1.245758e-08, -1.359058e-08, -1.50344e-08,
  -4.626294e-09, -5.683824e-09, -6.532793e-09, -7.182778e-09, -7.553118e-09, 
    -8.023932e-09, -8.482844e-09, -9.064243e-09, -9.386778e-09, 
    -9.660032e-09, -9.982575e-09, -1.059191e-08, -1.114683e-08, 
    -1.212506e-08, -1.279424e-08,
  -3.446344e-09, -4.809364e-09, -5.681405e-09, -6.594216e-09, -7.141203e-09, 
    -7.597031e-09, -7.986525e-09, -8.437337e-09, -8.967286e-09, 
    -9.289331e-09, -9.5748e-09, -9.903187e-09, -1.02828e-08, -1.075079e-08, 
    -1.137777e-08,
  -2.053937e-09, -3.613921e-09, -4.848239e-09, -5.73664e-09, -6.478686e-09, 
    -7.088127e-09, -7.584284e-09, -8.021511e-09, -8.361059e-09, -8.74901e-09, 
    -9.05224e-09, -9.34381e-09, -9.605511e-09, -9.910878e-09, -1.026548e-08,
  -1.651948e-09, -2.237895e-09, -3.666544e-09, -4.895238e-09, -5.793672e-09, 
    -6.363357e-09, -6.855952e-09, -7.3686e-09, -7.857357e-09, -8.280946e-09, 
    -8.616861e-09, -8.924932e-09, -9.154364e-09, -9.401395e-09, -9.598637e-09,
  -1.693481e-09, -1.715777e-09, -2.296443e-09, -3.614122e-09, -4.766414e-09, 
    -5.836172e-09, -6.368821e-09, -6.736935e-09, -7.040259e-09, 
    -7.453655e-09, -7.766143e-09, -8.216626e-09, -8.419545e-09, 
    -8.725782e-09, -8.847074e-09,
  -5.937718e-09, -7.149047e-09, -8.383024e-09, -9.462859e-09, -1.079028e-08, 
    -1.204851e-08, -1.268344e-08, -1.325957e-08, -1.428702e-08, 
    -1.594174e-08, -1.745392e-08, -1.903197e-08, -2.046053e-08, 
    -2.150372e-08, -2.237213e-08,
  -4.949606e-09, -6.422998e-09, -7.605853e-09, -8.749857e-09, -9.905819e-09, 
    -1.13503e-08, -1.249456e-08, -1.30136e-08, -1.350364e-08, -1.444983e-08, 
    -1.580092e-08, -1.708257e-08, -1.868865e-08, -2.027505e-08, -2.152004e-08,
  -4.311916e-09, -5.678328e-09, -6.942666e-09, -8.049268e-09, -9.142408e-09, 
    -1.048395e-08, -1.187187e-08, -1.282865e-08, -1.322114e-08, 
    -1.361175e-08, -1.439646e-08, -1.539267e-08, -1.66417e-08, -1.816175e-08, 
    -1.973081e-08,
  -3.906097e-09, -4.919257e-09, -6.293058e-09, -7.431649e-09, -8.518377e-09, 
    -9.767842e-09, -1.114493e-08, -1.239231e-08, -1.311222e-08, -1.32467e-08, 
    -1.35539e-08, -1.401184e-08, -1.477968e-08, -1.575996e-08, -1.698112e-08,
  -3.750243e-09, -4.472756e-09, -5.635171e-09, -6.861378e-09, -7.981885e-09, 
    -9.163657e-09, -1.041767e-08, -1.174714e-08, -1.284076e-08, -1.30812e-08, 
    -1.30825e-08, -1.312144e-08, -1.345036e-08, -1.395923e-08, -1.467481e-08,
  -3.650053e-09, -4.226993e-09, -5.144696e-09, -6.302349e-09, -7.428234e-09, 
    -8.702159e-09, -9.948318e-09, -1.107751e-08, -1.228964e-08, 
    -1.300275e-08, -1.298498e-08, -1.275498e-08, -1.261973e-08, 
    -1.270445e-08, -1.287809e-08,
  -3.494712e-09, -4.092845e-09, -4.787885e-09, -5.867381e-09, -6.97084e-09, 
    -8.027845e-09, -9.391835e-09, -1.061004e-08, -1.166107e-08, 
    -1.248291e-08, -1.276131e-08, -1.259389e-08, -1.241129e-08, 
    -1.222174e-08, -1.210776e-08,
  -3.333928e-09, -3.870199e-09, -4.471314e-09, -5.39497e-09, -6.531376e-09, 
    -7.64854e-09, -8.923283e-09, -1.013268e-08, -1.123564e-08, -1.212234e-08, 
    -1.251271e-08, -1.239235e-08, -1.2173e-08, -1.194551e-08, -1.176331e-08,
  -3.215626e-09, -3.643723e-09, -4.267795e-09, -4.965973e-09, -5.99275e-09, 
    -6.999529e-09, -8.435264e-09, -9.752909e-09, -1.072936e-08, 
    -1.156218e-08, -1.209772e-08, -1.220775e-08, -1.208748e-08, 
    -1.185066e-08, -1.163639e-08,
  -2.971465e-09, -3.543255e-09, -4.041019e-09, -4.623151e-09, -5.626011e-09, 
    -6.64261e-09, -7.836475e-09, -9.349391e-09, -1.062639e-08, -1.140409e-08, 
    -1.173981e-08, -1.18487e-08, -1.178499e-08, -1.157192e-08, -1.13785e-08,
  -4.253027e-09, -4.775387e-09, -5.464732e-09, -6.346916e-09, -7.279609e-09, 
    -8.634008e-09, -9.799503e-09, -1.121337e-08, -1.287015e-08, 
    -1.405215e-08, -1.490882e-08, -1.556649e-08, -1.600482e-08, 
    -1.629459e-08, -1.657815e-08,
  -3.667676e-09, -4.00153e-09, -4.484609e-09, -5.225529e-09, -5.988601e-09, 
    -7.04184e-09, -8.158028e-09, -9.480706e-09, -1.111738e-08, -1.277168e-08, 
    -1.422025e-08, -1.500446e-08, -1.559381e-08, -1.596909e-08, -1.616474e-08,
  -3.365328e-09, -3.537462e-09, -3.866799e-09, -4.302438e-09, -4.922058e-09, 
    -5.7351e-09, -6.745276e-09, -7.947887e-09, -9.476007e-09, -1.110713e-08, 
    -1.283725e-08, -1.418396e-08, -1.498037e-08, -1.555729e-08, -1.589264e-08,
  -3.191979e-09, -3.232036e-09, -3.537628e-09, -3.869049e-09, -4.217395e-09, 
    -4.800571e-09, -5.636863e-09, -6.694115e-09, -8.023314e-09, 
    -9.656756e-09, -1.132411e-08, -1.286269e-08, -1.420553e-08, 
    -1.491516e-08, -1.537803e-08,
  -2.944603e-09, -2.984277e-09, -3.315126e-09, -3.630679e-09, -3.901055e-09, 
    -4.232129e-09, -4.821447e-09, -5.696542e-09, -6.842698e-09, 
    -8.196043e-09, -9.906834e-09, -1.151097e-08, -1.30269e-08, -1.415845e-08, 
    -1.506158e-08,
  -2.822387e-09, -2.750117e-09, -3.057749e-09, -3.443787e-09, -3.728869e-09, 
    -3.999574e-09, -4.372195e-09, -4.946168e-09, -5.957646e-09, 
    -7.231315e-09, -8.690856e-09, -1.023674e-08, -1.175831e-08, 
    -1.297652e-08, -1.389582e-08,
  -2.65852e-09, -2.5827e-09, -2.820368e-09, -3.184285e-09, -3.49477e-09, 
    -3.761423e-09, -4.004455e-09, -4.364254e-09, -5.161133e-09, -6.41208e-09, 
    -7.85727e-09, -9.253926e-09, -1.076563e-08, -1.208559e-08, -1.309734e-08,
  -2.524279e-09, -2.447054e-09, -2.58036e-09, -2.968704e-09, -3.248214e-09, 
    -3.505132e-09, -3.717154e-09, -3.968318e-09, -4.602939e-09, 
    -5.796589e-09, -7.251159e-09, -8.695343e-09, -1.008324e-08, 
    -1.137475e-08, -1.248154e-08,
  -2.433781e-09, -2.317003e-09, -2.462633e-09, -2.696932e-09, -2.936178e-09, 
    -3.105372e-09, -3.455053e-09, -3.854515e-09, -4.383796e-09, 
    -5.352391e-09, -6.700649e-09, -8.184823e-09, -9.677559e-09, 
    -1.107316e-08, -1.235342e-08,
  -2.469319e-09, -2.316504e-09, -2.388763e-09, -2.4965e-09, -2.664908e-09, 
    -2.93316e-09, -3.242381e-09, -3.777377e-09, -4.301582e-09, -5.119992e-09, 
    -6.359238e-09, -7.909295e-09, -9.30549e-09, -1.107375e-08, -1.249746e-08,
  -6.996689e-09, -7.35678e-09, -7.829844e-09, -8.499737e-09, -9.264479e-09, 
    -1.006288e-08, -1.084813e-08, -1.146279e-08, -1.193678e-08, 
    -1.236622e-08, -1.270751e-08, -1.298841e-08, -1.324196e-08, -1.34565e-08, 
    -1.370954e-08,
  -5.97589e-09, -6.394537e-09, -6.783077e-09, -7.268791e-09, -7.88833e-09, 
    -8.577042e-09, -9.367142e-09, -1.001659e-08, -1.062663e-08, 
    -1.118858e-08, -1.169798e-08, -1.222035e-08, -1.252928e-08, 
    -1.271981e-08, -1.292093e-08,
  -4.725752e-09, -5.238792e-09, -5.682212e-09, -6.099725e-09, -6.595238e-09, 
    -7.144345e-09, -7.889165e-09, -8.589478e-09, -9.287061e-09, 
    -9.886135e-09, -1.047595e-08, -1.104569e-08, -1.161562e-08, 
    -1.194514e-08, -1.224674e-08,
  -3.720021e-09, -4.163641e-09, -4.673677e-09, -5.117322e-09, -5.537122e-09, 
    -5.96716e-09, -6.491967e-09, -7.152809e-09, -7.814395e-09, -8.465217e-09, 
    -9.177082e-09, -9.668974e-09, -1.020872e-08, -1.077611e-08, -1.130737e-08,
  -3.118068e-09, -3.37522e-09, -3.856365e-09, -4.370034e-09, -4.754964e-09, 
    -5.106029e-09, -5.495572e-09, -5.991297e-09, -6.624247e-09, 
    -7.160161e-09, -7.82673e-09, -8.48945e-09, -9.075801e-09, -9.756213e-09, 
    -1.040425e-08,
  -2.810591e-09, -2.965645e-09, -3.221392e-09, -3.719759e-09, -4.206946e-09, 
    -4.552221e-09, -4.898038e-09, -5.195048e-09, -5.675957e-09, 
    -6.106637e-09, -6.681277e-09, -7.336352e-09, -8.112404e-09, 
    -8.859445e-09, -9.550533e-09,
  -2.466902e-09, -2.685006e-09, -2.846699e-09, -3.172846e-09, -3.679329e-09, 
    -4.062274e-09, -4.406743e-09, -4.737674e-09, -5.062208e-09, 
    -5.363685e-09, -5.909449e-09, -6.55527e-09, -7.368399e-09, -8.051299e-09, 
    -8.777871e-09,
  -2.197298e-09, -2.335377e-09, -2.504855e-09, -2.810659e-09, -3.273892e-09, 
    -3.712592e-09, -3.945942e-09, -4.130833e-09, -4.488975e-09, 
    -4.792644e-09, -5.363332e-09, -5.903623e-09, -6.731818e-09, 
    -7.292338e-09, -7.885931e-09,
  -2.052538e-09, -2.061481e-09, -2.211548e-09, -2.49304e-09, -2.89969e-09, 
    -3.362614e-09, -3.642748e-09, -3.682729e-09, -3.856467e-09, 
    -4.222471e-09, -4.820992e-09, -5.356712e-09, -6.001025e-09, 
    -6.450289e-09, -6.920132e-09,
  -1.982346e-09, -1.983528e-09, -2.068284e-09, -2.312586e-09, -2.629076e-09, 
    -2.91527e-09, -3.154726e-09, -3.387138e-09, -3.587122e-09, -3.993492e-09, 
    -4.408698e-09, -4.921832e-09, -5.317892e-09, -5.636093e-09, -6.021742e-09,
  -1.48056e-08, -1.528233e-08, -1.567544e-08, -1.603586e-08, -1.617972e-08, 
    -1.623365e-08, -1.61556e-08, -1.59913e-08, -1.561968e-08, -1.529294e-08, 
    -1.486065e-08, -1.445066e-08, -1.418111e-08, -1.370739e-08, -1.30264e-08,
  -1.231834e-08, -1.314131e-08, -1.370899e-08, -1.422645e-08, -1.445448e-08, 
    -1.460363e-08, -1.46135e-08, -1.446195e-08, -1.419065e-08, -1.38973e-08, 
    -1.359669e-08, -1.325129e-08, -1.277422e-08, -1.212808e-08, -1.136912e-08,
  -9.581093e-09, -1.067617e-08, -1.143132e-08, -1.204302e-08, -1.249433e-08, 
    -1.271187e-08, -1.280339e-08, -1.275658e-08, -1.258214e-08, -1.23484e-08, 
    -1.203195e-08, -1.16794e-08, -1.120736e-08, -1.056021e-08, -9.865825e-09,
  -6.991707e-09, -7.837579e-09, -8.735019e-09, -9.509253e-09, -1.008503e-08, 
    -1.04875e-08, -1.073009e-08, -1.077086e-08, -1.070401e-08, -1.051848e-08, 
    -1.025707e-08, -9.922092e-09, -9.484819e-09, -8.930559e-09, -8.429995e-09,
  -5.602077e-09, -5.866244e-09, -6.290295e-09, -6.87197e-09, -7.426722e-09, 
    -7.858427e-09, -8.158574e-09, -8.335251e-09, -8.385456e-09, 
    -8.310141e-09, -8.166657e-09, -7.93054e-09, -7.668552e-09, -7.376781e-09, 
    -7.148396e-09,
  -4.893514e-09, -4.962969e-09, -5.087126e-09, -5.285622e-09, -5.547193e-09, 
    -5.812058e-09, -6.009435e-09, -6.135483e-09, -6.196203e-09, 
    -6.218225e-09, -6.206661e-09, -6.188005e-09, -6.211922e-09, 
    -6.155805e-09, -6.091087e-09,
  -4.610272e-09, -4.640694e-09, -4.641616e-09, -4.640593e-09, -4.678471e-09, 
    -4.680478e-09, -4.709766e-09, -4.757878e-09, -4.791784e-09, 
    -4.814276e-09, -4.862798e-09, -4.917026e-09, -4.958567e-09, 
    -4.993193e-09, -5.014015e-09,
  -4.154737e-09, -4.317877e-09, -4.35791e-09, -4.311695e-09, -4.238482e-09, 
    -4.201862e-09, -4.112889e-09, -4.107725e-09, -4.080063e-09, 
    -4.120646e-09, -4.15588e-09, -4.170991e-09, -4.133748e-09, -4.123914e-09, 
    -4.100638e-09,
  -3.105113e-09, -3.369374e-09, -3.499211e-09, -3.543985e-09, -3.572996e-09, 
    -3.630565e-09, -3.715396e-09, -3.768623e-09, -3.76626e-09, -3.766573e-09, 
    -3.694169e-09, -3.611925e-09, -3.47887e-09, -3.380408e-09, -3.309381e-09,
  -1.606919e-09, -1.881219e-09, -2.052198e-09, -2.211169e-09, -2.319912e-09, 
    -2.51166e-09, -2.704099e-09, -2.88408e-09, -2.89933e-09, -2.898166e-09, 
    -2.880926e-09, -2.812132e-09, -2.741337e-09, -2.665111e-09, -2.615257e-09,
  -9.32925e-09, -9.808974e-09, -1.037231e-08, -1.090624e-08, -1.157764e-08, 
    -1.225756e-08, -1.2934e-08, -1.36852e-08, -1.443583e-08, -1.515208e-08, 
    -1.59095e-08, -1.673684e-08, -1.755622e-08, -1.865014e-08, -1.981356e-08,
  -8.881153e-09, -9.518843e-09, -1.001236e-08, -1.046973e-08, -1.091551e-08, 
    -1.143338e-08, -1.205737e-08, -1.270011e-08, -1.334313e-08, 
    -1.412017e-08, -1.487944e-08, -1.567003e-08, -1.642162e-08, -1.72204e-08, 
    -1.809635e-08,
  -7.23828e-09, -8.575584e-09, -9.572672e-09, -1.008337e-08, -1.054296e-08, 
    -1.09291e-08, -1.133642e-08, -1.18815e-08, -1.239425e-08, -1.298006e-08, 
    -1.366171e-08, -1.431441e-08, -1.508016e-08, -1.588154e-08, -1.6618e-08,
  -5.974229e-09, -7.016849e-09, -8.19639e-09, -9.303669e-09, -1.002725e-08, 
    -1.055005e-08, -1.092726e-08, -1.132046e-08, -1.169782e-08, 
    -1.211802e-08, -1.261983e-08, -1.312677e-08, -1.372022e-08, 
    -1.433302e-08, -1.494003e-08,
  -5.771239e-09, -6.046822e-09, -6.800692e-09, -7.798953e-09, -8.958399e-09, 
    -9.911369e-09, -1.044704e-08, -1.079966e-08, -1.117968e-08, 
    -1.157321e-08, -1.196122e-08, -1.237672e-08, -1.283367e-08, 
    -1.319503e-08, -1.347197e-08,
  -5.894391e-09, -5.888193e-09, -6.161556e-09, -6.574115e-09, -7.414009e-09, 
    -8.527861e-09, -9.577259e-09, -1.033391e-08, -1.066887e-08, 
    -1.092762e-08, -1.122356e-08, -1.149493e-08, -1.178775e-08, 
    -1.197364e-08, -1.216174e-08,
  -6.296593e-09, -6.026233e-09, -5.987074e-09, -6.149889e-09, -6.441019e-09, 
    -7.083911e-09, -8.001778e-09, -9.002762e-09, -9.837367e-09, 
    -1.021387e-08, -1.035061e-08, -1.046668e-08, -1.05867e-08, -1.071697e-08, 
    -1.090908e-08,
  -6.08843e-09, -6.553181e-09, -6.475077e-09, -6.136227e-09, -6.127487e-09, 
    -6.330092e-09, -6.757132e-09, -7.527648e-09, -8.379142e-09, -9.09798e-09, 
    -9.462477e-09, -9.506985e-09, -9.562175e-09, -9.735613e-09, -9.981757e-09,
  -5.232863e-09, -5.945527e-09, -6.640202e-09, -6.883396e-09, -6.526018e-09, 
    -6.348601e-09, -6.353138e-09, -6.617309e-09, -7.149417e-09, 
    -7.850133e-09, -8.468218e-09, -9.067755e-09, -9.257918e-09, 
    -9.453188e-09, -9.660867e-09,
  -3.893422e-09, -5.020956e-09, -5.775314e-09, -6.430829e-09, -6.900467e-09, 
    -6.90251e-09, -6.680851e-09, -6.579551e-09, -6.646133e-09, -6.908227e-09, 
    -7.378692e-09, -7.899869e-09, -8.572641e-09, -9.128206e-09, -9.479088e-09,
  -3.96031e-09, -4.454698e-09, -5.081609e-09, -5.879849e-09, -6.817707e-09, 
    -7.819328e-09, -8.824406e-09, -9.730867e-09, -1.013704e-08, 
    -1.016517e-08, -1.005e-08, -1.011936e-08, -1.035964e-08, -1.058679e-08, 
    -1.07817e-08,
  -3.435783e-09, -3.922549e-09, -4.44653e-09, -5.136138e-09, -5.846098e-09, 
    -6.645457e-09, -7.437206e-09, -8.369019e-09, -9.352663e-09, 
    -9.887514e-09, -1.029865e-08, -1.051397e-08, -1.062676e-08, 
    -1.071499e-08, -1.062469e-08,
  -3.002128e-09, -3.331198e-09, -3.745344e-09, -4.308663e-09, -4.99781e-09, 
    -5.756175e-09, -6.491248e-09, -7.22187e-09, -8.123743e-09, -9.095882e-09, 
    -9.819089e-09, -1.050228e-08, -1.093404e-08, -1.122409e-08, -1.114358e-08,
  -2.647088e-09, -2.97639e-09, -3.304234e-09, -3.710657e-09, -4.24403e-09, 
    -4.975605e-09, -5.773901e-09, -6.444147e-09, -7.139455e-09, 
    -7.984403e-09, -8.874172e-09, -9.68269e-09, -1.057598e-08, -1.122781e-08, 
    -1.165217e-08,
  -2.364928e-09, -2.626646e-09, -2.965328e-09, -3.311835e-09, -3.694335e-09, 
    -4.204493e-09, -4.945084e-09, -5.805718e-09, -6.493085e-09, 
    -7.156987e-09, -7.952509e-09, -8.76436e-09, -9.701641e-09, -1.072877e-08, 
    -1.149002e-08,
  -2.104316e-09, -2.285015e-09, -2.57528e-09, -2.957118e-09, -3.34534e-09, 
    -3.73042e-09, -4.246514e-09, -4.986658e-09, -5.863821e-09, -6.59452e-09, 
    -7.357257e-09, -8.088134e-09, -8.952257e-09, -9.949448e-09, -1.094045e-08,
  -1.86906e-09, -2.017772e-09, -2.24567e-09, -2.574802e-09, -2.946935e-09, 
    -3.362429e-09, -3.821554e-09, -4.383105e-09, -5.070903e-09, 
    -5.899248e-09, -6.738026e-09, -7.563139e-09, -8.342592e-09, 
    -9.167111e-09, -1.003415e-08,
  -1.658235e-09, -1.878176e-09, -2.075133e-09, -2.357122e-09, -2.653898e-09, 
    -2.993799e-09, -3.412047e-09, -3.955691e-09, -4.584889e-09, 
    -5.284159e-09, -6.094564e-09, -6.968958e-09, -7.853673e-09, 
    -8.583356e-09, -9.193955e-09,
  -1.31522e-09, -1.580946e-09, -1.800397e-09, -2.081435e-09, -2.355268e-09, 
    -2.626432e-09, -2.985137e-09, -3.464371e-09, -4.115381e-09, 
    -4.835159e-09, -5.618675e-09, -6.452701e-09, -7.298831e-09, 
    -8.006888e-09, -8.54124e-09,
  -1.130568e-09, -1.292871e-09, -1.4812e-09, -1.687675e-09, -1.858143e-09, 
    -2.147334e-09, -2.529863e-09, -2.979236e-09, -3.554987e-09, 
    -4.300035e-09, -5.121525e-09, -5.950845e-09, -6.693457e-09, 
    -7.316136e-09, -7.818201e-09,
  -2.486527e-09, -2.515509e-09, -2.514636e-09, -2.644561e-09, -2.886847e-09, 
    -3.279166e-09, -3.88071e-09, -4.34918e-09, -4.819616e-09, -5.465403e-09, 
    -6.189404e-09, -6.881197e-09, -7.238688e-09, -7.449021e-09, -7.783082e-09,
  -2.548262e-09, -2.675601e-09, -2.696362e-09, -2.618163e-09, -2.568544e-09, 
    -2.602481e-09, -2.828311e-09, -3.212901e-09, -3.743598e-09, 
    -4.140188e-09, -4.560554e-09, -5.073034e-09, -5.628601e-09, 
    -6.155452e-09, -6.619805e-09,
  -2.403655e-09, -2.406117e-09, -2.36662e-09, -2.337738e-09, -2.354198e-09, 
    -2.3981e-09, -2.434848e-09, -2.564864e-09, -2.824116e-09, -3.25448e-09, 
    -3.695495e-09, -4.049958e-09, -4.422197e-09, -4.93707e-09, -5.467616e-09,
  -2.104743e-09, -2.115794e-09, -2.072549e-09, -2.020945e-09, -1.989388e-09, 
    -2.039808e-09, -2.13146e-09, -2.236559e-09, -2.393726e-09, -2.607859e-09, 
    -2.961031e-09, -3.360238e-09, -3.752495e-09, -4.162386e-09, -4.666311e-09,
  -1.758566e-09, -1.729155e-09, -1.80231e-09, -1.815661e-09, -1.748122e-09, 
    -1.74869e-09, -1.819897e-09, -1.914354e-09, -2.044577e-09, -2.230107e-09, 
    -2.460091e-09, -2.781713e-09, -3.116903e-09, -3.455631e-09, -3.869896e-09,
  -1.564231e-09, -1.591555e-09, -1.647001e-09, -1.631277e-09, -1.498419e-09, 
    -1.436727e-09, -1.471839e-09, -1.52011e-09, -1.639371e-09, -1.832324e-09, 
    -2.084542e-09, -2.37893e-09, -2.703669e-09, -3.003273e-09, -3.307617e-09,
  -1.424928e-09, -1.562839e-09, -1.702692e-09, -1.68065e-09, -1.467575e-09, 
    -1.453633e-09, -1.496864e-09, -1.546006e-09, -1.57533e-09, -1.611859e-09, 
    -1.731327e-09, -1.993705e-09, -2.328128e-09, -2.69274e-09, -3.079877e-09,
  -1.145359e-09, -1.434353e-09, -1.560097e-09, -1.15318e-09, -9.631717e-10, 
    -8.719967e-10, -9.483681e-10, -1.244821e-09, -1.467075e-09, 
    -1.522007e-09, -1.556918e-09, -1.658406e-09, -1.945889e-09, 
    -2.302015e-09, -2.728313e-09,
  -4.944921e-10, -5.086554e-10, -4.537565e-10, -2.208888e-10, -4.445144e-10, 
    -6.256634e-10, -6.856254e-10, -8.974128e-10, -9.646877e-10, 
    -1.126042e-09, -1.356302e-09, -1.479717e-09, -1.637045e-09, 
    -1.980325e-09, -2.406411e-09,
  -3.346883e-10, -2.349096e-10, -1.068135e-10, -2.039781e-11, -1.447754e-10, 
    -4.604113e-10, -5.491553e-10, -7.31574e-10, -8.459711e-10, -9.417241e-10, 
    -1.061111e-09, -1.260505e-09, -1.447052e-09, -1.700264e-09, -2.202031e-09,
  -1.031227e-09, -1.035222e-09, -1.121389e-09, -1.304897e-09, -1.577252e-09, 
    -1.894231e-09, -2.25267e-09, -2.673621e-09, -3.0248e-09, -3.567484e-09, 
    -4.931878e-09, -6.77975e-09, -9.103463e-09, -1.037425e-08, -1.116974e-08,
  -6.701366e-10, -6.293999e-10, -5.992886e-10, -6.507586e-10, -8.086454e-10, 
    -1.057608e-09, -1.368964e-09, -1.71562e-09, -2.127359e-09, -2.522868e-09, 
    -3.016124e-09, -3.631892e-09, -4.681909e-09, -6.382942e-09, -8.262483e-09,
  -6.352507e-10, -5.349071e-10, -4.07621e-10, -3.423625e-10, -3.388632e-10, 
    -4.795362e-10, -7.135156e-10, -1.006416e-09, -1.317338e-09, 
    -1.652279e-09, -2.065934e-09, -2.573123e-09, -3.125806e-09, 
    -3.798471e-09, -4.716182e-09,
  -5.686424e-10, -4.42345e-10, -3.179221e-10, -1.845063e-10, -1.568509e-10, 
    -1.695426e-10, -2.909837e-10, -4.607847e-10, -6.69548e-10, -9.33328e-10, 
    -1.247751e-09, -1.67909e-09, -2.192552e-09, -2.713423e-09, -3.194593e-09,
  -4.428261e-10, -4.922149e-10, -4.466611e-10, -5.338184e-10, -5.544276e-10, 
    -4.966771e-10, -4.741458e-10, -5.06569e-10, -5.792186e-10, -6.531181e-10, 
    -7.194983e-10, -8.7054e-10, -1.161591e-09, -1.568477e-09, -2.148218e-09,
  -4.646396e-10, -5.083035e-10, -5.988283e-10, -6.038838e-10, -6.134561e-10, 
    -6.280628e-10, -7.007306e-10, -7.98505e-10, -9.175057e-10, -9.914596e-10, 
    -9.936438e-10, -9.163096e-10, -8.613362e-10, -1.036532e-09, -1.313041e-09,
  -4.645255e-10, -3.292826e-10, -3.670527e-10, -1.943964e-10, -3.860727e-11, 
    7.882323e-11, 1.036354e-10, 1.899966e-11, -1.407646e-10, -3.889866e-10, 
    -7.1023e-10, -9.372044e-10, -1.090287e-09, -1.091067e-09, -1.19164e-09,
  -3.372723e-10, 9.57917e-12, 1.342761e-10, 4.533174e-10, 7.252405e-10, 
    7.30119e-10, 6.071225e-10, 4.968204e-10, 4.083918e-10, 3.174126e-10, 
    8.481229e-11, -2.215477e-10, -6.345952e-10, -1.029663e-09, -1.305318e-09,
  -2.919373e-10, -7.155024e-10, -6.318612e-10, -4.887171e-10, -3.495287e-10, 
    -2.262957e-10, -4.764087e-11, 1.270988e-10, 1.537649e-10, 2.229165e-10, 
    2.75471e-10, 1.638052e-10, -8.702899e-11, -4.668426e-10, -9.104302e-10,
  -5.805191e-10, -5.397367e-10, -3.855855e-10, -5.632717e-10, -5.65673e-10, 
    -5.10436e-10, -3.309149e-10, -1.828888e-10, 1.040646e-10, 1.987027e-10, 
    1.800108e-10, 1.023186e-10, -9.619211e-12, -1.224349e-10, -4.18562e-10,
  -2.452609e-09, -2.425353e-09, -2.452163e-09, -2.500613e-09, -2.563152e-09, 
    -2.6052e-09, -2.590185e-09, -2.541812e-09, -2.455839e-09, -2.370755e-09, 
    -2.319818e-09, -2.317917e-09, -2.279185e-09, -2.238162e-09, -2.026609e-09,
  -1.338796e-09, -1.351774e-09, -1.384911e-09, -1.392231e-09, -1.352306e-09, 
    -1.309352e-09, -1.248174e-09, -1.188686e-09, -1.094525e-09, -1.06387e-09, 
    -1.088547e-09, -1.019254e-09, -8.47973e-10, -7.01482e-10, -7.784072e-10,
  -8.432393e-10, -8.372399e-10, -8.621748e-10, -8.817919e-10, -8.806864e-10, 
    -8.160669e-10, -7.257942e-10, -6.197004e-10, -5.285538e-10, -4.53349e-10, 
    -3.439808e-10, -2.086188e-10, -1.659184e-10, -4.320431e-10, -5.073144e-10,
  -3.93396e-10, -3.813935e-10, -3.965532e-10, -3.982432e-10, -4.066085e-10, 
    -4.484334e-10, -4.558448e-10, -4.465473e-10, -4.307153e-10, -4.06974e-10, 
    -3.82285e-10, -3.307553e-10, -2.297367e-10, -3.552499e-10, -3.921134e-10,
  -1.935496e-10, -1.832376e-10, -2.039195e-10, -2.277638e-10, -3.107185e-10, 
    -4.430092e-10, -5.262043e-10, -5.899535e-10, -6.580293e-10, 
    -7.270817e-10, -8.250902e-10, -8.583724e-10, -7.464283e-10, 
    -5.908923e-10, -4.617326e-10,
  -1.406909e-10, -1.459593e-10, -2.020471e-10, -2.578027e-10, -3.845652e-10, 
    -4.989284e-10, -6.18448e-10, -7.088006e-10, -7.664288e-10, -8.264728e-10, 
    -8.993701e-10, -1.04452e-09, -1.107443e-09, -1.064806e-09, -9.007728e-10,
  -2.210822e-10, -2.722619e-10, -3.877041e-10, -4.454732e-10, -5.481222e-10, 
    -6.742987e-10, -7.239743e-10, -7.174357e-10, -6.86132e-10, -6.311658e-10, 
    -6.724293e-10, -6.930718e-10, -7.803928e-10, -8.915094e-10, -9.734471e-10,
  -3.721291e-10, -4.088971e-10, -4.775776e-10, -4.082412e-10, -3.968409e-10, 
    -3.682173e-10, -3.783988e-10, -3.450753e-10, -3.570644e-10, 
    -2.911661e-10, -2.407949e-10, -2.487884e-10, -2.586809e-10, 
    -3.613401e-10, -5.363767e-10,
  -3.392664e-10, -3.598667e-10, -3.281677e-10, -3.046017e-10, -2.09819e-10, 
    -1.11683e-10, -9.136363e-11, -8.137248e-11, -1.064583e-10, -1.669124e-10, 
    -1.901255e-10, -2.198546e-10, -2.19748e-10, -2.331216e-10, -3.051427e-10,
  -2.92475e-10, -2.659408e-10, -2.689107e-10, -2.641104e-10, -2.656468e-10, 
    -2.732092e-10, -2.706984e-10, -1.979238e-10, -1.203232e-10, 
    -2.359503e-10, -2.833551e-10, -3.83023e-10, -3.997271e-10, -3.072975e-10, 
    -2.446574e-10,
  -8.0507e-09, -9.386285e-09, -1.094989e-08, -1.263856e-08, -1.424199e-08, 
    -1.555003e-08, -1.655616e-08, -1.735691e-08, -1.805916e-08, 
    -1.849919e-08, -1.880705e-08, -1.885406e-08, -1.875584e-08, 
    -1.849491e-08, -1.810478e-08,
  -5.092514e-09, -5.894047e-09, -6.823573e-09, -7.822814e-09, -8.880245e-09, 
    -1.007709e-08, -1.130815e-08, -1.230858e-08, -1.311002e-08, -1.37223e-08, 
    -1.412548e-08, -1.432565e-08, -1.431018e-08, -1.409417e-08, -1.369934e-08,
  -3.18989e-09, -3.621174e-09, -4.148097e-09, -4.731243e-09, -5.374252e-09, 
    -6.059661e-09, -6.796246e-09, -7.54282e-09, -8.297833e-09, -8.876849e-09, 
    -9.307768e-09, -9.534072e-09, -9.558626e-09, -9.404857e-09, -9.082879e-09,
  -2.314592e-09, -2.437142e-09, -2.665551e-09, -2.948137e-09, -3.26021e-09, 
    -3.58905e-09, -3.950927e-09, -4.309337e-09, -4.695584e-09, -5.029293e-09, 
    -5.33808e-09, -5.509375e-09, -5.558677e-09, -5.442023e-09, -5.179509e-09,
  -1.788852e-09, -1.782809e-09, -1.840461e-09, -1.936021e-09, -2.046606e-09, 
    -2.166892e-09, -2.299905e-09, -2.430328e-09, -2.553206e-09, -2.64974e-09, 
    -2.716086e-09, -2.732016e-09, -2.711601e-09, -2.618092e-09, -2.472148e-09,
  -1.460893e-09, -1.43903e-09, -1.418777e-09, -1.436024e-09, -1.462082e-09, 
    -1.489102e-09, -1.518266e-09, -1.547546e-09, -1.567504e-09, 
    -1.577127e-09, -1.558135e-09, -1.517568e-09, -1.458258e-09, 
    -1.379124e-09, -1.298488e-09,
  -1.142283e-09, -1.156643e-09, -1.138323e-09, -1.126653e-09, -1.112778e-09, 
    -1.099691e-09, -1.081092e-09, -1.068757e-09, -1.050855e-09, 
    -1.036925e-09, -1.006286e-09, -9.708835e-10, -9.222883e-10, 
    -8.887384e-10, -8.387712e-10,
  -8.585548e-10, -8.646875e-10, -8.68098e-10, -8.78526e-10, -8.763196e-10, 
    -8.803613e-10, -8.626647e-10, -8.238379e-10, -7.744514e-10, 
    -7.207632e-10, -6.723239e-10, -6.24875e-10, -5.929418e-10, -5.562764e-10, 
    -5.297561e-10,
  -5.299821e-10, -5.125157e-10, -5.202555e-10, -5.283155e-10, -5.220826e-10, 
    -5.181708e-10, -5.037581e-10, -4.795835e-10, -4.451829e-10, 
    -4.105799e-10, -3.959348e-10, -3.720472e-10, -3.3353e-10, -2.886714e-10, 
    -2.555251e-10,
  -2.623786e-10, -2.396841e-10, -2.347274e-10, -2.571477e-10, -2.921517e-10, 
    -3.329945e-10, -3.716999e-10, -3.674546e-10, -4.202232e-10, 
    -4.709979e-10, -4.967763e-10, -4.615851e-10, -4.05481e-10, -3.443516e-10, 
    -3.103403e-10,
  -1.877334e-08, -1.94284e-08, -1.990456e-08, -1.889737e-08, -1.763543e-08, 
    -1.680657e-08, -1.642904e-08, -1.594136e-08, -1.537613e-08, 
    -1.510162e-08, -1.518372e-08, -1.560755e-08, -1.625505e-08, 
    -1.703373e-08, -1.784007e-08,
  -1.942897e-08, -1.907002e-08, -1.935613e-08, -2.001546e-08, -1.973166e-08, 
    -1.87637e-08, -1.797297e-08, -1.744325e-08, -1.712772e-08, -1.649585e-08, 
    -1.623555e-08, -1.647257e-08, -1.701852e-08, -1.774432e-08, -1.85574e-08,
  -1.840425e-08, -1.875665e-08, -1.889159e-08, -1.911188e-08, -1.943003e-08, 
    -1.915564e-08, -1.858984e-08, -1.797974e-08, -1.741533e-08, 
    -1.765357e-08, -1.803447e-08, -1.841174e-08, -1.881597e-08, 
    -1.918437e-08, -1.948685e-08,
  -1.582826e-08, -1.730744e-08, -1.78959e-08, -1.797384e-08, -1.858905e-08, 
    -1.87416e-08, -1.821386e-08, -1.767805e-08, -1.761532e-08, -1.77665e-08, 
    -1.808871e-08, -1.859624e-08, -1.914134e-08, -1.960832e-08, -1.976538e-08,
  -1.265932e-08, -1.445699e-08, -1.619285e-08, -1.728193e-08, -1.751023e-08, 
    -1.7489e-08, -1.749427e-08, -1.725163e-08, -1.678556e-08, -1.688428e-08, 
    -1.717354e-08, -1.763511e-08, -1.797416e-08, -1.836224e-08, -1.861002e-08,
  -8.742014e-09, -1.079842e-08, -1.272183e-08, -1.435821e-08, -1.572677e-08, 
    -1.658869e-08, -1.675012e-08, -1.659355e-08, -1.627687e-08, 
    -1.593288e-08, -1.589746e-08, -1.620513e-08, -1.650359e-08, 
    -1.685829e-08, -1.719016e-08,
  -5.203899e-09, -7.017253e-09, -8.843474e-09, -1.06837e-08, -1.231583e-08, 
    -1.348765e-08, -1.441201e-08, -1.494448e-08, -1.523493e-08, 
    -1.542405e-08, -1.530671e-08, -1.532057e-08, -1.527972e-08, 
    -1.519347e-08, -1.502326e-08,
  -3.042389e-09, -4.001652e-09, -5.538655e-09, -7.105804e-09, -8.672756e-09, 
    -1.012107e-08, -1.126659e-08, -1.213991e-08, -1.272267e-08, -1.30716e-08, 
    -1.325962e-08, -1.328666e-08, -1.318982e-08, -1.298176e-08, -1.262276e-08,
  -2.30086e-09, -2.607733e-09, -3.237691e-09, -4.215577e-09, -5.485337e-09, 
    -6.779474e-09, -7.990322e-09, -8.999144e-09, -9.782553e-09, 
    -1.029797e-08, -1.054679e-08, -1.068915e-08, -1.060548e-08, 
    -1.037857e-08, -9.95108e-09,
  -1.453579e-09, -1.77894e-09, -2.1793e-09, -2.670191e-09, -3.282518e-09, 
    -4.098044e-09, -4.988757e-09, -5.895421e-09, -6.717127e-09, 
    -7.386844e-09, -7.810818e-09, -7.98035e-09, -7.998032e-09, -7.803122e-09, 
    -7.506991e-09,
  -1.315836e-08, -1.331216e-08, -1.328643e-08, -1.318035e-08, -1.293046e-08, 
    -1.270853e-08, -1.264062e-08, -1.24995e-08, -1.243374e-08, -1.235065e-08, 
    -1.211299e-08, -1.181162e-08, -1.160305e-08, -1.132642e-08, -1.099925e-08,
  -1.331607e-08, -1.341806e-08, -1.351347e-08, -1.350618e-08, -1.337088e-08, 
    -1.327542e-08, -1.325692e-08, -1.311342e-08, -1.295591e-08, 
    -1.273965e-08, -1.244623e-08, -1.19544e-08, -1.141694e-08, -1.092222e-08, 
    -1.066856e-08,
  -1.409525e-08, -1.381845e-08, -1.363957e-08, -1.35776e-08, -1.344625e-08, 
    -1.336591e-08, -1.326139e-08, -1.309672e-08, -1.282074e-08, 
    -1.240214e-08, -1.208388e-08, -1.187907e-08, -1.169226e-08, 
    -1.164682e-08, -1.17272e-08,
  -1.403854e-08, -1.413614e-08, -1.417496e-08, -1.397764e-08, -1.374033e-08, 
    -1.356198e-08, -1.34457e-08, -1.316484e-08, -1.27645e-08, -1.239308e-08, 
    -1.214154e-08, -1.204555e-08, -1.200365e-08, -1.216724e-08, -1.225467e-08,
  -1.302114e-08, -1.354941e-08, -1.399193e-08, -1.418211e-08, -1.417532e-08, 
    -1.394621e-08, -1.376169e-08, -1.363727e-08, -1.333452e-08, -1.2901e-08, 
    -1.265654e-08, -1.262053e-08, -1.278362e-08, -1.29989e-08, -1.307891e-08,
  -1.18177e-08, -1.236264e-08, -1.294285e-08, -1.360788e-08, -1.401559e-08, 
    -1.446446e-08, -1.453607e-08, -1.436336e-08, -1.417419e-08, 
    -1.392138e-08, -1.362762e-08, -1.353726e-08, -1.376064e-08, 
    -1.390087e-08, -1.420211e-08,
  -1.054312e-08, -1.147008e-08, -1.193039e-08, -1.261892e-08, -1.326333e-08, 
    -1.392201e-08, -1.464324e-08, -1.525021e-08, -1.541386e-08, 
    -1.532395e-08, -1.535376e-08, -1.54201e-08, -1.57409e-08, -1.622563e-08, 
    -1.713319e-08,
  -8.297772e-09, -9.543573e-09, -1.05872e-08, -1.161834e-08, -1.246366e-08, 
    -1.323357e-08, -1.406833e-08, -1.484654e-08, -1.572365e-08, 
    -1.637183e-08, -1.69063e-08, -1.731882e-08, -1.810123e-08, -1.862104e-08, 
    -1.903996e-08,
  -5.662102e-09, -6.670202e-09, -7.820468e-09, -9.09533e-09, -1.046757e-08, 
    -1.164544e-08, -1.275804e-08, -1.381182e-08, -1.494134e-08, 
    -1.594833e-08, -1.67683e-08, -1.744369e-08, -1.785004e-08, -1.822547e-08, 
    -1.810932e-08,
  -3.267964e-09, -3.891301e-09, -4.652182e-09, -5.567486e-09, -6.598066e-09, 
    -7.868708e-09, -9.123934e-09, -1.046724e-08, -1.167861e-08, 
    -1.287372e-08, -1.385944e-08, -1.467047e-08, -1.51431e-08, -1.537353e-08, 
    -1.490604e-08,
  -1.601236e-08, -1.822413e-08, -1.955765e-08, -2.03213e-08, -2.084104e-08, 
    -2.126741e-08, -2.1604e-08, -2.192409e-08, -2.208817e-08, -2.216408e-08, 
    -2.209431e-08, -2.189163e-08, -2.162336e-08, -2.133526e-08, -2.08935e-08,
  -1.395453e-08, -1.512108e-08, -1.681423e-08, -1.839445e-08, -1.938989e-08, 
    -1.999348e-08, -2.025935e-08, -2.035305e-08, -2.04304e-08, -2.045794e-08, 
    -2.047679e-08, -2.037684e-08, -2.016869e-08, -1.968463e-08, -1.883323e-08,
  -1.305774e-08, -1.339488e-08, -1.397165e-08, -1.517984e-08, -1.661958e-08, 
    -1.80217e-08, -1.887053e-08, -1.918567e-08, -1.917521e-08, -1.915303e-08, 
    -1.900109e-08, -1.881711e-08, -1.832495e-08, -1.756304e-08, -1.674526e-08,
  -1.371208e-08, -1.332115e-08, -1.348312e-08, -1.387665e-08, -1.447423e-08, 
    -1.529119e-08, -1.624644e-08, -1.713832e-08, -1.76371e-08, -1.772632e-08, 
    -1.753359e-08, -1.712893e-08, -1.654578e-08, -1.595644e-08, -1.540203e-08,
  -1.419994e-08, -1.41734e-08, -1.39651e-08, -1.40211e-08, -1.423261e-08, 
    -1.454688e-08, -1.495338e-08, -1.544328e-08, -1.577239e-08, 
    -1.599028e-08, -1.587179e-08, -1.561273e-08, -1.529956e-08, 
    -1.499352e-08, -1.488504e-08,
  -1.366961e-08, -1.419247e-08, -1.440628e-08, -1.427742e-08, -1.424181e-08, 
    -1.421036e-08, -1.418663e-08, -1.426732e-08, -1.433573e-08, -1.43788e-08, 
    -1.438479e-08, -1.43094e-08, -1.420479e-08, -1.416473e-08, -1.426524e-08,
  -1.184325e-08, -1.268804e-08, -1.362796e-08, -1.417081e-08, -1.441626e-08, 
    -1.429462e-08, -1.409922e-08, -1.397526e-08, -1.384556e-08, 
    -1.381395e-08, -1.385868e-08, -1.382718e-08, -1.386404e-08, 
    -1.389726e-08, -1.407278e-08,
  -1.029882e-08, -1.07697e-08, -1.142888e-08, -1.206833e-08, -1.286466e-08, 
    -1.353831e-08, -1.393139e-08, -1.410773e-08, -1.412635e-08, 
    -1.417873e-08, -1.420473e-08, -1.422208e-08, -1.414753e-08, 
    -1.408256e-08, -1.39723e-08,
  -1.020255e-08, -1.02303e-08, -1.052225e-08, -1.089104e-08, -1.144115e-08, 
    -1.206562e-08, -1.272583e-08, -1.334216e-08, -1.38596e-08, -1.426255e-08, 
    -1.441807e-08, -1.445191e-08, -1.427837e-08, -1.386574e-08, -1.345944e-08,
  -9.845957e-09, -9.751449e-09, -9.708423e-09, -9.902113e-09, -1.016029e-08, 
    -1.064079e-08, -1.106095e-08, -1.15458e-08, -1.195443e-08, -1.225273e-08, 
    -1.229684e-08, -1.223706e-08, -1.199506e-08, -1.155288e-08, -1.112787e-08,
  -2.785351e-08, -2.727912e-08, -2.489546e-08, -2.28722e-08, -2.053258e-08, 
    -1.895929e-08, -1.854217e-08, -1.871303e-08, -1.889057e-08, 
    -1.919079e-08, -1.958523e-08, -2.013994e-08, -2.074026e-08, 
    -2.151132e-08, -2.214115e-08,
  -2.530285e-08, -2.682362e-08, -2.696824e-08, -2.581878e-08, -2.375832e-08, 
    -2.191514e-08, -2.040321e-08, -1.964904e-08, -1.94707e-08, -1.959373e-08, 
    -1.9883e-08, -2.034441e-08, -2.077514e-08, -2.128838e-08, -2.18195e-08,
  -2.157488e-08, -2.351395e-08, -2.527173e-08, -2.640097e-08, -2.663772e-08, 
    -2.519288e-08, -2.353938e-08, -2.206972e-08, -2.115273e-08, 
    -2.072571e-08, -2.065829e-08, -2.092648e-08, -2.126867e-08, 
    -2.151126e-08, -2.16706e-08,
  -1.803299e-08, -1.947019e-08, -2.1319e-08, -2.308998e-08, -2.448082e-08, 
    -2.539275e-08, -2.57121e-08, -2.500945e-08, -2.393978e-08, -2.289439e-08, 
    -2.232876e-08, -2.192619e-08, -2.187196e-08, -2.170251e-08, -2.151895e-08,
  -1.518772e-08, -1.608477e-08, -1.721559e-08, -1.874712e-08, -2.044887e-08, 
    -2.199814e-08, -2.313701e-08, -2.400059e-08, -2.451198e-08, 
    -2.448193e-08, -2.404221e-08, -2.335412e-08, -2.268946e-08, 
    -2.212483e-08, -2.151223e-08,
  -1.308297e-08, -1.331882e-08, -1.373333e-08, -1.438507e-08, -1.526045e-08, 
    -1.633724e-08, -1.754935e-08, -1.890113e-08, -2.010923e-08, 
    -2.105184e-08, -2.148041e-08, -2.158141e-08, -2.136948e-08, 
    -2.091556e-08, -2.043867e-08,
  -1.302214e-08, -1.275379e-08, -1.243458e-08, -1.233089e-08, -1.236662e-08, 
    -1.257889e-08, -1.290292e-08, -1.334008e-08, -1.386845e-08, 
    -1.447634e-08, -1.508955e-08, -1.556193e-08, -1.579743e-08, 
    -1.586685e-08, -1.579792e-08,
  -1.435934e-08, -1.413873e-08, -1.388345e-08, -1.361108e-08, -1.326444e-08, 
    -1.293938e-08, -1.259535e-08, -1.226927e-08, -1.213601e-08, 
    -1.217283e-08, -1.228669e-08, -1.242637e-08, -1.249073e-08, 
    -1.264034e-08, -1.272333e-08,
  -1.348871e-08, -1.386508e-08, -1.411221e-08, -1.427336e-08, -1.43762e-08, 
    -1.428645e-08, -1.419688e-08, -1.395517e-08, -1.36679e-08, -1.345549e-08, 
    -1.326265e-08, -1.315609e-08, -1.310594e-08, -1.316906e-08, -1.328466e-08,
  -9.818397e-09, -1.064312e-08, -1.136356e-08, -1.180902e-08, -1.231464e-08, 
    -1.267846e-08, -1.330642e-08, -1.35626e-08, -1.365962e-08, -1.370843e-08, 
    -1.364616e-08, -1.361573e-08, -1.356911e-08, -1.350172e-08, -1.342186e-08,
  -1.572747e-08, -1.442487e-08, -1.358511e-08, -1.28437e-08, -1.249852e-08, 
    -1.262916e-08, -1.259384e-08, -1.302154e-08, -1.328517e-08, 
    -1.360854e-08, -1.466723e-08, -1.605007e-08, -1.78292e-08, -1.957355e-08, 
    -2.081498e-08,
  -2.044261e-08, -1.866683e-08, -1.584659e-08, -1.421403e-08, -1.351594e-08, 
    -1.320903e-08, -1.303035e-08, -1.29439e-08, -1.316867e-08, -1.334672e-08, 
    -1.368699e-08, -1.470235e-08, -1.59964e-08, -1.799052e-08, -1.941262e-08,
  -2.350845e-08, -2.379518e-08, -2.18656e-08, -1.845315e-08, -1.574166e-08, 
    -1.446561e-08, -1.369491e-08, -1.348755e-08, -1.348703e-08, 
    -1.368785e-08, -1.392884e-08, -1.427403e-08, -1.501596e-08, 
    -1.615377e-08, -1.789118e-08,
  -2.322896e-08, -2.49796e-08, -2.564046e-08, -2.572912e-08, -2.362219e-08, 
    -1.939413e-08, -1.696712e-08, -1.508589e-08, -1.432335e-08, 
    -1.403263e-08, -1.398262e-08, -1.425647e-08, -1.468298e-08, 
    -1.544763e-08, -1.647625e-08,
  -2.319387e-08, -2.56898e-08, -2.727952e-08, -2.786351e-08, -2.826664e-08, 
    -2.809754e-08, -2.596653e-08, -2.282797e-08, -1.910499e-08, 
    -1.691961e-08, -1.57041e-08, -1.491962e-08, -1.474528e-08, -1.493446e-08, 
    -1.543814e-08,
  -1.979462e-08, -2.188956e-08, -2.414313e-08, -2.635723e-08, -2.804805e-08, 
    -2.904007e-08, -2.933965e-08, -2.924665e-08, -2.895586e-08, 
    -2.662347e-08, -2.402825e-08, -2.100772e-08, -1.8933e-08, -1.718219e-08, 
    -1.653062e-08,
  -1.64793e-08, -1.758618e-08, -1.918226e-08, -2.061889e-08, -2.214199e-08, 
    -2.342883e-08, -2.48555e-08, -2.600366e-08, -2.665996e-08, -2.690761e-08, 
    -2.694335e-08, -2.670434e-08, -2.611937e-08, -2.518864e-08, -2.37357e-08,
  -1.477236e-08, -1.512992e-08, -1.58479e-08, -1.664305e-08, -1.755544e-08, 
    -1.842988e-08, -1.933907e-08, -2.018266e-08, -2.103081e-08, 
    -2.192638e-08, -2.264856e-08, -2.32276e-08, -2.365332e-08, -2.388693e-08, 
    -2.392199e-08,
  -1.220354e-08, -1.261535e-08, -1.316566e-08, -1.368092e-08, -1.434054e-08, 
    -1.496949e-08, -1.561696e-08, -1.632814e-08, -1.692772e-08, 
    -1.758489e-08, -1.809307e-08, -1.854671e-08, -1.888838e-08, 
    -1.915144e-08, -1.936453e-08,
  -7.437438e-09, -7.953028e-09, -8.552377e-09, -9.173769e-09, -9.76013e-09, 
    -1.042733e-08, -1.115489e-08, -1.184036e-08, -1.25288e-08, -1.310805e-08, 
    -1.368359e-08, -1.407039e-08, -1.436392e-08, -1.452119e-08, -1.448826e-08,
  -7.586243e-09, -7.468509e-09, -7.534488e-09, -7.627462e-09, -7.803024e-09, 
    -8.128265e-09, -8.434847e-09, -8.831107e-09, -9.353504e-09, 
    -9.945571e-09, -1.045902e-08, -1.128957e-08, -1.244993e-08, 
    -1.429618e-08, -1.673565e-08,
  -8.269746e-09, -8.128776e-09, -8.066772e-09, -8.122622e-09, -8.154182e-09, 
    -8.296886e-09, -8.56125e-09, -8.837991e-09, -9.216872e-09, -9.715094e-09, 
    -1.012723e-08, -1.060289e-08, -1.132024e-08, -1.23333e-08, -1.412308e-08,
  -8.829396e-09, -8.872886e-09, -8.738714e-09, -8.624553e-09, -8.641623e-09, 
    -8.659641e-09, -8.781699e-09, -9.017223e-09, -9.283363e-09, 
    -9.716047e-09, -1.010371e-08, -1.049403e-08, -1.088721e-08, 
    -1.145033e-08, -1.233506e-08,
  -9.454798e-09, -9.516918e-09, -9.477183e-09, -9.445237e-09, -9.156245e-09, 
    -9.081269e-09, -9.11384e-09, -9.282342e-09, -9.475795e-09, -9.756103e-09, 
    -1.015009e-08, -1.056396e-08, -1.087054e-08, -1.125163e-08, -1.164886e-08,
  -1.048453e-08, -1.04834e-08, -1.054798e-08, -1.066242e-08, -1.067366e-08, 
    -1.029471e-08, -9.959089e-09, -9.811212e-09, -9.85076e-09, -9.970525e-09, 
    -1.020707e-08, -1.053628e-08, -1.085839e-08, -1.114967e-08, -1.157451e-08,
  -1.241362e-08, -1.162298e-08, -1.194369e-08, -1.243281e-08, -1.284408e-08, 
    -1.318731e-08, -1.32221e-08, -1.281669e-08, -1.243168e-08, -1.206491e-08, 
    -1.188619e-08, -1.184943e-08, -1.17374e-08, -1.166395e-08, -1.179901e-08,
  -1.488838e-08, -1.415113e-08, -1.34418e-08, -1.350853e-08, -1.398268e-08, 
    -1.487824e-08, -1.567938e-08, -1.635179e-08, -1.639066e-08, 
    -1.622779e-08, -1.56636e-08, -1.542158e-08, -1.531756e-08, -1.506683e-08, 
    -1.466067e-08,
  -1.688009e-08, -1.630061e-08, -1.596045e-08, -1.535794e-08, -1.47569e-08, 
    -1.484664e-08, -1.552091e-08, -1.632461e-08, -1.744068e-08, 
    -1.837227e-08, -1.882533e-08, -1.87829e-08, -1.848144e-08, -1.840706e-08, 
    -1.836919e-08,
  -1.621453e-08, -1.676129e-08, -1.699066e-08, -1.72563e-08, -1.713736e-08, 
    -1.683857e-08, -1.66923e-08, -1.658594e-08, -1.684801e-08, -1.740189e-08, 
    -1.815477e-08, -1.904568e-08, -1.991889e-08, -2.054367e-08, -2.094714e-08,
  -1.237768e-08, -1.372654e-08, -1.450857e-08, -1.510588e-08, -1.59523e-08, 
    -1.626448e-08, -1.687575e-08, -1.7285e-08, -1.736345e-08, -1.73062e-08, 
    -1.723512e-08, -1.73475e-08, -1.765246e-08, -1.812343e-08, -1.863454e-08,
  -8.523554e-09, -8.589023e-09, -8.762695e-09, -8.997728e-09, -9.220091e-09, 
    -9.456594e-09, -9.649094e-09, -9.909481e-09, -1.022992e-08, 
    -1.047878e-08, -1.076869e-08, -1.099359e-08, -1.123119e-08, 
    -1.118993e-08, -1.112441e-08,
  -7.982558e-09, -7.995759e-09, -8.184297e-09, -8.419327e-09, -8.599531e-09, 
    -8.700447e-09, -8.829209e-09, -8.914002e-09, -9.092802e-09, 
    -9.296459e-09, -9.591393e-09, -9.828312e-09, -1.019918e-08, 
    -1.067041e-08, -1.097516e-08,
  -7.861042e-09, -7.773967e-09, -7.836104e-09, -7.989287e-09, -8.146777e-09, 
    -8.191356e-09, -8.211821e-09, -8.196358e-09, -8.172166e-09, 
    -8.207043e-09, -8.366992e-09, -8.574077e-09, -8.885917e-09, 
    -9.253345e-09, -9.849035e-09,
  -7.957262e-09, -7.754932e-09, -7.73889e-09, -7.725617e-09, -7.751947e-09, 
    -7.775629e-09, -7.733131e-09, -7.655513e-09, -7.567491e-09, 
    -7.458933e-09, -7.451639e-09, -7.525228e-09, -7.725088e-09, 
    -7.917451e-09, -8.237497e-09,
  -8.567358e-09, -8.259698e-09, -8.073628e-09, -7.947555e-09, -7.828294e-09, 
    -7.745262e-09, -7.695806e-09, -7.565903e-09, -7.434691e-09, 
    -7.287435e-09, -7.182693e-09, -7.090872e-09, -7.125821e-09, 
    -7.215707e-09, -7.360436e-09,
  -9.17877e-09, -8.994713e-09, -8.70476e-09, -8.367634e-09, -8.16368e-09, 
    -7.968413e-09, -7.773068e-09, -7.62432e-09, -7.486538e-09, -7.373478e-09, 
    -7.255526e-09, -7.171434e-09, -7.138509e-09, -7.163731e-09, -7.188612e-09,
  -1.010357e-08, -1.009487e-08, -9.849524e-09, -9.605656e-09, -9.358098e-09, 
    -9.122152e-09, -8.970582e-09, -8.745981e-09, -8.420936e-09, 
    -8.116634e-09, -7.795075e-09, -7.559113e-09, -7.4331e-09, -7.402462e-09, 
    -7.418548e-09,
  -1.045205e-08, -1.063961e-08, -1.064998e-08, -1.046445e-08, -1.034276e-08, 
    -1.023779e-08, -1.017944e-08, -1.004555e-08, -9.843276e-09, 
    -9.686903e-09, -9.582143e-09, -9.47562e-09, -9.365674e-09, -9.208443e-09, 
    -9.049783e-09,
  -9.354562e-09, -1.017178e-08, -1.064091e-08, -1.108065e-08, -1.13399e-08, 
    -1.166762e-08, -1.197493e-08, -1.223567e-08, -1.23569e-08, -1.227064e-08, 
    -1.194184e-08, -1.16443e-08, -1.134344e-08, -1.11283e-08, -1.096446e-08,
  -7.786288e-09, -8.569236e-09, -9.284466e-09, -9.901934e-09, -1.06502e-08, 
    -1.13658e-08, -1.208682e-08, -1.278904e-08, -1.370182e-08, -1.446327e-08, 
    -1.504822e-08, -1.536974e-08, -1.537145e-08, -1.498528e-08, -1.452875e-08,
  -1.035781e-08, -1.07487e-08, -1.148984e-08, -1.242467e-08, -1.285752e-08, 
    -1.33889e-08, -1.37854e-08, -1.411792e-08, -1.418499e-08, -1.421413e-08, 
    -1.420267e-08, -1.411824e-08, -1.401029e-08, -1.37292e-08, -1.369957e-08,
  -9.384148e-09, -9.452425e-09, -9.665426e-09, -1.028189e-08, -1.101212e-08, 
    -1.159444e-08, -1.217875e-08, -1.275454e-08, -1.326442e-08, 
    -1.364531e-08, -1.390785e-08, -1.404842e-08, -1.417487e-08, -1.42083e-08, 
    -1.415344e-08,
  -9.132743e-09, -8.975886e-09, -8.947308e-09, -8.903293e-09, -9.264373e-09, 
    -9.895569e-09, -1.054573e-08, -1.111426e-08, -1.169543e-08, 
    -1.226901e-08, -1.275884e-08, -1.316443e-08, -1.343271e-08, 
    -1.363479e-08, -1.373535e-08,
  -9.716532e-09, -9.355557e-09, -8.974797e-09, -8.736499e-09, -8.536548e-09, 
    -8.55116e-09, -8.897418e-09, -9.436222e-09, -9.993374e-09, -1.053318e-08, 
    -1.10017e-08, -1.148767e-08, -1.19359e-08, -1.228703e-08, -1.255963e-08,
  -1.012794e-08, -1.00404e-08, -9.745914e-09, -9.293345e-09, -8.798781e-09, 
    -8.422623e-09, -8.234256e-09, -8.322075e-09, -8.577679e-09, -8.92006e-09, 
    -9.366442e-09, -9.771657e-09, -1.015269e-08, -1.049345e-08, -1.080141e-08,
  -9.880205e-09, -9.966681e-09, -1.003421e-08, -9.962083e-09, -9.6716e-09, 
    -9.186582e-09, -8.739664e-09, -8.36993e-09, -8.270335e-09, -8.281781e-09, 
    -8.40746e-09, -8.577755e-09, -8.794674e-09, -9.005081e-09, -9.20496e-09,
  -9.263675e-09, -9.604268e-09, -9.61618e-09, -9.660804e-09, -9.727948e-09, 
    -9.667083e-09, -9.374909e-09, -9.05032e-09, -8.786804e-09, -8.552441e-09, 
    -8.432002e-09, -8.368304e-09, -8.343965e-09, -8.329041e-09, -8.321575e-09,
  -8.167831e-09, -8.777279e-09, -9.18261e-09, -9.355381e-09, -9.463046e-09, 
    -9.456349e-09, -9.487052e-09, -9.399924e-09, -9.336512e-09, 
    -9.157012e-09, -8.924199e-09, -8.678081e-09, -8.474614e-09, 
    -8.363883e-09, -8.278552e-09,
  -6.619744e-09, -7.285369e-09, -8.023531e-09, -8.642596e-09, -9.023836e-09, 
    -9.177933e-09, -9.16809e-09, -9.285066e-09, -9.30839e-09, -9.324534e-09, 
    -9.266489e-09, -9.104781e-09, -8.925813e-09, -8.760722e-09, -8.672218e-09,
  -5.05481e-09, -5.698594e-09, -6.412084e-09, -7.185533e-09, -7.898945e-09, 
    -8.498393e-09, -8.727437e-09, -8.795773e-09, -9.015515e-09, 
    -9.254312e-09, -9.397575e-09, -9.469756e-09, -9.412826e-09, 
    -9.358311e-09, -9.299153e-09,
  -1.389687e-08, -1.428026e-08, -1.406962e-08, -1.432169e-08, -1.401386e-08, 
    -1.37037e-08, -1.389375e-08, -1.420538e-08, -1.449454e-08, -1.476354e-08, 
    -1.485537e-08, -1.452208e-08, -1.419226e-08, -1.434981e-08, -1.455679e-08,
  -1.268993e-08, -1.314932e-08, -1.390811e-08, -1.374106e-08, -1.410006e-08, 
    -1.422843e-08, -1.41445e-08, -1.406736e-08, -1.409174e-08, -1.438783e-08, 
    -1.477106e-08, -1.499831e-08, -1.487436e-08, -1.46613e-08, -1.442785e-08,
  -1.165115e-08, -1.224843e-08, -1.268235e-08, -1.36512e-08, -1.353091e-08, 
    -1.396975e-08, -1.430254e-08, -1.43274e-08, -1.431251e-08, -1.434284e-08, 
    -1.455863e-08, -1.484754e-08, -1.473454e-08, -1.458479e-08, -1.449278e-08,
  -1.048359e-08, -1.153698e-08, -1.205288e-08, -1.239933e-08, -1.291841e-08, 
    -1.31324e-08, -1.343169e-08, -1.404299e-08, -1.429851e-08, -1.440872e-08, 
    -1.456163e-08, -1.489665e-08, -1.527729e-08, -1.545468e-08, -1.534939e-08,
  -8.426341e-09, -1.024647e-08, -1.155459e-08, -1.205873e-08, -1.229606e-08, 
    -1.257641e-08, -1.24909e-08, -1.263138e-08, -1.317918e-08, -1.366246e-08, 
    -1.386312e-08, -1.415625e-08, -1.434524e-08, -1.457391e-08, -1.468143e-08,
  -6.178776e-09, -7.920333e-09, -9.986878e-09, -1.143665e-08, -1.198402e-08, 
    -1.234719e-08, -1.226717e-08, -1.212359e-08, -1.200254e-08, 
    -1.230076e-08, -1.255603e-08, -1.297634e-08, -1.312238e-08, 
    -1.331496e-08, -1.343315e-08,
  -4.074215e-09, -5.528345e-09, -7.420207e-09, -9.50614e-09, -1.108123e-08, 
    -1.196941e-08, -1.22402e-08, -1.203145e-08, -1.1809e-08, -1.167196e-08, 
    -1.184904e-08, -1.188183e-08, -1.220677e-08, -1.216001e-08, -1.213232e-08,
  -2.797163e-09, -3.791371e-09, -5.126615e-09, -6.890072e-09, -8.828984e-09, 
    -1.065868e-08, -1.182811e-08, -1.2031e-08, -1.177404e-08, -1.146775e-08, 
    -1.132451e-08, -1.140478e-08, -1.152606e-08, -1.164803e-08, -1.163361e-08,
  -1.903461e-09, -2.365459e-09, -3.320079e-09, -4.640559e-09, -6.307547e-09, 
    -8.167826e-09, -1.01431e-08, -1.152272e-08, -1.208602e-08, -1.158714e-08, 
    -1.131053e-08, -1.11573e-08, -1.117841e-08, -1.124999e-08, -1.136672e-08,
  -1.673942e-09, -1.785715e-09, -2.085498e-09, -2.862584e-09, -3.845642e-09, 
    -5.412366e-09, -7.376556e-09, -9.371793e-09, -1.100607e-08, 
    -1.190667e-08, -1.169617e-08, -1.1225e-08, -1.08985e-08, -1.086114e-08, 
    -1.090187e-08,
  -4.554447e-09, -6.022688e-09, -7.969177e-09, -9.315591e-09, -1.042454e-08, 
    -1.123382e-08, -1.173549e-08, -1.19108e-08, -1.225572e-08, -1.21939e-08, 
    -1.149096e-08, -9.653957e-09, -8.105029e-09, -7.853416e-09, -8.335136e-09,
  -3.418549e-09, -4.504332e-09, -6.066452e-09, -8.26103e-09, -9.657763e-09, 
    -1.087021e-08, -1.149447e-08, -1.199864e-08, -1.239876e-08, 
    -1.219689e-08, -1.172517e-08, -1.167628e-08, -1.034148e-08, 
    -8.662786e-09, -8.466199e-09,
  -2.715023e-09, -3.522933e-09, -4.778193e-09, -6.529189e-09, -8.8459e-09, 
    -1.024052e-08, -1.120426e-08, -1.181527e-08, -1.241649e-08, 
    -1.277405e-08, -1.247456e-08, -1.154727e-08, -1.083881e-08, 
    -1.060312e-08, -1.119049e-08,
  -2.308973e-09, -2.797639e-09, -3.80469e-09, -5.306028e-09, -7.352326e-09, 
    -9.76145e-09, -1.092662e-08, -1.161915e-08, -1.211152e-08, -1.257441e-08, 
    -1.275059e-08, -1.253097e-08, -1.187805e-08, -1.135803e-08, -1.200594e-08,
  -1.909055e-09, -2.349169e-09, -3.045325e-09, -4.23504e-09, -6.05825e-09, 
    -8.325559e-09, -1.062971e-08, -1.154592e-08, -1.195933e-08, 
    -1.240356e-08, -1.261778e-08, -1.202416e-08, -1.232975e-08, 
    -1.274202e-08, -1.354438e-08,
  -1.682193e-09, -1.973031e-09, -2.568392e-09, -3.438763e-09, -4.871177e-09, 
    -7.055514e-09, -9.466483e-09, -1.135756e-08, -1.199381e-08, -1.22586e-08, 
    -1.269186e-08, -1.249338e-08, -1.225122e-08, -1.303061e-08, -1.348692e-08,
  -1.684076e-09, -1.777791e-09, -2.120968e-09, -2.755782e-09, -3.85729e-09, 
    -5.725376e-09, -8.110231e-09, -1.060672e-08, -1.187149e-08, 
    -1.245294e-08, -1.25982e-08, -1.231751e-08, -1.29911e-08, -1.369664e-08, 
    -1.375006e-08,
  -1.694939e-09, -1.773723e-09, -1.884525e-09, -2.321738e-09, -2.945887e-09, 
    -4.460237e-09, -6.501506e-09, -9.254827e-09, -1.138366e-08, -1.24087e-08, 
    -1.277685e-08, -1.25919e-08, -1.271558e-08, -1.308479e-08, -1.343567e-08,
  -1.609811e-09, -1.650625e-09, -1.793297e-09, -2.022945e-09, -2.491652e-09, 
    -3.313757e-09, -4.977804e-09, -7.427407e-09, -9.992535e-09, 
    -1.229482e-08, -1.304464e-08, -1.285489e-08, -1.272728e-08, 
    -1.265575e-08, -1.339759e-08,
  -1.421048e-09, -1.558037e-09, -1.653832e-09, -1.76232e-09, -2.07018e-09, 
    -2.608674e-09, -3.487126e-09, -5.578439e-09, -8.227754e-09, 
    -1.092066e-08, -1.280998e-08, -1.317135e-08, -1.28528e-08, -1.286287e-08, 
    -1.361615e-08,
  -6.136935e-09, -6.531402e-09, -7.068591e-09, -7.520558e-09, -8.054228e-09, 
    -8.733471e-09, -1.008025e-08, -1.005863e-08, -9.837937e-09, 
    -1.040711e-08, -1.085815e-08, -1.121075e-08, -1.163423e-08, 
    -1.191484e-08, -1.169307e-08,
  -6.13821e-09, -6.306648e-09, -6.699624e-09, -7.277406e-09, -8.02063e-09, 
    -8.616849e-09, -8.8852e-09, -9.853951e-09, -1.003578e-08, -1.045036e-08, 
    -1.141931e-08, -1.201435e-08, -1.224567e-08, -1.216304e-08, -1.14959e-08,
  -6.032889e-09, -6.178285e-09, -6.463096e-09, -6.974717e-09, -7.515003e-09, 
    -8.452691e-09, -8.842767e-09, -9.24266e-09, -9.570032e-09, -1.099468e-08, 
    -1.170045e-08, -1.19711e-08, -1.218343e-08, -1.200172e-08, -1.158745e-08,
  -5.667493e-09, -5.900616e-09, -6.065178e-09, -6.627169e-09, -7.169496e-09, 
    -8.057795e-09, -8.786122e-09, -9.152572e-09, -9.191765e-09, 
    -1.060215e-08, -1.215259e-08, -1.194043e-08, -1.188938e-08, 
    -1.170329e-08, -1.156758e-08,
  -4.934475e-09, -5.328857e-09, -5.651594e-09, -6.004029e-09, -6.465841e-09, 
    -7.262211e-09, -8.012653e-09, -9.031307e-09, -9.113836e-09, 
    -9.604658e-09, -1.182448e-08, -1.207583e-08, -1.194898e-08, -1.16288e-08, 
    -1.15796e-08,
  -4.343364e-09, -4.616398e-09, -4.978684e-09, -5.422256e-09, -5.786587e-09, 
    -6.298274e-09, -7.063673e-09, -8.254047e-09, -8.91074e-09, -9.034111e-09, 
    -1.118071e-08, -1.214558e-08, -1.189955e-08, -1.18781e-08, -1.131616e-08,
  -3.89481e-09, -4.134659e-09, -4.440039e-09, -4.765481e-09, -5.158667e-09, 
    -5.597971e-09, -6.090991e-09, -7.157899e-09, -8.28917e-09, -8.545558e-09, 
    -1.043671e-08, -1.191423e-08, -1.177605e-08, -1.19719e-08, -1.136696e-08,
  -3.476915e-09, -3.670188e-09, -3.941816e-09, -4.183542e-09, -4.522324e-09, 
    -4.944817e-09, -5.395246e-09, -6.163274e-09, -7.261307e-09, 
    -8.163759e-09, -9.62783e-09, -1.145874e-08, -1.178005e-08, -1.186527e-08, 
    -1.1775e-08,
  -2.981984e-09, -3.200665e-09, -3.484776e-09, -3.701371e-09, -3.948924e-09, 
    -4.279095e-09, -4.630171e-09, -5.353489e-09, -6.257773e-09, 
    -7.407633e-09, -8.877236e-09, -1.055168e-08, -1.144551e-08, 
    -1.181662e-08, -1.217913e-08,
  -2.441872e-09, -2.724355e-09, -3.009138e-09, -3.204669e-09, -3.405338e-09, 
    -3.722567e-09, -4.03183e-09, -4.548769e-09, -5.346336e-09, -6.487411e-09, 
    -7.928246e-09, -9.728215e-09, -1.10989e-08, -1.166407e-08, -1.241006e-08,
  -3.55741e-09, -4.224914e-09, -5.051503e-09, -5.846912e-09, -6.421325e-09, 
    -6.978634e-09, -7.408895e-09, -7.673773e-09, -7.759706e-09, -7.78073e-09, 
    -7.676365e-09, -7.578458e-09, -7.458793e-09, -7.485563e-09, -7.614706e-09,
  -2.731796e-09, -3.3419e-09, -4.048977e-09, -4.803684e-09, -5.569586e-09, 
    -6.191576e-09, -6.711462e-09, -7.164186e-09, -7.406741e-09, 
    -7.413492e-09, -7.2955e-09, -7.217103e-09, -7.338365e-09, -7.458818e-09, 
    -7.595107e-09,
  -2.201755e-09, -2.548088e-09, -3.165817e-09, -3.883935e-09, -4.63905e-09, 
    -5.381527e-09, -6.027076e-09, -6.610257e-09, -6.953658e-09, 
    -6.975697e-09, -6.808667e-09, -6.845965e-09, -7.04549e-09, -7.213518e-09, 
    -7.300081e-09,
  -2.000798e-09, -2.166683e-09, -2.481815e-09, -3.08785e-09, -3.791352e-09, 
    -4.545794e-09, -5.393217e-09, -6.027913e-09, -6.548957e-09, 
    -6.643443e-09, -6.840551e-09, -6.774035e-09, -6.781201e-09, 
    -6.927386e-09, -7.120619e-09,
  -1.936309e-09, -2.01118e-09, -2.170565e-09, -2.54411e-09, -3.139361e-09, 
    -3.772993e-09, -4.691322e-09, -5.606982e-09, -6.117685e-09, 
    -6.406875e-09, -6.812908e-09, -6.818401e-09, -6.497687e-09, 
    -6.582198e-09, -7.316536e-09,
  -1.983568e-09, -1.978697e-09, -2.051292e-09, -2.270335e-09, -2.714508e-09, 
    -3.254062e-09, -3.921636e-09, -5.055177e-09, -5.971062e-09, 
    -6.250767e-09, -6.609874e-09, -6.891439e-09, -6.45758e-09, -6.599678e-09, 
    -7.333267e-09,
  -2.051487e-09, -2.081182e-09, -2.069142e-09, -2.17312e-09, -2.42568e-09, 
    -2.897231e-09, -3.415819e-09, -4.337495e-09, -5.748013e-09, 
    -6.180944e-09, -6.459989e-09, -6.982187e-09, -6.764765e-09, 
    -7.016335e-09, -7.87859e-09,
  -2.060376e-09, -2.227305e-09, -2.222148e-09, -2.249549e-09, -2.374079e-09, 
    -2.690065e-09, -3.159812e-09, -3.750796e-09, -5.058661e-09, 
    -6.080439e-09, -6.379629e-09, -7.095454e-09, -7.176399e-09, 
    -7.473727e-09, -8.964904e-09,
  -2.09147e-09, -2.201843e-09, -2.316264e-09, -2.371801e-09, -2.462057e-09, 
    -2.669898e-09, -3.018509e-09, -3.442612e-09, -4.341243e-09, 
    -5.598431e-09, -6.533675e-09, -7.376796e-09, -7.595212e-09, 
    -8.213389e-09, -1.005743e-08,
  -2.153458e-09, -2.295728e-09, -2.37334e-09, -2.428926e-09, -2.492019e-09, 
    -2.733038e-09, -3.11771e-09, -3.401614e-09, -4.029875e-09, -5.098715e-09, 
    -6.162046e-09, -7.660645e-09, -7.945062e-09, -8.860196e-09, -1.123004e-08,
  -2.579374e-09, -3.290577e-09, -4.116768e-09, -5.070314e-09, -6.078655e-09, 
    -7.275922e-09, -8.185599e-09, -8.935682e-09, -9.322474e-09, 
    -9.482378e-09, -9.50515e-09, -9.535167e-09, -9.559713e-09, -9.676888e-09, 
    -9.898327e-09,
  -2.136473e-09, -2.671364e-09, -3.323298e-09, -4.196427e-09, -5.079134e-09, 
    -6.039415e-09, -7.096396e-09, -8.034864e-09, -8.921557e-09, 
    -9.411272e-09, -9.50477e-09, -9.521496e-09, -9.500646e-09, -9.498817e-09, 
    -9.537604e-09,
  -1.800988e-09, -2.222318e-09, -2.747786e-09, -3.466162e-09, -4.306285e-09, 
    -5.21558e-09, -6.155241e-09, -7.097012e-09, -8.002464e-09, -8.882719e-09, 
    -9.428515e-09, -9.582736e-09, -9.554266e-09, -9.574123e-09, -9.546237e-09,
  -1.592739e-09, -1.907854e-09, -2.334341e-09, -2.900086e-09, -3.631445e-09, 
    -4.503211e-09, -5.435089e-09, -6.4108e-09, -7.157436e-09, -8.091437e-09, 
    -8.81248e-09, -9.37874e-09, -9.562774e-09, -9.568318e-09, -9.606447e-09,
  -1.415663e-09, -1.689051e-09, -2.061693e-09, -2.510372e-09, -3.133834e-09, 
    -3.862644e-09, -4.713898e-09, -5.714022e-09, -6.570836e-09, 
    -7.246938e-09, -8.082211e-09, -8.650782e-09, -9.166446e-09, 
    -9.436906e-09, -9.486672e-09,
  -1.493081e-09, -1.485252e-09, -1.772082e-09, -2.189103e-09, -2.739004e-09, 
    -3.471597e-09, -4.187645e-09, -4.942137e-09, -5.912705e-09, 
    -6.725509e-09, -7.347009e-09, -8.038885e-09, -8.418518e-09, 
    -8.921793e-09, -9.085088e-09,
  -1.505569e-09, -1.48512e-09, -1.587417e-09, -1.906629e-09, -2.329556e-09, 
    -3.011291e-09, -3.850577e-09, -4.516423e-09, -5.274716e-09, 
    -6.086212e-09, -6.815039e-09, -7.463417e-09, -8.005877e-09, 
    -8.459371e-09, -8.768382e-09,
  -1.531682e-09, -1.551482e-09, -1.529376e-09, -1.71332e-09, -2.052474e-09, 
    -2.50104e-09, -3.384067e-09, -4.15519e-09, -4.928787e-09, -5.635445e-09, 
    -6.332941e-09, -6.866672e-09, -7.490967e-09, -7.920808e-09, -8.16445e-09,
  -1.641541e-09, -1.514743e-09, -1.552029e-09, -1.593208e-09, -1.849843e-09, 
    -2.172792e-09, -2.793848e-09, -3.671513e-09, -4.519023e-09, 
    -5.235738e-09, -5.913584e-09, -6.370696e-09, -7.157907e-09, 
    -7.403215e-09, -8.221551e-09,
  -1.902529e-09, -1.654364e-09, -1.584952e-09, -1.581988e-09, -1.678081e-09, 
    -1.969022e-09, -2.439908e-09, -3.14369e-09, -4.008758e-09, -4.75301e-09, 
    -5.369739e-09, -5.968916e-09, -6.552044e-09, -7.147556e-09, -7.965113e-09,
  -2.963344e-09, -3.319592e-09, -4.068773e-09, -4.757698e-09, -5.475868e-09, 
    -6.286638e-09, -7.243015e-09, -7.981015e-09, -8.898756e-09, 
    -9.564977e-09, -1.006996e-08, -1.043238e-08, -1.072191e-08, 
    -1.099986e-08, -1.107381e-08,
  -2.48889e-09, -2.715265e-09, -3.105268e-09, -3.85839e-09, -4.556356e-09, 
    -5.401987e-09, -6.260277e-09, -7.239738e-09, -7.933926e-09, 
    -8.821248e-09, -9.391859e-09, -1.009063e-08, -1.04834e-08, -1.069547e-08, 
    -1.083496e-08,
  -2.116771e-09, -2.33168e-09, -2.54647e-09, -2.998116e-09, -3.682712e-09, 
    -4.461602e-09, -5.33009e-09, -6.276437e-09, -7.307313e-09, -7.993879e-09, 
    -8.687596e-09, -9.324202e-09, -9.95318e-09, -1.043157e-08, -1.06744e-08,
  -1.785879e-09, -1.945184e-09, -2.164408e-09, -2.427864e-09, -2.894523e-09, 
    -3.59094e-09, -4.445396e-09, -5.349494e-09, -6.31373e-09, -7.438117e-09, 
    -8.055754e-09, -8.54935e-09, -9.146324e-09, -9.784999e-09, -1.022558e-08,
  -1.606993e-09, -1.690112e-09, -1.846724e-09, -2.022928e-09, -2.31119e-09, 
    -2.802315e-09, -3.479633e-09, -4.440765e-09, -5.363511e-09, 
    -6.387411e-09, -7.459724e-09, -8.078047e-09, -8.478901e-09, 
    -8.911973e-09, -9.497944e-09,
  -1.455186e-09, -1.540498e-09, -1.615125e-09, -1.771917e-09, -1.908959e-09, 
    -2.229118e-09, -2.700436e-09, -3.430842e-09, -4.394095e-09, 
    -5.370678e-09, -6.362794e-09, -7.28136e-09, -7.864422e-09, -8.258632e-09, 
    -8.622903e-09,
  -1.430211e-09, -1.438807e-09, -1.48324e-09, -1.540972e-09, -1.669198e-09, 
    -1.814736e-09, -2.142414e-09, -2.664596e-09, -3.423382e-09, 
    -4.300946e-09, -5.294711e-09, -6.260851e-09, -7.071733e-09, -7.59723e-09, 
    -8.011303e-09,
  -1.572526e-09, -1.469925e-09, -1.439347e-09, -1.46403e-09, -1.490444e-09, 
    -1.601832e-09, -1.739005e-09, -2.113465e-09, -2.666517e-09, 
    -3.401194e-09, -4.148994e-09, -5.041242e-09, -6.068873e-09, 
    -6.756372e-09, -7.278267e-09,
  -1.754677e-09, -1.528907e-09, -1.497966e-09, -1.475326e-09, -1.49179e-09, 
    -1.485181e-09, -1.54321e-09, -1.676994e-09, -2.110715e-09, -2.70022e-09, 
    -3.418356e-09, -3.963851e-09, -4.85037e-09, -5.717125e-09, -6.320749e-09,
  -2.00782e-09, -1.733404e-09, -1.532531e-09, -1.47507e-09, -1.446353e-09, 
    -1.521657e-09, -1.489278e-09, -1.49627e-09, -1.629559e-09, -2.058878e-09, 
    -2.762942e-09, -3.34589e-09, -3.87901e-09, -4.682021e-09, -5.365442e-09,
  -4.859695e-09, -5.304619e-09, -5.788982e-09, -6.154553e-09, -6.49458e-09, 
    -6.767563e-09, -7.102803e-09, -7.449022e-09, -7.832911e-09, 
    -8.197843e-09, -8.576999e-09, -8.844312e-09, -9.361266e-09, 
    -1.005652e-08, -1.075914e-08,
  -4.13754e-09, -4.686066e-09, -5.198129e-09, -5.594476e-09, -5.938246e-09, 
    -6.234283e-09, -6.573838e-09, -6.868369e-09, -7.246357e-09, 
    -7.739257e-09, -8.216769e-09, -8.652244e-09, -8.945391e-09, 
    -9.509619e-09, -1.045864e-08,
  -3.4796e-09, -4.018544e-09, -4.618609e-09, -5.104016e-09, -5.47221e-09, 
    -5.779907e-09, -6.119949e-09, -6.43425e-09, -6.772753e-09, -7.193874e-09, 
    -7.797539e-09, -8.315086e-09, -8.7087e-09, -9.004704e-09, -9.948551e-09,
  -2.720446e-09, -3.300953e-09, -3.895444e-09, -4.519002e-09, -5.026229e-09, 
    -5.368368e-09, -5.679318e-09, -6.028347e-09, -6.342733e-09, 
    -6.682916e-09, -7.208029e-09, -7.901347e-09, -8.548871e-09, 
    -8.760772e-09, -9.321401e-09,
  -2.043073e-09, -2.589552e-09, -3.213999e-09, -3.818957e-09, -4.467371e-09, 
    -4.986021e-09, -5.349493e-09, -5.658603e-09, -6.029306e-09, 
    -6.310734e-09, -6.599406e-09, -7.205279e-09, -8.074049e-09, 
    -8.688056e-09, -8.929227e-09,
  -1.448898e-09, -1.917559e-09, -2.477039e-09, -3.141434e-09, -3.804617e-09, 
    -4.458959e-09, -4.948022e-09, -5.295537e-09, -5.562805e-09, 
    -6.006283e-09, -6.280779e-09, -6.601725e-09, -7.37678e-09, -8.364196e-09, 
    -8.722114e-09,
  -1.07868e-09, -1.397662e-09, -1.818592e-09, -2.359771e-09, -3.106047e-09, 
    -3.832652e-09, -4.4786e-09, -4.860609e-09, -5.216733e-09, -5.528588e-09, 
    -6.036755e-09, -6.361727e-09, -6.826346e-09, -7.918846e-09, -8.584978e-09,
  -8.466602e-10, -1.060718e-09, -1.349599e-09, -1.788876e-09, -2.327858e-09, 
    -3.098222e-09, -3.923091e-09, -4.495667e-09, -4.811294e-09, 
    -5.101857e-09, -5.494252e-09, -5.979273e-09, -6.472322e-09, 
    -7.408534e-09, -8.350786e-09,
  -7.265044e-10, -8.369552e-10, -1.07711e-09, -1.38633e-09, -1.849309e-09, 
    -2.346466e-09, -3.10251e-09, -3.983923e-09, -4.498446e-09, -4.768701e-09, 
    -5.131324e-09, -5.55896e-09, -5.950447e-09, -6.764812e-09, -7.973336e-09,
  -8.432491e-10, -7.880645e-10, -8.547894e-10, -1.111197e-09, -1.426446e-09, 
    -1.962375e-09, -2.461079e-09, -3.250985e-09, -4.073985e-09, 
    -4.345607e-09, -4.675303e-09, -5.191783e-09, -5.596029e-09, 
    -6.053656e-09, -7.096479e-09,
  -9.885976e-10, -1.193867e-09, -1.582174e-09, -2.191967e-09, -2.816408e-09, 
    -3.627912e-09, -4.734598e-09, -6.116339e-09, -7.546121e-09, 
    -8.668754e-09, -9.615203e-09, -1.031974e-08, -1.094323e-08, 
    -1.149728e-08, -1.199319e-08,
  -8.540512e-10, -1.013609e-09, -1.232616e-09, -1.685105e-09, -2.299926e-09, 
    -3.042928e-09, -3.901689e-09, -5.045552e-09, -6.368067e-09, 
    -7.751839e-09, -8.949137e-09, -9.832632e-09, -1.051965e-08, 
    -1.105519e-08, -1.141439e-08,
  -7.580523e-10, -8.689901e-10, -1.03206e-09, -1.339974e-09, -1.847313e-09, 
    -2.537991e-09, -3.322405e-09, -4.237145e-09, -5.377363e-09, 
    -6.728395e-09, -8.153958e-09, -9.315213e-09, -1.006689e-08, 
    -1.063442e-08, -1.102814e-08,
  -7.070528e-10, -7.603596e-10, -8.705143e-10, -1.081059e-09, -1.482699e-09, 
    -2.089366e-09, -2.874684e-09, -3.711957e-09, -4.677774e-09, 
    -5.881425e-09, -7.284734e-09, -8.696693e-09, -9.652932e-09, 
    -1.027821e-08, -1.072166e-08,
  -7.386067e-10, -7.211429e-10, -7.98154e-10, -9.449521e-10, -1.221482e-09, 
    -1.727921e-09, -2.441483e-09, -3.305432e-09, -4.182934e-09, 
    -5.248712e-09, -6.51312e-09, -7.976797e-09, -9.147413e-09, -9.947258e-09, 
    -1.042329e-08,
  -9.052809e-10, -7.435966e-10, -7.466663e-10, -8.669788e-10, -1.05653e-09, 
    -1.437682e-09, -2.069995e-09, -2.948314e-09, -3.824277e-09, 
    -4.802357e-09, -5.885936e-09, -7.31414e-09, -8.636571e-09, -9.669714e-09, 
    -1.025291e-08,
  -9.553012e-10, -9.272238e-10, -7.776446e-10, -8.334047e-10, -9.720881e-10, 
    -1.237612e-09, -1.740924e-09, -2.598233e-09, -3.524335e-09, -4.50527e-09, 
    -5.515093e-09, -6.735414e-09, -8.114468e-09, -9.261707e-09, -1.006175e-08,
  -8.917466e-10, -9.124749e-10, -8.995695e-10, -8.240896e-10, -9.415502e-10, 
    -1.145196e-09, -1.526108e-09, -2.276766e-09, -3.243644e-09, 
    -4.239836e-09, -5.293949e-09, -6.408458e-09, -7.71666e-09, -8.8578e-09, 
    -9.687107e-09,
  -7.962285e-10, -8.734752e-10, -8.889305e-10, -9.016518e-10, -8.984168e-10, 
    -1.051449e-09, -1.347142e-09, -2.018517e-09, -3.00051e-09, -4.047469e-09, 
    -5.167407e-09, -6.234967e-09, -7.39516e-09, -8.493727e-09, -9.296983e-09,
  -6.862735e-10, -7.471474e-10, -8.66594e-10, -8.89293e-10, -9.346486e-10, 
    -1.025924e-09, -1.230601e-09, -1.732407e-09, -2.72663e-09, -3.867455e-09, 
    -5.06365e-09, -6.194097e-09, -7.295214e-09, -8.349191e-09, -9.078946e-09,
  -2.868332e-09, -3.225982e-09, -3.550686e-09, -3.881758e-09, -4.257814e-09, 
    -4.704302e-09, -5.335961e-09, -6.495409e-09, -8.024686e-09, 
    -9.342108e-09, -1.064539e-08, -1.200259e-08, -1.328059e-08, 
    -1.435778e-08, -1.499771e-08,
  -2.068916e-09, -2.408397e-09, -2.742667e-09, -3.063084e-09, -3.365846e-09, 
    -3.687452e-09, -4.091147e-09, -4.667611e-09, -5.767234e-09, 
    -7.223058e-09, -8.710426e-09, -1.029648e-08, -1.182906e-08, 
    -1.327944e-08, -1.436692e-08,
  -1.509688e-09, -1.734016e-09, -1.985541e-09, -2.276495e-09, -2.582799e-09, 
    -2.876013e-09, -3.174359e-09, -3.531903e-09, -4.097716e-09, -5.23052e-09, 
    -6.681288e-09, -8.316424e-09, -1.016565e-08, -1.192896e-08, -1.3536e-08,
  -1.402145e-09, -1.410362e-09, -1.522777e-09, -1.692919e-09, -1.936811e-09, 
    -2.174635e-09, -2.425066e-09, -2.6813e-09, -3.042302e-09, -3.664181e-09, 
    -4.772452e-09, -6.373306e-09, -8.218659e-09, -1.01864e-08, -1.20454e-08,
  -1.377862e-09, -1.286229e-09, -1.292084e-09, -1.348956e-09, -1.462065e-09, 
    -1.639437e-09, -1.829316e-09, -2.008571e-09, -2.239608e-09, 
    -2.626398e-09, -3.350048e-09, -4.592181e-09, -6.316294e-09, -8.43584e-09, 
    -1.054696e-08,
  -1.440873e-09, -1.310266e-09, -1.1968e-09, -1.168038e-09, -1.186161e-09, 
    -1.259252e-09, -1.396537e-09, -1.538537e-09, -1.701227e-09, -1.9067e-09, 
    -2.344468e-09, -3.321266e-09, -4.823788e-09, -6.790199e-09, -9.26238e-09,
  -1.416333e-09, -1.398916e-09, -1.271773e-09, -1.142995e-09, -1.052902e-09, 
    -1.030127e-09, -1.080717e-09, -1.194019e-09, -1.343384e-09, 
    -1.485267e-09, -1.751476e-09, -2.446785e-09, -3.800548e-09, 
    -5.637174e-09, -8.202832e-09,
  -1.313964e-09, -1.390891e-09, -1.344126e-09, -1.165454e-09, -1.056293e-09, 
    -9.879432e-10, -9.617319e-10, -1.035501e-09, -1.145761e-09, 
    -1.312938e-09, -1.511597e-09, -1.959209e-09, -3.075144e-09, 
    -4.886784e-09, -7.475922e-09,
  -1.18617e-09, -1.296353e-09, -1.334346e-09, -1.233856e-09, -1.016498e-09, 
    -9.337439e-10, -8.944616e-10, -8.936021e-10, -9.442316e-10, 
    -1.062809e-09, -1.3489e-09, -1.72971e-09, -2.695618e-09, -4.394294e-09, 
    -6.94787e-09,
  -9.694542e-10, -1.186945e-09, -1.27191e-09, -1.300815e-09, -1.235614e-09, 
    -1.080054e-09, -1.019436e-09, -1.041043e-09, -1.018363e-09, 
    -1.063813e-09, -1.179959e-09, -1.550258e-09, -2.469945e-09, 
    -4.117898e-09, -6.630473e-09,
  -1.086765e-08, -1.147582e-08, -1.196013e-08, -1.192184e-08, -1.152395e-08, 
    -1.14906e-08, -1.157084e-08, -1.208251e-08, -1.252617e-08, -1.275613e-08, 
    -1.26941e-08, -1.271157e-08, -1.262828e-08, -1.260461e-08, -1.26235e-08,
  -9.415331e-09, -1.051491e-08, -1.105709e-08, -1.16075e-08, -1.176621e-08, 
    -1.149492e-08, -1.109951e-08, -1.06142e-08, -1.039621e-08, -1.067796e-08, 
    -1.103417e-08, -1.136199e-08, -1.141583e-08, -1.140402e-08, -1.154282e-08,
  -7.681787e-09, -8.87305e-09, -9.875035e-09, -1.062201e-08, -1.133512e-08, 
    -1.158662e-08, -1.147334e-08, -1.123834e-08, -1.080615e-08, 
    -1.056513e-08, -1.017041e-08, -9.865205e-09, -9.856507e-09, 
    -1.005231e-08, -1.024091e-08,
  -6.555769e-09, -7.490288e-09, -8.516213e-09, -9.390991e-09, -1.005292e-08, 
    -1.070722e-08, -1.113605e-08, -1.132542e-08, -1.140453e-08, 
    -1.123115e-08, -1.085202e-08, -1.024946e-08, -9.864711e-09, 
    -9.718031e-09, -9.737816e-09,
  -5.147487e-09, -6.32911e-09, -7.238417e-09, -8.118779e-09, -8.974455e-09, 
    -9.601052e-09, -1.041604e-08, -1.099233e-08, -1.13051e-08, -1.129094e-08, 
    -1.101971e-08, -1.051934e-08, -1.017663e-08, -9.943217e-09, -9.810138e-09,
  -3.904018e-09, -5.042897e-09, -6.146758e-09, -6.922749e-09, -7.722281e-09, 
    -8.471108e-09, -9.251425e-09, -1.003096e-08, -1.045508e-08, 
    -1.067001e-08, -1.078891e-08, -1.0668e-08, -1.03877e-08, -1.011553e-08, 
    -9.835817e-09,
  -2.733271e-09, -3.793709e-09, -5.001377e-09, -5.956724e-09, -6.460273e-09, 
    -7.120179e-09, -7.870142e-09, -8.509461e-09, -9.049356e-09, 
    -9.571145e-09, -1.012034e-08, -1.046762e-08, -1.042229e-08, 
    -1.018755e-08, -9.63883e-09,
  -1.911198e-09, -2.608714e-09, -3.726524e-09, -4.919145e-09, -5.515892e-09, 
    -5.914626e-09, -6.528253e-09, -7.23776e-09, -7.927816e-09, -8.77203e-09, 
    -9.393327e-09, -9.85237e-09, -9.993821e-09, -9.887799e-09, -9.37208e-09,
  -1.300279e-09, -1.688805e-09, -2.548582e-09, -3.745895e-09, -4.932748e-09, 
    -5.109155e-09, -5.417316e-09, -6.100568e-09, -6.810078e-09, 
    -8.041841e-09, -8.922489e-09, -9.274658e-09, -9.361867e-09, 
    -9.281345e-09, -8.828218e-09,
  -1.166873e-09, -1.265268e-09, -1.558959e-09, -2.533566e-09, -4.004062e-09, 
    -4.611322e-09, -4.671325e-09, -5.035093e-09, -6.029345e-09, 
    -7.391896e-09, -8.198976e-09, -8.555126e-09, -8.816815e-09, 
    -8.978359e-09, -8.671267e-09,
  -1.47189e-08, -1.611702e-08, -1.72884e-08, -1.823846e-08, -1.802917e-08, 
    -1.668829e-08, -1.525124e-08, -1.404964e-08, -1.381968e-08, 
    -1.398584e-08, -1.45516e-08, -1.526413e-08, -1.603821e-08, -1.66042e-08, 
    -1.681841e-08,
  -1.370325e-08, -1.510955e-08, -1.621657e-08, -1.741089e-08, -1.806151e-08, 
    -1.756502e-08, -1.714712e-08, -1.660387e-08, -1.635128e-08, 
    -1.626879e-08, -1.65637e-08, -1.695615e-08, -1.746042e-08, -1.784079e-08, 
    -1.835581e-08,
  -1.264369e-08, -1.439724e-08, -1.552254e-08, -1.643207e-08, -1.735444e-08, 
    -1.732743e-08, -1.718249e-08, -1.705139e-08, -1.693226e-08, 
    -1.701511e-08, -1.70603e-08, -1.736735e-08, -1.789724e-08, -1.853354e-08, 
    -1.911686e-08,
  -1.149008e-08, -1.33539e-08, -1.495902e-08, -1.579629e-08, -1.670289e-08, 
    -1.682236e-08, -1.670665e-08, -1.655776e-08, -1.64304e-08, -1.62331e-08, 
    -1.600149e-08, -1.577831e-08, -1.582116e-08, -1.621578e-08, -1.687908e-08,
  -1.018423e-08, -1.220022e-08, -1.412496e-08, -1.538664e-08, -1.56367e-08, 
    -1.609886e-08, -1.609373e-08, -1.556268e-08, -1.555186e-08, 
    -1.519602e-08, -1.513506e-08, -1.488511e-08, -1.484218e-08, 
    -1.483919e-08, -1.51887e-08,
  -8.891523e-09, -1.09068e-08, -1.302499e-08, -1.490598e-08, -1.516374e-08, 
    -1.538533e-08, -1.537977e-08, -1.520175e-08, -1.483381e-08, 
    -1.456827e-08, -1.417319e-08, -1.408384e-08, -1.373235e-08, 
    -1.383627e-08, -1.397623e-08,
  -7.347456e-09, -9.687673e-09, -1.168725e-08, -1.388813e-08, -1.509527e-08, 
    -1.497115e-08, -1.488159e-08, -1.487151e-08, -1.435275e-08, 
    -1.383786e-08, -1.354766e-08, -1.348078e-08, -1.350686e-08, -1.35257e-08, 
    -1.373996e-08,
  -5.618861e-09, -8.289251e-09, -1.054642e-08, -1.222708e-08, -1.410607e-08, 
    -1.440385e-08, -1.448088e-08, -1.43789e-08, -1.388121e-08, -1.325358e-08, 
    -1.286949e-08, -1.315685e-08, -1.339955e-08, -1.329266e-08, -1.286528e-08,
  -3.775095e-09, -6.480007e-09, -9.497938e-09, -1.136271e-08, -1.290746e-08, 
    -1.37202e-08, -1.398087e-08, -1.352841e-08, -1.301104e-08, -1.224934e-08, 
    -1.162977e-08, -1.162235e-08, -1.067076e-08, -9.914063e-09, -9.410476e-09,
  -2.580272e-09, -4.667097e-09, -7.81126e-09, -1.026765e-08, -1.198303e-08, 
    -1.326318e-08, -1.345932e-08, -1.294927e-08, -1.197482e-08, 
    -1.097325e-08, -1.126002e-08, -1.014528e-08, -9.331329e-09, -8.57766e-09, 
    -8.232752e-09,
  -1.198299e-08, -1.222305e-08, -1.301499e-08, -1.383799e-08, -1.464173e-08, 
    -1.540008e-08, -1.616915e-08, -1.646897e-08, -1.668182e-08, 
    -1.628804e-08, -1.589508e-08, -1.531243e-08, -1.479323e-08, -1.43875e-08, 
    -1.414512e-08,
  -1.197874e-08, -1.216846e-08, -1.257834e-08, -1.349239e-08, -1.457946e-08, 
    -1.546696e-08, -1.653577e-08, -1.69975e-08, -1.714415e-08, -1.693791e-08, 
    -1.652656e-08, -1.616302e-08, -1.575201e-08, -1.533451e-08, -1.490798e-08,
  -1.197168e-08, -1.209853e-08, -1.24735e-08, -1.286957e-08, -1.399581e-08, 
    -1.511058e-08, -1.616336e-08, -1.712743e-08, -1.773849e-08, 
    -1.812022e-08, -1.816552e-08, -1.829111e-08, -1.816926e-08, 
    -1.815179e-08, -1.789122e-08,
  -1.168007e-08, -1.210383e-08, -1.250529e-08, -1.275824e-08, -1.350546e-08, 
    -1.460678e-08, -1.570214e-08, -1.672036e-08, -1.748657e-08, 
    -1.800558e-08, -1.842998e-08, -1.875532e-08, -1.903109e-08, 
    -1.917006e-08, -1.918542e-08,
  -1.105911e-08, -1.19359e-08, -1.240924e-08, -1.282993e-08, -1.334873e-08, 
    -1.41408e-08, -1.533645e-08, -1.626973e-08, -1.702229e-08, -1.765363e-08, 
    -1.825275e-08, -1.852243e-08, -1.871678e-08, -1.853164e-08, -1.833685e-08,
  -1.04543e-08, -1.13801e-08, -1.234802e-08, -1.273291e-08, -1.317385e-08, 
    -1.386322e-08, -1.456099e-08, -1.560901e-08, -1.65445e-08, -1.76449e-08, 
    -1.803355e-08, -1.843037e-08, -1.8028e-08, -1.765904e-08, -1.703437e-08,
  -9.80221e-09, -1.057849e-08, -1.188776e-08, -1.269759e-08, -1.304668e-08, 
    -1.380002e-08, -1.449325e-08, -1.564591e-08, -1.654191e-08, 
    -1.719878e-08, -1.745674e-08, -1.737677e-08, -1.643126e-08, 
    -1.617672e-08, -1.560251e-08,
  -8.932751e-09, -9.942959e-09, -1.098391e-08, -1.206714e-08, -1.282059e-08, 
    -1.368986e-08, -1.463894e-08, -1.56595e-08, -1.613921e-08, -1.671147e-08, 
    -1.665704e-08, -1.592015e-08, -1.526401e-08, -1.449819e-08, -1.348455e-08,
  -7.927311e-09, -9.118215e-09, -1.028874e-08, -1.145871e-08, -1.252125e-08, 
    -1.323951e-08, -1.460299e-08, -1.514325e-08, -1.54951e-08, -1.594624e-08, 
    -1.554704e-08, -1.527482e-08, -1.366499e-08, -1.241594e-08, -1.120515e-08,
  -6.769428e-09, -8.231194e-09, -9.358956e-09, -1.057112e-08, -1.21049e-08, 
    -1.329099e-08, -1.488143e-08, -1.489176e-08, -1.514282e-08, 
    -1.516181e-08, -1.482112e-08, -1.443388e-08, -1.30018e-08, -1.11975e-08, 
    -1.019916e-08,
  -1.078483e-08, -1.105142e-08, -1.128972e-08, -1.14855e-08, -1.155684e-08, 
    -1.162674e-08, -1.165394e-08, -1.172217e-08, -1.189565e-08, 
    -1.217107e-08, -1.251691e-08, -1.291829e-08, -1.326191e-08, 
    -1.369689e-08, -1.423481e-08,
  -1.089604e-08, -1.101648e-08, -1.128323e-08, -1.145294e-08, -1.140743e-08, 
    -1.142438e-08, -1.147462e-08, -1.155432e-08, -1.179722e-08, 
    -1.213049e-08, -1.26467e-08, -1.321915e-08, -1.396451e-08, -1.448409e-08, 
    -1.501903e-08,
  -1.128696e-08, -1.115432e-08, -1.133497e-08, -1.157529e-08, -1.153793e-08, 
    -1.138205e-08, -1.140706e-08, -1.156968e-08, -1.196104e-08, 
    -1.252093e-08, -1.342646e-08, -1.414844e-08, -1.497218e-08, 
    -1.552831e-08, -1.594863e-08,
  -1.102859e-08, -1.144311e-08, -1.148732e-08, -1.156342e-08, -1.155048e-08, 
    -1.137955e-08, -1.143359e-08, -1.179351e-08, -1.230608e-08, 
    -1.339098e-08, -1.421362e-08, -1.494467e-08, -1.531176e-08, 
    -1.552569e-08, -1.533062e-08,
  -1.00277e-08, -1.097148e-08, -1.144354e-08, -1.153027e-08, -1.152374e-08, 
    -1.156649e-08, -1.16554e-08, -1.210884e-08, -1.337514e-08, -1.413297e-08, 
    -1.467525e-08, -1.542453e-08, -1.590596e-08, -1.539771e-08, -1.485644e-08,
  -9.187246e-09, -1.020963e-08, -1.111595e-08, -1.141791e-08, -1.146231e-08, 
    -1.169365e-08, -1.179582e-08, -1.285346e-08, -1.437244e-08, 
    -1.395266e-08, -1.514896e-08, -1.626347e-08, -1.48124e-08, -1.356173e-08, 
    -1.28838e-08,
  -8.151353e-09, -9.328606e-09, -1.059249e-08, -1.132425e-08, -1.156247e-08, 
    -1.179912e-08, -1.198476e-08, -1.325306e-08, -1.434755e-08, 
    -1.357731e-08, -1.56241e-08, -1.492121e-08, -1.177062e-08, -1.058755e-08, 
    -1.048172e-08,
  -7.268044e-09, -8.440116e-09, -9.76674e-09, -1.081589e-08, -1.143234e-08, 
    -1.18853e-08, -1.247357e-08, -1.324466e-08, -1.359085e-08, -1.332137e-08, 
    -1.480557e-08, -1.363908e-08, -1.098985e-08, -1.052061e-08, -1.130874e-08,
  -6.585755e-09, -7.631408e-09, -9.057357e-09, -1.040684e-08, -1.125103e-08, 
    -1.149046e-08, -1.243915e-08, -1.34982e-08, -1.348776e-08, -1.336551e-08, 
    -1.395182e-08, -1.291548e-08, -1.256395e-08, -1.262702e-08, -1.398229e-08,
  -5.886606e-09, -7.087369e-09, -8.252858e-09, -9.622771e-09, -1.091305e-08, 
    -1.181234e-08, -1.243422e-08, -1.339518e-08, -1.332829e-08, 
    -1.392492e-08, -1.357423e-08, -1.346231e-08, -1.561104e-08, 
    -1.443263e-08, -1.349064e-08,
  -1.102783e-08, -1.163493e-08, -1.235903e-08, -1.262632e-08, -1.226219e-08, 
    -1.125828e-08, -1.109424e-08, -1.133039e-08, -1.153746e-08, 
    -1.192725e-08, -1.268088e-08, -1.44057e-08, -1.476463e-08, -1.545996e-08, 
    -1.648209e-08,
  -1.008469e-08, -1.104432e-08, -1.176761e-08, -1.226323e-08, -1.237479e-08, 
    -1.258281e-08, -1.214805e-08, -1.172182e-08, -1.1355e-08, -1.151076e-08, 
    -1.13918e-08, -1.189448e-08, -1.331885e-08, -1.424165e-08, -1.487583e-08,
  -8.387127e-09, -9.772685e-09, -1.057786e-08, -1.119293e-08, -1.178734e-08, 
    -1.20433e-08, -1.223081e-08, -1.236394e-08, -1.181612e-08, -1.161271e-08, 
    -1.13158e-08, -1.154984e-08, -1.20683e-08, -1.313436e-08, -1.42266e-08,
  -6.542572e-09, -8.056627e-09, -9.435282e-09, -1.026724e-08, -1.111188e-08, 
    -1.166147e-08, -1.165296e-08, -1.203168e-08, -1.186919e-08, 
    -1.197569e-08, -1.203052e-08, -1.208098e-08, -1.227694e-08, 
    -1.253305e-08, -1.308073e-08,
  -5.019085e-09, -6.211552e-09, -7.676787e-09, -8.961536e-09, -1.023752e-08, 
    -1.112538e-08, -1.120236e-08, -1.149214e-08, -1.166171e-08, 
    -1.147779e-08, -1.186979e-08, -1.232509e-08, -1.24794e-08, -1.261028e-08, 
    -1.263046e-08,
  -4.000264e-09, -4.713594e-09, -5.904439e-09, -7.300272e-09, -8.751126e-09, 
    -1.028805e-08, -1.097975e-08, -1.107901e-08, -1.156972e-08, 
    -1.165874e-08, -1.162975e-08, -1.164816e-08, -1.190595e-08, -1.2612e-08, 
    -1.298621e-08,
  -3.263098e-09, -3.801296e-09, -4.584906e-09, -5.678773e-09, -7.089021e-09, 
    -8.827309e-09, -1.040672e-08, -1.068701e-08, -1.132701e-08, 
    -1.175103e-08, -1.161071e-08, -1.15095e-08, -1.138706e-08, -1.209806e-08, 
    -1.242486e-08,
  -2.629038e-09, -3.113729e-09, -3.738966e-09, -4.611729e-09, -5.70111e-09, 
    -7.264569e-09, -9.256381e-09, -1.036035e-08, -1.109766e-08, 
    -1.162796e-08, -1.150944e-08, -1.129027e-08, -1.143074e-08, 
    -1.152117e-08, -1.241358e-08,
  -2.309495e-09, -2.531825e-09, -3.027359e-09, -3.768886e-09, -4.792305e-09, 
    -5.971007e-09, -7.913397e-09, -9.597692e-09, -1.069458e-08, 
    -1.148884e-08, -1.158859e-08, -1.144902e-08, -1.147218e-08, 
    -1.147779e-08, -1.251732e-08,
  -2.092608e-09, -2.174724e-09, -2.507768e-09, -3.088295e-09, -3.867548e-09, 
    -5.012084e-09, -6.666803e-09, -8.685602e-09, -1.020745e-08, 
    -1.115696e-08, -1.154974e-08, -1.153712e-08, -1.1999e-08, -1.237439e-08, 
    -1.337373e-08,
  -4.973361e-09, -5.462895e-09, -6.046703e-09, -6.929755e-09, -7.887342e-09, 
    -8.795908e-09, -9.513472e-09, -1.04507e-08, -1.124832e-08, -1.191254e-08, 
    -1.31242e-08, -1.415921e-08, -1.430304e-08, -1.459135e-08, -1.528771e-08,
  -4.248356e-09, -4.73604e-09, -5.295087e-09, -6.075056e-09, -7.050878e-09, 
    -8.004723e-09, -8.816646e-09, -9.778435e-09, -1.057341e-08, 
    -1.125741e-08, -1.19387e-08, -1.307426e-08, -1.403639e-08, -1.487382e-08, 
    -1.510618e-08,
  -3.822434e-09, -4.215603e-09, -4.628735e-09, -5.259108e-09, -6.101911e-09, 
    -7.091304e-09, -8.050831e-09, -9.102343e-09, -1.004518e-08, 
    -1.082237e-08, -1.132492e-08, -1.211844e-08, -1.314236e-08, 
    -1.421976e-08, -1.522618e-08,
  -3.61067e-09, -3.832211e-09, -4.110386e-09, -4.539281e-09, -5.259849e-09, 
    -6.156261e-09, -7.28372e-09, -8.273808e-09, -9.237629e-09, -1.014369e-08, 
    -1.086299e-08, -1.155317e-08, -1.237143e-08, -1.325645e-08, -1.432753e-08,
  -3.449186e-09, -3.712191e-09, -3.822141e-09, -4.191809e-09, -4.707904e-09, 
    -5.351467e-09, -6.516783e-09, -7.370105e-09, -8.117586e-09, 
    -9.177658e-09, -1.026579e-08, -1.095265e-08, -1.180058e-08, 
    -1.247337e-08, -1.31497e-08,
  -3.382835e-09, -3.508084e-09, -3.630493e-09, -3.82111e-09, -4.210579e-09, 
    -4.763288e-09, -5.619318e-09, -6.664218e-09, -7.287532e-09, 
    -8.148033e-09, -9.214703e-09, -1.018972e-08, -1.111625e-08, 
    -1.191502e-08, -1.241809e-08,
  -3.420235e-09, -3.554341e-09, -3.591176e-09, -3.626945e-09, -3.869763e-09, 
    -4.324204e-09, -4.973074e-09, -5.862378e-09, -6.70576e-09, -7.497013e-09, 
    -8.483661e-09, -9.304973e-09, -1.030113e-08, -1.133893e-08, -1.202716e-08,
  -2.952557e-09, -3.310727e-09, -3.51841e-09, -3.536777e-09, -3.579439e-09, 
    -4.039493e-09, -4.574944e-09, -5.349491e-09, -6.112004e-09, 
    -6.949594e-09, -7.90754e-09, -8.626198e-09, -9.571805e-09, -1.058239e-08, 
    -1.153799e-08,
  -2.288759e-09, -2.677914e-09, -3.085775e-09, -3.317675e-09, -3.415363e-09, 
    -3.650283e-09, -4.209809e-09, -4.771713e-09, -5.804515e-09, -6.49873e-09, 
    -7.457322e-09, -8.06468e-09, -8.928042e-09, -9.857184e-09, -1.086061e-08,
  -1.646891e-09, -2.024084e-09, -2.409414e-09, -2.797269e-09, -2.972564e-09, 
    -3.245431e-09, -3.868343e-09, -4.353435e-09, -5.132859e-09, 
    -6.102623e-09, -6.991163e-09, -7.775523e-09, -8.42632e-09, -9.356004e-09, 
    -1.027793e-08,
  -3.166317e-09, -3.394895e-09, -3.571812e-09, -3.691989e-09, -3.922115e-09, 
    -4.245668e-09, -4.667578e-09, -5.055143e-09, -5.395211e-09, 
    -5.642141e-09, -5.918563e-09, -6.369142e-09, -6.916959e-09, 
    -7.443491e-09, -8.058448e-09,
  -2.360996e-09, -2.630547e-09, -2.932136e-09, -3.216588e-09, -3.465632e-09, 
    -3.718915e-09, -4.014892e-09, -4.416116e-09, -4.922797e-09, 
    -5.393785e-09, -5.657577e-09, -5.989213e-09, -6.587115e-09, 
    -7.326767e-09, -8.160937e-09,
  -1.857065e-09, -2.116261e-09, -2.371868e-09, -2.681706e-09, -3.035286e-09, 
    -3.355359e-09, -3.679606e-09, -4.041079e-09, -4.472537e-09, 
    -4.975167e-09, -5.471819e-09, -5.860883e-09, -6.271919e-09, 
    -6.982049e-09, -8.149827e-09,
  -1.420197e-09, -1.631657e-09, -1.860318e-09, -2.141283e-09, -2.449328e-09, 
    -2.794607e-09, -3.202228e-09, -3.678929e-09, -4.197866e-09, 
    -4.712214e-09, -5.14286e-09, -5.704837e-09, -6.262309e-09, -6.932458e-09, 
    -7.977464e-09,
  -1.113732e-09, -1.33882e-09, -1.565305e-09, -1.820257e-09, -2.105504e-09, 
    -2.420442e-09, -2.766042e-09, -3.162846e-09, -3.678103e-09, 
    -4.375631e-09, -4.923615e-09, -5.38889e-09, -6.094863e-09, -6.935116e-09, 
    -8.050204e-09,
  -8.081089e-10, -9.837213e-10, -1.226096e-09, -1.49924e-09, -1.822735e-09, 
    -2.163494e-09, -2.496155e-09, -2.874211e-09, -3.270275e-09, 
    -3.875915e-09, -4.579481e-09, -5.133989e-09, -5.77806e-09, -6.771058e-09, 
    -7.963853e-09,
  -6.218966e-10, -7.677982e-10, -9.475032e-10, -1.177734e-09, -1.490766e-09, 
    -1.864112e-09, -2.256011e-09, -2.630041e-09, -3.012667e-09, 
    -3.496742e-09, -4.153504e-09, -4.849183e-09, -5.466374e-09, 
    -6.440969e-09, -7.769066e-09,
  -5.640948e-10, -6.537628e-10, -7.471733e-10, -9.156759e-10, -1.200155e-09, 
    -1.573109e-09, -1.982626e-09, -2.421255e-09, -2.826555e-09, 
    -3.270414e-09, -3.808344e-09, -4.481767e-09, -5.206495e-09, 
    -6.098329e-09, -7.476713e-09,
  -4.917102e-10, -5.79946e-10, -6.824126e-10, -7.745417e-10, -9.679436e-10, 
    -1.295276e-09, -1.682104e-09, -2.124977e-09, -2.597763e-09, 
    -3.098536e-09, -3.613795e-09, -4.214882e-09, -4.866904e-09, 
    -5.662869e-09, -7.103483e-09,
  -2.968648e-10, -4.106391e-10, -6.197083e-10, -7.976138e-10, -9.296369e-10, 
    -1.105325e-09, -1.429383e-09, -1.849324e-09, -2.35049e-09, -2.871405e-09, 
    -3.448488e-09, -4.021965e-09, -4.693028e-09, -5.324388e-09, -6.565009e-09,
  -4.133331e-09, -4.503541e-09, -4.917388e-09, -5.4272e-09, -5.836799e-09, 
    -6.365768e-09, -6.676194e-09, -6.972823e-09, -7.2102e-09, -7.410926e-09, 
    -7.715665e-09, -7.916404e-09, -8.163183e-09, -8.147221e-09, -8.237016e-09,
  -2.520276e-09, -2.87042e-09, -3.266321e-09, -3.745201e-09, -4.21025e-09, 
    -4.713509e-09, -5.16216e-09, -5.549337e-09, -5.937247e-09, -6.254397e-09, 
    -6.568933e-09, -6.934918e-09, -7.199044e-09, -7.338542e-09, -7.476141e-09,
  -1.54859e-09, -1.723567e-09, -1.953567e-09, -2.245654e-09, -2.636843e-09, 
    -3.080002e-09, -3.616573e-09, -4.10163e-09, -4.592362e-09, -5.058159e-09, 
    -5.467171e-09, -5.909333e-09, -6.306884e-09, -6.621051e-09, -6.865889e-09,
  -1.04016e-09, -1.145188e-09, -1.268595e-09, -1.414312e-09, -1.596074e-09, 
    -1.845003e-09, -2.17687e-09, -2.614821e-09, -3.107858e-09, -3.658221e-09, 
    -4.197808e-09, -4.731299e-09, -5.307551e-09, -5.741556e-09, -6.12074e-09,
  -6.903838e-10, -7.707277e-10, -8.715502e-10, -9.771349e-10, -1.097497e-09, 
    -1.239411e-09, -1.422413e-09, -1.657101e-09, -2.008786e-09, 
    -2.405121e-09, -2.930588e-09, -3.508955e-09, -4.166095e-09, 
    -4.752289e-09, -5.268687e-09,
  -3.858477e-10, -4.401031e-10, -5.195822e-10, -5.9533e-10, -6.903789e-10, 
    -7.92352e-10, -9.30626e-10, -1.100855e-09, -1.334833e-09, -1.617869e-09, 
    -1.998951e-09, -2.461971e-09, -3.157272e-09, -3.820892e-09, -4.477035e-09,
  -2.249748e-10, -2.322567e-10, -2.413447e-10, -2.843758e-10, -3.621348e-10, 
    -4.655341e-10, -5.788411e-10, -7.152459e-10, -8.84426e-10, -1.078307e-09, 
    -1.33651e-09, -1.710365e-09, -2.253343e-09, -2.992484e-09, -3.69912e-09,
  -2.27289e-10, -2.165592e-10, -2.069672e-10, -1.427004e-10, -1.518288e-10, 
    -2.242519e-10, -3.364572e-10, -4.816434e-10, -6.588525e-10, 
    -8.520432e-10, -1.023788e-09, -1.277999e-09, -1.670595e-09, 
    -2.289514e-09, -3.007331e-09,
  -2.679201e-10, -2.977552e-10, -2.857823e-10, -1.711233e-10, -1.070813e-10, 
    -9.026613e-11, -1.252699e-10, -2.336262e-10, -3.90068e-10, -6.074197e-10, 
    -8.389672e-10, -1.016858e-09, -1.255448e-09, -1.739588e-09, -2.414412e-09,
  -1.695167e-10, -1.783686e-10, -8.519615e-11, -1.734514e-10, -1.75205e-10, 
    -1.384109e-10, -9.5943e-11, -9.053087e-11, -1.940897e-10, -3.506983e-10, 
    -5.862374e-10, -8.315458e-10, -1.030694e-09, -1.365358e-09, -1.968419e-09,
  -2.973892e-09, -3.18e-09, -3.41038e-09, -3.724603e-09, -4.142727e-09, 
    -4.701188e-09, -5.386618e-09, -6.135417e-09, -6.78899e-09, -7.395545e-09, 
    -7.883678e-09, -8.451031e-09, -9.096195e-09, -9.626731e-09, -9.135385e-09,
  -2.584123e-09, -2.739043e-09, -2.913128e-09, -3.103648e-09, -3.328156e-09, 
    -3.632507e-09, -3.984868e-09, -4.464418e-09, -4.905735e-09, 
    -5.471009e-09, -5.987836e-09, -6.582204e-09, -7.099723e-09, 
    -7.971173e-09, -8.138741e-09,
  -2.179822e-09, -2.357258e-09, -2.52091e-09, -2.66761e-09, -2.827846e-09, 
    -3.014179e-09, -3.243721e-09, -3.552022e-09, -3.897215e-09, 
    -4.284823e-09, -4.733276e-09, -5.365221e-09, -5.575693e-09, 
    -5.877543e-09, -6.611137e-09,
  -1.589391e-09, -1.875419e-09, -2.12767e-09, -2.328411e-09, -2.475937e-09, 
    -2.647148e-09, -2.826185e-09, -3.079511e-09, -3.38664e-09, -3.680038e-09, 
    -4.096169e-09, -4.579839e-09, -5.259457e-09, -4.990263e-09, -4.41515e-09,
  -9.210915e-10, -1.246364e-09, -1.589475e-09, -1.904561e-09, -2.144757e-09, 
    -2.33029e-09, -2.533559e-09, -2.711645e-09, -2.990768e-09, -3.233044e-09, 
    -3.599985e-09, -3.940518e-09, -5.183156e-09, -5.295198e-09, -4.170605e-09,
  -5.402274e-10, -6.760115e-10, -9.427722e-10, -1.266686e-09, -1.610565e-09, 
    -1.903592e-09, -2.208373e-09, -2.403146e-09, -2.691652e-09, 
    -2.884257e-09, -3.258465e-09, -3.490289e-09, -4.188241e-09, 
    -5.667609e-09, -4.673183e-09,
  -4.300833e-10, -4.653136e-10, -5.311301e-10, -6.59567e-10, -9.538422e-10, 
    -1.283032e-09, -1.667994e-09, -1.898623e-09, -2.240064e-09, 
    -2.453941e-09, -2.823825e-09, -3.145077e-09, -3.211055e-09, 
    -4.174334e-09, -5.155904e-09,
  -3.233898e-10, -3.423553e-10, -3.559564e-10, -3.999067e-10, -5.072636e-10, 
    -6.954426e-10, -1.044454e-09, -1.362018e-09, -1.731029e-09, 
    -2.050841e-09, -2.404712e-09, -2.758753e-09, -2.956108e-09, 
    -3.264775e-09, -4.145033e-09,
  -2.691333e-10, -3.020144e-10, -3.036339e-10, -3.38693e-10, -4.136281e-10, 
    -4.965578e-10, -6.542371e-10, -9.024939e-10, -1.227372e-09, 
    -1.592129e-09, -2.030814e-09, -2.379491e-09, -2.74822e-09, -2.986813e-09, 
    -3.600972e-09,
  -8.466319e-11, -1.857604e-10, -2.613182e-10, -3.341114e-10, -3.902786e-10, 
    -4.285717e-10, -5.018828e-10, -6.254787e-10, -8.564451e-10, 
    -1.157725e-09, -1.563812e-09, -1.976685e-09, -2.369078e-09, 
    -2.692607e-09, -3.153209e-09,
  -2.906104e-09, -2.98226e-09, -3.140946e-09, -3.35218e-09, -3.625809e-09, 
    -4.081562e-09, -4.826086e-09, -6.119284e-09, -8.370365e-09, 
    -1.076261e-08, -1.283667e-08, -1.453155e-08, -1.572622e-08, 
    -1.659424e-08, -1.781546e-08,
  -2.57394e-09, -2.746955e-09, -2.885458e-09, -3.021492e-09, -3.157727e-09, 
    -3.369944e-09, -3.72741e-09, -4.223982e-09, -5.198445e-09, -6.806072e-09, 
    -8.958887e-09, -1.1097e-08, -1.28424e-08, -1.40709e-08, -1.51206e-08,
  -1.973106e-09, -2.335339e-09, -2.572726e-09, -2.755353e-09, -2.889775e-09, 
    -2.992501e-09, -3.186815e-09, -3.416571e-09, -3.802056e-09, 
    -4.521592e-09, -5.672294e-09, -7.492892e-09, -9.374515e-09, 
    -1.116317e-08, -1.249066e-08,
  -1.309849e-09, -1.665047e-09, -2.051765e-09, -2.40979e-09, -2.633351e-09, 
    -2.792162e-09, -2.909103e-09, -3.099612e-09, -3.267788e-09, 
    -3.582116e-09, -4.03465e-09, -5.010321e-09, -6.391589e-09, -8.00573e-09, 
    -9.632056e-09,
  -8.869412e-10, -1.059406e-09, -1.348232e-09, -1.74102e-09, -2.20561e-09, 
    -2.509425e-09, -2.704212e-09, -2.868131e-09, -3.035901e-09, 
    -3.209168e-09, -3.398487e-09, -3.809593e-09, -4.496118e-09, 
    -5.644039e-09, -6.890796e-09,
  -6.915472e-10, -7.604071e-10, -9.085904e-10, -1.109747e-09, -1.476526e-09, 
    -1.971246e-09, -2.375981e-09, -2.679326e-09, -2.875138e-09, 
    -3.046534e-09, -3.165891e-09, -3.423203e-09, -3.674968e-09, 
    -4.491666e-09, -5.254091e-09,
  -5.351256e-10, -5.949099e-10, -6.796627e-10, -7.931729e-10, -9.569191e-10, 
    -1.28612e-09, -1.727343e-09, -2.198258e-09, -2.571829e-09, -2.875941e-09, 
    -3.044664e-09, -3.281264e-09, -3.451611e-09, -3.8291e-09, -4.561063e-09,
  -4.37094e-10, -4.631637e-10, -5.189329e-10, -6.086414e-10, -6.972806e-10, 
    -8.708308e-10, -1.18148e-09, -1.614488e-09, -2.086926e-09, -2.500267e-09, 
    -2.807387e-09, -3.052936e-09, -3.310528e-09, -3.454465e-09, -4.001019e-09,
  -3.934717e-10, -4.257004e-10, -4.099484e-10, -4.641817e-10, -5.394157e-10, 
    -6.291566e-10, -7.761886e-10, -1.094686e-09, -1.562633e-09, 
    -2.088398e-09, -2.486932e-09, -2.769458e-09, -3.123739e-09, 
    -3.294281e-09, -3.532776e-09,
  -3.375776e-10, -4.492097e-10, -4.798302e-10, -4.407095e-10, -4.836843e-10, 
    -5.384591e-10, -6.17581e-10, -7.625967e-10, -1.069309e-09, -1.574514e-09, 
    -2.108538e-09, -2.463932e-09, -2.824599e-09, -3.167629e-09, -3.343606e-09,
  -5.732913e-09, -5.964425e-09, -6.272638e-09, -6.726358e-09, -7.352714e-09, 
    -8.12767e-09, -8.883206e-09, -9.736344e-09, -1.042482e-08, -1.100405e-08, 
    -1.143653e-08, -1.17667e-08, -1.215069e-08, -1.249229e-08, -1.285758e-08,
  -5.295395e-09, -5.498541e-09, -5.769317e-09, -6.032844e-09, -6.381153e-09, 
    -6.839353e-09, -7.429468e-09, -8.138824e-09, -8.897295e-09, 
    -9.621838e-09, -1.02693e-08, -1.083523e-08, -1.123741e-08, -1.17111e-08, 
    -1.206605e-08,
  -4.753458e-09, -5.003666e-09, -5.283064e-09, -5.55477e-09, -5.803665e-09, 
    -6.069429e-09, -6.392611e-09, -6.837985e-09, -7.381277e-09, 
    -8.054204e-09, -8.748078e-09, -9.483364e-09, -1.007946e-08, 
    -1.060446e-08, -1.116404e-08,
  -3.942206e-09, -4.320318e-09, -4.660178e-09, -4.967158e-09, -5.279339e-09, 
    -5.555561e-09, -5.773682e-09, -6.057857e-09, -6.350997e-09, 
    -6.742704e-09, -7.277336e-09, -7.881482e-09, -8.559263e-09, 
    -9.175407e-09, -9.817088e-09,
  -3.07932e-09, -3.496186e-09, -3.882166e-09, -4.244092e-09, -4.596957e-09, 
    -4.954215e-09, -5.239418e-09, -5.490559e-09, -5.711208e-09, 
    -5.933792e-09, -6.175341e-09, -6.537592e-09, -7.007935e-09, 
    -7.567303e-09, -8.218418e-09,
  -2.272983e-09, -2.667082e-09, -3.013983e-09, -3.35615e-09, -3.717442e-09, 
    -4.124588e-09, -4.554922e-09, -4.92602e-09, -5.205212e-09, -5.394542e-09, 
    -5.556624e-09, -5.664949e-09, -5.9051e-09, -6.237157e-09, -6.741145e-09,
  -1.711442e-09, -1.90487e-09, -2.169952e-09, -2.509749e-09, -2.845439e-09, 
    -3.201894e-09, -3.59747e-09, -4.041427e-09, -4.479542e-09, -4.844965e-09, 
    -5.069594e-09, -5.153166e-09, -5.231216e-09, -5.354708e-09, -5.630251e-09,
  -1.370198e-09, -1.431064e-09, -1.5371e-09, -1.749052e-09, -2.053594e-09, 
    -2.3979e-09, -2.796061e-09, -3.166477e-09, -3.580604e-09, -4.00027e-09, 
    -4.398169e-09, -4.627568e-09, -4.728938e-09, -4.816477e-09, -4.933881e-09,
  -1.240424e-09, -1.255394e-09, -1.260202e-09, -1.295395e-09, -1.416298e-09, 
    -1.65499e-09, -1.984398e-09, -2.390851e-09, -2.833671e-09, -3.239403e-09, 
    -3.642651e-09, -3.965669e-09, -4.184028e-09, -4.370612e-09, -4.508677e-09,
  -1.068395e-09, -1.147326e-09, -1.1959e-09, -1.162729e-09, -1.186331e-09, 
    -1.262803e-09, -1.395805e-09, -1.619889e-09, -2.00541e-09, -2.460593e-09, 
    -2.910502e-09, -3.325331e-09, -3.643514e-09, -3.942163e-09, -4.161472e-09,
  -4.085503e-09, -4.319152e-09, -4.492388e-09, -4.651044e-09, -4.756297e-09, 
    -4.870454e-09, -5.034083e-09, -5.251374e-09, -5.505315e-09, 
    -5.795266e-09, -6.143893e-09, -6.489708e-09, -6.8379e-09, -7.196035e-09, 
    -7.522443e-09,
  -3.310832e-09, -3.547648e-09, -3.794293e-09, -3.934861e-09, -4.049379e-09, 
    -4.151683e-09, -4.292037e-09, -4.416898e-09, -4.614724e-09, 
    -4.882935e-09, -5.231885e-09, -5.587033e-09, -5.990281e-09, 
    -6.417935e-09, -6.821884e-09,
  -2.827634e-09, -3.015114e-09, -3.241056e-09, -3.427784e-09, -3.577263e-09, 
    -3.690755e-09, -3.817512e-09, -3.924547e-09, -4.090634e-09, 
    -4.337366e-09, -4.647871e-09, -4.968241e-09, -5.352391e-09, 
    -5.789837e-09, -6.218567e-09,
  -2.465117e-09, -2.696941e-09, -2.881665e-09, -3.046708e-09, -3.204619e-09, 
    -3.362324e-09, -3.515514e-09, -3.638987e-09, -3.791607e-09, -4.03202e-09, 
    -4.302059e-09, -4.615632e-09, -4.987621e-09, -5.386988e-09, -5.798805e-09,
  -2.087292e-09, -2.368381e-09, -2.626873e-09, -2.790034e-09, -2.918614e-09, 
    -3.025632e-09, -3.181233e-09, -3.346857e-09, -3.554395e-09, 
    -3.834064e-09, -4.113571e-09, -4.425468e-09, -4.78387e-09, -5.161227e-09, 
    -5.529951e-09,
  -1.799305e-09, -2.051338e-09, -2.338163e-09, -2.566649e-09, -2.75229e-09, 
    -2.868806e-09, -2.963112e-09, -3.098994e-09, -3.286378e-09, 
    -3.567252e-09, -3.892802e-09, -4.260007e-09, -4.645378e-09, 
    -5.012157e-09, -5.369703e-09,
  -1.575354e-09, -1.776771e-09, -2.043149e-09, -2.323734e-09, -2.564936e-09, 
    -2.757749e-09, -2.90087e-09, -3.016192e-09, -3.13363e-09, -3.342688e-09, 
    -3.629583e-09, -3.990002e-09, -4.397267e-09, -4.78787e-09, -5.168442e-09,
  -1.462236e-09, -1.625824e-09, -1.786968e-09, -2.031145e-09, -2.30182e-09, 
    -2.600736e-09, -2.850526e-09, -3.045396e-09, -3.187551e-09, 
    -3.320314e-09, -3.54021e-09, -3.84089e-09, -4.218949e-09, -4.612446e-09, 
    -4.988125e-09,
  -1.324398e-09, -1.52207e-09, -1.719928e-09, -1.898885e-09, -2.1173e-09, 
    -2.324127e-09, -2.65277e-09, -2.944192e-09, -3.192725e-09, -3.413529e-09, 
    -3.569961e-09, -3.780928e-09, -4.066765e-09, -4.460608e-09, -4.851588e-09,
  -1.219851e-09, -1.340731e-09, -1.553556e-09, -1.716993e-09, -1.944142e-09, 
    -2.185354e-09, -2.43415e-09, -2.748798e-09, -3.048654e-09, -3.362565e-09, 
    -3.640199e-09, -3.90455e-09, -4.106045e-09, -4.35011e-09, -4.674624e-09,
  -2.140411e-08, -2.158864e-08, -2.189861e-08, -2.20794e-08, -2.235178e-08, 
    -2.240879e-08, -2.279364e-08, -2.318414e-08, -2.334279e-08, 
    -2.343894e-08, -2.327097e-08, -2.296073e-08, -2.265221e-08, -2.18752e-08, 
    -2.066429e-08,
  -1.974761e-08, -1.980081e-08, -2.006187e-08, -2.033368e-08, -2.066699e-08, 
    -2.065875e-08, -2.051953e-08, -2.046322e-08, -2.021555e-08, 
    -2.002272e-08, -1.965027e-08, -1.938738e-08, -1.903989e-08, 
    -1.842178e-08, -1.736287e-08,
  -1.741209e-08, -1.806435e-08, -1.832271e-08, -1.850918e-08, -1.864624e-08, 
    -1.866831e-08, -1.847734e-08, -1.821054e-08, -1.779683e-08, 
    -1.739093e-08, -1.672223e-08, -1.594245e-08, -1.524496e-08, 
    -1.413001e-08, -1.307409e-08,
  -1.503913e-08, -1.57008e-08, -1.630649e-08, -1.645055e-08, -1.650155e-08, 
    -1.631773e-08, -1.62121e-08, -1.592428e-08, -1.55188e-08, -1.496146e-08, 
    -1.41822e-08, -1.335183e-08, -1.231965e-08, -1.122799e-08, -1.014023e-08,
  -1.213418e-08, -1.274352e-08, -1.319066e-08, -1.351997e-08, -1.369221e-08, 
    -1.360053e-08, -1.337301e-08, -1.302814e-08, -1.258141e-08, 
    -1.203064e-08, -1.130994e-08, -1.047876e-08, -9.485785e-09, 
    -8.335934e-09, -7.185345e-09,
  -9.258481e-09, -9.797883e-09, -1.01246e-08, -1.045129e-08, -1.055915e-08, 
    -1.052418e-08, -1.036043e-08, -1.005347e-08, -9.601943e-09, 
    -9.089418e-09, -8.393004e-09, -7.6816e-09, -6.833844e-09, -5.796978e-09, 
    -5.029572e-09,
  -6.888838e-09, -7.371582e-09, -7.593639e-09, -7.841626e-09, -7.897453e-09, 
    -7.871072e-09, -7.729798e-09, -7.476965e-09, -7.099369e-09, 
    -6.664314e-09, -6.105185e-09, -5.584437e-09, -4.662929e-09, 
    -3.932699e-09, -3.224161e-09,
  -5.234201e-09, -5.601791e-09, -5.784849e-09, -5.917576e-09, -5.947261e-09, 
    -5.862435e-09, -5.739833e-09, -5.459932e-09, -5.174773e-09, 
    -4.708013e-09, -4.375527e-09, -3.77816e-09, -3.22148e-09, -2.651007e-09, 
    -2.13598e-09,
  -3.474243e-09, -3.778202e-09, -3.976641e-09, -4.109546e-09, -4.136437e-09, 
    -4.061429e-09, -3.902119e-09, -3.693281e-09, -3.4369e-09, -3.131551e-09, 
    -2.831861e-09, -2.456755e-09, -2.205057e-09, -1.596218e-09, -1.441098e-09,
  -1.997146e-09, -2.254054e-09, -2.425594e-09, -2.536634e-09, -2.564193e-09, 
    -2.551509e-09, -2.460085e-09, -2.331467e-09, -2.208556e-09, -2.09139e-09, 
    -1.923419e-09, -1.776033e-09, -1.533432e-09, -8.606785e-10, -1.004645e-09,
  -1.190775e-08, -1.177466e-08, -1.159968e-08, -1.131411e-08, -1.107979e-08, 
    -1.069737e-08, -1.027412e-08, -9.864936e-09, -9.504978e-09, 
    -9.221182e-09, -8.918986e-09, -8.801136e-09, -8.90493e-09, -9.078383e-09, 
    -9.432202e-09,
  -1.205011e-08, -1.204679e-08, -1.189388e-08, -1.157316e-08, -1.129692e-08, 
    -1.103535e-08, -1.070901e-08, -1.03449e-08, -9.925257e-09, -9.513378e-09, 
    -9.288931e-09, -9.158026e-09, -9.182325e-09, -9.368146e-09, -9.665024e-09,
  -1.288881e-08, -1.268193e-08, -1.253057e-08, -1.232051e-08, -1.215352e-08, 
    -1.191738e-08, -1.162018e-08, -1.134979e-08, -1.109587e-08, -1.05928e-08, 
    -1.018325e-08, -9.892104e-09, -9.778987e-09, -9.942458e-09, -1.026681e-08,
  -1.416791e-08, -1.410122e-08, -1.384984e-08, -1.349122e-08, -1.323996e-08, 
    -1.302776e-08, -1.265167e-08, -1.225649e-08, -1.193973e-08, 
    -1.160236e-08, -1.129569e-08, -1.09397e-08, -1.060271e-08, -1.031813e-08, 
    -1.006526e-08,
  -1.405815e-08, -1.471298e-08, -1.523767e-08, -1.508061e-08, -1.485842e-08, 
    -1.44179e-08, -1.394314e-08, -1.35291e-08, -1.33046e-08, -1.320527e-08, 
    -1.321642e-08, -1.325743e-08, -1.330738e-08, -1.332095e-08, -1.319024e-08,
  -1.458908e-08, -1.501137e-08, -1.600069e-08, -1.616055e-08, -1.617372e-08, 
    -1.605086e-08, -1.585446e-08, -1.571331e-08, -1.557053e-08, 
    -1.558821e-08, -1.566443e-08, -1.589249e-08, -1.599179e-08, 
    -1.609464e-08, -1.595549e-08,
  -1.310603e-08, -1.420474e-08, -1.478336e-08, -1.546191e-08, -1.582977e-08, 
    -1.59847e-08, -1.624752e-08, -1.666839e-08, -1.743724e-08, -1.825586e-08, 
    -1.919421e-08, -1.984786e-08, -2.037379e-08, -2.068854e-08, -2.077115e-08,
  -1.184139e-08, -1.278256e-08, -1.344018e-08, -1.393491e-08, -1.4497e-08, 
    -1.499942e-08, -1.581399e-08, -1.651754e-08, -1.694446e-08, 
    -1.710161e-08, -1.744118e-08, -1.761263e-08, -1.753662e-08, 
    -1.720444e-08, -1.67382e-08,
  -1.161594e-08, -1.202984e-08, -1.246131e-08, -1.270848e-08, -1.310517e-08, 
    -1.361964e-08, -1.393406e-08, -1.423322e-08, -1.414921e-08, 
    -1.394543e-08, -1.385344e-08, -1.311207e-08, -1.231786e-08, 
    -1.177647e-08, -1.141786e-08,
  -1.143426e-08, -1.149007e-08, -1.138829e-08, -1.148885e-08, -1.160443e-08, 
    -1.202223e-08, -1.236817e-08, -1.254219e-08, -1.231653e-08, 
    -1.219276e-08, -1.130437e-08, -1.047279e-08, -9.957716e-09, 
    -9.675645e-09, -9.687832e-09,
  -1.209947e-08, -1.325956e-08, -1.42589e-08, -1.549413e-08, -1.656593e-08, 
    -1.767479e-08, -1.850294e-08, -1.931689e-08, -1.979446e-08, 
    -2.006532e-08, -2.005386e-08, -2.001918e-08, -1.993489e-08, 
    -1.985691e-08, -1.989752e-08,
  -1.052174e-08, -1.189063e-08, -1.30692e-08, -1.42348e-08, -1.520364e-08, 
    -1.625985e-08, -1.722605e-08, -1.805171e-08, -1.867496e-08, 
    -1.903216e-08, -1.903044e-08, -1.88071e-08, -1.856717e-08, -1.832322e-08, 
    -1.822636e-08,
  -8.665082e-09, -1.038533e-08, -1.167218e-08, -1.293855e-08, -1.405825e-08, 
    -1.500945e-08, -1.590825e-08, -1.666941e-08, -1.726335e-08, -1.75185e-08, 
    -1.746053e-08, -1.722075e-08, -1.697251e-08, -1.671939e-08, -1.652609e-08,
  -7.263811e-09, -8.760792e-09, -1.027272e-08, -1.159715e-08, -1.278005e-08, 
    -1.389096e-08, -1.481471e-08, -1.553394e-08, -1.600582e-08, 
    -1.616339e-08, -1.603248e-08, -1.584145e-08, -1.557083e-08, 
    -1.529211e-08, -1.501948e-08,
  -6.443369e-09, -7.387146e-09, -8.77005e-09, -1.028577e-08, -1.154461e-08, 
    -1.274779e-08, -1.361964e-08, -1.423846e-08, -1.453184e-08, 
    -1.466285e-08, -1.451848e-08, -1.437464e-08, -1.398415e-08, 
    -1.371406e-08, -1.347142e-08,
  -6.617403e-09, -6.759215e-09, -7.567547e-09, -8.864093e-09, -1.032072e-08, 
    -1.164574e-08, -1.26131e-08, -1.327217e-08, -1.348745e-08, -1.356186e-08, 
    -1.354754e-08, -1.323083e-08, -1.295887e-08, -1.287584e-08, -1.295647e-08,
  -6.964237e-09, -6.916472e-09, -7.262507e-09, -8.11547e-09, -9.268567e-09, 
    -1.035693e-08, -1.139216e-08, -1.178103e-08, -1.213479e-08, 
    -1.250142e-08, -1.283251e-08, -1.290274e-08, -1.317668e-08, 
    -1.371206e-08, -1.427254e-08,
  -7.391282e-09, -7.182392e-09, -7.244201e-09, -7.760554e-09, -8.614849e-09, 
    -9.473361e-09, -1.029145e-08, -1.078982e-08, -1.161796e-08, 
    -1.296149e-08, -1.33961e-08, -1.380145e-08, -1.43277e-08, -1.457803e-08, 
    -1.452137e-08,
  -7.808374e-09, -7.631636e-09, -7.875723e-09, -8.009434e-09, -8.370667e-09, 
    -8.934529e-09, -9.7043e-09, -1.08796e-08, -1.22416e-08, -1.353268e-08, 
    -1.404278e-08, -1.438443e-08, -1.43522e-08, -1.371345e-08, -1.228002e-08,
  -8.126645e-09, -8.012922e-09, -8.102633e-09, -8.450538e-09, -8.615447e-09, 
    -9.054123e-09, -1.060863e-08, -1.190156e-08, -1.313588e-08, -1.502e-08, 
    -1.45252e-08, -1.346033e-08, -1.245793e-08, -9.966377e-09, -8.420179e-09,
  -1.047388e-08, -1.100492e-08, -1.148496e-08, -1.207761e-08, -1.250105e-08, 
    -1.267995e-08, -1.272631e-08, -1.27065e-08, -1.254239e-08, -1.269324e-08, 
    -1.298111e-08, -1.331837e-08, -1.374501e-08, -1.436849e-08, -1.496987e-08,
  -9.791785e-09, -1.033561e-08, -1.086392e-08, -1.147245e-08, -1.190496e-08, 
    -1.215575e-08, -1.232707e-08, -1.208019e-08, -1.193352e-08, 
    -1.177879e-08, -1.177409e-08, -1.18241e-08, -1.213429e-08, -1.245728e-08, 
    -1.285698e-08,
  -9.229328e-09, -9.581932e-09, -1.000659e-08, -1.052775e-08, -1.089733e-08, 
    -1.122968e-08, -1.105825e-08, -1.080579e-08, -1.040396e-08, 
    -9.907018e-09, -9.638226e-09, -1.00111e-08, -1.045793e-08, -1.085654e-08, 
    -1.104993e-08,
  -8.858007e-09, -9.007186e-09, -9.260359e-09, -9.480376e-09, -9.798899e-09, 
    -9.75653e-09, -9.630282e-09, -9.13541e-09, -8.62066e-09, -8.366388e-09, 
    -9.007621e-09, -9.951597e-09, -1.030336e-08, -1.023372e-08, -1.042653e-08,
  -8.488987e-09, -8.655046e-09, -8.751968e-09, -8.742916e-09, -8.66271e-09, 
    -8.382703e-09, -8.204012e-09, -7.670747e-09, -7.706669e-09, 
    -8.357169e-09, -9.415438e-09, -9.8867e-09, -9.404355e-09, -9.430186e-09, 
    -9.544955e-09,
  -8.396573e-09, -8.271895e-09, -8.276845e-09, -8.222623e-09, -7.88e-09, 
    -7.694569e-09, -7.455705e-09, -7.356318e-09, -7.886258e-09, -8.52988e-09, 
    -9.098887e-09, -9.417908e-09, -8.745351e-09, -9.324613e-09, -9.027851e-09,
  -8.609637e-09, -8.317657e-09, -8.065098e-09, -7.9359e-09, -7.675635e-09, 
    -7.600127e-09, -7.522184e-09, -7.491779e-09, -7.921999e-09, 
    -8.383059e-09, -9.351192e-09, -9.251893e-09, -9.226778e-09, 
    -9.355526e-09, -9.656829e-09,
  -9.066896e-09, -8.575168e-09, -8.284727e-09, -8.058649e-09, -7.846657e-09, 
    -7.797361e-09, -7.727619e-09, -7.646952e-09, -8.123975e-09, -8.76897e-09, 
    -9.714816e-09, -9.385668e-09, -9.468947e-09, -9.751541e-09, -9.776679e-09,
  -9.581406e-09, -9.003267e-09, -8.623707e-09, -8.387498e-09, -8.177617e-09, 
    -8.037524e-09, -7.946091e-09, -7.898979e-09, -8.449796e-09, 
    -8.942418e-09, -9.759109e-09, -9.021865e-09, -1.039899e-08, 
    -1.082191e-08, -1.152235e-08,
  -9.968228e-09, -9.681145e-09, -9.232931e-09, -9.015001e-09, -8.624974e-09, 
    -8.475566e-09, -8.318117e-09, -8.38524e-09, -8.75303e-09, -9.279391e-09, 
    -9.580241e-09, -9.577721e-09, -1.210451e-08, -1.34037e-08, -9.862981e-09,
  -1.096263e-08, -1.090069e-08, -1.099096e-08, -1.118305e-08, -1.141335e-08, 
    -1.184437e-08, -1.208779e-08, -1.235137e-08, -1.246908e-08, 
    -1.243721e-08, -1.229758e-08, -1.177214e-08, -1.112008e-08, 
    -1.051219e-08, -1.009602e-08,
  -1.050129e-08, -1.036376e-08, -1.040578e-08, -1.061115e-08, -1.087404e-08, 
    -1.132496e-08, -1.146318e-08, -1.189072e-08, -1.197327e-08, 
    -1.200189e-08, -1.148016e-08, -1.094657e-08, -1.040922e-08, 
    -1.006066e-08, -9.846835e-09,
  -1.024334e-08, -1.012419e-08, -1.00939e-08, -1.031834e-08, -1.056621e-08, 
    -1.074623e-08, -1.123614e-08, -1.139402e-08, -1.150833e-08, 
    -1.119778e-08, -1.059251e-08, -1.012133e-08, -9.951065e-09, 
    -1.004471e-08, -1.004245e-08,
  -9.926383e-09, -9.946799e-09, -1.003521e-08, -1.013524e-08, -1.041932e-08, 
    -1.05607e-08, -1.079462e-08, -1.088704e-08, -1.090087e-08, -1.046277e-08, 
    -1.009908e-08, -9.919972e-09, -1.001623e-08, -1.017003e-08, -1.012051e-08,
  -9.907782e-09, -9.849289e-09, -9.930398e-09, -9.972094e-09, -1.014663e-08, 
    -1.034204e-08, -1.037665e-08, -1.052483e-08, -1.044456e-08, 
    -1.004473e-08, -9.911852e-09, -9.934987e-09, -1.00945e-08, -1.009572e-08, 
    -9.871543e-09,
  -9.900318e-09, -9.952601e-09, -1.002352e-08, -9.994096e-09, -9.963504e-09, 
    -1.006338e-08, -1.02126e-08, -1.034492e-08, -9.969671e-09, -9.821678e-09, 
    -9.664999e-09, -9.682283e-09, -9.963253e-09, -1.000993e-08, -1.014806e-08,
  -9.975323e-09, -9.970899e-09, -9.977008e-09, -1.004319e-08, -9.952282e-09, 
    -9.852373e-09, -9.987202e-09, -9.859197e-09, -9.582312e-09, 
    -9.496091e-09, -9.606906e-09, -9.790712e-09, -1.021766e-08, 
    -1.042816e-08, -1.074496e-08,
  -1.016928e-08, -1.015386e-08, -1.008692e-08, -1.009717e-08, -9.894655e-09, 
    -9.782434e-09, -9.605899e-09, -9.434493e-09, -9.201091e-09, 
    -9.513073e-09, -9.498732e-09, -1.003194e-08, -1.0481e-08, -1.062458e-08, 
    -1.039507e-08,
  -1.015509e-08, -1.03789e-08, -1.045643e-08, -1.035335e-08, -1.017523e-08, 
    -9.942153e-09, -9.859057e-09, -9.641924e-09, -9.814574e-09, 
    -9.722382e-09, -1.0084e-08, -1.052925e-08, -1.067046e-08, -1.015924e-08, 
    -8.99256e-09,
  -9.65408e-09, -9.984014e-09, -1.006066e-08, -1.002331e-08, -9.946842e-09, 
    -9.955651e-09, -9.781862e-09, -9.862349e-09, -9.897938e-09, 
    -1.011237e-08, -1.055674e-08, -1.049041e-08, -9.945828e-09, 
    -8.514307e-09, -7.220991e-09,
  -1.599977e-08, -1.606922e-08, -1.609722e-08, -1.601e-08, -1.599118e-08, 
    -1.584453e-08, -1.570509e-08, -1.532749e-08, -1.488621e-08, 
    -1.439531e-08, -1.388282e-08, -1.34982e-08, -1.30495e-08, -1.259572e-08, 
    -1.22274e-08,
  -1.492985e-08, -1.502606e-08, -1.518714e-08, -1.520185e-08, -1.522078e-08, 
    -1.503943e-08, -1.484231e-08, -1.446784e-08, -1.407464e-08, 
    -1.361542e-08, -1.318449e-08, -1.276941e-08, -1.229063e-08, 
    -1.189806e-08, -1.166142e-08,
  -1.357468e-08, -1.390832e-08, -1.41065e-08, -1.419044e-08, -1.42156e-08, 
    -1.410845e-08, -1.391983e-08, -1.359368e-08, -1.325945e-08, 
    -1.285069e-08, -1.257259e-08, -1.211293e-08, -1.171138e-08, 
    -1.137432e-08, -1.102707e-08,
  -1.193252e-08, -1.252516e-08, -1.275671e-08, -1.293368e-08, -1.301037e-08, 
    -1.30085e-08, -1.294695e-08, -1.277719e-08, -1.251158e-08, -1.233416e-08, 
    -1.203995e-08, -1.153107e-08, -1.117639e-08, -1.089527e-08, -1.062136e-08,
  -1.039529e-08, -1.098726e-08, -1.145543e-08, -1.170849e-08, -1.191049e-08, 
    -1.202607e-08, -1.20642e-08, -1.197382e-08, -1.182561e-08, -1.171722e-08, 
    -1.134578e-08, -1.098407e-08, -1.070707e-08, -1.044867e-08, -1.033544e-08,
  -9.2932e-09, -9.834079e-09, -1.026015e-08, -1.061751e-08, -1.090919e-08, 
    -1.112054e-08, -1.125581e-08, -1.122899e-08, -1.122849e-08, 
    -1.104711e-08, -1.078029e-08, -1.061795e-08, -1.036696e-08, -1.04164e-08, 
    -1.028839e-08,
  -8.380654e-09, -8.937704e-09, -9.3782e-09, -9.782647e-09, -1.009627e-08, 
    -1.033135e-08, -1.048369e-08, -1.057232e-08, -1.064033e-08, 
    -1.053621e-08, -1.050523e-08, -1.029064e-08, -1.020555e-08, 
    -1.005053e-08, -9.758588e-09,
  -7.615127e-09, -8.164154e-09, -8.653081e-09, -9.161921e-09, -9.560059e-09, 
    -9.884615e-09, -1.005666e-08, -1.023771e-08, -1.027834e-08, 
    -1.027278e-08, -1.001461e-08, -9.868747e-09, -9.859635e-09, 
    -9.460043e-09, -8.89587e-09,
  -6.910794e-09, -7.506106e-09, -8.074044e-09, -8.664793e-09, -9.085913e-09, 
    -9.469238e-09, -9.639685e-09, -9.857888e-09, -9.827256e-09, 
    -9.618399e-09, -9.565202e-09, -9.709861e-09, -9.245913e-09, 
    -8.480204e-09, -7.371286e-09,
  -6.008861e-09, -6.738202e-09, -7.439064e-09, -8.015197e-09, -8.610709e-09, 
    -8.988578e-09, -9.161742e-09, -9.321986e-09, -9.326033e-09, 
    -9.353384e-09, -9.528057e-09, -9.076042e-09, -8.044394e-09, 
    -6.861315e-09, -5.87456e-09,
  -2.536837e-08, -2.489102e-08, -2.409243e-08, -2.345807e-08, -2.312604e-08, 
    -2.279278e-08, -2.253528e-08, -2.236531e-08, -2.226833e-08, 
    -2.219211e-08, -2.216913e-08, -2.210079e-08, -2.198309e-08, 
    -2.182723e-08, -2.16507e-08,
  -2.511678e-08, -2.454996e-08, -2.40152e-08, -2.333656e-08, -2.298349e-08, 
    -2.280263e-08, -2.263243e-08, -2.243282e-08, -2.226023e-08, 
    -2.209766e-08, -2.19486e-08, -2.177464e-08, -2.165026e-08, -2.133546e-08, 
    -2.079798e-08,
  -2.338623e-08, -2.337678e-08, -2.326725e-08, -2.296343e-08, -2.243316e-08, 
    -2.202494e-08, -2.16783e-08, -2.129595e-08, -2.103481e-08, -2.072527e-08, 
    -2.028187e-08, -1.966243e-08, -1.884658e-08, -1.780862e-08, -1.657037e-08,
  -2.046547e-08, -2.107315e-08, -2.119174e-08, -2.100084e-08, -2.075357e-08, 
    -2.03063e-08, -1.969122e-08, -1.909334e-08, -1.836552e-08, -1.758618e-08, 
    -1.663817e-08, -1.551844e-08, -1.42514e-08, -1.283779e-08, -1.143491e-08,
  -1.575514e-08, -1.754385e-08, -1.849209e-08, -1.866741e-08, -1.83129e-08, 
    -1.783723e-08, -1.7206e-08, -1.63956e-08, -1.543317e-08, -1.430314e-08, 
    -1.299958e-08, -1.152638e-08, -9.977486e-09, -8.610004e-09, -7.551057e-09,
  -1.220208e-08, -1.416637e-08, -1.549115e-08, -1.629767e-08, -1.627511e-08, 
    -1.559486e-08, -1.47429e-08, -1.360747e-08, -1.222767e-08, -1.074426e-08, 
    -9.173432e-09, -7.778001e-09, -6.721453e-09, -5.986383e-09, -5.505628e-09,
  -8.745607e-09, -1.017339e-08, -1.108777e-08, -1.158421e-08, -1.171396e-08, 
    -1.147911e-08, -1.092918e-08, -9.915754e-09, -8.704146e-09, 
    -7.450504e-09, -6.391776e-09, -5.595813e-09, -5.025944e-09, 
    -4.662447e-09, -4.486304e-09,
  -5.403297e-09, -6.475003e-09, -7.247871e-09, -7.792996e-09, -8.188976e-09, 
    -8.11111e-09, -7.550742e-09, -6.801264e-09, -6.021986e-09, -5.276324e-09, 
    -4.611056e-09, -4.147476e-09, -3.979749e-09, -4.004236e-09, -4.122032e-09,
  -3.241983e-09, -3.770845e-09, -4.374529e-09, -4.856025e-09, -5.094747e-09, 
    -5.058672e-09, -4.765369e-09, -4.363256e-09, -3.971107e-09, 
    -3.625384e-09, -3.459403e-09, -3.514245e-09, -3.694947e-09, 
    -3.933299e-09, -4.293022e-09,
  -2.584672e-09, -2.506095e-09, -2.512648e-09, -2.608312e-09, -2.703555e-09, 
    -2.829828e-09, -2.791079e-09, -2.785544e-09, -2.84895e-09, -2.96141e-09, 
    -3.182412e-09, -3.433804e-09, -3.788075e-09, -4.169664e-09, -4.490192e-09,
  -1.969419e-08, -1.876453e-08, -1.716534e-08, -1.595715e-08, -1.533976e-08, 
    -1.504888e-08, -1.447923e-08, -1.360221e-08, -1.269599e-08, 
    -1.182971e-08, -1.120838e-08, -1.097332e-08, -1.140176e-08, 
    -1.213072e-08, -1.300839e-08,
  -1.928703e-08, -1.957037e-08, -1.887275e-08, -1.74141e-08, -1.608161e-08, 
    -1.527314e-08, -1.475728e-08, -1.433243e-08, -1.382771e-08, 
    -1.299457e-08, -1.213746e-08, -1.168439e-08, -1.14523e-08, -1.174397e-08, 
    -1.251475e-08,
  -1.627595e-08, -1.78456e-08, -1.901521e-08, -1.873416e-08, -1.755286e-08, 
    -1.648631e-08, -1.583635e-08, -1.532209e-08, -1.494908e-08, 
    -1.458253e-08, -1.408379e-08, -1.3512e-08, -1.313705e-08, -1.292134e-08, 
    -1.312516e-08,
  -1.351549e-08, -1.504445e-08, -1.701694e-08, -1.892492e-08, -1.932513e-08, 
    -1.837486e-08, -1.717017e-08, -1.656488e-08, -1.622666e-08, 
    -1.591417e-08, -1.564276e-08, -1.537173e-08, -1.502889e-08, 
    -1.476891e-08, -1.430979e-08,
  -1.077059e-08, -1.220233e-08, -1.389191e-08, -1.603181e-08, -1.804276e-08, 
    -1.970882e-08, -1.983259e-08, -1.924525e-08, -1.854784e-08, 
    -1.804271e-08, -1.775253e-08, -1.729039e-08, -1.675265e-08, 
    -1.609984e-08, -1.527703e-08,
  -8.129309e-09, -9.382657e-09, -1.094628e-08, -1.243334e-08, -1.452897e-08, 
    -1.675693e-08, -1.881787e-08, -2.030096e-08, -2.110922e-08, -2.10227e-08, 
    -2.052357e-08, -1.968397e-08, -1.841418e-08, -1.693103e-08, -1.538763e-08,
  -5.879826e-09, -6.956825e-09, -8.04443e-09, -9.476697e-09, -1.079193e-08, 
    -1.269045e-08, -1.467809e-08, -1.669668e-08, -1.836287e-08, 
    -1.966682e-08, -2.030895e-08, -1.979233e-08, -1.869945e-08, 
    -1.707163e-08, -1.544316e-08,
  -4.405246e-09, -5.016314e-09, -5.718626e-09, -6.681554e-09, -7.727631e-09, 
    -8.901764e-09, -1.028718e-08, -1.185853e-08, -1.319273e-08, 
    -1.427362e-08, -1.526837e-08, -1.600024e-08, -1.65773e-08, -1.657424e-08, 
    -1.584941e-08,
  -3.365675e-09, -3.580086e-09, -3.950829e-09, -4.471194e-09, -5.120103e-09, 
    -5.826653e-09, -6.511798e-09, -7.227617e-09, -8.13778e-09, -9.110142e-09, 
    -1.023429e-08, -1.11327e-08, -1.182636e-08, -1.225105e-08, -1.246159e-08,
  -2.9589e-09, -2.962924e-09, -3.102921e-09, -3.324413e-09, -3.600967e-09, 
    -3.868738e-09, -4.078788e-09, -4.421838e-09, -4.83568e-09, -5.434196e-09, 
    -6.057181e-09, -6.788649e-09, -7.494572e-09, -8.128669e-09, -8.593156e-09,
  -1.443274e-08, -1.557697e-08, -1.656003e-08, -1.754826e-08, -1.820791e-08, 
    -1.869008e-08, -1.899569e-08, -1.903949e-08, -1.905916e-08, 
    -1.872787e-08, -1.829678e-08, -1.781782e-08, -1.733466e-08, 
    -1.671576e-08, -1.609055e-08,
  -1.239726e-08, -1.366044e-08, -1.483526e-08, -1.590839e-08, -1.691943e-08, 
    -1.768591e-08, -1.830801e-08, -1.850773e-08, -1.855651e-08, 
    -1.849358e-08, -1.819649e-08, -1.781738e-08, -1.736455e-08, 
    -1.697843e-08, -1.638943e-08,
  -1.046504e-08, -1.145136e-08, -1.244408e-08, -1.350294e-08, -1.46075e-08, 
    -1.562596e-08, -1.647552e-08, -1.709265e-08, -1.73952e-08, -1.74258e-08, 
    -1.739353e-08, -1.719369e-08, -1.692175e-08, -1.658966e-08, -1.619621e-08,
  -9.210233e-09, -9.994754e-09, -1.065984e-08, -1.138264e-08, -1.227244e-08, 
    -1.324498e-08, -1.429125e-08, -1.518149e-08, -1.582442e-08, 
    -1.609416e-08, -1.621063e-08, -1.623199e-08, -1.61837e-08, -1.607943e-08, 
    -1.596459e-08,
  -8.604265e-09, -9.026339e-09, -9.515588e-09, -9.997626e-09, -1.043138e-08, 
    -1.100885e-08, -1.169567e-08, -1.256951e-08, -1.336563e-08, 
    -1.401602e-08, -1.439961e-08, -1.459489e-08, -1.476567e-08, 
    -1.484207e-08, -1.489901e-08,
  -8.218831e-09, -8.483434e-09, -8.806714e-09, -9.093492e-09, -9.434557e-09, 
    -9.723826e-09, -1.013384e-08, -1.059767e-08, -1.117205e-08, 
    -1.174139e-08, -1.226532e-08, -1.269978e-08, -1.302425e-08, 
    -1.322697e-08, -1.346695e-08,
  -7.896651e-09, -8.083701e-09, -8.208421e-09, -8.403897e-09, -8.595459e-09, 
    -8.830957e-09, -9.049466e-09, -9.32361e-09, -9.636929e-09, -1.004883e-08, 
    -1.0436e-08, -1.088184e-08, -1.128085e-08, -1.175793e-08, -1.21932e-08,
  -7.311856e-09, -7.704049e-09, -7.872142e-09, -7.987637e-09, -8.06995e-09, 
    -8.186121e-09, -8.288116e-09, -8.388579e-09, -8.529581e-09, 
    -8.701778e-09, -8.920857e-09, -9.208072e-09, -9.452485e-09, 
    -9.918096e-09, -1.045252e-08,
  -6.260413e-09, -6.912208e-09, -7.315204e-09, -7.609001e-09, -7.725602e-09, 
    -7.776055e-09, -7.809287e-09, -7.855928e-09, -7.925722e-09, 
    -7.952202e-09, -8.01086e-09, -8.109939e-09, -8.227986e-09, -8.590301e-09, 
    -8.785729e-09,
  -4.861248e-09, -5.564445e-09, -6.257688e-09, -6.713027e-09, -7.070323e-09, 
    -7.260558e-09, -7.348799e-09, -7.3494e-09, -7.378703e-09, -7.400192e-09, 
    -7.399965e-09, -7.446289e-09, -7.41864e-09, -7.665935e-09, -7.638096e-09,
  -7.378517e-09, -7.763559e-09, -8.099593e-09, -8.445082e-09, -8.77045e-09, 
    -9.110646e-09, -9.69604e-09, -1.057819e-08, -1.153069e-08, -1.248196e-08, 
    -1.335825e-08, -1.402975e-08, -1.45909e-08, -1.51165e-08, -1.567201e-08,
  -6.647753e-09, -7.060712e-09, -7.472535e-09, -7.86509e-09, -8.216291e-09, 
    -8.582658e-09, -8.995685e-09, -9.716985e-09, -1.063159e-08, 
    -1.161598e-08, -1.255018e-08, -1.343645e-08, -1.405008e-08, 
    -1.458243e-08, -1.51558e-08,
  -5.907443e-09, -6.339616e-09, -6.791221e-09, -7.264289e-09, -7.672081e-09, 
    -8.083911e-09, -8.46605e-09, -8.977683e-09, -9.763853e-09, -1.073982e-08, 
    -1.163568e-08, -1.246023e-08, -1.315497e-08, -1.371003e-08, -1.42261e-08,
  -5.206243e-09, -5.656079e-09, -6.132863e-09, -6.627586e-09, -7.090662e-09, 
    -7.541894e-09, -8.00143e-09, -8.422163e-09, -8.953437e-09, -9.763418e-09, 
    -1.065647e-08, -1.144574e-08, -1.212244e-08, -1.265446e-08, -1.313808e-08,
  -4.594923e-09, -5.053832e-09, -5.531737e-09, -6.046491e-09, -6.521445e-09, 
    -6.987245e-09, -7.471614e-09, -7.958573e-09, -8.455549e-09, 
    -9.035682e-09, -9.762915e-09, -1.045204e-08, -1.107688e-08, 
    -1.159192e-08, -1.19915e-08,
  -3.783741e-09, -4.358859e-09, -4.881304e-09, -5.456884e-09, -5.981182e-09, 
    -6.491748e-09, -6.955764e-09, -7.414923e-09, -7.872748e-09, 
    -8.415623e-09, -9.004425e-09, -9.544052e-09, -1.005304e-08, -1.04727e-08, 
    -1.075265e-08,
  -2.881427e-09, -3.479162e-09, -4.123998e-09, -4.752648e-09, -5.38365e-09, 
    -5.962818e-09, -6.519525e-09, -7.010861e-09, -7.433271e-09, 
    -7.906806e-09, -8.420193e-09, -8.889102e-09, -9.288519e-09, 
    -9.624882e-09, -9.875845e-09,
  -2.059127e-09, -2.551888e-09, -3.182317e-09, -3.93232e-09, -4.638167e-09, 
    -5.308646e-09, -5.947547e-09, -6.532611e-09, -7.025512e-09, 
    -7.526737e-09, -7.97289e-09, -8.480971e-09, -8.956426e-09, -9.21981e-09, 
    -9.532164e-09,
  -1.684018e-09, -1.869572e-09, -2.284293e-09, -2.948952e-09, -3.76232e-09, 
    -4.560807e-09, -5.296217e-09, -5.966714e-09, -6.564773e-09, 
    -7.135994e-09, -7.633759e-09, -8.125144e-09, -8.570697e-09, 
    -8.969637e-09, -9.154101e-09,
  -1.655527e-09, -1.668377e-09, -1.762476e-09, -2.087192e-09, -2.663705e-09, 
    -3.537366e-09, -4.404756e-09, -5.271377e-09, -6.042667e-09, 
    -6.656597e-09, -7.30745e-09, -7.855069e-09, -8.261591e-09, -8.784173e-09, 
    -8.981851e-09,
  -2.659239e-09, -3.000771e-09, -3.493729e-09, -4.138744e-09, -4.927128e-09, 
    -5.803142e-09, -6.775351e-09, -7.775146e-09, -8.821915e-09, 
    -9.930658e-09, -1.095469e-08, -1.205831e-08, -1.321114e-08, 
    -1.429774e-08, -1.509394e-08,
  -1.852275e-09, -2.137665e-09, -2.455338e-09, -2.842131e-09, -3.337587e-09, 
    -3.947545e-09, -4.725633e-09, -5.619975e-09, -6.581971e-09, 
    -7.640484e-09, -8.694095e-09, -9.738288e-09, -1.075448e-08, 
    -1.172622e-08, -1.260975e-08,
  -1.479819e-09, -1.617107e-09, -1.777033e-09, -1.993782e-09, -2.297223e-09, 
    -2.702682e-09, -3.240011e-09, -3.908298e-09, -4.6438e-09, -5.481792e-09, 
    -6.454755e-09, -7.511405e-09, -8.563648e-09, -9.585997e-09, -1.05148e-08,
  -1.279909e-09, -1.315651e-09, -1.410627e-09, -1.519758e-09, -1.683618e-09, 
    -1.913114e-09, -2.261299e-09, -2.711293e-09, -3.282784e-09, 
    -3.956607e-09, -4.742197e-09, -5.649114e-09, -6.61401e-09, -7.657045e-09, 
    -8.617788e-09,
  -1.255183e-09, -1.168757e-09, -1.194708e-09, -1.275586e-09, -1.356221e-09, 
    -1.464598e-09, -1.625469e-09, -1.875146e-09, -2.218848e-09, 
    -2.746452e-09, -3.403546e-09, -4.223272e-09, -5.125324e-09, 
    -6.104129e-09, -7.112349e-09,
  -1.52715e-09, -1.363739e-09, -1.260837e-09, -1.242766e-09, -1.27606e-09, 
    -1.332916e-09, -1.394217e-09, -1.5003e-09, -1.629497e-09, -1.908113e-09, 
    -2.39026e-09, -3.085911e-09, -3.857592e-09, -4.725571e-09, -5.718426e-09,
  -2.02627e-09, -1.871066e-09, -1.664003e-09, -1.458869e-09, -1.363064e-09, 
    -1.345526e-09, -1.363637e-09, -1.411251e-09, -1.439176e-09, 
    -1.531877e-09, -1.829821e-09, -2.362418e-09, -3.075586e-09, 
    -3.826075e-09, -4.706754e-09,
  -2.469085e-09, -2.394882e-09, -2.25195e-09, -2.003251e-09, -1.748884e-09, 
    -1.583817e-09, -1.462479e-09, -1.457305e-09, -1.443335e-09, 
    -1.432278e-09, -1.564627e-09, -1.878067e-09, -2.425912e-09, 
    -3.122399e-09, -3.960965e-09,
  -2.648773e-09, -2.65163e-09, -2.600676e-09, -2.420109e-09, -2.176233e-09, 
    -1.954229e-09, -1.782452e-09, -1.635321e-09, -1.566414e-09, 
    -1.473849e-09, -1.45841e-09, -1.595077e-09, -1.969272e-09, -2.558022e-09, 
    -3.33104e-09,
  -2.36952e-09, -2.541173e-09, -2.556938e-09, -2.597175e-09, -2.427555e-09, 
    -2.254064e-09, -2.125893e-09, -1.971098e-09, -1.793414e-09, 
    -1.604782e-09, -1.462651e-09, -1.446897e-09, -1.660299e-09, -2.13461e-09, 
    -2.818996e-09,
  -3.377449e-09, -3.757368e-09, -4.290985e-09, -5.101607e-09, -6.133443e-09, 
    -7.266532e-09, -8.384893e-09, -9.438609e-09, -1.056432e-08, 
    -1.189267e-08, -1.368245e-08, -1.571815e-08, -1.83501e-08, -2.122266e-08, 
    -2.421376e-08,
  -2.366588e-09, -2.723056e-09, -3.164624e-09, -3.645786e-09, -4.233555e-09, 
    -4.954205e-09, -5.87913e-09, -6.974883e-09, -8.170411e-09, -9.28685e-09, 
    -1.061049e-08, -1.203209e-08, -1.372312e-08, -1.583332e-08, -1.85748e-08,
  -1.783118e-09, -1.939389e-09, -2.197011e-09, -2.550769e-09, -2.924418e-09, 
    -3.369509e-09, -3.912523e-09, -4.646873e-09, -5.648559e-09, 
    -6.805862e-09, -8.04834e-09, -9.284362e-09, -1.060019e-08, -1.197501e-08, 
    -1.368246e-08,
  -1.503857e-09, -1.599542e-09, -1.698362e-09, -1.831087e-09, -2.049312e-09, 
    -2.346637e-09, -2.678623e-09, -3.124666e-09, -3.785817e-09, -4.66563e-09, 
    -5.697206e-09, -6.871712e-09, -8.10005e-09, -9.346864e-09, -1.058444e-08,
  -1.354485e-09, -1.332111e-09, -1.281519e-09, -1.297798e-09, -1.425044e-09, 
    -1.641519e-09, -1.915501e-09, -2.236098e-09, -2.63542e-09, -3.174862e-09, 
    -3.858892e-09, -4.656914e-09, -5.761746e-09, -7.069238e-09, -8.41137e-09,
  -1.415998e-09, -1.337848e-09, -1.25072e-09, -1.186819e-09, -1.191683e-09, 
    -1.263013e-09, -1.429462e-09, -1.72502e-09, -1.979849e-09, -2.196202e-09, 
    -2.590236e-09, -2.906254e-09, -3.490728e-09, -4.465562e-09, -5.826756e-09,
  -2.021135e-09, -1.753642e-09, -1.597944e-09, -1.475697e-09, -1.343615e-09, 
    -1.301854e-09, -1.299573e-09, -1.381997e-09, -1.641e-09, -1.785107e-09, 
    -1.845985e-09, -1.937486e-09, -2.152986e-09, -2.803598e-09, -3.72343e-09,
  -2.545715e-09, -2.518734e-09, -2.292431e-09, -2.055014e-09, -1.824398e-09, 
    -1.678089e-09, -1.572528e-09, -1.507786e-09, -1.451541e-09, 
    -1.577915e-09, -1.722587e-09, -1.715125e-09, -1.62879e-09, -1.611574e-09, 
    -2.107101e-09,
  -2.593152e-09, -2.61632e-09, -2.6358e-09, -2.530795e-09, -2.422254e-09, 
    -2.329594e-09, -2.268143e-09, -2.151187e-09, -1.909633e-09, 
    -1.737583e-09, -1.696032e-09, -1.922551e-09, -1.886411e-09, 
    -1.647968e-09, -1.390549e-09,
  -2.32487e-09, -2.455689e-09, -2.490463e-09, -2.548e-09, -2.452716e-09, 
    -2.486932e-09, -2.498631e-09, -2.506142e-09, -2.429995e-09, 
    -2.363446e-09, -2.185883e-09, -2.062814e-09, -2.048832e-09, -2.02225e-09, 
    -1.854109e-09,
  -2.206294e-09, -2.478075e-09, -2.916933e-09, -3.533903e-09, -4.40594e-09, 
    -5.444054e-09, -6.942404e-09, -8.72843e-09, -1.054732e-08, -1.365151e-08, 
    -1.755426e-08, -2.13817e-08, -2.289897e-08, -2.256575e-08, -2.122059e-08,
  -1.989641e-09, -2.137621e-09, -2.358129e-09, -2.743206e-09, -3.298089e-09, 
    -4.115792e-09, -5.051549e-09, -6.354679e-09, -7.729002e-09, 
    -9.509182e-09, -1.20105e-08, -1.543277e-08, -1.946117e-08, -2.213311e-08, 
    -2.330013e-08,
  -1.786103e-09, -1.842683e-09, -1.934754e-09, -2.110872e-09, -2.465845e-09, 
    -3.019064e-09, -3.789367e-09, -4.729376e-09, -5.886014e-09, 
    -7.151768e-09, -8.63784e-09, -1.066187e-08, -1.36758e-08, -1.767014e-08, 
    -2.07046e-08,
  -1.454712e-09, -1.572152e-09, -1.557555e-09, -1.649826e-09, -1.811106e-09, 
    -2.164659e-09, -2.706301e-09, -3.429843e-09, -4.344012e-09, 
    -5.486505e-09, -6.732416e-09, -8.105389e-09, -9.76794e-09, -1.217882e-08, 
    -1.576077e-08,
  -1.159298e-09, -1.204975e-09, -1.166305e-09, -1.153739e-09, -1.225113e-09, 
    -1.426248e-09, -1.910555e-09, -2.560425e-09, -3.30086e-09, -4.152205e-09, 
    -5.239044e-09, -6.361367e-09, -7.621283e-09, -9.196667e-09, -1.118701e-08,
  -1.001064e-09, -1.057742e-09, -1.082588e-09, -9.997414e-10, -9.758963e-10, 
    -9.886501e-10, -1.161217e-09, -1.633117e-09, -2.36901e-09, -3.199846e-09, 
    -4.12608e-09, -5.109037e-09, -6.121147e-09, -7.327976e-09, -8.840796e-09,
  -1.018651e-09, -1.094838e-09, -1.172206e-09, -1.197551e-09, -1.039929e-09, 
    -1.003307e-09, -1.011031e-09, -1.197335e-09, -1.591787e-09, 
    -2.222411e-09, -3.060412e-09, -4.100852e-09, -5.112609e-09, -5.922e-09, 
    -7.148124e-09,
  -1.098018e-09, -1.215109e-09, -1.391383e-09, -1.600009e-09, -1.585675e-09, 
    -1.386623e-09, -1.199316e-09, -1.108504e-09, -1.220818e-09, 
    -1.625014e-09, -2.218253e-09, -3.012384e-09, -4.080951e-09, 
    -5.129865e-09, -5.984511e-09,
  -1.163816e-09, -1.24894e-09, -1.418822e-09, -1.642492e-09, -1.944144e-09, 
    -1.945262e-09, -1.743692e-09, -1.521171e-09, -1.318164e-09, 
    -1.306206e-09, -1.653431e-09, -2.204321e-09, -3.07787e-09, -4.060249e-09, 
    -5.104376e-09,
  -1.152402e-09, -1.297569e-09, -1.397814e-09, -1.510622e-09, -1.722023e-09, 
    -1.976401e-09, -1.919743e-09, -1.821835e-09, -1.700225e-09, 
    -1.528223e-09, -1.48188e-09, -1.705061e-09, -2.272847e-09, -3.141122e-09, 
    -4.083304e-09,
  -3.399987e-09, -3.586642e-09, -3.690388e-09, -3.720495e-09, -3.881685e-09, 
    -3.904509e-09, -4.06533e-09, -3.694394e-09, -3.991851e-09, -4.665688e-09, 
    -5.958268e-09, -7.514798e-09, -9.459774e-09, -1.144173e-08, -1.344923e-08,
  -2.652165e-09, -2.930685e-09, -3.163525e-09, -3.462381e-09, -3.592896e-09, 
    -3.906612e-09, -4.197076e-09, -3.952692e-09, -3.839346e-09, 
    -4.125563e-09, -4.492683e-09, -5.386839e-09, -6.774733e-09, 
    -8.649474e-09, -1.067618e-08,
  -1.94215e-09, -2.000529e-09, -2.129845e-09, -2.456768e-09, -2.860203e-09, 
    -3.083132e-09, -3.619186e-09, -3.670721e-09, -3.440166e-09, 
    -3.393078e-09, -3.497422e-09, -4.005534e-09, -4.829312e-09, 
    -6.127132e-09, -7.922966e-09,
  -1.40919e-09, -1.413365e-09, -1.349785e-09, -1.576756e-09, -1.902901e-09, 
    -2.198211e-09, -2.445345e-09, -2.817e-09, -2.963969e-09, -3.001235e-09, 
    -3.02598e-09, -3.222752e-09, -3.628025e-09, -4.391323e-09, -5.609337e-09,
  -1.147039e-09, -1.174664e-09, -1.153662e-09, -1.179583e-09, -1.341173e-09, 
    -1.512819e-09, -1.65688e-09, -1.949224e-09, -2.250782e-09, -2.589901e-09, 
    -2.717242e-09, -2.865536e-09, -3.047374e-09, -3.336716e-09, -4.060058e-09,
  -1.092996e-09, -1.093511e-09, -1.191474e-09, -1.103822e-09, -1.077187e-09, 
    -1.160576e-09, -1.230324e-09, -1.411402e-09, -1.605361e-09, 
    -1.779376e-09, -2.107932e-09, -2.422738e-09, -2.688769e-09, 
    -2.915131e-09, -3.23357e-09,
  -1.039513e-09, -1.029972e-09, -1.060063e-09, -1.102652e-09, -9.356912e-10, 
    -9.171581e-10, -1.011438e-09, -1.149498e-09, -1.301003e-09, 
    -1.392676e-09, -1.591265e-09, -1.863727e-09, -2.179091e-09, 
    -2.461325e-09, -2.729776e-09,
  -9.644938e-10, -1.020235e-09, -9.72681e-10, -8.547684e-10, -7.168684e-10, 
    -5.183112e-10, -5.863968e-10, -7.035059e-10, -8.829111e-10, 
    -1.051463e-09, -1.22663e-09, -1.416369e-09, -1.684506e-09, -1.984614e-09, 
    -2.290766e-09,
  -7.517104e-10, -8.638483e-10, -9.025539e-10, -9.215851e-10, -6.88359e-10, 
    -4.584082e-10, -3.940878e-10, -6.229201e-10, -8.045078e-10, 
    -9.342876e-10, -1.031956e-09, -1.077059e-09, -1.252481e-09, 
    -1.543462e-09, -1.866697e-09,
  -6.979243e-10, -7.367324e-10, -9.010306e-10, -9.932409e-10, -9.076724e-10, 
    -7.628488e-10, -5.336658e-10, -4.30182e-10, -5.91084e-10, -7.868089e-10, 
    -8.27598e-10, -8.917196e-10, -9.130791e-10, -1.080477e-09, -1.3902e-09,
  -6.733905e-09, -7.68528e-09, -8.923186e-09, -1.020617e-08, -1.132032e-08, 
    -1.226743e-08, -1.302713e-08, -1.308957e-08, -1.235656e-08, 
    -1.207491e-08, -1.072917e-08, -9.04641e-09, -7.386488e-09, -6.483571e-09, 
    -6.228706e-09,
  -4.081077e-09, -4.677102e-09, -5.396211e-09, -6.225653e-09, -7.17886e-09, 
    -8.362201e-09, -9.643488e-09, -1.129064e-08, -1.207165e-08, 
    -1.210339e-08, -1.136898e-08, -9.775714e-09, -8.649407e-09, 
    -7.399672e-09, -6.573033e-09,
  -2.91366e-09, -3.165897e-09, -3.538926e-09, -4.012327e-09, -4.556335e-09, 
    -5.297871e-09, -6.133339e-09, -7.454092e-09, -8.960651e-09, 
    -9.833167e-09, -1.019347e-08, -9.646699e-09, -8.109147e-09, -6.8649e-09, 
    -6.009765e-09,
  -2.366129e-09, -2.454014e-09, -2.602449e-09, -2.825187e-09, -3.122727e-09, 
    -3.491371e-09, -3.999714e-09, -4.566603e-09, -5.44863e-09, -6.661701e-09, 
    -7.65951e-09, -8.290412e-09, -7.929147e-09, -6.583244e-09, -5.3289e-09,
  -2.054245e-09, -2.174336e-09, -2.23691e-09, -2.301003e-09, -2.41315e-09, 
    -2.590004e-09, -2.844498e-09, -3.18442e-09, -3.609984e-09, -4.101144e-09, 
    -5.133572e-09, -6.114947e-09, -7.092248e-09, -6.928788e-09, -5.979647e-09,
  -1.624759e-09, -1.789753e-09, -1.912666e-09, -1.989565e-09, -2.046926e-09, 
    -2.12238e-09, -2.228671e-09, -2.410279e-09, -2.709555e-09, -3.011982e-09, 
    -3.450905e-09, -4.416413e-09, -5.410705e-09, -6.239262e-09, -6.352138e-09,
  -1.09864e-09, -1.301942e-09, -1.468019e-09, -1.583108e-09, -1.685614e-09, 
    -1.775288e-09, -1.845832e-09, -1.948628e-09, -2.092669e-09, 
    -2.333661e-09, -2.654968e-09, -3.068828e-09, -3.872445e-09, 
    -4.694752e-09, -5.473954e-09,
  -5.14047e-10, -7.33927e-10, -9.264483e-10, -1.087208e-09, -1.222207e-09, 
    -1.357135e-09, -1.505862e-09, -1.652503e-09, -1.761069e-09, 
    -1.934265e-09, -2.200638e-09, -2.505526e-09, -2.884682e-09, 
    -3.541608e-09, -4.189038e-09,
  -1.265652e-10, -2.440435e-10, -3.844932e-10, -5.733976e-10, -7.453747e-10, 
    -9.074423e-10, -1.100263e-09, -1.32227e-09, -1.495559e-09, -1.61175e-09, 
    -1.755293e-09, -2.005601e-09, -2.323054e-09, -2.746811e-09, -3.278745e-09,
  1.016978e-11, -1.020131e-10, -1.736878e-10, -2.726185e-10, -3.881258e-10, 
    -5.564509e-10, -8.363489e-10, -1.031087e-09, -1.158173e-09, 
    -1.321892e-09, -1.42302e-09, -1.592362e-09, -1.859019e-09, -2.197781e-09, 
    -2.582906e-09,
  -6.059494e-09, -6.275822e-09, -6.575724e-09, -6.988932e-09, -7.682267e-09, 
    -8.488624e-09, -9.57133e-09, -1.064008e-08, -1.147764e-08, -1.177076e-08, 
    -1.226953e-08, -1.321153e-08, -1.425452e-08, -1.569373e-08, -1.742712e-08,
  -5.254485e-09, -5.74137e-09, -6.136632e-09, -6.468284e-09, -6.862585e-09, 
    -7.477651e-09, -8.348895e-09, -9.423218e-09, -1.078049e-08, 
    -1.201828e-08, -1.274678e-08, -1.328577e-08, -1.400667e-08, 
    -1.482695e-08, -1.575643e-08,
  -3.783289e-09, -4.534018e-09, -5.245978e-09, -5.794797e-09, -6.211113e-09, 
    -6.620258e-09, -7.172508e-09, -7.950394e-09, -9.039024e-09, 
    -1.045863e-08, -1.189768e-08, -1.319668e-08, -1.43326e-08, -1.504846e-08, 
    -1.560977e-08,
  -2.106789e-09, -2.887661e-09, -3.684133e-09, -4.527462e-09, -5.271578e-09, 
    -5.850091e-09, -6.323356e-09, -6.809779e-09, -7.406189e-09, 
    -8.267541e-09, -9.551095e-09, -1.101015e-08, -1.259664e-08, 
    -1.409413e-08, -1.54649e-08,
  -1.10656e-09, -1.592694e-09, -2.194634e-09, -2.938491e-09, -3.786879e-09, 
    -4.644026e-09, -5.394252e-09, -5.986114e-09, -6.460446e-09, 
    -6.895383e-09, -7.465888e-09, -8.347492e-09, -9.540253e-09, 
    -1.110951e-08, -1.255156e-08,
  -5.977812e-10, -8.759058e-10, -1.268056e-09, -1.771985e-09, -2.36845e-09, 
    -3.144718e-09, -4.003134e-09, -4.8807e-09, -5.637683e-09, -6.176355e-09, 
    -6.558107e-09, -6.916118e-09, -7.404356e-09, -8.190471e-09, -9.273482e-09,
  -4.135392e-10, -5.784756e-10, -8.167821e-10, -1.125037e-09, -1.565683e-09, 
    -2.06615e-09, -2.625781e-09, -3.357623e-09, -4.238388e-09, -5.14062e-09, 
    -5.900509e-09, -6.353615e-09, -6.620018e-09, -6.850112e-09, -7.230041e-09,
  -2.33941e-10, -3.747083e-10, -5.125075e-10, -7.018234e-10, -9.399282e-10, 
    -1.318724e-09, -1.82178e-09, -2.412849e-09, -3.034394e-09, -3.737195e-09, 
    -4.527354e-09, -5.353984e-09, -5.995704e-09, -6.435114e-09, -6.565846e-09,
  1.890896e-11, -8.725159e-11, -2.209312e-10, -3.802059e-10, -5.531484e-10, 
    -7.686228e-10, -1.039313e-09, -1.40273e-09, -1.917543e-09, -2.54925e-09, 
    -3.306479e-09, -4.102779e-09, -4.87608e-09, -5.451097e-09, -5.982108e-09,
  2.053025e-10, 2.25672e-10, 2.183335e-10, 1.615882e-10, 2.628229e-11, 
    -1.97861e-10, -5.63887e-10, -9.054242e-10, -1.216686e-09, -1.664987e-09, 
    -2.105156e-09, -2.728958e-09, -3.452483e-09, -4.309209e-09, -5.011602e-09,
  -3.498334e-09, -3.795133e-09, -4.459673e-09, -5.243749e-09, -5.681565e-09, 
    -5.346027e-09, -4.378015e-09, -4.294607e-09, -5.175573e-09, 
    -6.944992e-09, -9.672992e-09, -1.240623e-08, -1.415248e-08, 
    -1.584804e-08, -1.76122e-08,
  -2.995459e-09, -3.328579e-09, -3.648276e-09, -4.240804e-09, -4.888447e-09, 
    -5.603684e-09, -5.543989e-09, -4.596504e-09, -4.358094e-09, 
    -5.006814e-09, -6.557821e-09, -8.991157e-09, -1.152304e-08, 
    -1.339769e-08, -1.545993e-08,
  -2.431117e-09, -2.801869e-09, -3.154907e-09, -3.527028e-09, -4.071183e-09, 
    -4.711425e-09, -5.390217e-09, -5.269874e-09, -4.473951e-09, -4.33924e-09, 
    -5.020953e-09, -6.488324e-09, -8.830233e-09, -1.104146e-08, -1.303116e-08,
  -1.845739e-09, -2.176561e-09, -2.560417e-09, -2.993542e-09, -3.403233e-09, 
    -3.965961e-09, -4.634788e-09, -5.210647e-09, -5.07534e-09, -4.473285e-09, 
    -4.446069e-09, -5.125443e-09, -6.59156e-09, -8.619764e-09, -1.074038e-08,
  -1.35501e-09, -1.605248e-09, -1.91513e-09, -2.320963e-09, -2.767493e-09, 
    -3.261769e-09, -3.853983e-09, -4.639341e-09, -5.173129e-09, 
    -5.028737e-09, -4.56159e-09, -4.699193e-09, -5.577881e-09, -7.011408e-09, 
    -8.70237e-09,
  -9.292723e-10, -1.128648e-09, -1.374282e-09, -1.6789e-09, -2.065481e-09, 
    -2.571404e-09, -3.076168e-09, -3.721933e-09, -4.537311e-09, 
    -5.102248e-09, -5.145868e-09, -4.917122e-09, -5.155448e-09, 
    -6.052342e-09, -7.272534e-09,
  -6.65651e-10, -7.461073e-10, -9.365718e-10, -1.168078e-09, -1.444141e-09, 
    -1.836888e-09, -2.374557e-09, -2.914224e-09, -3.658053e-09, 
    -4.428158e-09, -5.042875e-09, -5.315005e-09, -5.195815e-09, 
    -5.481791e-09, -6.337159e-09,
  -5.054072e-10, -5.547844e-10, -6.527213e-10, -8.252194e-10, -1.014788e-09, 
    -1.24222e-09, -1.599377e-09, -2.102314e-09, -2.66098e-09, -3.456329e-09, 
    -4.313106e-09, -4.990979e-09, -5.309091e-09, -5.37902e-09, -5.799387e-09,
  -5.984793e-10, -5.765982e-10, -5.665005e-10, -6.4465e-10, -8.043066e-10, 
    -9.823281e-10, -1.20332e-09, -1.525447e-09, -1.981359e-09, -2.529047e-09, 
    -3.247163e-09, -4.111661e-09, -4.84903e-09, -5.212849e-09, -5.589826e-09,
  -6.798875e-10, -6.663837e-10, -6.783711e-10, -6.625019e-10, -7.068138e-10, 
    -8.381697e-10, -1.051001e-09, -1.262712e-09, -1.531718e-09, 
    -1.995127e-09, -2.555294e-09, -3.192452e-09, -3.990684e-09, 
    -4.740386e-09, -5.238229e-09,
  -3.322401e-09, -3.499933e-09, -3.62579e-09, -3.567045e-09, -3.824957e-09, 
    -4.394656e-09, -4.830243e-09, -4.783221e-09, -5.100559e-09, 
    -6.198063e-09, -7.669077e-09, -9.397183e-09, -1.143248e-08, 
    -1.268668e-08, -1.322229e-08,
  -2.740706e-09, -2.944181e-09, -3.168636e-09, -3.295791e-09, -3.424781e-09, 
    -3.690167e-09, -4.267508e-09, -4.643196e-09, -4.456929e-09, 
    -4.490685e-09, -5.137897e-09, -6.238212e-09, -8.235922e-09, 
    -1.068141e-08, -1.211981e-08,
  -2.402245e-09, -2.566509e-09, -2.76044e-09, -2.975793e-09, -3.126048e-09, 
    -3.382922e-09, -3.747551e-09, -4.371619e-09, -4.649286e-09, 
    -4.134266e-09, -4.047173e-09, -4.332495e-09, -5.325935e-09, 
    -7.409722e-09, -1.048771e-08,
  -1.853528e-09, -2.025613e-09, -2.176479e-09, -2.395121e-09, -2.64563e-09, 
    -2.910608e-09, -3.27263e-09, -3.812147e-09, -4.491784e-09, -4.772814e-09, 
    -4.128177e-09, -3.814571e-09, -3.956092e-09, -4.834131e-09, -6.807389e-09,
  -1.371727e-09, -1.562921e-09, -1.732714e-09, -1.935142e-09, -2.17946e-09, 
    -2.425672e-09, -2.705856e-09, -3.118531e-09, -3.808334e-09, 
    -4.613483e-09, -4.68702e-09, -3.926594e-09, -3.369766e-09, -3.428461e-09, 
    -4.470223e-09,
  -1.003193e-09, -1.120386e-09, -1.317173e-09, -1.536819e-09, -1.755896e-09, 
    -2.006492e-09, -2.251767e-09, -2.535982e-09, -3.032713e-09, 
    -3.879497e-09, -4.715258e-09, -4.536589e-09, -3.612379e-09, 
    -3.000065e-09, -3.306308e-09,
  -8.449021e-10, -8.86078e-10, -9.619502e-10, -1.152681e-09, -1.384283e-09, 
    -1.633232e-09, -1.893664e-09, -2.149474e-09, -2.444406e-09, 
    -3.017886e-09, -3.974799e-09, -4.623833e-09, -4.412169e-09, 
    -3.543743e-09, -3.136368e-09,
  -7.249455e-10, -7.61021e-10, -7.955919e-10, -8.675054e-10, -1.026757e-09, 
    -1.258595e-09, -1.538655e-09, -1.838906e-09, -2.103185e-09, 
    -2.469957e-09, -3.04178e-09, -3.989571e-09, -4.601605e-09, -4.385091e-09, 
    -3.655414e-09,
  -6.458894e-10, -6.362448e-10, -6.610045e-10, -6.789599e-10, -7.9182e-10, 
    -8.986736e-10, -1.123853e-09, -1.446709e-09, -1.771374e-09, 
    -2.110227e-09, -2.492175e-09, -3.092595e-09, -4.017841e-09, 
    -4.552422e-09, -4.562787e-09,
  -7.418786e-10, -6.944776e-10, -6.032497e-10, -5.802187e-10, -5.74535e-10, 
    -6.295069e-10, -7.580147e-10, -1.015338e-09, -1.354986e-09, 
    -1.733647e-09, -2.116566e-09, -2.489717e-09, -3.209269e-09, 
    -4.047687e-09, -4.521136e-09,
  -9.592508e-09, -1.067708e-08, -1.171497e-08, -1.239738e-08, -1.267899e-08, 
    -1.262051e-08, -1.210079e-08, -1.140183e-08, -1.156371e-08, 
    -1.225137e-08, -1.331231e-08, -1.448219e-08, -1.567287e-08, 
    -1.654391e-08, -1.747596e-08,
  -6.606706e-09, -7.893344e-09, -9.023448e-09, -1.008007e-08, -1.099846e-08, 
    -1.168147e-08, -1.185214e-08, -1.170471e-08, -1.107276e-08, 
    -1.092379e-08, -1.137318e-08, -1.231605e-08, -1.340869e-08, 
    -1.427593e-08, -1.513811e-08,
  -4.367023e-09, -5.041896e-09, -6.052318e-09, -7.305764e-09, -8.562909e-09, 
    -9.644931e-09, -1.049845e-08, -1.099917e-08, -1.088884e-08, 
    -1.045166e-08, -1.019906e-08, -1.048248e-08, -1.123724e-08, 
    -1.220715e-08, -1.305281e-08,
  -3.649034e-09, -3.940414e-09, -4.383746e-09, -5.004288e-09, -5.934383e-09, 
    -7.116063e-09, -8.334971e-09, -9.287395e-09, -9.933527e-09, 
    -1.011429e-08, -9.805004e-09, -9.553196e-09, -9.675161e-09, 
    -9.968096e-09, -1.063221e-08,
  -2.911075e-09, -3.183816e-09, -3.522588e-09, -3.965032e-09, -4.473686e-09, 
    -5.131221e-09, -6.0177e-09, -7.021296e-09, -7.905189e-09, -8.562087e-09, 
    -9.033847e-09, -9.244161e-09, -9.062752e-09, -9.005441e-09, -8.991417e-09,
  -2.224716e-09, -2.478955e-09, -2.802625e-09, -3.224535e-09, -3.645711e-09, 
    -4.068159e-09, -4.562261e-09, -5.119163e-09, -5.794835e-09, 
    -6.552023e-09, -7.298754e-09, -7.936563e-09, -8.352107e-09, 
    -8.338773e-09, -8.377503e-09,
  -1.836982e-09, -1.958631e-09, -2.18348e-09, -2.53345e-09, -2.957063e-09, 
    -3.334043e-09, -3.699322e-09, -4.051177e-09, -4.432495e-09, 
    -4.907272e-09, -5.555273e-09, -6.330949e-09, -6.970508e-09, -7.32557e-09, 
    -7.573614e-09,
  -1.737014e-09, -1.753274e-09, -1.841452e-09, -1.999623e-09, -2.290006e-09, 
    -2.64424e-09, -2.992252e-09, -3.31648e-09, -3.605301e-09, -3.911194e-09, 
    -4.262575e-09, -4.793292e-09, -5.457371e-09, -6.10871e-09, -6.535403e-09,
  -1.550683e-09, -1.544684e-09, -1.605327e-09, -1.710575e-09, -1.847906e-09, 
    -2.108231e-09, -2.365716e-09, -2.642809e-09, -2.935606e-09, 
    -3.251716e-09, -3.536328e-09, -3.817673e-09, -4.220829e-09, 
    -4.700564e-09, -5.305805e-09,
  -1.246319e-09, -1.30796e-09, -1.36457e-09, -1.435409e-09, -1.543498e-09, 
    -1.732994e-09, -1.981011e-09, -2.208052e-09, -2.405238e-09, 
    -2.648094e-09, -2.943801e-09, -3.194288e-09, -3.499282e-09, 
    -3.834847e-09, -4.2048e-09,
  -7.218603e-09, -7.238998e-09, -7.279933e-09, -7.427654e-09, -7.60505e-09, 
    -7.885171e-09, -8.292105e-09, -8.691485e-09, -8.544492e-09, 
    -8.197344e-09, -8.075109e-09, -8.11992e-09, -8.554192e-09, -9.114569e-09, 
    -9.688745e-09,
  -6.580942e-09, -6.625327e-09, -6.727797e-09, -6.849144e-09, -7.008255e-09, 
    -7.233545e-09, -7.612533e-09, -8.119013e-09, -8.633539e-09, 
    -8.716502e-09, -8.382815e-09, -8.193027e-09, -8.327748e-09, -8.67728e-09, 
    -9.306605e-09,
  -6.066502e-09, -6.138361e-09, -6.256407e-09, -6.352405e-09, -6.503746e-09, 
    -6.735356e-09, -7.050455e-09, -7.459971e-09, -8.033721e-09, 
    -8.578517e-09, -8.810058e-09, -8.605473e-09, -8.339298e-09, 
    -8.438043e-09, -8.853482e-09,
  -5.470548e-09, -5.46206e-09, -5.522861e-09, -5.675674e-09, -5.888003e-09, 
    -6.126729e-09, -6.405722e-09, -6.846622e-09, -7.350987e-09, 
    -7.930165e-09, -8.536317e-09, -8.875253e-09, -8.783157e-09, 
    -8.618226e-09, -8.560868e-09,
  -4.767465e-09, -4.760953e-09, -4.786318e-09, -4.976739e-09, -5.188995e-09, 
    -5.494244e-09, -5.809621e-09, -6.190409e-09, -6.697349e-09, 
    -7.323547e-09, -8.020211e-09, -8.723597e-09, -9.013537e-09, 
    -9.016305e-09, -8.80877e-09,
  -4.053651e-09, -4.010424e-09, -3.99763e-09, -4.082511e-09, -4.265002e-09, 
    -4.596402e-09, -5.0298e-09, -5.480022e-09, -5.989973e-09, -6.565547e-09, 
    -7.353166e-09, -8.171923e-09, -8.986135e-09, -9.24554e-09, -9.238677e-09,
  -3.794574e-09, -3.632945e-09, -3.633878e-09, -3.516934e-09, -3.49592e-09, 
    -3.665606e-09, -3.9748e-09, -4.435847e-09, -4.997215e-09, -5.717406e-09, 
    -6.485572e-09, -7.451495e-09, -8.333631e-09, -9.200272e-09, -9.449939e-09,
  -3.478201e-09, -3.495704e-09, -3.454658e-09, -3.271056e-09, -3.096815e-09, 
    -3.11516e-09, -3.29617e-09, -3.548256e-09, -3.942828e-09, -4.519138e-09, 
    -5.285459e-09, -6.304143e-09, -7.429191e-09, -8.489763e-09, -9.246922e-09,
  -3.043815e-09, -3.288626e-09, -3.319393e-09, -3.134195e-09, -2.877969e-09, 
    -2.735645e-09, -2.84255e-09, -3.017703e-09, -3.265987e-09, -3.654098e-09, 
    -4.222023e-09, -4.937728e-09, -6.040163e-09, -7.305129e-09, -8.457514e-09,
  -2.630435e-09, -2.95996e-09, -3.19793e-09, -3.433e-09, -3.282246e-09, 
    -2.883939e-09, -2.801819e-09, -2.795767e-09, -2.745874e-09, 
    -2.977858e-09, -3.336738e-09, -4.042874e-09, -4.850694e-09, 
    -5.867425e-09, -7.223006e-09,
  -1.34976e-08, -1.362988e-08, -1.372881e-08, -1.375006e-08, -1.369743e-08, 
    -1.356805e-08, -1.337707e-08, -1.314041e-08, -1.288104e-08, 
    -1.260757e-08, -1.233195e-08, -1.208549e-08, -1.186394e-08, -1.17213e-08, 
    -1.162508e-08,
  -1.085142e-08, -1.105105e-08, -1.121482e-08, -1.133606e-08, -1.140624e-08, 
    -1.140515e-08, -1.137102e-08, -1.131276e-08, -1.123985e-08, -1.11364e-08, 
    -1.100943e-08, -1.087124e-08, -1.075974e-08, -1.071058e-08, -1.065172e-08,
  -8.576577e-09, -8.829288e-09, -9.020592e-09, -9.194038e-09, -9.343791e-09, 
    -9.447122e-09, -9.516735e-09, -9.5587e-09, -9.558803e-09, -9.531629e-09, 
    -9.479379e-09, -9.398445e-09, -9.325634e-09, -9.283625e-09, -9.252052e-09,
  -6.265025e-09, -6.570632e-09, -6.835159e-09, -7.067242e-09, -7.28165e-09, 
    -7.449906e-09, -7.585822e-09, -7.694174e-09, -7.743036e-09, 
    -7.840968e-09, -7.933672e-09, -7.981932e-09, -8.054615e-09, 
    -8.132036e-09, -8.259301e-09,
  -4.144136e-09, -4.427657e-09, -4.729647e-09, -4.996674e-09, -5.251203e-09, 
    -5.451634e-09, -5.625257e-09, -5.782073e-09, -5.980953e-09, 
    -6.229818e-09, -6.439648e-09, -6.568042e-09, -6.70449e-09, -6.787284e-09, 
    -6.897436e-09,
  -2.723052e-09, -2.937631e-09, -3.172433e-09, -3.432744e-09, -3.701024e-09, 
    -3.954939e-09, -4.201091e-09, -4.449609e-09, -4.767295e-09, 
    -5.050329e-09, -5.230139e-09, -5.365343e-09, -5.350858e-09, -5.42108e-09, 
    -5.491644e-09,
  -1.996547e-09, -2.12815e-09, -2.290369e-09, -2.458184e-09, -2.64056e-09, 
    -2.84743e-09, -3.086624e-09, -3.379899e-09, -3.639502e-09, -3.861283e-09, 
    -4.042978e-09, -4.181463e-09, -4.201495e-09, -4.343989e-09, -4.417164e-09,
  -1.66688e-09, -1.727166e-09, -1.817748e-09, -1.913386e-09, -2.057461e-09, 
    -2.201791e-09, -2.423582e-09, -2.647727e-09, -2.896261e-09, 
    -3.217346e-09, -3.385243e-09, -3.455045e-09, -3.516039e-09, 
    -3.689577e-09, -3.841797e-09,
  -1.43026e-09, -1.519398e-09, -1.661482e-09, -1.72662e-09, -1.809261e-09, 
    -1.948599e-09, -2.091616e-09, -2.289016e-09, -2.379184e-09, 
    -2.691416e-09, -2.82064e-09, -2.898046e-09, -3.012722e-09, -3.122966e-09, 
    -3.260405e-09,
  -1.074265e-09, -1.215134e-09, -1.348038e-09, -1.497741e-09, -1.609141e-09, 
    -1.768725e-09, -1.90015e-09, -2.085869e-09, -2.282659e-09, -2.598318e-09, 
    -3.001096e-09, -3.430915e-09, -3.235107e-09, -3.171502e-09, -3.317018e-09,
  -1.230002e-08, -1.281963e-08, -1.335566e-08, -1.380938e-08, -1.426472e-08, 
    -1.462316e-08, -1.491428e-08, -1.514934e-08, -1.537446e-08, 
    -1.559031e-08, -1.576589e-08, -1.589216e-08, -1.596313e-08, 
    -1.596697e-08, -1.591378e-08,
  -1.028754e-08, -1.09386e-08, -1.160671e-08, -1.218402e-08, -1.272794e-08, 
    -1.318227e-08, -1.361326e-08, -1.395271e-08, -1.419522e-08, -1.43756e-08, 
    -1.450276e-08, -1.459284e-08, -1.463459e-08, -1.465765e-08, -1.463071e-08,
  -7.701392e-09, -8.630741e-09, -9.460532e-09, -1.017331e-08, -1.082623e-08, 
    -1.140214e-08, -1.190183e-08, -1.232257e-08, -1.269677e-08, 
    -1.297198e-08, -1.316721e-08, -1.3296e-08, -1.335483e-08, -1.336774e-08, 
    -1.333145e-08,
  -4.833914e-09, -5.716742e-09, -6.633548e-09, -7.583131e-09, -8.464815e-09, 
    -9.220544e-09, -9.868224e-09, -1.041576e-08, -1.090084e-08, 
    -1.128835e-08, -1.160665e-08, -1.184066e-08, -1.199225e-08, 
    -1.206716e-08, -1.206936e-08,
  -2.588903e-09, -3.128469e-09, -3.772474e-09, -4.512682e-09, -5.339306e-09, 
    -6.207069e-09, -7.077862e-09, -7.891556e-09, -8.589388e-09, 
    -9.156421e-09, -9.605172e-09, -9.968943e-09, -1.023424e-08, 
    -1.040715e-08, -1.053811e-08,
  -1.537082e-09, -1.782986e-09, -2.085379e-09, -2.467021e-09, -2.928892e-09, 
    -3.469164e-09, -4.097824e-09, -4.791467e-09, -5.553575e-09, 
    -6.278755e-09, -6.957584e-09, -7.502419e-09, -7.967859e-09, 
    -8.259472e-09, -8.498882e-09,
  -1.089826e-09, -1.215656e-09, -1.356458e-09, -1.523379e-09, -1.727244e-09, 
    -1.978646e-09, -2.298682e-09, -2.674096e-09, -3.128376e-09, 
    -3.644814e-09, -4.232843e-09, -4.814241e-09, -5.385716e-09, 
    -5.868503e-09, -6.344244e-09,
  -8.050663e-10, -8.97133e-10, -9.988769e-10, -1.106091e-09, -1.224698e-09, 
    -1.351277e-09, -1.498874e-09, -1.666644e-09, -1.871937e-09, -2.12101e-09, 
    -2.419782e-09, -2.763026e-09, -3.149649e-09, -3.581734e-09, -4.099221e-09,
  -6.880698e-10, -7.324669e-10, -7.870816e-10, -8.578455e-10, -9.445087e-10, 
    -1.044248e-09, -1.151667e-09, -1.268394e-09, -1.391266e-09, -1.5203e-09, 
    -1.661159e-09, -1.817681e-09, -1.978366e-09, -2.149154e-09, -2.473472e-09,
  -6.345698e-10, -6.731987e-10, -7.171626e-10, -7.644818e-10, -8.106515e-10, 
    -8.659277e-10, -9.430656e-10, -1.02358e-09, -1.124288e-09, -1.228233e-09, 
    -1.32471e-09, -1.416999e-09, -1.503517e-09, -1.619188e-09, -1.757903e-09,
  -1.254191e-08, -1.327265e-08, -1.393184e-08, -1.448046e-08, -1.498423e-08, 
    -1.530778e-08, -1.547177e-08, -1.555678e-08, -1.54681e-08, -1.532239e-08, 
    -1.525107e-08, -1.530246e-08, -1.54087e-08, -1.556451e-08, -1.568958e-08,
  -1.018428e-08, -1.102888e-08, -1.185374e-08, -1.258774e-08, -1.332252e-08, 
    -1.404047e-08, -1.466384e-08, -1.514079e-08, -1.564078e-08, 
    -1.600464e-08, -1.617403e-08, -1.616077e-08, -1.608093e-08, 
    -1.594293e-08, -1.57861e-08,
  -7.210741e-09, -7.930744e-09, -8.895655e-09, -9.874102e-09, -1.077367e-08, 
    -1.166951e-08, -1.258856e-08, -1.340052e-08, -1.414466e-08, 
    -1.480321e-08, -1.537875e-08, -1.584097e-08, -1.614313e-08, 
    -1.629369e-08, -1.631288e-08,
  -4.704692e-09, -5.193658e-09, -5.731035e-09, -6.48316e-09, -7.356013e-09, 
    -8.316221e-09, -9.365048e-09, -1.034481e-08, -1.135191e-08, 
    -1.226172e-08, -1.308249e-08, -1.377862e-08, -1.441026e-08, 
    -1.492717e-08, -1.532647e-08,
  -2.759468e-09, -2.979745e-09, -3.264882e-09, -3.651153e-09, -4.183307e-09, 
    -4.817561e-09, -5.6667e-09, -6.636433e-09, -7.677988e-09, -8.704872e-09, 
    -9.65711e-09, -1.050079e-08, -1.130292e-08, -1.202604e-08, -1.267657e-08,
  -1.889594e-09, -1.972165e-09, -2.043693e-09, -2.148436e-09, -2.311877e-09, 
    -2.56247e-09, -2.94255e-09, -3.455579e-09, -4.067108e-09, -4.913929e-09, 
    -5.841865e-09, -6.822009e-09, -7.734957e-09, -8.639252e-09, -9.490187e-09,
  -1.140222e-09, -1.228731e-09, -1.311089e-09, -1.400619e-09, -1.447916e-09, 
    -1.516852e-09, -1.660497e-09, -1.873673e-09, -2.148378e-09, 
    -2.459604e-09, -2.832421e-09, -3.344382e-09, -4.056343e-09, 
    -4.926913e-09, -5.881994e-09,
  -4.854013e-10, -5.629172e-10, -6.407381e-10, -7.441001e-10, -8.225854e-10, 
    -8.89489e-10, -9.711741e-10, -1.078681e-09, -1.228588e-09, -1.418941e-09, 
    -1.647589e-09, -1.878032e-09, -2.135238e-09, -2.494816e-09, -3.011846e-09,
  -2.172487e-10, -2.716831e-10, -3.363526e-10, -4.12347e-10, -4.807354e-10, 
    -5.4454e-10, -5.966792e-10, -6.571635e-10, -7.336568e-10, -8.202466e-10, 
    -9.279969e-10, -1.090635e-09, -1.300806e-09, -1.51656e-09, -1.769898e-09,
  -1.395069e-10, -1.297915e-10, -1.564943e-10, -1.688889e-10, -2.019651e-10, 
    -2.824668e-10, -3.806971e-10, -4.709364e-10, -5.450657e-10, 
    -6.212698e-10, -6.86979e-10, -7.56025e-10, -8.390122e-10, -9.408178e-10, 
    -1.089088e-09,
  -7.068944e-09, -7.372901e-09, -7.705752e-09, -8.064488e-09, -8.352423e-09, 
    -8.774793e-09, -9.232502e-09, -9.66414e-09, -1.015948e-08, -1.05583e-08, 
    -1.108072e-08, -1.161162e-08, -1.205082e-08, -1.251598e-08, -1.303415e-08,
  -6.830619e-09, -7.245559e-09, -7.578532e-09, -7.9422e-09, -8.203946e-09, 
    -8.510626e-09, -8.89907e-09, -9.279499e-09, -9.656165e-09, -1.00829e-08, 
    -1.055206e-08, -1.106908e-08, -1.157788e-08, -1.206926e-08, -1.264023e-08,
  -6.411981e-09, -6.919965e-09, -7.284469e-09, -7.642783e-09, -7.976102e-09, 
    -8.230615e-09, -8.605321e-09, -9.008272e-09, -9.401865e-09, 
    -9.749895e-09, -1.010993e-08, -1.041226e-08, -1.083838e-08, 
    -1.136465e-08, -1.199209e-08,
  -5.971186e-09, -6.432115e-09, -6.910285e-09, -7.344357e-09, -7.810292e-09, 
    -8.08523e-09, -8.319634e-09, -8.668866e-09, -9.119862e-09, -9.581924e-09, 
    -9.97946e-09, -1.036221e-08, -1.069452e-08, -1.101957e-08, -1.143572e-08,
  -5.501538e-09, -5.863253e-09, -6.332248e-09, -6.736073e-09, -7.235862e-09, 
    -7.625904e-09, -7.883396e-09, -8.011154e-09, -8.259777e-09, 
    -8.723713e-09, -9.358468e-09, -9.924841e-09, -1.046492e-08, 
    -1.083812e-08, -1.116006e-08,
  -5.190819e-09, -5.493699e-09, -5.847295e-09, -6.149259e-09, -6.504216e-09, 
    -6.874437e-09, -7.217514e-09, -7.498792e-09, -7.596118e-09, 
    -7.813834e-09, -8.229549e-09, -8.90647e-09, -9.56027e-09, -1.019748e-08, 
    -1.070364e-08,
  -4.910997e-09, -5.117267e-09, -5.326952e-09, -5.579824e-09, -5.916748e-09, 
    -6.19095e-09, -6.584755e-09, -6.720829e-09, -7.118377e-09, -7.298259e-09, 
    -7.428492e-09, -7.804465e-09, -8.457689e-09, -9.215657e-09, -9.81823e-09,
  -4.217581e-09, -4.34967e-09, -4.441873e-09, -4.557484e-09, -4.710576e-09, 
    -4.845151e-09, -5.035784e-09, -5.565516e-09, -6.060589e-09, -6.35458e-09, 
    -6.596005e-09, -6.717912e-09, -6.936826e-09, -7.465525e-09, -8.101308e-09,
  -3.401747e-09, -3.500917e-09, -3.552355e-09, -3.63076e-09, -3.625708e-09, 
    -3.716239e-09, -3.952204e-09, -4.303107e-09, -4.553232e-09, 
    -4.913954e-09, -5.295656e-09, -5.527445e-09, -5.48624e-09, -5.519709e-09, 
    -5.900887e-09,
  -2.431888e-09, -2.603461e-09, -2.692702e-09, -2.689589e-09, -2.517191e-09, 
    -2.500012e-09, -2.789903e-09, -3.062236e-09, -3.128166e-09, 
    -3.301871e-09, -3.612632e-09, -3.857844e-09, -3.908184e-09, 
    -3.859765e-09, -3.982735e-09,
  -2.889922e-09, -2.862837e-09, -2.812885e-09, -2.775172e-09, -2.697052e-09, 
    -2.657667e-09, -2.557283e-09, -2.517916e-09, -2.482448e-09, 
    -2.521419e-09, -2.575866e-09, -2.620876e-09, -2.697861e-09, 
    -2.844475e-09, -3.124936e-09,
  -2.556767e-09, -2.553689e-09, -2.566662e-09, -2.522725e-09, -2.483448e-09, 
    -2.443838e-09, -2.415026e-09, -2.352266e-09, -2.383111e-09, 
    -2.404073e-09, -2.493249e-09, -2.586076e-09, -2.67413e-09, -2.772993e-09, 
    -2.910773e-09,
  -2.446822e-09, -2.429572e-09, -2.433361e-09, -2.444174e-09, -2.397681e-09, 
    -2.297156e-09, -2.231894e-09, -2.216232e-09, -2.262971e-09, 
    -2.348339e-09, -2.392213e-09, -2.465788e-09, -2.543876e-09, 
    -2.639758e-09, -2.783888e-09,
  -2.482667e-09, -2.407583e-09, -2.37274e-09, -2.380955e-09, -2.440209e-09, 
    -2.525871e-09, -2.471744e-09, -2.355096e-09, -2.318753e-09, 
    -2.408565e-09, -2.530777e-09, -2.614576e-09, -2.697508e-09, 
    -2.765173e-09, -2.776469e-09,
  -2.817544e-09, -2.672428e-09, -2.565297e-09, -2.493723e-09, -2.486944e-09, 
    -2.573899e-09, -2.735609e-09, -2.858736e-09, -2.845475e-09, 
    -2.784835e-09, -2.707411e-09, -2.741338e-09, -2.929018e-09, 
    -3.123913e-09, -3.272236e-09,
  -3.270472e-09, -3.253171e-09, -3.107268e-09, -2.957991e-09, -2.81479e-09, 
    -2.779542e-09, -2.878902e-09, -3.086639e-09, -3.256801e-09, 
    -3.401672e-09, -3.381857e-09, -3.159555e-09, -3.141424e-09, 
    -3.302424e-09, -3.558016e-09,
  -3.455834e-09, -3.666696e-09, -3.741667e-09, -3.719499e-09, -3.619827e-09, 
    -3.472321e-09, -3.320668e-09, -3.382811e-09, -3.620158e-09, -3.84761e-09, 
    -4.062087e-09, -4.102374e-09, -3.973208e-09, -3.743239e-09, -3.822403e-09,
  -3.135418e-09, -3.552399e-09, -3.960888e-09, -4.215598e-09, -4.2545e-09, 
    -4.170647e-09, -4.092128e-09, -3.951878e-09, -3.897211e-09, 
    -4.067516e-09, -4.410148e-09, -4.640768e-09, -4.736915e-09, 
    -4.799957e-09, -4.639733e-09,
  -2.739152e-09, -3.077689e-09, -3.586313e-09, -4.077407e-09, -4.405438e-09, 
    -4.527175e-09, -4.706844e-09, -4.596542e-09, -4.536748e-09, 
    -4.622791e-09, -4.637238e-09, -4.797871e-09, -5.081922e-09, 
    -5.360405e-09, -5.522395e-09,
  -2.5059e-09, -2.674414e-09, -2.969875e-09, -3.345355e-09, -3.765706e-09, 
    -4.130433e-09, -4.6275e-09, -5.16537e-09, -5.240764e-09, -5.136101e-09, 
    -4.999551e-09, -5.146951e-09, -5.379665e-09, -5.506065e-09, -5.691816e-09,
  -2.590589e-09, -2.639684e-09, -2.716708e-09, -2.837155e-09, -2.951688e-09, 
    -3.091567e-09, -3.290853e-09, -3.543791e-09, -3.829739e-09, 
    -4.116928e-09, -4.406245e-09, -4.723468e-09, -5.064518e-09, 
    -5.412693e-09, -5.744618e-09,
  -1.6297e-09, -1.670967e-09, -1.763833e-09, -1.903129e-09, -2.047682e-09, 
    -2.234892e-09, -2.426682e-09, -2.612336e-09, -2.795894e-09, 
    -2.969044e-09, -3.139581e-09, -3.340062e-09, -3.577536e-09, 
    -3.866755e-09, -4.195053e-09,
  -1.217502e-09, -1.245423e-09, -1.3463e-09, -1.484055e-09, -1.64866e-09, 
    -1.817129e-09, -1.979188e-09, -2.146435e-09, -2.285967e-09, 
    -2.411898e-09, -2.527208e-09, -2.65604e-09, -2.811118e-09, -2.994648e-09, 
    -3.201938e-09,
  -9.238886e-10, -9.529824e-10, -1.030163e-09, -1.167355e-09, -1.333415e-09, 
    -1.481017e-09, -1.632315e-09, -1.785218e-09, -1.923344e-09, 
    -2.046032e-09, -2.165675e-09, -2.292623e-09, -2.428917e-09, 
    -2.556897e-09, -2.690941e-09,
  -7.721261e-10, -8.080847e-10, -8.75174e-10, -9.887972e-10, -1.11517e-09, 
    -1.234522e-09, -1.356331e-09, -1.487413e-09, -1.615887e-09, 
    -1.744386e-09, -1.875724e-09, -2.028294e-09, -2.181396e-09, 
    -2.320271e-09, -2.424593e-09,
  -6.730229e-10, -6.971473e-10, -7.434166e-10, -8.235684e-10, -9.304621e-10, 
    -1.0291e-09, -1.1303e-09, -1.238002e-09, -1.357664e-09, -1.484185e-09, 
    -1.620032e-09, -1.790232e-09, -1.959106e-09, -2.102113e-09, -2.209352e-09,
  -6.536194e-10, -6.653294e-10, -6.883233e-10, -7.285479e-10, -8.000191e-10, 
    -8.854492e-10, -9.534417e-10, -1.03675e-09, -1.140167e-09, -1.254081e-09, 
    -1.396295e-09, -1.58322e-09, -1.770474e-09, -1.91389e-09, -2.02105e-09,
  -6.914971e-10, -6.821438e-10, -6.887018e-10, -6.985653e-10, -7.314414e-10, 
    -7.812072e-10, -8.444133e-10, -9.124121e-10, -1.000596e-09, -1.0925e-09, 
    -1.224178e-09, -1.426935e-09, -1.641094e-09, -1.80352e-09, -1.903234e-09,
  -7.096515e-10, -6.808403e-10, -6.736628e-10, -6.630589e-10, -6.74524e-10, 
    -7.047023e-10, -7.562551e-10, -8.302341e-10, -9.050566e-10, 
    -9.880906e-10, -1.087959e-09, -1.263007e-09, -1.516356e-09, 
    -1.742735e-09, -1.93259e-09,
  -6.934874e-10, -6.806634e-10, -6.532561e-10, -6.467559e-10, -6.317047e-10, 
    -6.568038e-10, -7.115195e-10, -7.821065e-10, -8.639605e-10, 
    -9.515231e-10, -1.065184e-09, -1.221433e-09, -1.436868e-09, 
    -1.722395e-09, -1.949997e-09,
  -1.482696e-08, -1.592575e-08, -1.712942e-08, -1.806014e-08, -1.861557e-08, 
    -1.905217e-08, -1.929822e-08, -1.911137e-08, -1.87135e-08, -1.818405e-08, 
    -1.769866e-08, -1.709427e-08, -1.655893e-08, -1.596512e-08, -1.537482e-08,
  -1.197691e-08, -1.307617e-08, -1.400162e-08, -1.494989e-08, -1.557843e-08, 
    -1.595814e-08, -1.614328e-08, -1.609731e-08, -1.584307e-08, 
    -1.549947e-08, -1.504219e-08, -1.451555e-08, -1.392746e-08, 
    -1.327596e-08, -1.267497e-08,
  -9.28912e-09, -1.003375e-08, -1.080004e-08, -1.153699e-08, -1.213191e-08, 
    -1.251414e-08, -1.275193e-08, -1.280125e-08, -1.271034e-08, 
    -1.252535e-08, -1.222193e-08, -1.181065e-08, -1.125859e-08, 
    -1.075494e-08, -1.028647e-08,
  -6.940414e-09, -7.441594e-09, -7.965635e-09, -8.436534e-09, -8.827684e-09, 
    -9.153423e-09, -9.337946e-09, -9.432514e-09, -9.380374e-09, 
    -9.256694e-09, -9.030193e-09, -8.713879e-09, -8.395122e-09, -8.05929e-09, 
    -7.708953e-09,
  -5.196201e-09, -5.708352e-09, -6.128467e-09, -6.463546e-09, -6.678698e-09, 
    -6.825162e-09, -6.888477e-09, -6.88878e-09, -6.822993e-09, -6.712908e-09, 
    -6.556635e-09, -6.39522e-09, -6.210672e-09, -5.99759e-09, -5.704428e-09,
  -3.899116e-09, -4.232938e-09, -4.546907e-09, -4.833762e-09, -5.048754e-09, 
    -5.195953e-09, -5.252017e-09, -5.237983e-09, -5.163169e-09, 
    -5.054439e-09, -4.918526e-09, -4.735985e-09, -4.519744e-09, 
    -4.253772e-09, -3.97557e-09,
  -3.320961e-09, -3.476245e-09, -3.612824e-09, -3.772748e-09, -3.902179e-09, 
    -4.014024e-09, -4.04881e-09, -4.032076e-09, -3.950776e-09, -3.853798e-09, 
    -3.718094e-09, -3.546531e-09, -3.313079e-09, -3.036696e-09, -2.81789e-09,
  -2.484238e-09, -2.68869e-09, -2.860131e-09, -2.985242e-09, -3.049943e-09, 
    -3.087267e-09, -3.086503e-09, -3.027202e-09, -2.977461e-09, 
    -2.902517e-09, -2.802771e-09, -2.658916e-09, -2.490395e-09, 
    -2.336081e-09, -2.193894e-09,
  -1.51041e-09, -1.758376e-09, -2.000298e-09, -2.206214e-09, -2.315709e-09, 
    -2.351871e-09, -2.380246e-09, -2.34683e-09, -2.293781e-09, -2.235834e-09, 
    -2.153178e-09, -2.074851e-09, -2.006636e-09, -1.941412e-09, -1.885534e-09,
  -1.050814e-09, -1.145969e-09, -1.278596e-09, -1.442939e-09, -1.541047e-09, 
    -1.628135e-09, -1.754952e-09, -1.817975e-09, -1.778165e-09, 
    -1.774348e-09, -1.73117e-09, -1.700976e-09, -1.674556e-09, -1.633898e-09, 
    -1.577269e-09,
  -9.032441e-09, -1.130996e-08, -1.442825e-08, -1.769959e-08, -2.019886e-08, 
    -2.286403e-08, -2.466279e-08, -2.554581e-08, -2.548719e-08, 
    -2.524491e-08, -2.508678e-08, -2.530101e-08, -2.545418e-08, 
    -2.554827e-08, -2.554894e-08,
  -7.291619e-09, -8.96114e-09, -1.125356e-08, -1.429745e-08, -1.73098e-08, 
    -1.995687e-08, -2.236387e-08, -2.405378e-08, -2.497746e-08, -2.50696e-08, 
    -2.461429e-08, -2.436027e-08, -2.447333e-08, -2.461845e-08, -2.462529e-08,
  -5.671587e-09, -6.93232e-09, -8.523227e-09, -1.079967e-08, -1.364561e-08, 
    -1.678208e-08, -1.957268e-08, -2.170191e-08, -2.32636e-08, -2.406233e-08, 
    -2.429904e-08, -2.411659e-08, -2.397818e-08, -2.385106e-08, -2.361191e-08,
  -4.910684e-09, -5.592881e-09, -6.639271e-09, -8.094803e-09, -1.011267e-08, 
    -1.267658e-08, -1.557062e-08, -1.824089e-08, -2.004322e-08, 
    -2.132335e-08, -2.201607e-08, -2.219906e-08, -2.217045e-08, 
    -2.189228e-08, -2.143649e-08,
  -5.088927e-09, -4.842495e-09, -5.276361e-09, -6.160686e-09, -7.44877e-09, 
    -9.294456e-09, -1.159787e-08, -1.423795e-08, -1.668931e-08, 
    -1.819801e-08, -1.911908e-08, -1.948863e-08, -1.959817e-08, 
    -1.938983e-08, -1.896845e-08,
  -7.196626e-09, -5.600598e-09, -4.823348e-09, -4.912801e-09, -5.498541e-09, 
    -6.387438e-09, -7.807644e-09, -9.719962e-09, -1.199319e-08, 
    -1.416133e-08, -1.569065e-08, -1.64015e-08, -1.663511e-08, -1.649878e-08, 
    -1.616142e-08,
  -8.443983e-09, -8.024771e-09, -6.8229e-09, -5.360812e-09, -4.888228e-09, 
    -5.157315e-09, -5.661855e-09, -6.455414e-09, -7.712802e-09, 
    -9.330561e-09, -1.112283e-08, -1.245653e-08, -1.327207e-08, 
    -1.342242e-08, -1.302626e-08,
  -7.031592e-09, -7.928551e-09, -8.19077e-09, -7.757151e-09, -6.577235e-09, 
    -5.451438e-09, -5.059801e-09, -5.306261e-09, -5.767931e-09, 
    -6.398682e-09, -7.135605e-09, -8.102782e-09, -8.732132e-09, 
    -9.090624e-09, -8.907839e-09,
  -4.161766e-09, -5.445466e-09, -6.732835e-09, -7.483523e-09, -7.595649e-09, 
    -7.40773e-09, -6.586981e-09, -5.748713e-09, -5.29642e-09, -5.359278e-09, 
    -5.545477e-09, -5.743853e-09, -5.85619e-09, -5.870517e-09, -5.807952e-09,
  -2.789029e-09, -3.10524e-09, -3.793631e-09, -4.870857e-09, -6.016771e-09, 
    -6.539912e-09, -6.925759e-09, -6.981814e-09, -6.659442e-09, 
    -6.165299e-09, -5.737173e-09, -5.468552e-09, -5.324804e-09, 
    -5.258901e-09, -5.229602e-09,
  -5.200595e-09, -5.883766e-09, -7.038942e-09, -8.573137e-09, -1.06313e-08, 
    -1.361109e-08, -1.687994e-08, -1.973554e-08, -2.174236e-08, 
    -2.414174e-08, -2.567581e-08, -2.63338e-08, -2.64977e-08, -2.653259e-08, 
    -2.680576e-08,
  -4.131553e-09, -4.540464e-09, -5.166479e-09, -6.132133e-09, -7.419156e-09, 
    -9.383041e-09, -1.25001e-08, -1.60045e-08, -1.913199e-08, -2.154596e-08, 
    -2.368666e-08, -2.47946e-08, -2.551743e-08, -2.633715e-08, -2.687956e-08,
  -3.782636e-09, -3.893077e-09, -4.151032e-09, -4.62026e-09, -5.404646e-09, 
    -6.520673e-09, -8.409015e-09, -1.138015e-08, -1.489151e-08, 
    -1.829766e-08, -2.119902e-08, -2.322814e-08, -2.437686e-08, 
    -2.519629e-08, -2.605006e-08,
  -3.846092e-09, -3.738306e-09, -3.747799e-09, -3.873136e-09, -4.200777e-09, 
    -4.790617e-09, -5.79985e-09, -7.538313e-09, -1.024748e-08, -1.367704e-08, 
    -1.716509e-08, -2.028302e-08, -2.244581e-08, -2.382569e-08, -2.486704e-08,
  -3.967441e-09, -3.876472e-09, -3.775686e-09, -3.720696e-09, -3.736228e-09, 
    -3.881595e-09, -4.308019e-09, -5.130973e-09, -6.596022e-09, -8.99905e-09, 
    -1.223796e-08, -1.582352e-08, -1.921687e-08, -2.160654e-08, -2.327116e-08,
  -4.126792e-09, -3.963192e-09, -3.854327e-09, -3.792187e-09, -3.791305e-09, 
    -3.777091e-09, -3.848994e-09, -4.114591e-09, -4.726113e-09, 
    -5.846176e-09, -7.722504e-09, -1.03862e-08, -1.377741e-08, -1.723512e-08, 
    -2.026152e-08,
  -4.845535e-09, -4.413913e-09, -4.050325e-09, -3.738094e-09, -3.641266e-09, 
    -3.689728e-09, -3.746706e-09, -3.854473e-09, -4.056295e-09, 
    -4.532983e-09, -5.394964e-09, -6.767203e-09, -8.734655e-09, 
    -1.134094e-08, -1.428992e-08,
  -5.621583e-09, -5.580297e-09, -5.221604e-09, -4.648532e-09, -3.957201e-09, 
    -3.616457e-09, -3.541414e-09, -3.607891e-09, -3.727565e-09, 
    -3.900589e-09, -4.263939e-09, -4.872313e-09, -5.8779e-09, -7.286223e-09, 
    -9.069547e-09,
  -5.650084e-09, -5.785097e-09, -5.938711e-09, -5.95723e-09, -5.686162e-09, 
    -4.974178e-09, -4.17994e-09, -3.666909e-09, -3.536025e-09, -3.552419e-09, 
    -3.694467e-09, -3.881233e-09, -4.252095e-09, -4.745912e-09, -5.502711e-09,
  -5.443852e-09, -5.638318e-09, -5.781173e-09, -5.909737e-09, -6.03768e-09, 
    -6.148992e-09, -6.096154e-09, -5.647558e-09, -4.847105e-09, 
    -4.193326e-09, -3.801186e-09, -3.679255e-09, -3.742123e-09, 
    -3.842116e-09, -4.023274e-09,
  -1.432762e-08, -1.576293e-08, -1.692976e-08, -1.840192e-08, -1.970139e-08, 
    -2.075918e-08, -2.13286e-08, -2.175897e-08, -2.188935e-08, -2.213908e-08, 
    -2.204808e-08, -2.189106e-08, -2.166575e-08, -2.160728e-08, -2.164299e-08,
  -1.071705e-08, -1.255007e-08, -1.41659e-08, -1.54156e-08, -1.661192e-08, 
    -1.795766e-08, -1.903175e-08, -2.005602e-08, -2.068658e-08, 
    -2.120954e-08, -2.15538e-08, -2.188437e-08, -2.197778e-08, -2.193494e-08, 
    -2.190226e-08,
  -7.571162e-09, -8.847599e-09, -1.04987e-08, -1.22588e-08, -1.383469e-08, 
    -1.517144e-08, -1.63642e-08, -1.756577e-08, -1.859295e-08, -1.954052e-08, 
    -2.028882e-08, -2.081443e-08, -2.130421e-08, -2.169294e-08, -2.197585e-08,
  -6.207772e-09, -6.661852e-09, -7.549146e-09, -8.728886e-09, -1.017277e-08, 
    -1.178482e-08, -1.328523e-08, -1.462697e-08, -1.588193e-08, -1.6949e-08, 
    -1.801727e-08, -1.895705e-08, -1.984755e-08, -2.05523e-08, -2.114281e-08,
  -5.362099e-09, -5.674649e-09, -6.005683e-09, -6.548246e-09, -7.358282e-09, 
    -8.396752e-09, -9.673829e-09, -1.106323e-08, -1.248245e-08, 
    -1.378044e-08, -1.502499e-08, -1.613174e-08, -1.717444e-08, 
    -1.826913e-08, -1.922623e-08,
  -4.853205e-09, -5.008057e-09, -5.247026e-09, -5.519831e-09, -5.87232e-09, 
    -6.371551e-09, -7.0587e-09, -7.955228e-09, -9.00833e-09, -1.017334e-08, 
    -1.140076e-08, -1.263069e-08, -1.384483e-08, -1.497052e-08, -1.615224e-08,
  -4.586135e-09, -4.657246e-09, -4.736598e-09, -4.91489e-09, -5.114848e-09, 
    -5.37049e-09, -5.690795e-09, -6.107516e-09, -6.681406e-09, -7.399117e-09, 
    -8.222686e-09, -9.132015e-09, -1.014195e-08, -1.120277e-08, -1.233414e-08,
  -4.317433e-09, -4.492412e-09, -4.565816e-09, -4.675018e-09, -4.749807e-09, 
    -4.832696e-09, -5.003913e-09, -5.216506e-09, -5.478342e-09, 
    -5.808068e-09, -6.248232e-09, -6.790382e-09, -7.392312e-09, 
    -8.051677e-09, -8.777915e-09,
  -3.939588e-09, -4.087258e-09, -4.284309e-09, -4.470808e-09, -4.617014e-09, 
    -4.686445e-09, -4.732303e-09, -4.774597e-09, -4.863437e-09, 
    -5.014605e-09, -5.194615e-09, -5.45056e-09, -5.753502e-09, -6.121526e-09, 
    -6.505405e-09,
  -3.617425e-09, -3.791433e-09, -3.954146e-09, -4.16419e-09, -4.337157e-09, 
    -4.489119e-09, -4.633415e-09, -4.714537e-09, -4.735742e-09, 
    -4.747644e-09, -4.787026e-09, -4.848399e-09, -4.955353e-09, 
    -5.104074e-09, -5.283457e-09,
  -1.648675e-08, -1.712975e-08, -1.783538e-08, -1.86931e-08, -1.948984e-08, 
    -2.036599e-08, -2.091784e-08, -2.113478e-08, -2.160845e-08, 
    -2.190551e-08, -2.205762e-08, -2.191949e-08, -2.16814e-08, -2.169715e-08, 
    -2.15159e-08,
  -1.48258e-08, -1.560078e-08, -1.631681e-08, -1.708288e-08, -1.789718e-08, 
    -1.883611e-08, -1.988825e-08, -2.061188e-08, -2.110167e-08, -2.17262e-08, 
    -2.204867e-08, -2.251206e-08, -2.218539e-08, -2.199016e-08, -2.165949e-08,
  -1.326362e-08, -1.387342e-08, -1.463646e-08, -1.53983e-08, -1.632511e-08, 
    -1.717734e-08, -1.816369e-08, -1.918623e-08, -1.996621e-08, 
    -2.075333e-08, -2.14325e-08, -2.212832e-08, -2.251353e-08, -2.250237e-08, 
    -2.234373e-08,
  -1.192379e-08, -1.24734e-08, -1.305178e-08, -1.370064e-08, -1.450421e-08, 
    -1.540654e-08, -1.62993e-08, -1.728693e-08, -1.828527e-08, -1.926983e-08, 
    -2.01168e-08, -2.101044e-08, -2.174101e-08, -2.225901e-08, -2.248068e-08,
  -1.054995e-08, -1.108854e-08, -1.1579e-08, -1.215946e-08, -1.280993e-08, 
    -1.354396e-08, -1.439628e-08, -1.536044e-08, -1.626891e-08, 
    -1.727531e-08, -1.833167e-08, -1.932815e-08, -2.031993e-08, 
    -2.104749e-08, -2.167441e-08,
  -9.32492e-09, -9.742717e-09, -1.025913e-08, -1.076292e-08, -1.134457e-08, 
    -1.191565e-08, -1.258029e-08, -1.335896e-08, -1.42148e-08, -1.513675e-08, 
    -1.609939e-08, -1.715954e-08, -1.823921e-08, -1.932602e-08, -2.021159e-08,
  -7.94051e-09, -8.421975e-09, -8.925734e-09, -9.479987e-09, -1.002613e-08, 
    -1.05718e-08, -1.116988e-08, -1.175144e-08, -1.241149e-08, -1.316854e-08, 
    -1.398962e-08, -1.490771e-08, -1.58459e-08, -1.690433e-08, -1.797407e-08,
  -6.727933e-09, -7.149653e-09, -7.626264e-09, -8.018056e-09, -8.488358e-09, 
    -9.04667e-09, -9.62227e-09, -1.021594e-08, -1.083017e-08, -1.149278e-08, 
    -1.216459e-08, -1.290092e-08, -1.367994e-08, -1.454262e-08, -1.543448e-08,
  -5.978295e-09, -6.137665e-09, -6.416797e-09, -6.770186e-09, -7.116348e-09, 
    -7.507503e-09, -8.061672e-09, -8.590668e-09, -9.158803e-09, 
    -9.790351e-09, -1.045169e-08, -1.110149e-08, -1.179265e-08, 
    -1.249954e-08, -1.325882e-08,
  -5.278161e-09, -5.410768e-09, -5.510341e-09, -5.665374e-09, -5.841886e-09, 
    -6.075844e-09, -6.654143e-09, -7.127094e-09, -7.528453e-09, 
    -8.021434e-09, -8.584245e-09, -9.213008e-09, -9.874745e-09, 
    -1.052629e-08, -1.120822e-08,
  -1.663204e-08, -1.72749e-08, -1.788571e-08, -1.838988e-08, -1.865174e-08, 
    -1.876473e-08, -1.880369e-08, -1.861419e-08, -1.841733e-08, 
    -1.845845e-08, -1.861565e-08, -1.887626e-08, -1.920355e-08, 
    -1.950118e-08, -1.970534e-08,
  -1.48533e-08, -1.611158e-08, -1.688073e-08, -1.755392e-08, -1.806092e-08, 
    -1.844004e-08, -1.855948e-08, -1.855603e-08, -1.841337e-08, 
    -1.835689e-08, -1.836428e-08, -1.858557e-08, -1.893097e-08, 
    -1.925921e-08, -1.956415e-08,
  -1.270671e-08, -1.41711e-08, -1.557316e-08, -1.644255e-08, -1.715074e-08, 
    -1.767249e-08, -1.806092e-08, -1.819791e-08, -1.815591e-08, -1.81712e-08, 
    -1.809799e-08, -1.811005e-08, -1.848875e-08, -1.899779e-08, -1.934946e-08,
  -1.13144e-08, -1.238156e-08, -1.363456e-08, -1.497814e-08, -1.596573e-08, 
    -1.671616e-08, -1.720379e-08, -1.76402e-08, -1.778538e-08, -1.782547e-08, 
    -1.780765e-08, -1.770779e-08, -1.792764e-08, -1.845274e-08, -1.901194e-08,
  -1.005983e-08, -1.10534e-08, -1.200635e-08, -1.314314e-08, -1.438935e-08, 
    -1.548134e-08, -1.619786e-08, -1.678679e-08, -1.722015e-08, 
    -1.742068e-08, -1.758584e-08, -1.751317e-08, -1.758489e-08, 
    -1.788008e-08, -1.84148e-08,
  -9.026992e-09, -9.891941e-09, -1.070725e-08, -1.156313e-08, -1.264143e-08, 
    -1.382546e-08, -1.492994e-08, -1.563178e-08, -1.617211e-08, -1.64929e-08, 
    -1.67272e-08, -1.692801e-08, -1.710385e-08, -1.734512e-08, -1.77825e-08,
  -8.126352e-09, -8.928793e-09, -9.605617e-09, -1.034982e-08, -1.113531e-08, 
    -1.213858e-08, -1.328589e-08, -1.43036e-08, -1.507682e-08, -1.558644e-08, 
    -1.591881e-08, -1.619401e-08, -1.634067e-08, -1.649323e-08, -1.676435e-08,
  -6.927553e-09, -7.840744e-09, -8.592475e-09, -9.28294e-09, -1.001409e-08, 
    -1.073997e-08, -1.164306e-08, -1.271925e-08, -1.369968e-08, 
    -1.451874e-08, -1.508034e-08, -1.543135e-08, -1.560344e-08, -1.57174e-08, 
    -1.585294e-08,
  -5.957077e-09, -6.581842e-09, -7.393908e-09, -8.205131e-09, -8.964405e-09, 
    -9.649725e-09, -1.031411e-08, -1.108162e-08, -1.19952e-08, -1.288425e-08, 
    -1.374541e-08, -1.434979e-08, -1.474946e-08, -1.497735e-08, -1.510177e-08,
  -5.145341e-09, -5.710532e-09, -6.256672e-09, -6.978095e-09, -7.771957e-09, 
    -8.567556e-09, -9.239298e-09, -9.900339e-09, -1.062428e-08, 
    -1.135331e-08, -1.213392e-08, -1.286607e-08, -1.342995e-08, 
    -1.390652e-08, -1.415768e-08,
  -9.482736e-09, -1.038551e-08, -1.148874e-08, -1.270654e-08, -1.398389e-08, 
    -1.531306e-08, -1.647886e-08, -1.753534e-08, -1.827639e-08, 
    -1.877831e-08, -1.910941e-08, -1.935901e-08, -1.959522e-08, 
    -1.977135e-08, -1.987754e-08,
  -7.162122e-09, -8.025439e-09, -8.999879e-09, -1.001576e-08, -1.115685e-08, 
    -1.245823e-08, -1.380008e-08, -1.518504e-08, -1.648116e-08, 
    -1.745821e-08, -1.810346e-08, -1.855987e-08, -1.891364e-08, 
    -1.919146e-08, -1.935105e-08,
  -5.754677e-09, -6.336938e-09, -7.09749e-09, -7.97207e-09, -8.904466e-09, 
    -9.987367e-09, -1.114328e-08, -1.243191e-08, -1.376209e-08, 
    -1.511246e-08, -1.633834e-08, -1.72523e-08, -1.783053e-08, -1.830147e-08, 
    -1.86006e-08,
  -4.777314e-09, -5.180497e-09, -5.70558e-09, -6.400682e-09, -7.22741e-09, 
    -8.148104e-09, -9.12289e-09, -1.01431e-08, -1.142136e-08, -1.272872e-08, 
    -1.410169e-08, -1.541428e-08, -1.652686e-08, -1.730269e-08, -1.775258e-08,
  -4.119658e-09, -4.40718e-09, -4.758157e-09, -5.231942e-09, -5.882256e-09, 
    -6.703762e-09, -7.603772e-09, -8.417924e-09, -9.417118e-09, 
    -1.063392e-08, -1.194996e-08, -1.334722e-08, -1.464676e-08, 
    -1.589299e-08, -1.680007e-08,
  -3.648492e-09, -3.893431e-09, -4.127166e-09, -4.395033e-09, -4.838448e-09, 
    -5.460199e-09, -6.346665e-09, -7.310029e-09, -8.204312e-09, 
    -9.171495e-09, -1.025646e-08, -1.15234e-08, -1.287058e-08, -1.415186e-08, 
    -1.539715e-08,
  -3.196005e-09, -3.480149e-09, -3.690356e-09, -3.869203e-09, -4.127144e-09, 
    -4.548144e-09, -5.107337e-09, -5.941405e-09, -6.970792e-09, 
    -7.989789e-09, -9.00573e-09, -1.004819e-08, -1.128669e-08, -1.255707e-08, 
    -1.375847e-08,
  -2.567594e-09, -2.876809e-09, -3.194564e-09, -3.468206e-09, -3.734962e-09, 
    -4.077945e-09, -4.473257e-09, -5.007356e-09, -5.82256e-09, -6.803695e-09, 
    -7.882659e-09, -8.907641e-09, -9.985978e-09, -1.11794e-08, -1.23966e-08,
  -2.061713e-09, -2.217319e-09, -2.514688e-09, -2.899839e-09, -3.277617e-09, 
    -3.623909e-09, -3.99294e-09, -4.377849e-09, -4.921024e-09, -5.680568e-09, 
    -6.69818e-09, -7.745309e-09, -8.889029e-09, -9.997177e-09, -1.122449e-08,
  -1.976319e-09, -2.019607e-09, -2.088759e-09, -2.311783e-09, -2.650372e-09, 
    -3.118265e-09, -3.564017e-09, -3.977489e-09, -4.382949e-09, 
    -4.886996e-09, -5.646867e-09, -6.600627e-09, -7.724791e-09, 
    -8.886079e-09, -1.011035e-08,
  -1.077478e-08, -1.200555e-08, -1.343136e-08, -1.493006e-08, -1.64678e-08, 
    -1.79612e-08, -1.928052e-08, -2.047865e-08, -2.155489e-08, -2.245261e-08, 
    -2.307892e-08, -2.347904e-08, -2.386277e-08, -2.416977e-08, -2.436814e-08,
  -8.229468e-09, -9.210409e-09, -1.031326e-08, -1.151582e-08, -1.291148e-08, 
    -1.424203e-08, -1.569588e-08, -1.707585e-08, -1.841081e-08, 
    -1.958635e-08, -2.077419e-08, -2.168931e-08, -2.231462e-08, 
    -2.283098e-08, -2.325862e-08,
  -6.214427e-09, -6.942781e-09, -7.72503e-09, -8.624737e-09, -9.657201e-09, 
    -1.081536e-08, -1.210712e-08, -1.349427e-08, -1.493778e-08, 
    -1.628699e-08, -1.759958e-08, -1.889205e-08, -2.007839e-08, 
    -2.101246e-08, -2.166021e-08,
  -4.940274e-09, -5.45458e-09, -6.006968e-09, -6.626037e-09, -7.354492e-09, 
    -8.207257e-09, -9.191298e-09, -1.02502e-08, -1.135336e-08, -1.255806e-08, 
    -1.383357e-08, -1.512603e-08, -1.637419e-08, -1.76851e-08, -1.891959e-08,
  -4.097578e-09, -4.339963e-09, -4.662929e-09, -5.078116e-09, -5.568149e-09, 
    -6.202612e-09, -6.981689e-09, -7.79038e-09, -8.615826e-09, -9.514494e-09, 
    -1.060857e-08, -1.184922e-08, -1.305811e-08, -1.435177e-08, -1.551499e-08,
  -3.768471e-09, -3.869525e-09, -4.001258e-09, -4.191836e-09, -4.456261e-09, 
    -4.849962e-09, -5.381872e-09, -5.96924e-09, -6.551894e-09, -7.301427e-09, 
    -8.269761e-09, -9.275825e-09, -1.031316e-08, -1.148085e-08, -1.25692e-08,
  -3.58273e-09, -3.613714e-09, -3.643671e-09, -3.657807e-09, -3.733483e-09, 
    -3.944659e-09, -4.249301e-09, -4.677553e-09, -5.128069e-09, 
    -5.577319e-09, -6.213206e-09, -6.982013e-09, -7.861149e-09, 
    -8.884386e-09, -9.972432e-09,
  -3.359475e-09, -3.39707e-09, -3.42567e-09, -3.376867e-09, -3.302373e-09, 
    -3.352195e-09, -3.48645e-09, -3.712676e-09, -4.079923e-09, -4.437714e-09, 
    -4.79547e-09, -5.297583e-09, -5.912399e-09, -6.731633e-09, -7.641481e-09,
  -3.138056e-09, -3.139807e-09, -3.161716e-09, -3.153004e-09, -3.136248e-09, 
    -3.0808e-09, -3.111123e-09, -3.188652e-09, -3.307358e-09, -3.55553e-09, 
    -3.85411e-09, -4.191674e-09, -4.614749e-09, -5.118393e-09, -5.755708e-09,
  -2.910087e-09, -2.970036e-09, -2.964975e-09, -2.922843e-09, -2.847949e-09, 
    -2.860129e-09, -2.928791e-09, -2.986788e-09, -3.030701e-09, 
    -3.127935e-09, -3.249298e-09, -3.442866e-09, -3.735082e-09, -4.13394e-09, 
    -4.582767e-09,
  -1.756156e-08, -1.730707e-08, -1.636306e-08, -1.578095e-08, -1.509639e-08, 
    -1.488418e-08, -1.506253e-08, -1.564395e-08, -1.622335e-08, 
    -1.680063e-08, -1.751573e-08, -1.812641e-08, -1.85552e-08, -1.910153e-08, 
    -1.968981e-08,
  -1.68889e-08, -1.759873e-08, -1.746319e-08, -1.694446e-08, -1.616849e-08, 
    -1.592078e-08, -1.578944e-08, -1.598469e-08, -1.645402e-08, 
    -1.692969e-08, -1.744759e-08, -1.808004e-08, -1.853621e-08, 
    -1.900257e-08, -1.930989e-08,
  -1.55401e-08, -1.61869e-08, -1.664306e-08, -1.684102e-08, -1.673332e-08, 
    -1.628115e-08, -1.624973e-08, -1.649929e-08, -1.688328e-08, 
    -1.732956e-08, -1.772632e-08, -1.813712e-08, -1.850628e-08, 
    -1.890563e-08, -1.920531e-08,
  -1.490863e-08, -1.566459e-08, -1.617462e-08, -1.62573e-08, -1.64076e-08, 
    -1.649134e-08, -1.646248e-08, -1.652527e-08, -1.691998e-08, 
    -1.751435e-08, -1.808495e-08, -1.868242e-08, -1.905003e-08, 
    -1.927937e-08, -1.940254e-08,
  -1.383044e-08, -1.414622e-08, -1.487956e-08, -1.561533e-08, -1.576501e-08, 
    -1.578561e-08, -1.606345e-08, -1.648624e-08, -1.681615e-08, 
    -1.736383e-08, -1.781355e-08, -1.840063e-08, -1.893613e-08, 
    -1.946395e-08, -1.968777e-08,
  -1.201752e-08, -1.327103e-08, -1.380523e-08, -1.439082e-08, -1.498407e-08, 
    -1.536937e-08, -1.553248e-08, -1.579773e-08, -1.630496e-08, 
    -1.697645e-08, -1.769162e-08, -1.834205e-08, -1.890223e-08, 
    -1.936014e-08, -1.985914e-08,
  -8.14785e-09, -1.075605e-08, -1.249463e-08, -1.334873e-08, -1.390407e-08, 
    -1.431922e-08, -1.475511e-08, -1.505479e-08, -1.545455e-08, 
    -1.617416e-08, -1.699505e-08, -1.786371e-08, -1.862485e-08, 
    -1.935027e-08, -2.005609e-08,
  -5.334927e-09, -7.599637e-09, -9.977554e-09, -1.162212e-08, -1.245948e-08, 
    -1.295054e-08, -1.354287e-08, -1.410631e-08, -1.460472e-08, 
    -1.519541e-08, -1.602104e-08, -1.667708e-08, -1.733308e-08, 
    -1.818432e-08, -1.916132e-08,
  -4.34106e-09, -5.257271e-09, -7.166281e-09, -9.148552e-09, -1.057044e-08, 
    -1.129487e-08, -1.198526e-08, -1.270591e-08, -1.33861e-08, -1.387201e-08, 
    -1.403559e-08, -1.461478e-08, -1.556637e-08, -1.637952e-08, -1.695873e-08,
  -4.057974e-09, -4.420608e-09, -5.288941e-09, -6.898296e-09, -8.307699e-09, 
    -9.594377e-09, -1.036859e-08, -1.081031e-08, -1.128993e-08, 
    -1.185185e-08, -1.216471e-08, -1.251452e-08, -1.291478e-08, 
    -1.358174e-08, -1.425914e-08,
  -9.626056e-09, -1.098762e-08, -1.173072e-08, -1.24955e-08, -1.281153e-08, 
    -1.250352e-08, -1.211244e-08, -1.15882e-08, -1.094832e-08, -1.061496e-08, 
    -1.044944e-08, -1.052123e-08, -1.052778e-08, -1.063834e-08, -1.076413e-08,
  -8.778202e-09, -9.981471e-09, -1.10515e-08, -1.181498e-08, -1.22668e-08, 
    -1.236996e-08, -1.198598e-08, -1.155163e-08, -1.099293e-08, -1.05028e-08, 
    -1.006604e-08, -9.913604e-09, -1.001321e-08, -1.026516e-08, -1.044432e-08,
  -8.08343e-09, -8.9556e-09, -1.007874e-08, -1.119893e-08, -1.181372e-08, 
    -1.21027e-08, -1.196991e-08, -1.161875e-08, -1.101132e-08, -1.046733e-08, 
    -9.96209e-09, -9.609235e-09, -9.423142e-09, -9.57143e-09, -9.948103e-09,
  -7.505507e-09, -8.338419e-09, -9.336592e-09, -1.028172e-08, -1.132258e-08, 
    -1.178775e-08, -1.185075e-08, -1.157558e-08, -1.123753e-08, 
    -1.057561e-08, -9.968188e-09, -9.549764e-09, -9.224246e-09, 
    -9.039695e-09, -9.204165e-09,
  -6.821904e-09, -7.750582e-09, -8.799259e-09, -9.895975e-09, -1.075936e-08, 
    -1.161678e-08, -1.185594e-08, -1.159892e-08, -1.126261e-08, 
    -1.096643e-08, -1.032194e-08, -9.681728e-09, -9.296306e-09, 
    -9.004957e-09, -8.828738e-09,
  -5.728101e-09, -7.12381e-09, -8.092867e-09, -9.201407e-09, -1.033124e-08, 
    -1.119312e-08, -1.189083e-08, -1.188016e-08, -1.135435e-08, 
    -1.100611e-08, -1.073674e-08, -1.017661e-08, -9.611314e-09, 
    -9.131591e-09, -8.760584e-09,
  -4.887391e-09, -6.245313e-09, -7.680378e-09, -8.728169e-09, -9.730906e-09, 
    -1.083243e-08, -1.170126e-08, -1.229238e-08, -1.204627e-08, 
    -1.137756e-08, -1.09068e-08, -1.057442e-08, -1.015855e-08, -9.645596e-09, 
    -9.044824e-09,
  -4.473825e-09, -5.167387e-09, -6.761753e-09, -8.302124e-09, -9.381631e-09, 
    -1.046824e-08, -1.148847e-08, -1.229332e-08, -1.255837e-08, -1.21952e-08, 
    -1.155835e-08, -1.101978e-08, -1.059567e-08, -1.012343e-08, -9.59828e-09,
  -4.144916e-09, -4.548674e-09, -5.612546e-09, -7.439907e-09, -8.953079e-09, 
    -1.017873e-08, -1.134111e-08, -1.245198e-08, -1.303059e-08, 
    -1.298082e-08, -1.232401e-08, -1.181675e-08, -1.128726e-08, 
    -1.062292e-08, -9.944622e-09,
  -3.825773e-09, -4.197574e-09, -4.765394e-09, -6.267377e-09, -8.035732e-09, 
    -9.730138e-09, -1.098846e-08, -1.226506e-08, -1.307064e-08, 
    -1.363496e-08, -1.328342e-08, -1.24786e-08, -1.19673e-08, -1.144376e-08, 
    -1.082006e-08,
  -9.881183e-09, -1.101554e-08, -1.095457e-08, -1.172684e-08, -1.237945e-08, 
    -1.359914e-08, -1.481843e-08, -1.64778e-08, -1.827592e-08, -1.864906e-08, 
    -1.709269e-08, -1.572942e-08, -1.546116e-08, -1.548043e-08, -1.59725e-08,
  -8.659774e-09, -9.796916e-09, -1.05759e-08, -1.137783e-08, -1.247788e-08, 
    -1.218613e-08, -1.350982e-08, -1.487853e-08, -1.671745e-08, 
    -1.872433e-08, -1.897716e-08, -1.71957e-08, -1.603134e-08, -1.559884e-08, 
    -1.553118e-08,
  -7.074842e-09, -8.122714e-09, -9.326151e-09, -1.048444e-08, -1.208478e-08, 
    -1.241972e-08, -1.222573e-08, -1.346469e-08, -1.500347e-08, 
    -1.723508e-08, -1.886621e-08, -1.859471e-08, -1.721038e-08, 
    -1.632853e-08, -1.582285e-08,
  -6.064489e-09, -6.579135e-09, -7.686446e-09, -9.079353e-09, -1.071153e-08, 
    -1.228678e-08, -1.207064e-08, -1.243322e-08, -1.334574e-08, 
    -1.522904e-08, -1.75434e-08, -1.867073e-08, -1.816115e-08, -1.718004e-08, 
    -1.656155e-08,
  -5.224176e-09, -5.639278e-09, -6.242746e-09, -7.396673e-09, -9.224363e-09, 
    -1.108688e-08, -1.175813e-08, -1.187923e-08, -1.21575e-08, -1.313512e-08, 
    -1.563497e-08, -1.744201e-08, -1.82121e-08, -1.782867e-08, -1.721117e-08,
  -4.571658e-09, -4.977004e-09, -5.20849e-09, -5.930141e-09, -7.457365e-09, 
    -9.575415e-09, -1.110604e-08, -1.145496e-08, -1.161686e-08, 
    -1.175791e-08, -1.329857e-08, -1.593891e-08, -1.709402e-08, 
    -1.758752e-08, -1.747719e-08,
  -4.315562e-09, -4.535459e-09, -4.751196e-09, -4.992465e-09, -5.915912e-09, 
    -7.924978e-09, -9.907687e-09, -1.070529e-08, -1.130163e-08, 
    -1.136417e-08, -1.139844e-08, -1.37864e-08, -1.555158e-08, -1.656942e-08, 
    -1.697616e-08,
  -4.167608e-09, -4.232739e-09, -4.439402e-09, -4.610305e-09, -4.954e-09, 
    -6.268033e-09, -8.647678e-09, -9.84942e-09, -1.067147e-08, -1.115359e-08, 
    -1.0951e-08, -1.172545e-08, -1.369777e-08, -1.51409e-08, -1.597894e-08,
  -3.90512e-09, -3.952737e-09, -4.115694e-09, -4.339764e-09, -4.627235e-09, 
    -5.114443e-09, -6.964957e-09, -8.984921e-09, -9.703147e-09, 
    -1.047654e-08, -1.081699e-08, -1.076423e-08, -1.183404e-08, 
    -1.360024e-08, -1.475826e-08,
  -3.510804e-09, -3.756537e-09, -3.826636e-09, -4.076317e-09, -4.321818e-09, 
    -4.683315e-09, -5.588193e-09, -7.680114e-09, -8.920582e-09, 
    -9.700507e-09, -1.039069e-08, -1.03805e-08, -1.073298e-08, -1.212168e-08, 
    -1.351249e-08,
  -1.169241e-08, -1.254521e-08, -1.316329e-08, -1.362135e-08, -1.421633e-08, 
    -1.506139e-08, -1.678198e-08, -1.685857e-08, -1.622102e-08, 
    -1.345775e-08, -1.302474e-08, -1.334136e-08, -1.522666e-08, 
    -1.731811e-08, -1.820779e-08,
  -1.068159e-08, -1.132502e-08, -1.193363e-08, -1.237792e-08, -1.318686e-08, 
    -1.389277e-08, -1.455473e-08, -1.581661e-08, -1.561917e-08, 
    -1.435673e-08, -1.368557e-08, -1.352392e-08, -1.498771e-08, 
    -1.751464e-08, -1.870293e-08,
  -1.00142e-08, -1.030828e-08, -1.078943e-08, -1.145526e-08, -1.212574e-08, 
    -1.310213e-08, -1.329203e-08, -1.399373e-08, -1.487509e-08, 
    -1.468084e-08, -1.403935e-08, -1.396891e-08, -1.459445e-08, 
    -1.746593e-08, -1.846203e-08,
  -9.778226e-09, -9.855023e-09, -1.016037e-08, -1.065203e-08, -1.134296e-08, 
    -1.222524e-08, -1.262703e-08, -1.295797e-08, -1.362962e-08, 
    -1.395988e-08, -1.429827e-08, -1.448741e-08, -1.468118e-08, 
    -1.717889e-08, -1.848266e-08,
  -9.330728e-09, -9.573363e-09, -9.783467e-09, -1.01397e-08, -1.060503e-08, 
    -1.139138e-08, -1.213833e-08, -1.228802e-08, -1.279068e-08, 
    -1.313693e-08, -1.341628e-08, -1.485442e-08, -1.494456e-08, 
    -1.644947e-08, -1.766532e-08,
  -8.518321e-09, -8.863211e-09, -9.416198e-09, -9.789828e-09, -1.010265e-08, 
    -1.077717e-08, -1.138722e-08, -1.17629e-08, -1.220985e-08, -1.244675e-08, 
    -1.274142e-08, -1.399292e-08, -1.526876e-08, -1.619769e-08, -1.722984e-08,
  -7.615525e-09, -8.052609e-09, -8.42704e-09, -9.133073e-09, -9.519411e-09, 
    -1.009519e-08, -1.086856e-08, -1.14411e-08, -1.17109e-08, -1.210599e-08, 
    -1.221134e-08, -1.326512e-08, -1.476374e-08, -1.618328e-08, -1.675601e-08,
  -6.816104e-09, -7.374324e-09, -7.717344e-09, -8.278686e-09, -8.763425e-09, 
    -9.185575e-09, -1.000712e-08, -1.071987e-08, -1.128965e-08, 
    -1.178071e-08, -1.196844e-08, -1.242395e-08, -1.399834e-08, 
    -1.588321e-08, -1.670639e-08,
  -6.025411e-09, -6.53742e-09, -6.963845e-09, -7.455817e-09, -8.123412e-09, 
    -8.517439e-09, -9.02778e-09, -9.967547e-09, -1.048722e-08, -1.111148e-08, 
    -1.176494e-08, -1.225056e-08, -1.302814e-08, -1.510103e-08, -1.643158e-08,
  -5.241541e-09, -5.682312e-09, -6.211821e-09, -6.678287e-09, -7.143111e-09, 
    -7.644586e-09, -8.144699e-09, -9.055993e-09, -9.709601e-09, 
    -1.036437e-08, -1.108613e-08, -1.204943e-08, -1.246475e-08, -1.39631e-08, 
    -1.600326e-08,
  -5.78939e-09, -5.924553e-09, -6.002383e-09, -6.239016e-09, -6.480446e-09, 
    -6.942083e-09, -7.53878e-09, -8.253692e-09, -9.246146e-09, -9.957392e-09, 
    -1.068577e-08, -1.13605e-08, -1.194961e-08, -1.276064e-08, -1.285657e-08,
  -5.52338e-09, -5.715694e-09, -5.776505e-09, -5.950268e-09, -6.187802e-09, 
    -6.5586e-09, -7.192159e-09, -7.810306e-09, -8.704575e-09, -9.419142e-09, 
    -1.02649e-08, -1.11024e-08, -1.172197e-08, -1.261871e-08, -1.319774e-08,
  -5.092357e-09, -5.388993e-09, -5.523647e-09, -5.681509e-09, -5.918392e-09, 
    -6.244934e-09, -6.805411e-09, -7.487357e-09, -8.253179e-09, 
    -9.032352e-09, -9.828713e-09, -1.075042e-08, -1.131725e-08, 
    -1.252837e-08, -1.329815e-08,
  -4.580829e-09, -4.908597e-09, -5.182311e-09, -5.40432e-09, -5.673153e-09, 
    -6.004787e-09, -6.444334e-09, -7.093815e-09, -7.855216e-09, 
    -8.555423e-09, -9.459296e-09, -1.035027e-08, -1.11532e-08, -1.222683e-08, 
    -1.336499e-08,
  -4.054471e-09, -4.420355e-09, -4.840923e-09, -5.113187e-09, -5.427335e-09, 
    -5.778601e-09, -6.220639e-09, -6.764967e-09, -7.433067e-09, 
    -8.106248e-09, -8.991988e-09, -9.934913e-09, -1.087693e-08, 
    -1.210137e-08, -1.322307e-08,
  -3.390161e-09, -3.871536e-09, -4.409372e-09, -4.779793e-09, -5.11545e-09, 
    -5.460683e-09, -5.918538e-09, -6.487848e-09, -7.131086e-09, 
    -7.664116e-09, -8.579673e-09, -9.503816e-09, -1.066624e-08, 
    -1.160352e-08, -1.302674e-08,
  -2.746225e-09, -3.32181e-09, -3.921101e-09, -4.41912e-09, -4.794418e-09, 
    -5.147599e-09, -5.597251e-09, -6.188705e-09, -6.866463e-09, 
    -7.390546e-09, -8.042893e-09, -9.066874e-09, -1.02712e-08, -1.155167e-08, 
    -1.272626e-08,
  -2.115931e-09, -2.627294e-09, -3.32451e-09, -3.933992e-09, -4.334356e-09, 
    -4.724193e-09, -5.208741e-09, -5.807537e-09, -6.599513e-09, 
    -7.212938e-09, -7.742892e-09, -8.525838e-09, -9.729736e-09, 
    -1.096868e-08, -1.24838e-08,
  -1.702639e-09, -2.030091e-09, -2.587021e-09, -3.306067e-09, -3.852795e-09, 
    -4.279392e-09, -4.761801e-09, -5.335813e-09, -6.15153e-09, -6.998663e-09, 
    -7.596159e-09, -8.186026e-09, -9.224435e-09, -1.055382e-08, -1.18262e-08,
  -1.447511e-09, -1.673139e-09, -1.994678e-09, -2.554926e-09, -3.132337e-09, 
    -3.775233e-09, -4.383066e-09, -4.962967e-09, -5.694776e-09, 
    -6.585243e-09, -7.350337e-09, -7.892942e-09, -8.70648e-09, -1.006501e-08, 
    -1.132718e-08,
  -2.424583e-09, -1.984025e-09, -2.066489e-09, -2.187217e-09, -2.288402e-09, 
    -2.411878e-09, -2.534361e-09, -2.824484e-09, -3.065738e-09, 
    -3.421369e-09, -3.698873e-09, -4.086751e-09, -4.544427e-09, 
    -5.198789e-09, -5.862388e-09,
  -2.069121e-09, -1.889124e-09, -1.955722e-09, -1.866074e-09, -1.902553e-09, 
    -2.020826e-09, -2.249538e-09, -2.540824e-09, -2.841782e-09, 
    -3.083507e-09, -3.299995e-09, -3.578841e-09, -4.038508e-09, 
    -4.656583e-09, -5.390719e-09,
  -2.109691e-09, -2.19553e-09, -2.240284e-09, -2.156129e-09, -2.115385e-09, 
    -2.067711e-09, -1.955819e-09, -2.056725e-09, -2.394161e-09, -2.80208e-09, 
    -3.113194e-09, -3.396428e-09, -3.637683e-09, -4.210975e-09, -4.931632e-09,
  -1.703671e-09, -1.772134e-09, -1.834693e-09, -1.945977e-09, -1.952794e-09, 
    -2.070829e-09, -2.104744e-09, -2.001896e-09, -2.122532e-09, 
    -2.529647e-09, -2.912062e-09, -3.337751e-09, -3.544053e-09, 
    -3.878673e-09, -4.510798e-09,
  -1.291084e-09, -1.339391e-09, -1.420625e-09, -1.561548e-09, -1.551519e-09, 
    -1.806456e-09, -2.133861e-09, -2.257933e-09, -2.376328e-09, 
    -2.571924e-09, -2.835106e-09, -3.230016e-09, -3.635486e-09, -3.82649e-09, 
    -4.208867e-09,
  -9.549423e-10, -9.870069e-10, -1.061585e-09, -1.046176e-09, -1.187633e-09, 
    -1.468558e-09, -1.804604e-09, -2.170186e-09, -2.39688e-09, -2.723075e-09, 
    -2.984842e-09, -3.234921e-09, -3.574685e-09, -3.919701e-09, -4.162272e-09,
  -8.307248e-10, -8.543778e-10, -8.742404e-10, -6.816969e-10, -8.864949e-10, 
    -1.15396e-09, -1.393226e-09, -1.762666e-09, -2.126055e-09, -2.520835e-09, 
    -2.999886e-09, -3.356031e-09, -3.631755e-09, -3.932486e-09, -4.199621e-09,
  -5.505205e-10, -6.125978e-10, -6.894145e-10, -6.446633e-10, -6.353943e-10, 
    -8.35969e-10, -1.032935e-09, -1.311042e-09, -1.714741e-09, -2.128415e-09, 
    -2.71887e-09, -3.294194e-09, -3.69126e-09, -4.036339e-09, -4.214117e-09,
  -3.735306e-10, -4.266987e-10, -5.201279e-10, -5.333233e-10, -5.116037e-10, 
    -6.254878e-10, -8.116758e-10, -9.844068e-10, -1.240422e-09, -1.69702e-09, 
    -2.299791e-09, -3.046194e-09, -3.668418e-09, -4.092003e-09, -4.285833e-09,
  -1.774376e-10, -2.185157e-10, -2.286457e-10, -3.5081e-10, -3.296947e-10, 
    -4.497825e-10, -5.832727e-10, -8.449547e-10, -9.35765e-10, -1.222152e-09, 
    -1.801696e-09, -2.624683e-09, -3.473841e-09, -4.130043e-09, -4.349162e-09,
  -6.33338e-09, -6.587452e-09, -6.798222e-09, -7.002626e-09, -7.285473e-09, 
    -7.585987e-09, -7.932718e-09, -8.26511e-09, -8.593572e-09, -8.845891e-09, 
    -9.055472e-09, -9.223858e-09, -9.308752e-09, -9.257615e-09, -9.171531e-09,
  -5.056643e-09, -5.220011e-09, -5.357274e-09, -5.529545e-09, -5.680505e-09, 
    -5.885161e-09, -6.034632e-09, -6.205279e-09, -6.444591e-09, 
    -6.742964e-09, -7.082979e-09, -7.422875e-09, -7.723235e-09, 
    -7.843693e-09, -7.907329e-09,
  -4.745426e-09, -4.716097e-09, -4.691474e-09, -4.716509e-09, -4.708389e-09, 
    -4.77588e-09, -4.833402e-09, -4.879511e-09, -4.962056e-09, -5.115819e-09, 
    -5.372554e-09, -5.689374e-09, -5.993343e-09, -6.207705e-09, -6.348677e-09,
  -4.766923e-09, -4.632325e-09, -4.507754e-09, -4.408174e-09, -4.293465e-09, 
    -4.243972e-09, -4.181872e-09, -4.125731e-09, -4.057895e-09, 
    -4.084557e-09, -4.238422e-09, -4.434727e-09, -4.619313e-09, 
    -4.747563e-09, -4.899782e-09,
  -5.043371e-09, -4.848059e-09, -4.665768e-09, -4.494716e-09, -4.329257e-09, 
    -4.170884e-09, -4.063073e-09, -3.922252e-09, -3.780399e-09, 
    -3.676526e-09, -3.673007e-09, -3.716716e-09, -3.772814e-09, 
    -3.839365e-09, -3.981429e-09,
  -4.974528e-09, -4.813376e-09, -4.625769e-09, -4.467538e-09, -4.293273e-09, 
    -4.110543e-09, -3.883015e-09, -3.646425e-09, -3.459279e-09, -3.36079e-09, 
    -3.341396e-09, -3.32397e-09, -3.297682e-09, -3.30642e-09, -3.424989e-09,
  -4.427862e-09, -4.380472e-09, -4.253404e-09, -4.144494e-09, -4.047075e-09, 
    -3.986293e-09, -3.792873e-09, -3.551571e-09, -3.312729e-09, 
    -3.186305e-09, -3.066057e-09, -3.010319e-09, -2.966292e-09, 
    -2.983984e-09, -3.139335e-09,
  -3.588461e-09, -3.647744e-09, -3.594498e-09, -3.521521e-09, -3.502066e-09, 
    -3.46492e-09, -3.382247e-09, -3.244975e-09, -3.216164e-09, -3.137248e-09, 
    -3.080399e-09, -2.95191e-09, -2.822949e-09, -2.745642e-09, -2.854738e-09,
  -2.602655e-09, -2.681308e-09, -2.738576e-09, -2.798819e-09, -2.944451e-09, 
    -2.936751e-09, -2.930194e-09, -2.87675e-09, -2.925389e-09, -2.941106e-09, 
    -2.930563e-09, -2.884967e-09, -2.810796e-09, -2.720688e-09, -2.700784e-09,
  -1.658053e-09, -1.706432e-09, -1.77036e-09, -1.932111e-09, -2.136183e-09, 
    -2.297435e-09, -2.356854e-09, -2.323212e-09, -2.420592e-09, 
    -2.607611e-09, -2.663155e-09, -2.692953e-09, -2.713344e-09, 
    -2.687255e-09, -2.665187e-09,
  -1.404319e-08, -1.415144e-08, -1.434745e-08, -1.45841e-08, -1.47597e-08, 
    -1.49675e-08, -1.509092e-08, -1.516133e-08, -1.519194e-08, -1.518097e-08, 
    -1.518249e-08, -1.520285e-08, -1.526503e-08, -1.535808e-08, -1.54391e-08,
  -1.2706e-08, -1.28858e-08, -1.300262e-08, -1.322781e-08, -1.346257e-08, 
    -1.364545e-08, -1.379276e-08, -1.391305e-08, -1.395169e-08, 
    -1.393303e-08, -1.387896e-08, -1.377565e-08, -1.366355e-08, 
    -1.355619e-08, -1.350364e-08,
  -1.186759e-08, -1.190697e-08, -1.200188e-08, -1.21095e-08, -1.225815e-08, 
    -1.242412e-08, -1.259264e-08, -1.270934e-08, -1.279529e-08, 
    -1.277407e-08, -1.270681e-08, -1.25712e-08, -1.238512e-08, -1.215312e-08, 
    -1.192251e-08,
  -1.136973e-08, -1.138722e-08, -1.137668e-08, -1.137993e-08, -1.136955e-08, 
    -1.142739e-08, -1.151323e-08, -1.16259e-08, -1.169617e-08, -1.172672e-08, 
    -1.168484e-08, -1.156884e-08, -1.140738e-08, -1.117979e-08, -1.091144e-08,
  -1.034275e-08, -1.062403e-08, -1.077412e-08, -1.0811e-08, -1.074783e-08, 
    -1.067999e-08, -1.058668e-08, -1.062149e-08, -1.069537e-08, 
    -1.074229e-08, -1.074682e-08, -1.066282e-08, -1.056066e-08, 
    -1.040994e-08, -1.023691e-08,
  -9.228219e-09, -9.660615e-09, -9.949554e-09, -1.01198e-08, -1.014642e-08, 
    -1.010403e-08, -1.006147e-08, -9.964283e-09, -9.897881e-09, 
    -9.867668e-09, -9.922647e-09, -9.89756e-09, -9.809621e-09, -9.715969e-09, 
    -9.61127e-09,
  -7.88223e-09, -8.283077e-09, -8.704184e-09, -9.04982e-09, -9.258989e-09, 
    -9.30274e-09, -9.35619e-09, -9.385677e-09, -9.396325e-09, -9.37024e-09, 
    -9.394437e-09, -9.390091e-09, -9.332219e-09, -9.22197e-09, -9.136944e-09,
  -6.526097e-09, -6.876054e-09, -7.29148e-09, -7.690352e-09, -8.053891e-09, 
    -8.291827e-09, -8.441328e-09, -8.517352e-09, -8.61876e-09, -8.677199e-09, 
    -8.703247e-09, -8.754951e-09, -8.767044e-09, -8.705498e-09, -8.584419e-09,
  -5.471919e-09, -5.603263e-09, -5.85228e-09, -6.20625e-09, -6.614962e-09, 
    -6.981544e-09, -7.269477e-09, -7.455962e-09, -7.568553e-09, 
    -7.670562e-09, -7.719843e-09, -7.764863e-09, -7.803436e-09, 
    -7.832481e-09, -7.758701e-09,
  -4.787527e-09, -4.822434e-09, -4.88263e-09, -5.001545e-09, -5.232875e-09, 
    -5.605016e-09, -5.99863e-09, -6.264761e-09, -6.411019e-09, -6.536026e-09, 
    -6.635894e-09, -6.719804e-09, -6.770566e-09, -6.836964e-09, -6.874188e-09,
  -2.370204e-08, -2.346169e-08, -2.309774e-08, -2.25943e-08, -2.155302e-08, 
    -2.088027e-08, -2.077633e-08, -2.104099e-08, -2.152296e-08, 
    -2.170404e-08, -2.182271e-08, -2.169523e-08, -2.171728e-08, 
    -2.168791e-08, -2.189505e-08,
  -2.268451e-08, -2.25344e-08, -2.252544e-08, -2.236667e-08, -2.202861e-08, 
    -2.142537e-08, -2.097261e-08, -2.063946e-08, -2.074237e-08, 
    -2.093993e-08, -2.120126e-08, -2.134658e-08, -2.148011e-08, -2.14137e-08, 
    -2.151741e-08,
  -2.126234e-08, -2.131161e-08, -2.143155e-08, -2.151544e-08, -2.147188e-08, 
    -2.123481e-08, -2.102248e-08, -2.077883e-08, -2.066949e-08, 
    -2.065413e-08, -2.070747e-08, -2.079777e-08, -2.085453e-08, 
    -2.086953e-08, -2.079758e-08,
  -1.865137e-08, -1.941579e-08, -1.988213e-08, -2.017835e-08, -2.03964e-08, 
    -2.034632e-08, -2.02854e-08, -2.021424e-08, -2.023527e-08, -2.020354e-08, 
    -2.022937e-08, -2.029351e-08, -2.031681e-08, -2.036821e-08, -2.032002e-08,
  -1.568734e-08, -1.673402e-08, -1.756481e-08, -1.827942e-08, -1.86196e-08, 
    -1.884787e-08, -1.885028e-08, -1.883055e-08, -1.878521e-08, 
    -1.874316e-08, -1.877439e-08, -1.880298e-08, -1.891026e-08, 
    -1.896512e-08, -1.903127e-08,
  -1.349803e-08, -1.403119e-08, -1.486885e-08, -1.563605e-08, -1.628769e-08, 
    -1.667419e-08, -1.691328e-08, -1.695484e-08, -1.692851e-08, 
    -1.679137e-08, -1.665597e-08, -1.65708e-08, -1.652334e-08, -1.651543e-08, 
    -1.646156e-08,
  -1.191933e-08, -1.246658e-08, -1.280173e-08, -1.337602e-08, -1.392083e-08, 
    -1.433909e-08, -1.466324e-08, -1.482073e-08, -1.484552e-08, 
    -1.478589e-08, -1.463116e-08, -1.438733e-08, -1.414369e-08, 
    -1.394216e-08, -1.371451e-08,
  -1.06286e-08, -1.121817e-08, -1.150944e-08, -1.176431e-08, -1.206442e-08, 
    -1.238764e-08, -1.267523e-08, -1.277206e-08, -1.276835e-08, 
    -1.269502e-08, -1.257155e-08, -1.236497e-08, -1.211023e-08, 
    -1.181738e-08, -1.148882e-08,
  -9.64877e-09, -9.878042e-09, -1.037782e-08, -1.059428e-08, -1.080031e-08, 
    -1.091201e-08, -1.102618e-08, -1.115739e-08, -1.113745e-08, 
    -1.108909e-08, -1.098939e-08, -1.085325e-08, -1.061648e-08, 
    -1.035006e-08, -1.004517e-08,
  -8.664073e-09, -9.013719e-09, -9.228564e-09, -9.571239e-09, -9.610481e-09, 
    -9.782481e-09, -9.979199e-09, -9.957042e-09, -9.943417e-09, -9.876e-09, 
    -9.77847e-09, -9.644983e-09, -9.45497e-09, -9.239521e-09, -9.055151e-09,
  -1.809487e-08, -1.880708e-08, -1.970075e-08, -2.085639e-08, -2.231302e-08, 
    -2.400281e-08, -2.539667e-08, -2.54847e-08, -2.484834e-08, -2.421725e-08, 
    -2.382692e-08, -2.386202e-08, -2.366635e-08, -2.456974e-08, -2.416407e-08,
  -1.760906e-08, -1.885082e-08, -1.964357e-08, -2.046034e-08, -2.194039e-08, 
    -2.326159e-08, -2.475795e-08, -2.54342e-08, -2.509512e-08, -2.448837e-08, 
    -2.409344e-08, -2.380367e-08, -2.331511e-08, -2.336472e-08, -2.352514e-08,
  -1.733591e-08, -1.85203e-08, -1.946071e-08, -2.009615e-08, -2.137081e-08, 
    -2.273209e-08, -2.405869e-08, -2.513557e-08, -2.514327e-08, 
    -2.449855e-08, -2.411805e-08, -2.387383e-08, -2.340615e-08, 
    -2.313956e-08, -2.319564e-08,
  -1.677991e-08, -1.8157e-08, -1.936919e-08, -1.997492e-08, -2.091107e-08, 
    -2.237919e-08, -2.363394e-08, -2.455292e-08, -2.528929e-08, 
    -2.493419e-08, -2.440331e-08, -2.42691e-08, -2.39816e-08, -2.337607e-08, 
    -2.352458e-08,
  -1.59117e-08, -1.712847e-08, -1.884535e-08, -1.99357e-08, -2.054952e-08, 
    -2.180172e-08, -2.334064e-08, -2.438961e-08, -2.512797e-08, 
    -2.543915e-08, -2.501734e-08, -2.485983e-08, -2.47077e-08, -2.41935e-08, 
    -2.381522e-08,
  -1.58814e-08, -1.622091e-08, -1.749625e-08, -1.928362e-08, -2.039935e-08, 
    -2.139453e-08, -2.269146e-08, -2.398086e-08, -2.499044e-08, 
    -2.578735e-08, -2.560029e-08, -2.543876e-08, -2.531607e-08, 
    -2.503878e-08, -2.448103e-08,
  -1.584738e-08, -1.579183e-08, -1.633317e-08, -1.758376e-08, -1.948601e-08, 
    -2.090657e-08, -2.216217e-08, -2.345422e-08, -2.445545e-08, 
    -2.570691e-08, -2.620272e-08, -2.620792e-08, -2.592569e-08, 
    -2.566238e-08, -2.509261e-08,
  -1.566697e-08, -1.605009e-08, -1.608899e-08, -1.638229e-08, -1.773662e-08, 
    -1.968673e-08, -2.126389e-08, -2.255263e-08, -2.377106e-08, 
    -2.473102e-08, -2.575106e-08, -2.627795e-08, -2.627041e-08, 
    -2.597429e-08, -2.534144e-08,
  -1.446631e-08, -1.563831e-08, -1.624326e-08, -1.628399e-08, -1.640058e-08, 
    -1.77973e-08, -1.990475e-08, -2.138107e-08, -2.264201e-08, -2.379521e-08, 
    -2.471746e-08, -2.544054e-08, -2.575454e-08, -2.577069e-08, -2.540159e-08,
  -1.23951e-08, -1.400201e-08, -1.544463e-08, -1.630432e-08, -1.632622e-08, 
    -1.60054e-08, -1.758174e-08, -1.974471e-08, -2.113985e-08, -2.227431e-08, 
    -2.328651e-08, -2.424036e-08, -2.487939e-08, -2.5024e-08, -2.490968e-08,
  -1.502275e-08, -1.556787e-08, -1.618451e-08, -1.676853e-08, -1.781131e-08, 
    -1.896242e-08, -2.069811e-08, -2.175255e-08, -2.271918e-08, 
    -2.317008e-08, -2.395721e-08, -2.489557e-08, -2.569034e-08, 
    -2.574229e-08, -2.524376e-08,
  -1.462592e-08, -1.504538e-08, -1.561644e-08, -1.616084e-08, -1.690371e-08, 
    -1.803294e-08, -1.964933e-08, -2.110285e-08, -2.201191e-08, 
    -2.328825e-08, -2.370828e-08, -2.472418e-08, -2.537604e-08, 
    -2.582567e-08, -2.539703e-08,
  -1.426366e-08, -1.459117e-08, -1.511814e-08, -1.558632e-08, -1.611158e-08, 
    -1.695152e-08, -1.821505e-08, -2.013512e-08, -2.136255e-08, 
    -2.252076e-08, -2.340307e-08, -2.438794e-08, -2.541197e-08, 
    -2.582619e-08, -2.582125e-08,
  -1.373244e-08, -1.42955e-08, -1.464566e-08, -1.517011e-08, -1.555221e-08, 
    -1.615066e-08, -1.695458e-08, -1.853991e-08, -2.038507e-08, 
    -2.171561e-08, -2.297212e-08, -2.391952e-08, -2.489876e-08, -2.56728e-08, 
    -2.610624e-08,
  -1.298096e-08, -1.380504e-08, -1.433899e-08, -1.473591e-08, -1.51541e-08, 
    -1.553459e-08, -1.629879e-08, -1.710355e-08, -1.87845e-08, -2.048807e-08, 
    -2.19269e-08, -2.326067e-08, -2.448029e-08, -2.526968e-08, -2.586309e-08,
  -1.213545e-08, -1.301561e-08, -1.385645e-08, -1.437449e-08, -1.477883e-08, 
    -1.512147e-08, -1.563468e-08, -1.655128e-08, -1.741684e-08, 
    -1.906007e-08, -2.05822e-08, -2.203552e-08, -2.351613e-08, -2.464744e-08, 
    -2.568481e-08,
  -1.171793e-08, -1.215533e-08, -1.290523e-08, -1.369362e-08, -1.429696e-08, 
    -1.47324e-08, -1.502581e-08, -1.582404e-08, -1.676025e-08, -1.764029e-08, 
    -1.915684e-08, -2.039682e-08, -2.225441e-08, -2.35734e-08, -2.482209e-08,
  -1.132625e-08, -1.190661e-08, -1.228356e-08, -1.288548e-08, -1.347125e-08, 
    -1.42545e-08, -1.468157e-08, -1.525148e-08, -1.630005e-08, -1.699529e-08, 
    -1.798812e-08, -1.894889e-08, -2.015929e-08, -2.212232e-08, -2.352876e-08,
  -1.083753e-08, -1.150795e-08, -1.212359e-08, -1.249441e-08, -1.280736e-08, 
    -1.32766e-08, -1.387733e-08, -1.431083e-08, -1.530029e-08, -1.654902e-08, 
    -1.738758e-08, -1.82166e-08, -1.876836e-08, -1.989173e-08, -2.164115e-08,
  -1.06057e-08, -1.101906e-08, -1.167608e-08, -1.234741e-08, -1.252182e-08, 
    -1.295884e-08, -1.351081e-08, -1.386764e-08, -1.410228e-08, 
    -1.517554e-08, -1.662617e-08, -1.759839e-08, -1.829698e-08, -1.86396e-08, 
    -1.955371e-08,
  -1.440441e-08, -1.504863e-08, -1.569103e-08, -1.656605e-08, -1.744751e-08, 
    -1.790461e-08, -1.830439e-08, -1.82384e-08, -1.758137e-08, -1.719481e-08, 
    -1.71591e-08, -1.743419e-08, -1.814132e-08, -1.940394e-08, -2.065796e-08,
  -1.372333e-08, -1.445535e-08, -1.517483e-08, -1.591671e-08, -1.692951e-08, 
    -1.763263e-08, -1.796589e-08, -1.846537e-08, -1.80216e-08, -1.758938e-08, 
    -1.722514e-08, -1.732753e-08, -1.767821e-08, -1.870668e-08, -1.992651e-08,
  -1.284413e-08, -1.360916e-08, -1.446287e-08, -1.527033e-08, -1.621296e-08, 
    -1.726129e-08, -1.776134e-08, -1.821009e-08, -1.83576e-08, -1.795173e-08, 
    -1.755721e-08, -1.734344e-08, -1.757776e-08, -1.803592e-08, -1.93085e-08,
  -1.195907e-08, -1.273466e-08, -1.363851e-08, -1.454773e-08, -1.543303e-08, 
    -1.656426e-08, -1.743132e-08, -1.788845e-08, -1.836615e-08, 
    -1.824294e-08, -1.799702e-08, -1.757514e-08, -1.758971e-08, 
    -1.780055e-08, -1.868067e-08,
  -1.087985e-08, -1.183242e-08, -1.267579e-08, -1.377722e-08, -1.471678e-08, 
    -1.574032e-08, -1.690135e-08, -1.755912e-08, -1.806591e-08, 
    -1.825335e-08, -1.83082e-08, -1.798879e-08, -1.773116e-08, -1.774403e-08, 
    -1.812055e-08,
  -9.755998e-09, -1.089326e-08, -1.178582e-08, -1.282824e-08, -1.390313e-08, 
    -1.490233e-08, -1.616381e-08, -1.715036e-08, -1.775695e-08, 
    -1.813179e-08, -1.830419e-08, -1.836101e-08, -1.802079e-08, 
    -1.785338e-08, -1.788732e-08,
  -8.469988e-09, -9.857009e-09, -1.088076e-08, -1.191544e-08, -1.309705e-08, 
    -1.407548e-08, -1.519036e-08, -1.636892e-08, -1.726564e-08, 
    -1.784682e-08, -1.815598e-08, -1.846195e-08, -1.839453e-08, 
    -1.808461e-08, -1.798289e-08,
  -7.571416e-09, -8.771874e-09, -9.978065e-09, -1.103343e-08, -1.215089e-08, 
    -1.332734e-08, -1.442017e-08, -1.563863e-08, -1.659119e-08, 
    -1.733383e-08, -1.792148e-08, -1.822746e-08, -1.865991e-08, 
    -1.838676e-08, -1.818058e-08,
  -7.020423e-09, -7.728471e-09, -9.037862e-09, -1.027317e-08, -1.138274e-08, 
    -1.240638e-08, -1.347442e-08, -1.461932e-08, -1.592937e-08, 
    -1.676292e-08, -1.742128e-08, -1.806901e-08, -1.850149e-08, 
    -1.873337e-08, -1.84846e-08,
  -6.750105e-09, -7.194924e-09, -8.076475e-09, -9.405968e-09, -1.076475e-08, 
    -1.204322e-08, -1.284111e-08, -1.381365e-08, -1.485104e-08, 
    -1.612369e-08, -1.67656e-08, -1.754382e-08, -1.835755e-08, -1.876133e-08, 
    -1.889634e-08,
  -1.682706e-08, -1.7408e-08, -1.783968e-08, -1.827781e-08, -1.842475e-08, 
    -1.862682e-08, -1.895803e-08, -1.936008e-08, -2.038612e-08, 
    -2.070964e-08, -1.924991e-08, -1.762254e-08, -1.731922e-08, 
    -1.736993e-08, -1.802487e-08,
  -1.541867e-08, -1.621495e-08, -1.684774e-08, -1.733056e-08, -1.774962e-08, 
    -1.800894e-08, -1.853198e-08, -1.884966e-08, -1.9708e-08, -2.06079e-08, 
    -2.012414e-08, -1.858803e-08, -1.737539e-08, -1.741601e-08, -1.77531e-08,
  -1.346413e-08, -1.442695e-08, -1.537254e-08, -1.612515e-08, -1.680569e-08, 
    -1.718887e-08, -1.763856e-08, -1.823023e-08, -1.884649e-08, 
    -2.016126e-08, -2.065971e-08, -1.968644e-08, -1.797538e-08, 
    -1.720426e-08, -1.746648e-08,
  -1.123473e-08, -1.223165e-08, -1.33732e-08, -1.444032e-08, -1.542207e-08, 
    -1.62227e-08, -1.675791e-08, -1.738546e-08, -1.796259e-08, -1.904153e-08, 
    -2.046741e-08, -2.044728e-08, -1.947411e-08, -1.770869e-08, -1.731857e-08,
  -8.997915e-09, -9.98821e-09, -1.112704e-08, -1.240039e-08, -1.354623e-08, 
    -1.470625e-08, -1.555199e-08, -1.639694e-08, -1.706894e-08, 
    -1.797722e-08, -1.931235e-08, -2.01132e-08, -1.990474e-08, -1.89818e-08, 
    -1.767985e-08,
  -7.418283e-09, -8.065918e-09, -8.969866e-09, -1.015494e-08, -1.14722e-08, 
    -1.274986e-08, -1.386523e-08, -1.496785e-08, -1.601173e-08, -1.70336e-08, 
    -1.817414e-08, -1.951514e-08, -1.974705e-08, -1.947524e-08, -1.838725e-08,
  -6.41595e-09, -6.948571e-09, -7.552287e-09, -8.344919e-09, -9.467088e-09, 
    -1.083408e-08, -1.208529e-08, -1.325531e-08, -1.441468e-08, -1.56691e-08, 
    -1.706919e-08, -1.843258e-08, -1.935115e-08, -1.949181e-08, -1.889789e-08,
  -5.078324e-09, -5.782086e-09, -6.418382e-09, -7.105138e-09, -7.853346e-09, 
    -9.015232e-09, -1.03817e-08, -1.166178e-08, -1.297929e-08, -1.407799e-08, 
    -1.563781e-08, -1.704633e-08, -1.860903e-08, -1.913937e-08, -1.92153e-08,
  -4.07502e-09, -4.377556e-09, -5.060547e-09, -5.892313e-09, -6.748039e-09, 
    -7.623561e-09, -8.749585e-09, -9.990669e-09, -1.142191e-08, 
    -1.272183e-08, -1.404235e-08, -1.566342e-08, -1.716213e-08, 
    -1.858385e-08, -1.899911e-08,
  -3.786379e-09, -3.699443e-09, -3.852509e-09, -4.420003e-09, -5.301309e-09, 
    -6.486736e-09, -7.6685e-09, -8.683299e-09, -9.917982e-09, -1.127986e-08, 
    -1.263433e-08, -1.40626e-08, -1.563535e-08, -1.735398e-08, -1.842485e-08,
  -1.957922e-08, -1.985662e-08, -2.006239e-08, -2.020455e-08, -2.024965e-08, 
    -2.025374e-08, -2.022303e-08, -2.036752e-08, -2.049954e-08, 
    -2.068966e-08, -2.084568e-08, -2.088817e-08, -2.111906e-08, 
    -2.102366e-08, -2.032836e-08,
  -1.871854e-08, -1.912108e-08, -1.932435e-08, -1.951665e-08, -1.955922e-08, 
    -1.964777e-08, -1.977776e-08, -2.000439e-08, -2.016615e-08, 
    -2.026525e-08, -2.009362e-08, -1.985496e-08, -1.967967e-08, 
    -1.962532e-08, -1.983713e-08,
  -1.759644e-08, -1.820536e-08, -1.853845e-08, -1.868652e-08, -1.880609e-08, 
    -1.884831e-08, -1.892958e-08, -1.916898e-08, -1.945667e-08, 
    -1.974005e-08, -1.964776e-08, -1.945358e-08, -1.90665e-08, -1.869969e-08, 
    -1.857932e-08,
  -1.588185e-08, -1.65546e-08, -1.725684e-08, -1.778051e-08, -1.804734e-08, 
    -1.814773e-08, -1.825397e-08, -1.837337e-08, -1.840762e-08, -1.8617e-08, 
    -1.876563e-08, -1.894443e-08, -1.905297e-08, -1.863108e-08, -1.825378e-08,
  -1.412886e-08, -1.470579e-08, -1.542459e-08, -1.619199e-08, -1.673702e-08, 
    -1.710218e-08, -1.750555e-08, -1.766726e-08, -1.761997e-08, 
    -1.740248e-08, -1.74025e-08, -1.777292e-08, -1.829316e-08, -1.875918e-08, 
    -1.851416e-08,
  -1.191464e-08, -1.24644e-08, -1.327183e-08, -1.438422e-08, -1.523748e-08, 
    -1.5853e-08, -1.639533e-08, -1.672871e-08, -1.687944e-08, -1.695486e-08, 
    -1.683846e-08, -1.682511e-08, -1.717055e-08, -1.782589e-08, -1.850057e-08,
  -9.806206e-09, -1.020329e-08, -1.079299e-08, -1.162828e-08, -1.278416e-08, 
    -1.392269e-08, -1.477909e-08, -1.54286e-08, -1.580155e-08, -1.602416e-08, 
    -1.623652e-08, -1.64713e-08, -1.66337e-08, -1.685388e-08, -1.750169e-08,
  -8.428097e-09, -8.819681e-09, -9.268579e-09, -9.677361e-09, -1.02636e-08, 
    -1.111717e-08, -1.196477e-08, -1.303442e-08, -1.39007e-08, -1.452858e-08, 
    -1.500896e-08, -1.553529e-08, -1.598855e-08, -1.631373e-08, -1.653378e-08,
  -7.373164e-09, -7.470641e-09, -7.752422e-09, -8.115006e-09, -8.562146e-09, 
    -9.130813e-09, -9.816444e-09, -1.052916e-08, -1.14408e-08, -1.238126e-08, 
    -1.310343e-08, -1.38518e-08, -1.471953e-08, -1.549038e-08, -1.624653e-08,
  -6.385968e-09, -6.560167e-09, -6.637284e-09, -6.810412e-09, -6.915825e-09, 
    -7.381064e-09, -8.265546e-09, -8.981272e-09, -9.425548e-09, 
    -1.025392e-08, -1.111243e-08, -1.17947e-08, -1.267368e-08, -1.377721e-08, 
    -1.469523e-08,
  -2.00859e-08, -2.042131e-08, -2.105239e-08, -2.177191e-08, -2.240339e-08, 
    -2.297174e-08, -2.332657e-08, -2.37233e-08, -2.42107e-08, -2.423934e-08, 
    -2.456627e-08, -2.511665e-08, -2.540011e-08, -2.583302e-08, -2.68199e-08,
  -1.943524e-08, -1.99026e-08, -2.017891e-08, -2.066155e-08, -2.128875e-08, 
    -2.189047e-08, -2.256041e-08, -2.302945e-08, -2.372959e-08, 
    -2.410276e-08, -2.453776e-08, -2.492038e-08, -2.510884e-08, 
    -2.538422e-08, -2.58165e-08,
  -1.884245e-08, -1.937674e-08, -1.981611e-08, -2.004122e-08, -2.033928e-08, 
    -2.089255e-08, -2.156213e-08, -2.229048e-08, -2.295554e-08, 
    -2.361932e-08, -2.410776e-08, -2.463439e-08, -2.479013e-08, 
    -2.495176e-08, -2.549089e-08,
  -1.738873e-08, -1.811336e-08, -1.874102e-08, -1.931955e-08, -1.96575e-08, 
    -1.997866e-08, -2.051548e-08, -2.120697e-08, -2.207248e-08, 
    -2.292542e-08, -2.372076e-08, -2.428633e-08, -2.468563e-08, -2.47986e-08, 
    -2.538308e-08,
  -1.579456e-08, -1.640432e-08, -1.713364e-08, -1.789381e-08, -1.844443e-08, 
    -1.881336e-08, -1.918477e-08, -1.975326e-08, -2.044277e-08, 
    -2.130796e-08, -2.227412e-08, -2.317587e-08, -2.392149e-08, 
    -2.410219e-08, -2.445767e-08,
  -1.413912e-08, -1.471918e-08, -1.534436e-08, -1.610401e-08, -1.692969e-08, 
    -1.774582e-08, -1.815949e-08, -1.855192e-08, -1.900797e-08, 
    -1.958975e-08, -2.030692e-08, -2.105313e-08, -2.183357e-08, -2.22062e-08, 
    -2.260775e-08,
  -1.183471e-08, -1.267777e-08, -1.342543e-08, -1.416645e-08, -1.496739e-08, 
    -1.577004e-08, -1.662107e-08, -1.734529e-08, -1.793367e-08, 
    -1.835388e-08, -1.874628e-08, -1.89981e-08, -1.926308e-08, -1.971295e-08, 
    -2.020536e-08,
  -9.417924e-09, -1.035846e-08, -1.130451e-08, -1.213361e-08, -1.289669e-08, 
    -1.371677e-08, -1.445002e-08, -1.512307e-08, -1.584815e-08, 
    -1.650686e-08, -1.691068e-08, -1.715368e-08, -1.739077e-08, 
    -1.769773e-08, -1.781005e-08,
  -7.571945e-09, -8.112936e-09, -8.826909e-09, -9.623829e-09, -1.0462e-08, 
    -1.136429e-08, -1.228095e-08, -1.295926e-08, -1.349739e-08, 
    -1.403051e-08, -1.441343e-08, -1.490755e-08, -1.538658e-08, 
    -1.566378e-08, -1.599105e-08,
  -6.250741e-09, -6.665003e-09, -7.073895e-09, -7.565841e-09, -8.049653e-09, 
    -8.732349e-09, -9.734523e-09, -1.062915e-08, -1.127649e-08, 
    -1.200522e-08, -1.252199e-08, -1.310543e-08, -1.359288e-08, 
    -1.394296e-08, -1.430589e-08,
  -2.396853e-08, -2.283291e-08, -2.256184e-08, -2.084654e-08, -1.761856e-08, 
    -1.586565e-08, -1.807419e-08, -1.965718e-08, -2.047941e-08, 
    -2.083587e-08, -2.04975e-08, -2.083736e-08, -2.077126e-08, -2.142909e-08, 
    -2.232066e-08,
  -2.074366e-08, -2.122819e-08, -1.997334e-08, -1.70936e-08, -1.590462e-08, 
    -1.686232e-08, -1.83004e-08, -1.895774e-08, -1.926207e-08, -1.946129e-08, 
    -1.972247e-08, -1.983813e-08, -1.978212e-08, -2.04013e-08, -2.090039e-08,
  -1.84378e-08, -1.906185e-08, -1.823981e-08, -1.695335e-08, -1.656186e-08, 
    -1.76416e-08, -1.786071e-08, -1.755792e-08, -1.746955e-08, -1.783707e-08, 
    -1.804948e-08, -1.829993e-08, -1.870793e-08, -1.918195e-08, -1.971411e-08,
  -1.755168e-08, -1.824125e-08, -1.790836e-08, -1.750063e-08, -1.800583e-08, 
    -1.871504e-08, -1.874022e-08, -1.824173e-08, -1.807543e-08, 
    -1.838393e-08, -1.820955e-08, -1.788023e-08, -1.785432e-08, 
    -1.818151e-08, -1.855613e-08,
  -1.787613e-08, -1.853251e-08, -1.804857e-08, -1.764206e-08, -1.793398e-08, 
    -1.8429e-08, -1.856183e-08, -1.810745e-08, -1.834845e-08, -1.880656e-08, 
    -1.891099e-08, -1.851908e-08, -1.823924e-08, -1.806953e-08, -1.814182e-08,
  -1.790102e-08, -1.870884e-08, -1.907042e-08, -1.828097e-08, -1.708078e-08, 
    -1.646042e-08, -1.635263e-08, -1.627836e-08, -1.684433e-08, 
    -1.732803e-08, -1.755568e-08, -1.739377e-08, -1.737693e-08, 
    -1.746116e-08, -1.766635e-08,
  -1.750729e-08, -1.879791e-08, -2.000836e-08, -1.897567e-08, -1.702276e-08, 
    -1.626404e-08, -1.614253e-08, -1.549758e-08, -1.566213e-08, 
    -1.575624e-08, -1.621416e-08, -1.638821e-08, -1.63604e-08, -1.642288e-08, 
    -1.66447e-08,
  -1.623439e-08, -1.735406e-08, -1.804755e-08, -1.695306e-08, -1.628626e-08, 
    -1.676805e-08, -1.673437e-08, -1.641192e-08, -1.596897e-08, 
    -1.585206e-08, -1.619224e-08, -1.628655e-08, -1.645758e-08, 
    -1.639437e-08, -1.628488e-08,
  -1.456664e-08, -1.468826e-08, -1.487555e-08, -1.442685e-08, -1.434694e-08, 
    -1.518385e-08, -1.574721e-08, -1.59328e-08, -1.614388e-08, -1.612407e-08, 
    -1.620582e-08, -1.632721e-08, -1.648044e-08, -1.660579e-08, -1.674291e-08,
  -1.264981e-08, -1.246176e-08, -1.284951e-08, -1.267606e-08, -1.148696e-08, 
    -1.162662e-08, -1.261308e-08, -1.318023e-08, -1.360788e-08, 
    -1.409304e-08, -1.439632e-08, -1.479133e-08, -1.521021e-08, 
    -1.566861e-08, -1.608234e-08,
  -2.172681e-08, -2.061054e-08, -2.073044e-08, -1.928957e-08, -1.853359e-08, 
    -1.650324e-08, -1.432013e-08, -1.359758e-08, -1.296503e-08, 
    -1.193432e-08, -1.176253e-08, -1.212888e-08, -1.353125e-08, 
    -1.462608e-08, -1.632112e-08,
  -2.511442e-08, -2.364503e-08, -2.476111e-08, -2.193337e-08, -1.901673e-08, 
    -1.744827e-08, -1.799205e-08, -1.971137e-08, -1.939816e-08, 
    -1.665041e-08, -1.655044e-08, -1.699167e-08, -1.539039e-08, 
    -1.511534e-08, -1.635482e-08,
  -2.803882e-08, -2.693896e-08, -2.87027e-08, -2.51096e-08, -2.032488e-08, 
    -1.83513e-08, -1.951308e-08, -2.015889e-08, -1.780804e-08, -1.598945e-08, 
    -1.593606e-08, -1.692379e-08, -1.739643e-08, -1.674724e-08, -1.546922e-08,
  -3.038119e-08, -2.98017e-08, -2.94736e-08, -2.602864e-08, -2.362085e-08, 
    -2.15711e-08, -1.970779e-08, -1.825976e-08, -1.57362e-08, -1.467456e-08, 
    -1.519346e-08, -1.581541e-08, -1.687205e-08, -1.7607e-08, -1.767964e-08,
  -3.007668e-08, -3.114733e-08, -3.111292e-08, -2.916425e-08, -2.600265e-08, 
    -2.217861e-08, -1.920027e-08, -1.944103e-08, -1.76603e-08, -1.677118e-08, 
    -1.63146e-08, -1.633352e-08, -1.668174e-08, -1.706881e-08, -1.711497e-08,
  -3.083559e-08, -3.145848e-08, -3.109182e-08, -3.015436e-08, -2.675396e-08, 
    -2.209554e-08, -2.110071e-08, -2.054745e-08, -1.733738e-08, 
    -1.568547e-08, -1.516976e-08, -1.485086e-08, -1.449014e-08, -1.43014e-08, 
    -1.444044e-08,
  -2.988799e-08, -3.049518e-08, -3.099839e-08, -3.002938e-08, -2.59357e-08, 
    -2.226461e-08, -2.188225e-08, -2.0612e-08, -1.778786e-08, -1.656741e-08, 
    -1.550286e-08, -1.420738e-08, -1.39525e-08, -1.304366e-08, -1.29305e-08,
  -2.868914e-08, -2.939681e-08, -3.000952e-08, -2.924828e-08, -2.676147e-08, 
    -2.414851e-08, -2.268977e-08, -2.072649e-08, -1.864018e-08, 
    -1.750704e-08, -1.635517e-08, -1.529616e-08, -1.490666e-08, 
    -1.450524e-08, -1.381284e-08,
  -2.759842e-08, -2.841244e-08, -2.844819e-08, -2.823114e-08, -2.741174e-08, 
    -2.46219e-08, -2.243005e-08, -2.075015e-08, -1.873738e-08, -1.74773e-08, 
    -1.668329e-08, -1.572375e-08, -1.474559e-08, -1.494053e-08, -1.510784e-08,
  -2.562452e-08, -2.630627e-08, -2.68422e-08, -2.684699e-08, -2.593718e-08, 
    -2.341107e-08, -2.040605e-08, -1.898753e-08, -1.728465e-08, 
    -1.579111e-08, -1.470162e-08, -1.396477e-08, -1.31686e-08, -1.361611e-08, 
    -1.455918e-08,
  -8.875499e-09, -9.14531e-09, -9.013069e-09, -9.92562e-09, -1.162622e-08, 
    -1.269795e-08, -1.311708e-08, -1.238053e-08, -1.079382e-08, 
    -9.245188e-09, -8.820908e-09, -7.982546e-09, -7.43906e-09, -7.671938e-09, 
    -9.196886e-09,
  -9.91573e-09, -1.015697e-08, -1.132084e-08, -1.409838e-08, -1.51551e-08, 
    -1.477504e-08, -1.423723e-08, -1.349134e-08, -1.375752e-08, 
    -1.437741e-08, -1.240008e-08, -1.205731e-08, -1.443055e-08, 
    -1.621071e-08, -1.637271e-08,
  -1.087088e-08, -1.205062e-08, -1.52149e-08, -1.69971e-08, -1.748652e-08, 
    -1.720994e-08, -1.630208e-08, -1.711392e-08, -1.782359e-08, 
    -1.798693e-08, -1.770326e-08, -1.757439e-08, -1.749016e-08, -1.69936e-08, 
    -1.631442e-08,
  -1.284188e-08, -1.452532e-08, -1.764758e-08, -2.046472e-08, -2.124116e-08, 
    -2.043406e-08, -2.108143e-08, -2.051219e-08, -2.093381e-08, 
    -2.178454e-08, -2.118047e-08, -2.030107e-08, -1.867696e-08, 
    -1.678667e-08, -1.464302e-08,
  -1.427111e-08, -1.719522e-08, -2.271272e-08, -2.371931e-08, -2.368927e-08, 
    -2.430369e-08, -2.446768e-08, -2.471399e-08, -2.465272e-08, 
    -2.501619e-08, -2.276522e-08, -2.093963e-08, -1.797629e-08, 
    -1.575497e-08, -1.381427e-08,
  -1.594104e-08, -1.987928e-08, -2.410342e-08, -2.561358e-08, -2.600879e-08, 
    -2.599139e-08, -2.652586e-08, -2.66291e-08, -2.610554e-08, -2.480242e-08, 
    -2.377287e-08, -2.088561e-08, -1.735802e-08, -1.522954e-08, -1.457878e-08,
  -1.684444e-08, -2.167755e-08, -2.659277e-08, -2.634849e-08, -2.726029e-08, 
    -2.870449e-08, -2.970441e-08, -2.880397e-08, -2.75194e-08, -2.515132e-08, 
    -2.37863e-08, -2.194251e-08, -1.821108e-08, -1.622308e-08, -1.52541e-08,
  -1.730229e-08, -2.191955e-08, -2.65197e-08, -2.824669e-08, -2.952174e-08, 
    -3.201266e-08, -3.203037e-08, -3.217831e-08, -2.936278e-08, -2.67413e-08, 
    -2.443064e-08, -2.230441e-08, -1.840146e-08, -1.613011e-08, -1.507432e-08,
  -1.738364e-08, -2.136498e-08, -2.629729e-08, -2.856519e-08, -3.059982e-08, 
    -3.237717e-08, -3.338809e-08, -3.313743e-08, -3.12872e-08, -2.894886e-08, 
    -2.556265e-08, -2.289675e-08, -1.907227e-08, -1.673475e-08, -1.520888e-08,
  -1.646377e-08, -1.988734e-08, -2.52393e-08, -2.798318e-08, -3.164373e-08, 
    -3.319052e-08, -3.277771e-08, -3.301056e-08, -3.131523e-08, 
    -2.879304e-08, -2.507851e-08, -2.204347e-08, -1.925556e-08, 
    -1.707313e-08, -1.513724e-08,
  -7.000598e-09, -6.779155e-09, -6.507607e-09, -6.276448e-09, -6.030647e-09, 
    -5.762584e-09, -5.356365e-09, -4.820919e-09, -4.301386e-09, 
    -3.845124e-09, -3.484036e-09, -3.310438e-09, -3.39823e-09, -3.532239e-09, 
    -3.746151e-09,
  -6.69157e-09, -6.499651e-09, -6.286227e-09, -6.034788e-09, -5.762667e-09, 
    -5.498382e-09, -5.24048e-09, -5.016843e-09, -4.784519e-09, -4.455999e-09, 
    -4.151037e-09, -3.870952e-09, -3.620072e-09, -3.667169e-09, -3.950815e-09,
  -6.388942e-09, -6.138878e-09, -6.003549e-09, -5.848862e-09, -5.598848e-09, 
    -5.306809e-09, -5.003064e-09, -4.763398e-09, -4.631619e-09, 
    -4.540071e-09, -4.394802e-09, -4.325836e-09, -4.423341e-09, 
    -4.701606e-09, -5.187952e-09,
  -6.242418e-09, -6.037643e-09, -5.880637e-09, -5.707474e-09, -5.479499e-09, 
    -5.157582e-09, -4.830857e-09, -4.565485e-09, -4.360093e-09, 
    -4.334283e-09, -4.537876e-09, -5.024529e-09, -5.687863e-09, 
    -6.483648e-09, -7.082716e-09,
  -5.942281e-09, -5.887657e-09, -5.806056e-09, -5.673346e-09, -5.438848e-09, 
    -5.150344e-09, -4.831537e-09, -4.536945e-09, -4.38595e-09, -4.636421e-09, 
    -5.192334e-09, -6.471204e-09, -7.500984e-09, -7.891837e-09, -8.427619e-09,
  -5.683333e-09, -5.606987e-09, -5.586748e-09, -5.515839e-09, -5.435656e-09, 
    -5.189464e-09, -4.869151e-09, -4.763009e-09, -5.007989e-09, 
    -5.798733e-09, -7.058095e-09, -7.924484e-09, -8.584816e-09, 
    -1.019964e-08, -1.193188e-08,
  -5.432113e-09, -5.390254e-09, -5.296147e-09, -5.332148e-09, -5.311732e-09, 
    -5.246334e-09, -5.282746e-09, -5.486515e-09, -6.510654e-09, 
    -7.859761e-09, -8.67562e-09, -9.694365e-09, -1.161312e-08, -1.377305e-08, 
    -1.484267e-08,
  -5.188319e-09, -5.172662e-09, -5.118803e-09, -5.156052e-09, -5.230385e-09, 
    -5.381001e-09, -5.66297e-09, -6.923585e-09, -8.414163e-09, -9.491074e-09, 
    -1.049736e-08, -1.24752e-08, -1.517641e-08, -1.674286e-08, -1.602691e-08,
  -4.929651e-09, -4.878083e-09, -4.98519e-09, -5.104691e-09, -5.203389e-09, 
    -5.468946e-09, -6.606984e-09, -8.299301e-09, -9.614203e-09, 
    -1.100592e-08, -1.287719e-08, -1.543362e-08, -1.775236e-08, 
    -1.887728e-08, -1.839438e-08,
  -4.702814e-09, -4.670394e-09, -4.81386e-09, -4.935707e-09, -5.260059e-09, 
    -5.964031e-09, -7.494523e-09, -9.160972e-09, -1.08946e-08, -1.271397e-08, 
    -1.4854e-08, -1.74639e-08, -1.970438e-08, -2.100693e-08, -2.036573e-08,
  -8.036485e-09, -8.232653e-09, -8.308804e-09, -8.350637e-09, -8.247968e-09, 
    -8.036173e-09, -7.519354e-09, -6.90288e-09, -6.019639e-09, -5.349992e-09, 
    -4.904415e-09, -4.735516e-09, -4.695961e-09, -4.733263e-09, -4.816028e-09,
  -8.69082e-09, -8.735419e-09, -8.782581e-09, -8.888773e-09, -8.976522e-09, 
    -8.946182e-09, -8.889414e-09, -8.705755e-09, -8.486388e-09, 
    -7.984904e-09, -7.183147e-09, -6.304941e-09, -5.518111e-09, 
    -4.990069e-09, -4.709614e-09,
  -9.240643e-09, -9.179686e-09, -9.160578e-09, -9.208473e-09, -9.344244e-09, 
    -9.491536e-09, -9.574349e-09, -9.567386e-09, -9.486041e-09, 
    -9.387955e-09, -9.128589e-09, -8.716498e-09, -7.986418e-09, 
    -7.093874e-09, -6.233849e-09,
  -9.446297e-09, -9.535459e-09, -9.551501e-09, -9.532229e-09, -9.610881e-09, 
    -9.719119e-09, -9.864591e-09, -9.936537e-09, -1.000723e-08, 
    -1.000409e-08, -9.956503e-09, -9.821568e-09, -9.603959e-09, 
    -9.201662e-09, -8.68847e-09,
  -9.216106e-09, -9.534843e-09, -9.725429e-09, -9.81325e-09, -9.873357e-09, 
    -9.979202e-09, -1.007958e-08, -1.018551e-08, -1.023115e-08, 
    -1.028297e-08, -1.028381e-08, -1.028559e-08, -1.022247e-08, 
    -1.014393e-08, -9.988995e-09,
  -8.654589e-09, -9.060202e-09, -9.412455e-09, -9.717681e-09, -9.931941e-09, 
    -1.009862e-08, -1.025772e-08, -1.033468e-08, -1.041185e-08, 
    -1.043255e-08, -1.044547e-08, -1.038773e-08, -1.031567e-08, 
    -1.033038e-08, -1.035655e-08,
  -8.002215e-09, -8.421687e-09, -8.794207e-09, -9.224956e-09, -9.613177e-09, 
    -9.908427e-09, -1.017596e-08, -1.034107e-08, -1.046315e-08, 
    -1.049546e-08, -1.048708e-08, -1.042959e-08, -1.032538e-08, 
    -1.024717e-08, -1.027614e-08,
  -7.157558e-09, -7.627368e-09, -8.072083e-09, -8.47889e-09, -8.943911e-09, 
    -9.368757e-09, -9.745042e-09, -1.003009e-08, -1.021406e-08, 
    -1.032832e-08, -1.035179e-08, -1.031527e-08, -1.020886e-08, 
    -1.006596e-08, -9.946349e-09,
  -6.394985e-09, -6.779925e-09, -7.302968e-09, -7.780113e-09, -8.286566e-09, 
    -8.756834e-09, -9.19982e-09, -9.579024e-09, -9.846716e-09, -9.993639e-09, 
    -1.002981e-08, -9.931749e-09, -9.73013e-09, -9.444798e-09, -9.152046e-09,
  -5.513628e-09, -5.981481e-09, -6.356957e-09, -6.928173e-09, -7.428142e-09, 
    -8.005006e-09, -8.58161e-09, -9.020773e-09, -9.30141e-09, -9.441429e-09, 
    -9.422316e-09, -9.262501e-09, -8.989632e-09, -8.637051e-09, -8.263917e-09,
  -8.273863e-09, -8.738654e-09, -9.261615e-09, -9.756029e-09, -1.013656e-08, 
    -1.044574e-08, -1.07356e-08, -1.101998e-08, -1.125946e-08, -1.145908e-08, 
    -1.165751e-08, -1.188416e-08, -1.208184e-08, -1.225619e-08, -1.239428e-08,
  -7.031125e-09, -7.525243e-09, -8.009709e-09, -8.468498e-09, -8.876209e-09, 
    -9.241601e-09, -9.545723e-09, -9.803335e-09, -1.004097e-08, 
    -1.024179e-08, -1.040704e-08, -1.057164e-08, -1.071821e-08, -1.08557e-08, 
    -1.095484e-08,
  -6.105954e-09, -6.535435e-09, -6.950639e-09, -7.335226e-09, -7.713898e-09, 
    -8.062097e-09, -8.393248e-09, -8.662076e-09, -8.8992e-09, -9.103084e-09, 
    -9.275903e-09, -9.427032e-09, -9.548642e-09, -9.641463e-09, -9.688759e-09,
  -5.221806e-09, -5.629641e-09, -5.99563e-09, -6.325124e-09, -6.635178e-09, 
    -6.940421e-09, -7.238854e-09, -7.511299e-09, -7.74563e-09, -7.95901e-09, 
    -8.140834e-09, -8.294601e-09, -8.409481e-09, -8.479636e-09, -8.501772e-09,
  -4.50614e-09, -4.843215e-09, -5.149096e-09, -5.430898e-09, -5.691914e-09, 
    -5.942615e-09, -6.183909e-09, -6.427631e-09, -6.647356e-09, 
    -6.845225e-09, -7.011659e-09, -7.152793e-09, -7.253906e-09, -7.32244e-09, 
    -7.357498e-09,
  -3.982997e-09, -4.204746e-09, -4.452515e-09, -4.681598e-09, -4.89244e-09, 
    -5.070851e-09, -5.261333e-09, -5.44708e-09, -5.629966e-09, -5.791394e-09, 
    -5.940104e-09, -6.061937e-09, -6.150074e-09, -6.221766e-09, -6.282635e-09,
  -3.597425e-09, -3.780177e-09, -3.952088e-09, -4.144495e-09, -4.299987e-09, 
    -4.436154e-09, -4.562012e-09, -4.687864e-09, -4.812176e-09, 
    -4.942623e-09, -5.060979e-09, -5.161096e-09, -5.243215e-09, 
    -5.325271e-09, -5.391208e-09,
  -3.425602e-09, -3.539591e-09, -3.652491e-09, -3.745113e-09, -3.843208e-09, 
    -3.936959e-09, -4.019994e-09, -4.091128e-09, -4.157875e-09, 
    -4.240539e-09, -4.326667e-09, -4.419416e-09, -4.535266e-09, 
    -4.683725e-09, -4.858335e-09,
  -3.362666e-09, -3.466492e-09, -3.515032e-09, -3.587717e-09, -3.630307e-09, 
    -3.673929e-09, -3.717193e-09, -3.743833e-09, -3.792584e-09, 
    -3.880786e-09, -4.0097e-09, -4.172207e-09, -4.383983e-09, -4.653674e-09, 
    -4.966179e-09,
  -3.311959e-09, -3.399343e-09, -3.438383e-09, -3.481504e-09, -3.504207e-09, 
    -3.499629e-09, -3.631478e-09, -3.648491e-09, -3.682968e-09, -3.82303e-09, 
    -4.031932e-09, -4.300689e-09, -4.625949e-09, -4.994903e-09, -5.393299e-09,
  -5.107629e-09, -6.231999e-09, -7.675587e-09, -9.314404e-09, -1.108565e-08, 
    -1.289145e-08, -1.507731e-08, -1.695886e-08, -1.863052e-08, 
    -2.016267e-08, -2.047536e-08, -1.998338e-08, -1.998139e-08, 
    -2.022676e-08, -2.076006e-08,
  -4.341068e-09, -5.206162e-09, -6.440342e-09, -7.833984e-09, -9.581112e-09, 
    -1.122834e-08, -1.317544e-08, -1.493184e-08, -1.673704e-08, 
    -1.813603e-08, -1.960987e-08, -2.043124e-08, -2.014706e-08, 
    -1.980873e-08, -1.997316e-08,
  -3.77214e-09, -4.424404e-09, -5.293899e-09, -6.405228e-09, -7.964967e-09, 
    -9.593465e-09, -1.147506e-08, -1.32195e-08, -1.504753e-08, -1.652188e-08, 
    -1.788511e-08, -1.919255e-08, -2.017876e-08, -2.011295e-08, -1.978449e-08,
  -3.516449e-09, -3.920897e-09, -4.563095e-09, -5.337935e-09, -6.503901e-09, 
    -7.94576e-09, -9.697549e-09, -1.148612e-08, -1.326909e-08, -1.500173e-08, 
    -1.639045e-08, -1.771e-08, -1.89102e-08, -1.984239e-08, -1.999498e-08,
  -3.322238e-09, -3.569131e-09, -4.032073e-09, -4.611246e-09, -5.400883e-09, 
    -6.509771e-09, -7.966343e-09, -9.702015e-09, -1.140283e-08, 
    -1.311213e-08, -1.478609e-08, -1.6117e-08, -1.735195e-08, -1.860938e-08, 
    -1.945132e-08,
  -3.190826e-09, -3.364444e-09, -3.653417e-09, -4.080884e-09, -4.617726e-09, 
    -5.385604e-09, -6.424872e-09, -7.903833e-09, -9.579447e-09, 
    -1.122261e-08, -1.278505e-08, -1.446313e-08, -1.566689e-08, 
    -1.676543e-08, -1.783167e-08,
  -2.872279e-09, -3.165817e-09, -3.391734e-09, -3.732804e-09, -4.137378e-09, 
    -4.640121e-09, -5.324372e-09, -6.291315e-09, -7.658228e-09, 
    -9.215635e-09, -1.073516e-08, -1.224393e-08, -1.386883e-08, 
    -1.508907e-08, -1.602737e-08,
  -2.656735e-09, -2.870611e-09, -3.113444e-09, -3.384539e-09, -3.740829e-09, 
    -4.148704e-09, -4.641746e-09, -5.278761e-09, -6.176062e-09, -7.37825e-09, 
    -8.758161e-09, -1.005901e-08, -1.142654e-08, -1.296831e-08, -1.420411e-08,
  -2.630147e-09, -2.628715e-09, -2.825065e-09, -3.106756e-09, -3.401201e-09, 
    -3.724846e-09, -4.089527e-09, -4.549237e-09, -5.120663e-09, -5.9221e-09, 
    -6.995466e-09, -8.170583e-09, -9.246233e-09, -1.041403e-08, -1.178766e-08,
  -2.631805e-09, -2.575344e-09, -2.576147e-09, -2.756616e-09, -3.036523e-09, 
    -3.381781e-09, -3.691266e-09, -4.025239e-09, -4.404461e-09, 
    -4.889241e-09, -5.563375e-09, -6.452884e-09, -7.424012e-09, 
    -8.291141e-09, -9.269153e-09,
  -5.374817e-09, -6.175738e-09, -7.042209e-09, -7.82472e-09, -8.713558e-09, 
    -9.714308e-09, -1.056708e-08, -1.174477e-08, -1.27564e-08, -1.341631e-08, 
    -1.39824e-08, -1.415494e-08, -1.438557e-08, -1.472787e-08, -1.52054e-08,
  -4.919751e-09, -5.592929e-09, -6.409667e-09, -7.204782e-09, -7.969078e-09, 
    -8.962136e-09, -9.812275e-09, -1.082788e-08, -1.206364e-08, 
    -1.298982e-08, -1.385719e-08, -1.42711e-08, -1.448218e-08, -1.465279e-08, 
    -1.496852e-08,
  -4.543601e-09, -5.104272e-09, -5.794125e-09, -6.59928e-09, -7.265344e-09, 
    -8.223913e-09, -9.077024e-09, -1.000519e-08, -1.123778e-08, 
    -1.246012e-08, -1.351765e-08, -1.421285e-08, -1.4593e-08, -1.476131e-08, 
    -1.490613e-08,
  -4.284618e-09, -4.719185e-09, -5.302292e-09, -6.020602e-09, -6.717948e-09, 
    -7.495737e-09, -8.409061e-09, -9.201261e-09, -1.03273e-08, -1.16641e-08, 
    -1.311802e-08, -1.403394e-08, -1.467211e-08, -1.492063e-08, -1.506675e-08,
  -4.140798e-09, -4.527479e-09, -4.924034e-09, -5.508934e-09, -6.176105e-09, 
    -6.891863e-09, -7.692474e-09, -8.550434e-09, -9.427011e-09, 
    -1.068349e-08, -1.21833e-08, -1.358827e-08, -1.448892e-08, -1.509356e-08, 
    -1.525519e-08,
  -4.007177e-09, -4.305456e-09, -4.62346e-09, -5.084275e-09, -5.699496e-09, 
    -6.259341e-09, -6.890062e-09, -7.680833e-09, -8.657687e-09, 
    -9.689311e-09, -1.113679e-08, -1.265814e-08, -1.385549e-08, 
    -1.477525e-08, -1.543922e-08,
  -3.869093e-09, -4.029587e-09, -4.309985e-09, -4.634459e-09, -5.1984e-09, 
    -5.731708e-09, -6.193718e-09, -6.846682e-09, -7.71174e-09, -8.847386e-09, 
    -1.011186e-08, -1.16122e-08, -1.304515e-08, -1.432729e-08, -1.514161e-08,
  -3.811528e-09, -3.893432e-09, -4.049916e-09, -4.297304e-09, -4.633583e-09, 
    -5.100194e-09, -5.591836e-09, -6.169966e-09, -6.859528e-09, -7.74144e-09, 
    -9.06478e-09, -1.047163e-08, -1.191555e-08, -1.333265e-08, -1.487113e-08,
  -3.819389e-09, -3.731732e-09, -3.898691e-09, -4.09492e-09, -4.233887e-09, 
    -4.448588e-09, -4.775299e-09, -5.312002e-09, -5.963091e-09, 
    -6.688364e-09, -7.653122e-09, -9.070027e-09, -1.059722e-08, 
    -1.202787e-08, -1.354637e-08,
  -3.787494e-09, -3.703494e-09, -3.664582e-09, -3.78252e-09, -3.902924e-09, 
    -4.020208e-09, -4.164832e-09, -4.36628e-09, -4.861972e-09, -5.534062e-09, 
    -6.318877e-09, -7.467673e-09, -8.921022e-09, -1.048955e-08, -1.199715e-08,
  -2.532278e-09, -2.75693e-09, -3.093992e-09, -3.380403e-09, -3.524709e-09, 
    -3.845082e-09, -4.126357e-09, -4.478728e-09, -4.785017e-09, 
    -5.252798e-09, -5.814735e-09, -6.311601e-09, -6.606874e-09, 
    -6.770851e-09, -6.981169e-09,
  -2.468692e-09, -2.748229e-09, -3.087797e-09, -3.489281e-09, -3.778853e-09, 
    -3.985273e-09, -4.344034e-09, -4.736739e-09, -5.1791e-09, -5.600929e-09, 
    -6.087649e-09, -6.681266e-09, -7.061228e-09, -7.348737e-09, -7.47518e-09,
  -2.611024e-09, -2.769243e-09, -2.978388e-09, -3.295208e-09, -3.591085e-09, 
    -3.846484e-09, -4.226776e-09, -4.656653e-09, -5.167585e-09, -5.68048e-09, 
    -6.086879e-09, -6.611934e-09, -7.146314e-09, -7.541747e-09, -7.759276e-09,
  -2.52487e-09, -2.623881e-09, -2.810624e-09, -3.159454e-09, -3.499158e-09, 
    -3.798216e-09, -4.153551e-09, -4.570099e-09, -5.039316e-09, 
    -5.537282e-09, -6.031451e-09, -6.437302e-09, -6.945343e-09, 
    -7.480629e-09, -7.828022e-09,
  -2.462538e-09, -2.606681e-09, -2.77641e-09, -3.168765e-09, -3.55585e-09, 
    -3.865257e-09, -4.275885e-09, -4.727416e-09, -5.176066e-09, 
    -5.600614e-09, -5.997513e-09, -6.360068e-09, -6.831923e-09, 
    -7.388968e-09, -7.860102e-09,
  -2.422718e-09, -2.696231e-09, -2.928401e-09, -3.238718e-09, -3.688057e-09, 
    -4.127173e-09, -4.604086e-09, -5.087124e-09, -5.528791e-09, 
    -5.909497e-09, -6.35096e-09, -6.663026e-09, -7.084363e-09, -7.612449e-09, 
    -8.074543e-09,
  -2.441644e-09, -2.738349e-09, -3.100174e-09, -3.569548e-09, -4.010186e-09, 
    -4.55059e-09, -5.111577e-09, -5.569105e-09, -6.159471e-09, -6.673482e-09, 
    -7.09357e-09, -7.413156e-09, -7.73557e-09, -8.157357e-09, -8.56506e-09,
  -2.652113e-09, -2.986734e-09, -3.329348e-09, -3.864875e-09, -4.525153e-09, 
    -5.078147e-09, -5.569612e-09, -6.216345e-09, -6.829297e-09, 
    -7.464343e-09, -8.163423e-09, -8.568695e-09, -8.970283e-09, 
    -9.314957e-09, -9.548992e-09,
  -2.830461e-09, -3.188596e-09, -3.697537e-09, -4.251641e-09, -4.800063e-09, 
    -5.453422e-09, -6.290806e-09, -6.930792e-09, -7.838204e-09, 
    -8.582488e-09, -9.273486e-09, -9.704942e-09, -1.013668e-08, 
    -1.047992e-08, -1.069406e-08,
  -2.954766e-09, -3.224396e-09, -3.821356e-09, -4.484213e-09, -5.243175e-09, 
    -6.171472e-09, -6.917015e-09, -7.910558e-09, -8.611301e-09, 
    -9.319159e-09, -9.954828e-09, -1.053682e-08, -1.13459e-08, -1.183601e-08, 
    -1.227523e-08,
  -7.496547e-09, -7.498459e-09, -7.587196e-09, -7.665747e-09, -7.778825e-09, 
    -7.874228e-09, -7.906809e-09, -8.030526e-09, -8.22849e-09, -8.351709e-09, 
    -8.380519e-09, -8.314557e-09, -8.146354e-09, -7.9289e-09, -7.926648e-09,
  -7.252925e-09, -7.198287e-09, -7.216941e-09, -7.174103e-09, -7.112713e-09, 
    -7.082878e-09, -7.038996e-09, -7.074602e-09, -7.152455e-09, 
    -7.223956e-09, -7.168765e-09, -7.098456e-09, -6.949146e-09, 
    -6.804014e-09, -6.713812e-09,
  -7.163842e-09, -7.058194e-09, -6.922562e-09, -6.787575e-09, -6.684005e-09, 
    -6.598105e-09, -6.588269e-09, -6.587554e-09, -6.61261e-09, -6.611224e-09, 
    -6.494973e-09, -6.288009e-09, -6.040807e-09, -5.814385e-09, -5.665785e-09,
  -7.117336e-09, -6.973762e-09, -6.837721e-09, -6.655458e-09, -6.472911e-09, 
    -6.337622e-09, -6.288344e-09, -6.164233e-09, -6.11114e-09, -6.047691e-09, 
    -5.918193e-09, -5.741233e-09, -5.561063e-09, -5.375311e-09, -5.201768e-09,
  -7.148568e-09, -6.997647e-09, -6.793197e-09, -6.572025e-09, -6.375102e-09, 
    -6.187276e-09, -6.13054e-09, -6.054093e-09, -5.944554e-09, -5.746104e-09, 
    -5.50163e-09, -5.276122e-09, -5.074705e-09, -4.907983e-09, -4.77129e-09,
  -7.208503e-09, -6.98659e-09, -6.771221e-09, -6.495615e-09, -6.284691e-09, 
    -6.137497e-09, -5.946962e-09, -5.800822e-09, -5.572625e-09, 
    -5.286612e-09, -5.0336e-09, -4.780378e-09, -4.588002e-09, -4.393022e-09, 
    -4.246069e-09,
  -7.253663e-09, -6.970197e-09, -6.702887e-09, -6.446927e-09, -6.217175e-09, 
    -5.936614e-09, -5.724284e-09, -5.419747e-09, -5.105268e-09, 
    -4.792865e-09, -4.544494e-09, -4.281145e-09, -4.043445e-09, 
    -3.852901e-09, -3.69054e-09,
  -7.22506e-09, -6.927037e-09, -6.60974e-09, -6.268134e-09, -5.974487e-09, 
    -5.623877e-09, -5.287859e-09, -4.909992e-09, -4.557197e-09, 
    -4.172056e-09, -3.997916e-09, -3.822394e-09, -3.768137e-09, 
    -3.795242e-09, -3.907259e-09,
  -7.107878e-09, -6.873945e-09, -6.510331e-09, -6.153111e-09, -5.673787e-09, 
    -5.196512e-09, -4.729897e-09, -4.27072e-09, -3.831009e-09, -3.622151e-09, 
    -3.573564e-09, -3.612906e-09, -3.740845e-09, -3.942606e-09, -4.257859e-09,
  -6.844392e-09, -6.488162e-09, -6.194073e-09, -5.831443e-09, -5.172431e-09, 
    -4.655352e-09, -4.001004e-09, -3.619981e-09, -3.453956e-09, 
    -3.576046e-09, -4.012433e-09, -4.705608e-09, -5.295161e-09, 
    -5.902636e-09, -6.126095e-09,
  -3.763285e-09, -3.90571e-09, -4.085818e-09, -4.253626e-09, -4.315897e-09, 
    -4.343274e-09, -4.370776e-09, -4.404274e-09, -4.449074e-09, 
    -4.616692e-09, -5.048814e-09, -5.447283e-09, -5.741367e-09, 
    -6.062745e-09, -6.422431e-09,
  -3.800419e-09, -3.84843e-09, -3.932098e-09, -4.12067e-09, -4.321305e-09, 
    -4.458379e-09, -4.479856e-09, -4.593511e-09, -4.841229e-09, 
    -5.184414e-09, -5.587558e-09, -5.975993e-09, -6.342023e-09, 
    -6.635921e-09, -6.920155e-09,
  -3.721776e-09, -3.614014e-09, -3.584252e-09, -3.773303e-09, -4.125613e-09, 
    -4.403295e-09, -4.577617e-09, -4.727537e-09, -4.95864e-09, -5.352767e-09, 
    -5.88095e-09, -6.363094e-09, -6.805864e-09, -7.112937e-09, -7.417754e-09,
  -3.420997e-09, -3.414252e-09, -3.438716e-09, -3.551603e-09, -3.900951e-09, 
    -4.310345e-09, -4.646765e-09, -4.844905e-09, -5.086419e-09, 
    -5.474301e-09, -6.008572e-09, -6.569039e-09, -7.140836e-09, 
    -7.510454e-09, -7.798225e-09,
  -3.396199e-09, -3.627207e-09, -3.775681e-09, -3.863495e-09, -4.064004e-09, 
    -4.397174e-09, -4.781104e-09, -4.985601e-09, -5.1981e-09, -5.580747e-09, 
    -6.149524e-09, -6.681842e-09, -7.21153e-09, -7.586734e-09, -7.835697e-09,
  -3.27671e-09, -3.651005e-09, -3.847247e-09, -4.015287e-09, -4.316843e-09, 
    -4.662466e-09, -5.098438e-09, -5.394823e-09, -5.637941e-09, 
    -5.929445e-09, -6.392576e-09, -6.883829e-09, -7.429305e-09, 
    -7.874054e-09, -8.196333e-09,
  -3.738314e-09, -4.145576e-09, -4.248435e-09, -4.420953e-09, -4.637708e-09, 
    -4.9728e-09, -5.411864e-09, -5.735203e-09, -6.017859e-09, -6.420102e-09, 
    -6.915347e-09, -7.400203e-09, -7.943632e-09, -8.400311e-09, -8.733804e-09,
  -5.074264e-09, -5.358644e-09, -5.512761e-09, -5.797312e-09, -6.131296e-09, 
    -6.263503e-09, -6.475704e-09, -6.583203e-09, -6.831715e-09, 
    -7.211711e-09, -7.668613e-09, -8.113491e-09, -8.571337e-09, 
    -8.869639e-09, -9.075988e-09,
  -5.673826e-09, -6.047909e-09, -6.408651e-09, -6.804615e-09, -7.15706e-09, 
    -7.423433e-09, -7.72854e-09, -7.908442e-09, -8.162041e-09, -8.381632e-09, 
    -8.67228e-09, -8.880074e-09, -9.019472e-09, -9.046586e-09, -9.077365e-09,
  -6.862312e-09, -7.31771e-09, -7.697937e-09, -8.10296e-09, -8.465341e-09, 
    -8.921658e-09, -8.996964e-09, -9.08878e-09, -9.057501e-09, -9.083238e-09, 
    -8.963866e-09, -8.88857e-09, -8.875236e-09, -8.906327e-09, -8.872846e-09,
  -6.458603e-09, -6.340219e-09, -6.225094e-09, -6.053947e-09, -5.81276e-09, 
    -5.470699e-09, -5.111894e-09, -4.727085e-09, -4.368644e-09, 
    -4.042778e-09, -3.792896e-09, -3.639476e-09, -3.500073e-09, 
    -3.410842e-09, -3.3648e-09,
  -5.928787e-09, -5.919191e-09, -5.869096e-09, -5.644368e-09, -5.305787e-09, 
    -4.947118e-09, -4.58106e-09, -4.272422e-09, -4.04361e-09, -3.856913e-09, 
    -3.690612e-09, -3.531917e-09, -3.370215e-09, -3.238971e-09, -3.117592e-09,
  -5.644712e-09, -5.628535e-09, -5.448003e-09, -5.084924e-09, -4.798645e-09, 
    -4.525753e-09, -4.312311e-09, -4.162468e-09, -4.046029e-09, 
    -3.910921e-09, -3.777345e-09, -3.653774e-09, -3.517198e-09, 
    -3.384615e-09, -3.235096e-09,
  -5.164477e-09, -5.143655e-09, -4.946578e-09, -4.715712e-09, -4.571061e-09, 
    -4.452484e-09, -4.402123e-09, -4.344499e-09, -4.290376e-09, 
    -4.232734e-09, -4.203534e-09, -4.172568e-09, -4.137869e-09, 
    -4.051417e-09, -3.932264e-09,
  -4.91051e-09, -4.910002e-09, -4.810647e-09, -4.625919e-09, -4.482764e-09, 
    -4.438138e-09, -4.404349e-09, -4.380905e-09, -4.423283e-09, 
    -4.503645e-09, -4.640583e-09, -4.773196e-09, -4.848179e-09, 
    -4.884907e-09, -4.829247e-09,
  -4.790563e-09, -4.893326e-09, -4.841545e-09, -4.78212e-09, -4.680011e-09, 
    -4.536955e-09, -4.43868e-09, -4.409529e-09, -4.527893e-09, -4.65421e-09, 
    -4.890558e-09, -5.076465e-09, -5.311309e-09, -5.538116e-09, -5.710485e-09,
  -5.015952e-09, -5.107191e-09, -5.102672e-09, -5.144111e-09, -4.968796e-09, 
    -4.847923e-09, -4.601744e-09, -4.627682e-09, -4.657358e-09, 
    -4.738198e-09, -5.005091e-09, -5.243884e-09, -5.501576e-09, 
    -5.646527e-09, -5.786197e-09,
  -5.735056e-09, -5.960381e-09, -5.829007e-09, -5.901938e-09, -5.659279e-09, 
    -5.692782e-09, -5.625068e-09, -5.329805e-09, -5.373603e-09, 
    -5.288582e-09, -5.203898e-09, -5.237979e-09, -5.484122e-09, 
    -5.719148e-09, -5.843754e-09,
  -6.261469e-09, -6.675287e-09, -6.816947e-09, -7.250126e-09, -7.492228e-09, 
    -7.203557e-09, -7.102961e-09, -6.867038e-09, -6.747074e-09, 
    -6.715706e-09, -6.799892e-09, -6.710559e-09, -6.643024e-09, 
    -6.650382e-09, -6.734327e-09,
  -6.136398e-09, -6.897419e-09, -7.51251e-09, -8.327968e-09, -9.00515e-09, 
    -9.229189e-09, -9.079537e-09, -8.995339e-09, -8.731463e-09, 
    -8.448639e-09, -7.985814e-09, -7.829142e-09, -7.725891e-09, 
    -7.725111e-09, -7.881146e-09,
  -1.239573e-08, -1.270042e-08, -1.302056e-08, -1.322006e-08, -1.349715e-08, 
    -1.375965e-08, -1.398836e-08, -1.414204e-08, -1.425456e-08, 
    -1.429222e-08, -1.430018e-08, -1.42456e-08, -1.420126e-08, -1.418234e-08, 
    -1.423258e-08,
  -1.143221e-08, -1.163419e-08, -1.190559e-08, -1.22836e-08, -1.266366e-08, 
    -1.295082e-08, -1.321346e-08, -1.333133e-08, -1.33069e-08, -1.319992e-08, 
    -1.308335e-08, -1.298501e-08, -1.289487e-08, -1.28237e-08, -1.275752e-08,
  -1.077126e-08, -1.091013e-08, -1.112077e-08, -1.156627e-08, -1.193023e-08, 
    -1.221901e-08, -1.235025e-08, -1.235236e-08, -1.225802e-08, 
    -1.213136e-08, -1.198036e-08, -1.185922e-08, -1.173802e-08, 
    -1.165178e-08, -1.153298e-08,
  -9.855217e-09, -1.00674e-08, -1.043706e-08, -1.090917e-08, -1.129502e-08, 
    -1.148208e-08, -1.15222e-08, -1.144632e-08, -1.136907e-08, -1.124575e-08, 
    -1.110905e-08, -1.096095e-08, -1.080566e-08, -1.063905e-08, -1.048412e-08,
  -9.138231e-09, -9.379325e-09, -9.706945e-09, -1.016394e-08, -1.054518e-08, 
    -1.073472e-08, -1.076759e-08, -1.071297e-08, -1.063046e-08, 
    -1.048646e-08, -1.029251e-08, -1.00851e-08, -9.8518e-09, -9.59487e-09, 
    -9.334395e-09,
  -8.400644e-09, -8.724616e-09, -9.083338e-09, -9.478422e-09, -9.810014e-09, 
    -1.002266e-08, -1.013847e-08, -1.009178e-08, -9.949956e-09, -9.72515e-09, 
    -9.445886e-09, -9.145704e-09, -8.811075e-09, -8.456321e-09, -8.148929e-09,
  -7.724918e-09, -8.144646e-09, -8.500022e-09, -8.90059e-09, -9.268428e-09, 
    -9.471929e-09, -9.444427e-09, -9.31122e-09, -9.097104e-09, -8.845548e-09, 
    -8.531862e-09, -8.171727e-09, -7.849392e-09, -7.505325e-09, -7.232048e-09,
  -7.208939e-09, -7.698559e-09, -8.021223e-09, -8.489987e-09, -8.780695e-09, 
    -8.909927e-09, -8.834236e-09, -8.712773e-09, -8.4748e-09, -8.120455e-09, 
    -7.739425e-09, -7.28853e-09, -6.911111e-09, -6.645409e-09, -6.459391e-09,
  -6.819418e-09, -7.320569e-09, -7.777116e-09, -8.165225e-09, -8.325085e-09, 
    -8.293944e-09, -8.295936e-09, -8.113276e-09, -7.945251e-09, 
    -7.643468e-09, -7.422171e-09, -7.199775e-09, -6.940113e-09, 
    -6.696101e-09, -6.50824e-09,
  -6.67121e-09, -7.244817e-09, -7.645417e-09, -7.807412e-09, -7.998401e-09, 
    -8.109435e-09, -7.822112e-09, -7.723329e-09, -7.501254e-09, 
    -7.298668e-09, -7.049948e-09, -6.892523e-09, -6.856586e-09, 
    -6.807416e-09, -6.866367e-09,
  -9.530105e-09, -1.032002e-08, -1.130136e-08, -1.192888e-08, -1.241449e-08, 
    -1.255725e-08, -1.174616e-08, -1.186496e-08, -1.29937e-08, -1.430211e-08, 
    -1.556965e-08, -1.702968e-08, -1.798854e-08, -1.860737e-08, -1.936262e-08,
  -8.882445e-09, -9.689543e-09, -1.049877e-08, -1.133426e-08, -1.183802e-08, 
    -1.228664e-08, -1.241328e-08, -1.194416e-08, -1.22864e-08, -1.316932e-08, 
    -1.425826e-08, -1.548462e-08, -1.655651e-08, -1.777415e-08, -1.830321e-08,
  -7.980542e-09, -9.008177e-09, -9.977734e-09, -1.070989e-08, -1.129146e-08, 
    -1.168738e-08, -1.204163e-08, -1.213719e-08, -1.212505e-08, 
    -1.253233e-08, -1.324737e-08, -1.434777e-08, -1.521812e-08, 
    -1.640985e-08, -1.765006e-08,
  -7.37544e-09, -8.176465e-09, -9.296283e-09, -1.024831e-08, -1.077529e-08, 
    -1.122531e-08, -1.150786e-08, -1.198089e-08, -1.212675e-08, -1.22686e-08, 
    -1.266817e-08, -1.354938e-08, -1.440005e-08, -1.512418e-08, -1.639916e-08,
  -7.114783e-09, -7.602878e-09, -8.453923e-09, -9.571091e-09, -1.029827e-08, 
    -1.07703e-08, -1.102087e-08, -1.143884e-08, -1.18461e-08, -1.202898e-08, 
    -1.21442e-08, -1.272043e-08, -1.366685e-08, -1.438811e-08, -1.524127e-08,
  -6.820555e-09, -7.343709e-09, -7.873471e-09, -8.875759e-09, -9.790212e-09, 
    -1.040811e-08, -1.070491e-08, -1.101988e-08, -1.143601e-08, 
    -1.185805e-08, -1.207357e-08, -1.248304e-08, -1.322122e-08, 
    -1.402176e-08, -1.472315e-08,
  -6.357285e-09, -7.002107e-09, -7.518714e-09, -8.325895e-09, -9.314577e-09, 
    -1.002786e-08, -1.042192e-08, -1.067704e-08, -1.105975e-08, 
    -1.154503e-08, -1.1973e-08, -1.245161e-08, -1.299709e-08, -1.364156e-08, 
    -1.417697e-08,
  -5.850041e-09, -6.715628e-09, -7.238298e-09, -8.07311e-09, -9.077048e-09, 
    -9.888409e-09, -1.03542e-08, -1.064449e-08, -1.090065e-08, -1.14175e-08, 
    -1.198225e-08, -1.249156e-08, -1.288636e-08, -1.332442e-08, -1.373634e-08,
  -5.392726e-09, -6.43742e-09, -7.20024e-09, -7.976237e-09, -8.932182e-09, 
    -9.696175e-09, -1.032301e-08, -1.072693e-08, -1.103514e-08, 
    -1.145468e-08, -1.20535e-08, -1.25096e-08, -1.27169e-08, -1.297067e-08, 
    -1.329521e-08,
  -5.000285e-09, -6.161074e-09, -7.184872e-09, -8.122452e-09, -9.12524e-09, 
    -9.935927e-09, -1.031349e-08, -1.079222e-08, -1.119299e-08, 
    -1.156866e-08, -1.192424e-08, -1.229145e-08, -1.252788e-08, 
    -1.268885e-08, -1.281474e-08,
  -9.447945e-09, -9.633213e-09, -9.589009e-09, -9.626081e-09, -9.863832e-09, 
    -9.93759e-09, -1.012234e-08, -1.051157e-08, -1.100298e-08, -1.153584e-08, 
    -1.200414e-08, -1.248858e-08, -1.404528e-08, -1.550728e-08, -1.557216e-08,
  -9.278777e-09, -9.48445e-09, -9.551618e-09, -9.559354e-09, -9.698374e-09, 
    -9.850296e-09, -9.876674e-09, -1.010972e-08, -1.045958e-08, 
    -1.090396e-08, -1.145481e-08, -1.19794e-08, -1.25825e-08, -1.399871e-08, 
    -1.500721e-08,
  -9.137562e-09, -9.234098e-09, -9.381552e-09, -9.432064e-09, -9.542469e-09, 
    -9.75789e-09, -9.862467e-09, -9.865158e-09, -1.005374e-08, -1.044671e-08, 
    -1.081381e-08, -1.138566e-08, -1.179992e-08, -1.255073e-08, -1.380905e-08,
  -8.496568e-09, -8.826428e-09, -9.064839e-09, -9.247596e-09, -9.408568e-09, 
    -9.647357e-09, -9.832519e-09, -9.876965e-09, -9.750479e-09, 
    -1.025556e-08, -1.062623e-08, -1.094776e-08, -1.134426e-08, 
    -1.168064e-08, -1.268732e-08,
  -7.794576e-09, -8.111948e-09, -8.493806e-09, -8.921627e-09, -9.188451e-09, 
    -9.544087e-09, -9.75307e-09, -9.879692e-09, -9.753855e-09, -9.922966e-09, 
    -1.050074e-08, -1.08592e-08, -1.118617e-08, -1.13499e-08, -1.185652e-08,
  -7.07415e-09, -7.409221e-09, -7.765159e-09, -8.320504e-09, -8.81013e-09, 
    -9.313937e-09, -9.700607e-09, -9.887332e-09, -9.893857e-09, 
    -9.832646e-09, -1.016281e-08, -1.044124e-08, -1.083288e-08, 
    -1.122157e-08, -1.139176e-08,
  -6.429187e-09, -6.801628e-09, -7.125422e-09, -7.625859e-09, -8.197318e-09, 
    -8.847823e-09, -9.442307e-09, -9.753963e-09, -9.933302e-09, 
    -9.842997e-09, -9.961056e-09, -1.005059e-08, -1.030204e-08, 
    -1.072432e-08, -1.1195e-08,
  -5.88872e-09, -6.207036e-09, -6.549537e-09, -6.982483e-09, -7.568009e-09, 
    -8.274048e-09, -9.118112e-09, -9.516102e-09, -9.920713e-09, 
    -9.911417e-09, -9.914186e-09, -9.889559e-09, -9.859458e-09, 
    -1.023697e-08, -1.059235e-08,
  -5.23498e-09, -5.569805e-09, -5.981501e-09, -6.366346e-09, -6.904328e-09, 
    -7.496726e-09, -8.405292e-09, -9.123502e-09, -9.555277e-09, 
    -9.744237e-09, -9.815325e-09, -1.002422e-08, -9.937906e-09, 
    -9.911481e-09, -1.017879e-08,
  -4.579653e-09, -4.976768e-09, -5.334528e-09, -5.796157e-09, -6.350055e-09, 
    -7.024405e-09, -7.751349e-09, -8.607143e-09, -9.290819e-09, 
    -9.510047e-09, -9.577781e-09, -9.797969e-09, -9.976157e-09, -9.89008e-09, 
    -9.929638e-09,
  -1.084265e-08, -1.10316e-08, -1.090862e-08, -1.074087e-08, -1.058738e-08, 
    -1.039903e-08, -1.044948e-08, -1.06597e-08, -1.092534e-08, -1.099198e-08, 
    -1.124919e-08, -1.13929e-08, -1.140205e-08, -1.203937e-08, -1.330943e-08,
  -1.11655e-08, -1.141323e-08, -1.128908e-08, -1.105024e-08, -1.082585e-08, 
    -1.055389e-08, -1.03811e-08, -1.03086e-08, -1.038473e-08, -1.047674e-08, 
    -1.067713e-08, -1.104729e-08, -1.125558e-08, -1.144876e-08, -1.278281e-08,
  -1.107697e-08, -1.123222e-08, -1.120792e-08, -1.109147e-08, -1.091071e-08, 
    -1.068884e-08, -1.05242e-08, -1.030636e-08, -1.021595e-08, -1.024175e-08, 
    -1.026941e-08, -1.051338e-08, -1.087284e-08, -1.102547e-08, -1.201354e-08,
  -1.087534e-08, -1.095721e-08, -1.094295e-08, -1.088976e-08, -1.073071e-08, 
    -1.062209e-08, -1.05486e-08, -1.044488e-08, -1.024225e-08, -1.019885e-08, 
    -1.016108e-08, -1.01473e-08, -1.039383e-08, -1.058914e-08, -1.1096e-08,
  -1.050009e-08, -1.051362e-08, -1.0534e-08, -1.059021e-08, -1.055888e-08, 
    -1.053622e-08, -1.052503e-08, -1.045484e-08, -1.028706e-08, 
    -1.020496e-08, -1.013567e-08, -1.001823e-08, -1.00683e-08, -1.024552e-08, 
    -1.043284e-08,
  -1.021859e-08, -1.013988e-08, -1.014442e-08, -1.020013e-08, -1.029692e-08, 
    -1.044465e-08, -1.0435e-08, -1.048095e-08, -1.031712e-08, -1.023501e-08, 
    -1.009064e-08, -1.000918e-08, -9.879815e-09, -1.005783e-08, -1.011151e-08,
  -9.978919e-09, -9.925481e-09, -9.875488e-09, -9.912251e-09, -9.973685e-09, 
    -1.017605e-08, -1.027534e-08, -1.037816e-08, -1.040203e-08, 
    -1.038338e-08, -1.039729e-08, -1.021832e-08, -9.928585e-09, 
    -9.795769e-09, -9.99018e-09,
  -9.553375e-09, -9.535794e-09, -9.533351e-09, -9.586856e-09, -9.659801e-09, 
    -9.757112e-09, -9.904245e-09, -1.007866e-08, -1.027782e-08, 
    -1.033661e-08, -1.056653e-08, -1.046885e-08, -1.044291e-08, 
    -1.011132e-08, -1.005973e-08,
  -9.032979e-09, -9.05784e-09, -9.132767e-09, -9.182216e-09, -9.275592e-09, 
    -9.294355e-09, -9.36836e-09, -9.493426e-09, -9.849487e-09, -1.007589e-08, 
    -1.036803e-08, -1.045611e-08, -1.049156e-08, -1.031187e-08, -1.015117e-08,
  -8.428583e-09, -8.528183e-09, -8.647115e-09, -8.736466e-09, -8.811118e-09, 
    -8.90793e-09, -8.947048e-09, -9.013404e-09, -9.253835e-09, -9.571811e-09, 
    -1.000094e-08, -1.031881e-08, -1.045881e-08, -1.045227e-08, -1.01764e-08,
  -1.201982e-08, -1.221816e-08, -1.280908e-08, -1.288936e-08, -1.351865e-08, 
    -1.435657e-08, -1.520169e-08, -1.575361e-08, -1.577588e-08, 
    -1.547384e-08, -1.539298e-08, -1.531855e-08, -1.539247e-08, 
    -1.564303e-08, -1.599197e-08,
  -1.13757e-08, -1.170513e-08, -1.19541e-08, -1.223792e-08, -1.235473e-08, 
    -1.266935e-08, -1.321822e-08, -1.403393e-08, -1.497033e-08, -1.54278e-08, 
    -1.535123e-08, -1.51064e-08, -1.505033e-08, -1.507134e-08, -1.50991e-08,
  -1.078997e-08, -1.111202e-08, -1.138805e-08, -1.158965e-08, -1.173732e-08, 
    -1.192859e-08, -1.215643e-08, -1.256015e-08, -1.323847e-08, 
    -1.408517e-08, -1.496195e-08, -1.527431e-08, -1.512048e-08, -1.48937e-08, 
    -1.474478e-08,
  -1.064145e-08, -1.08046e-08, -1.118736e-08, -1.135535e-08, -1.134482e-08, 
    -1.126757e-08, -1.127185e-08, -1.143749e-08, -1.186339e-08, 
    -1.241446e-08, -1.321889e-08, -1.418762e-08, -1.499188e-08, 
    -1.525506e-08, -1.507722e-08,
  -1.020574e-08, -1.049344e-08, -1.070789e-08, -1.115082e-08, -1.146747e-08, 
    -1.147065e-08, -1.11948e-08, -1.097099e-08, -1.096597e-08, -1.132072e-08, 
    -1.176921e-08, -1.235476e-08, -1.313424e-08, -1.3937e-08, -1.46662e-08,
  -9.889274e-09, -9.837465e-09, -1.003727e-08, -1.03224e-08, -1.075123e-08, 
    -1.103008e-08, -1.112477e-08, -1.110679e-08, -1.093905e-08, 
    -1.096465e-08, -1.107646e-08, -1.139994e-08, -1.192995e-08, 
    -1.239423e-08, -1.304695e-08,
  -9.965631e-09, -9.779187e-09, -9.691588e-09, -9.764452e-09, -9.993698e-09, 
    -1.031766e-08, -1.052717e-08, -1.065327e-08, -1.073489e-08, -1.07073e-08, 
    -1.076211e-08, -1.088092e-08, -1.111767e-08, -1.147207e-08, -1.194819e-08,
  -1.00229e-08, -9.933975e-09, -9.762072e-09, -9.581189e-09, -9.536491e-09, 
    -9.758025e-09, -1.002007e-08, -1.022423e-08, -1.03662e-08, -1.045621e-08, 
    -1.045508e-08, -1.049178e-08, -1.0567e-08, -1.070625e-08, -1.10713e-08,
  -9.670652e-09, -9.835984e-09, -9.828752e-09, -9.728004e-09, -9.537994e-09, 
    -9.500298e-09, -9.697647e-09, -9.94262e-09, -1.010887e-08, -1.02692e-08, 
    -1.031256e-08, -1.032963e-08, -1.041284e-08, -1.045701e-08, -1.05826e-08,
  -8.802624e-09, -9.209425e-09, -9.491271e-09, -9.628287e-09, -9.607334e-09, 
    -9.584885e-09, -9.673271e-09, -9.818242e-09, -9.939089e-09, 
    -1.009213e-08, -1.019943e-08, -1.027335e-08, -1.035622e-08, 
    -1.047489e-08, -1.057562e-08,
  -1.36206e-08, -1.413774e-08, -1.479826e-08, -1.525953e-08, -1.565339e-08, 
    -1.58981e-08, -1.630401e-08, -1.672609e-08, -1.738319e-08, -1.814396e-08, 
    -1.861837e-08, -1.934065e-08, -2.004999e-08, -2.069308e-08, -2.117769e-08,
  -1.316991e-08, -1.35245e-08, -1.392078e-08, -1.443265e-08, -1.496476e-08, 
    -1.53694e-08, -1.58567e-08, -1.626374e-08, -1.656924e-08, -1.707046e-08, 
    -1.765038e-08, -1.807746e-08, -1.867413e-08, -1.92265e-08, -1.986534e-08,
  -1.243934e-08, -1.292155e-08, -1.33776e-08, -1.374968e-08, -1.427089e-08, 
    -1.46799e-08, -1.508821e-08, -1.566764e-08, -1.597792e-08, -1.628702e-08, 
    -1.67827e-08, -1.720709e-08, -1.763541e-08, -1.805452e-08, -1.845467e-08,
  -1.15057e-08, -1.211542e-08, -1.260702e-08, -1.320804e-08, -1.355442e-08, 
    -1.402952e-08, -1.439242e-08, -1.487098e-08, -1.542506e-08, 
    -1.565567e-08, -1.587551e-08, -1.627188e-08, -1.668021e-08, 
    -1.717548e-08, -1.761207e-08,
  -1.080083e-08, -1.127649e-08, -1.184453e-08, -1.247694e-08, -1.30333e-08, 
    -1.34471e-08, -1.388802e-08, -1.422157e-08, -1.469705e-08, -1.518877e-08, 
    -1.536658e-08, -1.551738e-08, -1.577403e-08, -1.609445e-08, -1.652825e-08,
  -9.82496e-09, -1.043156e-08, -1.088074e-08, -1.153593e-08, -1.228594e-08, 
    -1.284612e-08, -1.328634e-08, -1.370878e-08, -1.399644e-08, 
    -1.440973e-08, -1.483882e-08, -1.49573e-08, -1.517084e-08, -1.537636e-08, 
    -1.559379e-08,
  -8.868183e-09, -9.550799e-09, -1.012075e-08, -1.053994e-08, -1.124855e-08, 
    -1.198331e-08, -1.256336e-08, -1.308064e-08, -1.353464e-08, 
    -1.379093e-08, -1.41147e-08, -1.440861e-08, -1.454812e-08, -1.47433e-08, 
    -1.486081e-08,
  -8.480911e-09, -8.863348e-09, -9.41825e-09, -9.904912e-09, -1.028046e-08, 
    -1.095297e-08, -1.163378e-08, -1.221609e-08, -1.278974e-08, 
    -1.327223e-08, -1.356801e-08, -1.386625e-08, -1.405059e-08, 
    -1.410455e-08, -1.424189e-08,
  -8.014328e-09, -8.325213e-09, -8.646487e-09, -9.061919e-09, -9.633049e-09, 
    -1.005111e-08, -1.06678e-08, -1.129196e-08, -1.186116e-08, -1.241441e-08, 
    -1.27739e-08, -1.310605e-08, -1.337536e-08, -1.349858e-08, -1.358205e-08,
  -7.563869e-09, -7.938022e-09, -8.217632e-09, -8.520321e-09, -8.745634e-09, 
    -9.217947e-09, -9.800966e-09, -1.036439e-08, -1.075774e-08, 
    -1.129236e-08, -1.183353e-08, -1.222505e-08, -1.254519e-08, 
    -1.278806e-08, -1.292873e-08,
  -1.188828e-08, -1.20641e-08, -1.294055e-08, -1.368804e-08, -1.462557e-08, 
    -1.478764e-08, -1.532524e-08, -1.538855e-08, -1.586648e-08, 
    -1.677641e-08, -1.75028e-08, -1.814389e-08, -1.862477e-08, -1.927195e-08, 
    -1.994073e-08,
  -1.104012e-08, -1.125048e-08, -1.171516e-08, -1.238044e-08, -1.323877e-08, 
    -1.398188e-08, -1.430092e-08, -1.454918e-08, -1.468642e-08, -1.5125e-08, 
    -1.576936e-08, -1.665564e-08, -1.751641e-08, -1.817206e-08, -1.88631e-08,
  -1.100613e-08, -1.105081e-08, -1.104395e-08, -1.132279e-08, -1.186497e-08, 
    -1.26516e-08, -1.329017e-08, -1.360499e-08, -1.376059e-08, -1.390269e-08, 
    -1.437322e-08, -1.503013e-08, -1.599109e-08, -1.669268e-08, -1.732948e-08,
  -1.173419e-08, -1.142067e-08, -1.124876e-08, -1.107011e-08, -1.111755e-08, 
    -1.138445e-08, -1.198128e-08, -1.245252e-08, -1.269944e-08, 
    -1.287204e-08, -1.320122e-08, -1.363554e-08, -1.435075e-08, -1.51547e-08, 
    -1.584537e-08,
  -1.139456e-08, -1.170512e-08, -1.172365e-08, -1.154606e-08, -1.129544e-08, 
    -1.105119e-08, -1.117124e-08, -1.149962e-08, -1.175345e-08, 
    -1.205826e-08, -1.232493e-08, -1.265992e-08, -1.311414e-08, 
    -1.382103e-08, -1.443982e-08,
  -1.032662e-08, -1.123397e-08, -1.163492e-08, -1.184356e-08, -1.179674e-08, 
    -1.156323e-08, -1.121411e-08, -1.117583e-08, -1.136927e-08, 
    -1.153191e-08, -1.186468e-08, -1.214579e-08, -1.248102e-08, 
    -1.299447e-08, -1.353762e-08,
  -9.48588e-09, -1.01391e-08, -1.101938e-08, -1.150387e-08, -1.18128e-08, 
    -1.192379e-08, -1.185507e-08, -1.152576e-08, -1.145008e-08, 
    -1.155663e-08, -1.171535e-08, -1.201138e-08, -1.223606e-08, -1.25717e-08, 
    -1.301915e-08,
  -8.899399e-09, -9.35767e-09, -9.973273e-09, -1.083729e-08, -1.137571e-08, 
    -1.17654e-08, -1.201191e-08, -1.207761e-08, -1.19179e-08, -1.18018e-08, 
    -1.189119e-08, -1.211409e-08, -1.235243e-08, -1.248002e-08, -1.271021e-08,
  -8.621553e-09, -8.773888e-09, -9.12911e-09, -9.845535e-09, -1.070565e-08, 
    -1.135616e-08, -1.173374e-08, -1.202538e-08, -1.215176e-08, 
    -1.219017e-08, -1.216161e-08, -1.225377e-08, -1.252167e-08, 
    -1.273996e-08, -1.287378e-08,
  -8.154641e-09, -8.544516e-09, -8.691848e-09, -8.950489e-09, -9.55546e-09, 
    -1.058808e-08, -1.135192e-08, -1.18135e-08, -1.210037e-08, -1.216763e-08, 
    -1.238054e-08, -1.24587e-08, -1.255149e-08, -1.280072e-08, -1.298302e-08,
  -1.394335e-08, -1.572744e-08, -1.618161e-08, -1.62107e-08, -1.655217e-08, 
    -1.704455e-08, -1.77841e-08, -1.818513e-08, -1.845823e-08, -1.922968e-08, 
    -1.984549e-08, -2.112918e-08, -2.202193e-08, -2.315452e-08, -2.41062e-08,
  -1.433523e-08, -1.549635e-08, -1.655298e-08, -1.676565e-08, -1.672198e-08, 
    -1.697372e-08, -1.757861e-08, -1.821309e-08, -1.865756e-08, 
    -1.918976e-08, -1.987405e-08, -2.073223e-08, -2.18502e-08, -2.294145e-08, 
    -2.412022e-08,
  -1.342889e-08, -1.427621e-08, -1.593155e-08, -1.717798e-08, -1.746823e-08, 
    -1.729857e-08, -1.749618e-08, -1.814009e-08, -1.874623e-08, 
    -1.926445e-08, -1.976078e-08, -2.05978e-08, -2.160127e-08, -2.283306e-08, 
    -2.404968e-08,
  -1.355366e-08, -1.35779e-08, -1.450703e-08, -1.619047e-08, -1.747878e-08, 
    -1.798326e-08, -1.790422e-08, -1.819286e-08, -1.892924e-08, 
    -1.958285e-08, -1.996912e-08, -2.053432e-08, -2.156005e-08, 
    -2.265784e-08, -2.385264e-08,
  -1.255046e-08, -1.342062e-08, -1.375122e-08, -1.480591e-08, -1.637631e-08, 
    -1.762371e-08, -1.825197e-08, -1.837986e-08, -1.90202e-08, -1.973535e-08, 
    -2.029861e-08, -2.058892e-08, -2.12828e-08, -2.237134e-08, -2.354746e-08,
  -1.111428e-08, -1.262855e-08, -1.343073e-08, -1.395307e-08, -1.508946e-08, 
    -1.637108e-08, -1.753214e-08, -1.829953e-08, -1.875391e-08, 
    -1.966117e-08, -2.027019e-08, -2.068574e-08, -2.101063e-08, 
    -2.176487e-08, -2.278228e-08,
  -1.028739e-08, -1.145247e-08, -1.269586e-08, -1.336957e-08, -1.41466e-08, 
    -1.530905e-08, -1.626823e-08, -1.739269e-08, -1.814727e-08, 
    -1.891905e-08, -2.000928e-08, -2.043062e-08, -2.091732e-08, 
    -2.130462e-08, -2.202884e-08,
  -9.233101e-09, -1.029562e-08, -1.161439e-08, -1.280988e-08, -1.344458e-08, 
    -1.439965e-08, -1.550141e-08, -1.637235e-08, -1.73724e-08, -1.81555e-08, 
    -1.921458e-08, -2.02612e-08, -2.056719e-08, -2.105345e-08, -2.144453e-08,
  -8.092547e-09, -9.109816e-09, -1.02775e-08, -1.176364e-08, -1.295099e-08, 
    -1.355658e-08, -1.452973e-08, -1.55771e-08, -1.655189e-08, -1.737435e-08, 
    -1.833128e-08, -1.943903e-08, -2.040965e-08, -2.084405e-08, -2.118125e-08,
  -7.071971e-09, -8.118984e-09, -9.134127e-09, -1.030952e-08, -1.182322e-08, 
    -1.316184e-08, -1.380312e-08, -1.477444e-08, -1.578196e-08, 
    -1.679149e-08, -1.767451e-08, -1.859713e-08, -1.970234e-08, 
    -2.061508e-08, -2.103678e-08,
  -9.361046e-09, -9.816739e-09, -1.02643e-08, -1.082633e-08, -1.138641e-08, 
    -1.187416e-08, -1.239857e-08, -1.271494e-08, -1.272124e-08, 
    -1.240242e-08, -1.201144e-08, -1.179448e-08, -1.189338e-08, 
    -1.240978e-08, -1.337974e-08,
  -8.741002e-09, -9.237164e-09, -9.687498e-09, -1.011129e-08, -1.047175e-08, 
    -1.098605e-08, -1.145313e-08, -1.193461e-08, -1.230818e-08, 
    -1.246495e-08, -1.237752e-08, -1.210469e-08, -1.18288e-08, -1.184992e-08, 
    -1.207627e-08,
  -8.201537e-09, -8.67972e-09, -9.169851e-09, -9.623328e-09, -9.908452e-09, 
    -1.024896e-08, -1.069869e-08, -1.114685e-08, -1.157999e-08, 
    -1.194896e-08, -1.215263e-08, -1.223607e-08, -1.208461e-08, 
    -1.190111e-08, -1.191092e-08,
  -7.754304e-09, -8.209437e-09, -8.665395e-09, -9.136262e-09, -9.515025e-09, 
    -9.739399e-09, -1.011861e-08, -1.052483e-08, -1.088728e-08, 
    -1.127534e-08, -1.1604e-08, -1.180624e-08, -1.19356e-08, -1.187369e-08, 
    -1.187614e-08,
  -7.478733e-09, -7.786223e-09, -8.263823e-09, -8.709577e-09, -9.151211e-09, 
    -9.463268e-09, -9.763557e-09, -1.007141e-08, -1.035829e-08, 
    -1.060624e-08, -1.09492e-08, -1.120344e-08, -1.140002e-08, -1.158706e-08, 
    -1.160296e-08,
  -7.265218e-09, -7.452092e-09, -7.868099e-09, -8.355436e-09, -8.799231e-09, 
    -9.17444e-09, -9.529273e-09, -9.89191e-09, -1.006321e-08, -1.024931e-08, 
    -1.04407e-08, -1.069027e-08, -1.081776e-08, -1.106091e-08, -1.119517e-08,
  -7.043209e-09, -7.264491e-09, -7.528755e-09, -7.97973e-09, -8.49197e-09, 
    -8.92459e-09, -9.21515e-09, -9.611773e-09, -9.959422e-09, -1.005336e-08, 
    -1.017226e-08, -1.037992e-08, -1.054572e-08, -1.064294e-08, -1.079198e-08,
  -6.656272e-09, -7.014184e-09, -7.29421e-09, -7.645584e-09, -8.060103e-09, 
    -8.657543e-09, -9.10847e-09, -9.441172e-09, -9.765051e-09, -9.989853e-09, 
    -1.00866e-08, -1.017831e-08, -1.036117e-08, -1.048973e-08, -1.06075e-08,
  -6.353378e-09, -6.685856e-09, -7.038043e-09, -7.410961e-09, -7.836204e-09, 
    -8.23195e-09, -8.739246e-09, -9.251371e-09, -9.599063e-09, -9.876241e-09, 
    -9.977515e-09, -1.016105e-08, -1.030837e-08, -1.0394e-08, -1.049266e-08,
  -6.116376e-09, -6.362979e-09, -6.675504e-09, -7.070244e-09, -7.517678e-09, 
    -8.208365e-09, -8.61955e-09, -9.013006e-09, -9.43077e-09, -9.688224e-09, 
    -1.003975e-08, -1.010913e-08, -1.039147e-08, -1.058301e-08, -1.065319e-08,
  -1.360307e-08, -1.401712e-08, -1.413074e-08, -1.485105e-08, -1.542887e-08, 
    -1.610287e-08, -1.697822e-08, -1.771964e-08, -1.848877e-08, 
    -1.882317e-08, -1.838637e-08, -1.763e-08, -1.727548e-08, -1.784321e-08, 
    -1.92085e-08,
  -1.227923e-08, -1.27089e-08, -1.312559e-08, -1.345224e-08, -1.409371e-08, 
    -1.477515e-08, -1.573465e-08, -1.666707e-08, -1.733505e-08, -1.81338e-08, 
    -1.846965e-08, -1.825698e-08, -1.745693e-08, -1.687303e-08, -1.740984e-08,
  -1.041556e-08, -1.123269e-08, -1.190341e-08, -1.239814e-08, -1.286033e-08, 
    -1.339359e-08, -1.412196e-08, -1.520093e-08, -1.630069e-08, 
    -1.707343e-08, -1.783049e-08, -1.7982e-08, -1.804742e-08, -1.742841e-08, 
    -1.676766e-08,
  -8.531434e-09, -9.245505e-09, -1.00767e-08, -1.096461e-08, -1.163656e-08, 
    -1.226724e-08, -1.282517e-08, -1.350004e-08, -1.453579e-08, 
    -1.575952e-08, -1.684321e-08, -1.753386e-08, -1.769738e-08, 
    -1.772933e-08, -1.731305e-08,
  -7.546127e-09, -7.861377e-09, -8.342627e-09, -9.046018e-09, -9.927273e-09, 
    -1.078158e-08, -1.155271e-08, -1.221916e-08, -1.291946e-08, 
    -1.384842e-08, -1.508831e-08, -1.634874e-08, -1.708127e-08, 
    -1.744719e-08, -1.746633e-08,
  -7.303637e-09, -7.345485e-09, -7.471167e-09, -7.764166e-09, -8.291499e-09, 
    -9.061685e-09, -9.963412e-09, -1.083128e-08, -1.159744e-08, -1.23061e-08, 
    -1.318901e-08, -1.430323e-08, -1.562107e-08, -1.640862e-08, -1.687739e-08,
  -7.267531e-09, -7.220117e-09, -7.19168e-09, -7.226927e-09, -7.329615e-09, 
    -7.743096e-09, -8.372729e-09, -9.204734e-09, -1.009945e-08, -1.0859e-08, 
    -1.157998e-08, -1.235531e-08, -1.343866e-08, -1.469727e-08, -1.558624e-08,
  -7.386702e-09, -7.320013e-09, -7.220991e-09, -7.105832e-09, -7.055372e-09, 
    -7.109974e-09, -7.42654e-09, -7.896633e-09, -8.625568e-09, -9.466455e-09, 
    -1.026032e-08, -1.096258e-08, -1.16523e-08, -1.257234e-08, -1.367276e-08,
  -7.435847e-09, -7.350557e-09, -7.231948e-09, -7.158773e-09, -7.070343e-09, 
    -6.990872e-09, -7.014058e-09, -7.199862e-09, -7.544285e-09, 
    -8.101862e-09, -8.861639e-09, -9.667354e-09, -1.039445e-08, 
    -1.105467e-08, -1.17917e-08,
  -7.433173e-09, -7.429354e-09, -7.255961e-09, -7.163467e-09, -7.048747e-09, 
    -7.066097e-09, -7.063705e-09, -7.039088e-09, -7.142381e-09, 
    -7.367861e-09, -7.765631e-09, -8.376492e-09, -9.154571e-09, 
    -9.863633e-09, -1.047928e-08,
  -1.888933e-08, -1.896714e-08, -1.905716e-08, -1.860977e-08, -1.827615e-08, 
    -1.764753e-08, -1.68718e-08, -1.622357e-08, -1.652255e-08, -1.707312e-08, 
    -1.711756e-08, -1.715992e-08, -1.747173e-08, -1.773525e-08, -1.80567e-08,
  -1.632369e-08, -1.695802e-08, -1.757512e-08, -1.81421e-08, -1.811849e-08, 
    -1.805822e-08, -1.783149e-08, -1.728197e-08, -1.651263e-08, 
    -1.666532e-08, -1.71607e-08, -1.742704e-08, -1.758077e-08, -1.769535e-08, 
    -1.777229e-08,
  -1.308093e-08, -1.400908e-08, -1.50453e-08, -1.596715e-08, -1.684874e-08, 
    -1.737632e-08, -1.753272e-08, -1.764493e-08, -1.73324e-08, -1.669498e-08, 
    -1.672323e-08, -1.715075e-08, -1.758749e-08, -1.790119e-08, -1.797063e-08,
  -1.099614e-08, -1.153087e-08, -1.234482e-08, -1.337339e-08, -1.447575e-08, 
    -1.549751e-08, -1.645024e-08, -1.692565e-08, -1.732507e-08, -1.72781e-08, 
    -1.694586e-08, -1.692372e-08, -1.720298e-08, -1.763368e-08, -1.804204e-08,
  -9.892344e-09, -9.913257e-09, -1.019046e-08, -1.076951e-08, -1.173608e-08, 
    -1.295596e-08, -1.410858e-08, -1.529927e-08, -1.621726e-08, 
    -1.684059e-08, -1.715556e-08, -1.703644e-08, -1.719343e-08, 
    -1.737268e-08, -1.761605e-08,
  -1.017798e-08, -9.829709e-09, -9.627413e-09, -9.653827e-09, -9.907009e-09, 
    -1.060285e-08, -1.169982e-08, -1.290312e-08, -1.415067e-08, 
    -1.539718e-08, -1.625293e-08, -1.694355e-08, -1.71472e-08, -1.742726e-08, 
    -1.758934e-08,
  -1.124211e-08, -1.073896e-08, -1.015935e-08, -9.78548e-09, -9.498826e-09, 
    -9.460575e-09, -9.836911e-09, -1.066903e-08, -1.192449e-08, 
    -1.316341e-08, -1.446773e-08, -1.565017e-08, -1.656014e-08, 
    -1.722887e-08, -1.758456e-08,
  -1.205419e-08, -1.171291e-08, -1.116259e-08, -1.061009e-08, -1.001866e-08, 
    -9.607329e-09, -9.340031e-09, -9.365011e-09, -9.926934e-09, 
    -1.115065e-08, -1.239586e-08, -1.377328e-08, -1.503155e-08, 
    -1.610191e-08, -1.709208e-08,
  -1.277277e-08, -1.229314e-08, -1.19002e-08, -1.142775e-08, -1.094393e-08, 
    -1.030029e-08, -9.812426e-09, -9.339994e-09, -9.120957e-09, 
    -9.302869e-09, -1.025134e-08, -1.163845e-08, -1.31167e-08, -1.453115e-08, 
    -1.569571e-08,
  -1.261078e-08, -1.250077e-08, -1.215636e-08, -1.178581e-08, -1.140472e-08, 
    -1.104238e-08, -1.06553e-08, -1.01318e-08, -9.574292e-09, -9.200677e-09, 
    -9.039296e-09, -9.583742e-09, -1.081549e-08, -1.23644e-08, -1.397645e-08,
  -1.91252e-08, -1.927286e-08, -1.925502e-08, -1.927098e-08, -1.947586e-08, 
    -1.961981e-08, -1.967885e-08, -1.974347e-08, -1.975389e-08, 
    -1.965468e-08, -1.911478e-08, -1.823505e-08, -1.738188e-08, 
    -1.679294e-08, -1.675693e-08,
  -1.873565e-08, -1.891784e-08, -1.919823e-08, -1.936121e-08, -1.934351e-08, 
    -1.932501e-08, -1.940149e-08, -1.952044e-08, -1.964235e-08, 
    -1.981875e-08, -1.984943e-08, -1.953586e-08, -1.885004e-08, 
    -1.781211e-08, -1.692705e-08,
  -1.75102e-08, -1.773219e-08, -1.811592e-08, -1.83455e-08, -1.859406e-08, 
    -1.861569e-08, -1.864518e-08, -1.877785e-08, -1.893916e-08, 
    -1.914878e-08, -1.938711e-08, -1.95696e-08, -1.961017e-08, -1.925792e-08, 
    -1.847846e-08,
  -1.642881e-08, -1.647214e-08, -1.67043e-08, -1.69679e-08, -1.719843e-08, 
    -1.742835e-08, -1.761933e-08, -1.77886e-08, -1.797637e-08, -1.822404e-08, 
    -1.853418e-08, -1.882725e-08, -1.909217e-08, -1.92655e-08, -1.919773e-08,
  -1.534045e-08, -1.543214e-08, -1.537131e-08, -1.539828e-08, -1.544469e-08, 
    -1.553407e-08, -1.570467e-08, -1.590376e-08, -1.613411e-08, 
    -1.643129e-08, -1.677062e-08, -1.723422e-08, -1.769709e-08, 
    -1.816542e-08, -1.858072e-08,
  -1.478846e-08, -1.462075e-08, -1.449013e-08, -1.441297e-08, -1.42074e-08, 
    -1.406902e-08, -1.393532e-08, -1.391119e-08, -1.398139e-08, 
    -1.416859e-08, -1.44644e-08, -1.490548e-08, -1.550963e-08, -1.618262e-08, 
    -1.685371e-08,
  -1.514807e-08, -1.471856e-08, -1.429793e-08, -1.399263e-08, -1.374938e-08, 
    -1.34082e-08, -1.319029e-08, -1.296863e-08, -1.280459e-08, -1.272945e-08, 
    -1.278452e-08, -1.293573e-08, -1.326308e-08, -1.382317e-08, -1.458284e-08,
  -1.591668e-08, -1.548096e-08, -1.502468e-08, -1.463875e-08, -1.417802e-08, 
    -1.374921e-08, -1.330182e-08, -1.293461e-08, -1.261967e-08, 
    -1.240626e-08, -1.220923e-08, -1.213089e-08, -1.208764e-08, 
    -1.223272e-08, -1.260726e-08,
  -1.673652e-08, -1.622234e-08, -1.566521e-08, -1.526177e-08, -1.489568e-08, 
    -1.452446e-08, -1.416635e-08, -1.372638e-08, -1.327662e-08, 
    -1.284825e-08, -1.248825e-08, -1.212456e-08, -1.181472e-08, 
    -1.159446e-08, -1.159013e-08,
  -1.723096e-08, -1.700065e-08, -1.654101e-08, -1.606875e-08, -1.561846e-08, 
    -1.522343e-08, -1.502393e-08, -1.472794e-08, -1.437493e-08, 
    -1.404332e-08, -1.36122e-08, -1.317171e-08, -1.271389e-08, -1.224725e-08, 
    -1.186222e-08,
  -1.184312e-08, -1.260061e-08, -1.32032e-08, -1.3555e-08, -1.412043e-08, 
    -1.459037e-08, -1.50747e-08, -1.536095e-08, -1.572293e-08, -1.616725e-08, 
    -1.680721e-08, -1.745156e-08, -1.827645e-08, -1.926287e-08, -2.054074e-08,
  -1.19833e-08, -1.268241e-08, -1.332626e-08, -1.371518e-08, -1.422892e-08, 
    -1.473398e-08, -1.53601e-08, -1.57743e-08, -1.600361e-08, -1.634469e-08, 
    -1.689409e-08, -1.750147e-08, -1.824841e-08, -1.891966e-08, -2.022866e-08,
  -1.205334e-08, -1.278058e-08, -1.357179e-08, -1.399829e-08, -1.451598e-08, 
    -1.501288e-08, -1.556612e-08, -1.599317e-08, -1.620943e-08, 
    -1.650683e-08, -1.697435e-08, -1.754231e-08, -1.830381e-08, 
    -1.896588e-08, -1.969898e-08,
  -1.253312e-08, -1.312274e-08, -1.392318e-08, -1.448446e-08, -1.493439e-08, 
    -1.537999e-08, -1.602064e-08, -1.649975e-08, -1.669523e-08, 
    -1.686822e-08, -1.724218e-08, -1.767231e-08, -1.838229e-08, 
    -1.916353e-08, -1.954286e-08,
  -1.305449e-08, -1.363364e-08, -1.454786e-08, -1.517508e-08, -1.569974e-08, 
    -1.614552e-08, -1.670468e-08, -1.72895e-08, -1.759626e-08, -1.774151e-08, 
    -1.799249e-08, -1.825573e-08, -1.872306e-08, -1.950519e-08, -1.978797e-08,
  -1.366947e-08, -1.432407e-08, -1.52708e-08, -1.601457e-08, -1.652007e-08, 
    -1.688251e-08, -1.752272e-08, -1.812152e-08, -1.84624e-08, -1.859529e-08, 
    -1.877206e-08, -1.891365e-08, -1.925882e-08, -1.997675e-08, -2.026358e-08,
  -1.41738e-08, -1.496965e-08, -1.581354e-08, -1.663646e-08, -1.702888e-08, 
    -1.737138e-08, -1.787242e-08, -1.852099e-08, -1.889535e-08, 
    -1.899477e-08, -1.904984e-08, -1.921659e-08, -1.952034e-08, 
    -2.014137e-08, -2.06005e-08,
  -1.469373e-08, -1.542971e-08, -1.619414e-08, -1.697902e-08, -1.760202e-08, 
    -1.785504e-08, -1.846554e-08, -1.88792e-08, -1.925039e-08, -1.931995e-08, 
    -1.936492e-08, -1.940848e-08, -1.957825e-08, -1.989257e-08, -2.04186e-08,
  -1.500116e-08, -1.565934e-08, -1.654269e-08, -1.713558e-08, -1.755779e-08, 
    -1.79335e-08, -1.850084e-08, -1.923136e-08, -1.958334e-08, -1.962523e-08, 
    -1.945391e-08, -1.93068e-08, -1.938103e-08, -1.983781e-08, -2.044003e-08,
  -1.5015e-08, -1.569475e-08, -1.665603e-08, -1.742687e-08, -1.819458e-08, 
    -1.867633e-08, -1.977019e-08, -1.964635e-08, -1.977114e-08, -1.97052e-08, 
    -1.965266e-08, -1.974847e-08, -1.977642e-08, -1.978792e-08, -2.021676e-08,
  -3.360779e-09, -3.62136e-09, -3.879433e-09, -4.213411e-09, -4.512735e-09, 
    -4.872388e-09, -5.16108e-09, -5.657242e-09, -6.275623e-09, -7.003575e-09, 
    -7.597559e-09, -8.252984e-09, -8.86983e-09, -9.64783e-09, -1.053075e-08,
  -3.085629e-09, -3.417351e-09, -3.698597e-09, -3.990985e-09, -4.24918e-09, 
    -4.527998e-09, -4.830035e-09, -5.227933e-09, -5.735321e-09, 
    -6.413596e-09, -7.106018e-09, -7.737565e-09, -8.271665e-09, 
    -8.932941e-09, -9.62119e-09,
  -2.933898e-09, -3.244861e-09, -3.523562e-09, -3.78681e-09, -4.03341e-09, 
    -4.288815e-09, -4.590585e-09, -4.981558e-09, -5.415725e-09, -5.97407e-09, 
    -6.666559e-09, -7.436909e-09, -7.966789e-09, -8.520418e-09, -9.155988e-09,
  -2.864897e-09, -3.143047e-09, -3.416332e-09, -3.65976e-09, -3.869508e-09, 
    -4.130933e-09, -4.437817e-09, -4.841467e-09, -5.247864e-09, 
    -5.711295e-09, -6.279069e-09, -7.010684e-09, -7.651266e-09, 
    -8.160505e-09, -8.831223e-09,
  -2.827449e-09, -3.077303e-09, -3.331504e-09, -3.585463e-09, -3.804395e-09, 
    -4.130292e-09, -4.475344e-09, -4.878501e-09, -5.258648e-09, 
    -5.695486e-09, -6.191746e-09, -6.821331e-09, -7.42892e-09, -7.936405e-09, 
    -8.562459e-09,
  -2.822687e-09, -3.065376e-09, -3.34375e-09, -3.640822e-09, -3.927741e-09, 
    -4.267279e-09, -4.637884e-09, -5.015143e-09, -5.421529e-09, 
    -5.821397e-09, -6.280744e-09, -6.858347e-09, -7.398967e-09, 
    -7.919382e-09, -8.587348e-09,
  -2.830812e-09, -3.070492e-09, -3.424714e-09, -3.806626e-09, -4.096222e-09, 
    -4.492008e-09, -4.802499e-09, -5.236267e-09, -5.593e-09, -6.037026e-09, 
    -6.517554e-09, -7.002526e-09, -7.491858e-09, -8.034336e-09, -8.709203e-09,
  -2.865257e-09, -3.188349e-09, -3.565682e-09, -3.993511e-09, -4.400279e-09, 
    -4.785709e-09, -5.249403e-09, -5.439389e-09, -5.805495e-09, 
    -6.280008e-09, -6.765767e-09, -7.307249e-09, -7.837671e-09, 
    -8.440055e-09, -9.020309e-09,
  -2.914262e-09, -3.387043e-09, -3.8996e-09, -4.319329e-09, -4.735728e-09, 
    -5.086539e-09, -5.295822e-09, -5.752269e-09, -6.203905e-09, -6.75263e-09, 
    -7.23131e-09, -7.729724e-09, -8.286983e-09, -9.007637e-09, -9.697031e-09,
  -3.015704e-09, -3.669595e-09, -4.15301e-09, -4.599389e-09, -4.985556e-09, 
    -5.328644e-09, -6.058003e-09, -6.122443e-09, -6.651228e-09, 
    -7.217466e-09, -7.721683e-09, -8.252485e-09, -8.973181e-09, -9.70559e-09, 
    -1.028303e-08,
  -3.828187e-09, -3.715299e-09, -3.704793e-09, -3.647743e-09, -3.516418e-09, 
    -3.435756e-09, -3.389044e-09, -3.544771e-09, -3.812217e-09, 
    -4.093621e-09, -4.326489e-09, -4.785089e-09, -5.49613e-09, -6.271062e-09, 
    -6.784658e-09,
  -3.622872e-09, -3.474352e-09, -3.383788e-09, -3.341194e-09, -3.252964e-09, 
    -3.221745e-09, -3.19231e-09, -3.28639e-09, -3.473323e-09, -3.842962e-09, 
    -4.047862e-09, -4.309135e-09, -4.899134e-09, -5.721087e-09, -6.465433e-09,
  -3.615836e-09, -3.400903e-09, -3.25466e-09, -3.149514e-09, -3.069148e-09, 
    -3.052458e-09, -3.050757e-09, -3.132764e-09, -3.212705e-09, -3.49932e-09, 
    -3.828303e-09, -4.029596e-09, -4.414932e-09, -5.113132e-09, -5.991251e-09,
  -3.369035e-09, -3.151529e-09, -3.01679e-09, -2.922236e-09, -2.834126e-09, 
    -2.829251e-09, -2.889772e-09, -3.005796e-09, -3.150344e-09, 
    -3.286942e-09, -3.582393e-09, -3.822954e-09, -4.122741e-09, 
    -4.675342e-09, -5.506769e-09,
  -3.244037e-09, -2.997913e-09, -2.836989e-09, -2.73676e-09, -2.661787e-09, 
    -2.601946e-09, -2.674673e-09, -2.810501e-09, -3.043821e-09, 
    -3.187667e-09, -3.39077e-09, -3.619881e-09, -3.869126e-09, -4.295273e-09, 
    -5.052653e-09,
  -3.049162e-09, -2.808282e-09, -2.636227e-09, -2.520287e-09, -2.460809e-09, 
    -2.465059e-09, -2.565282e-09, -2.70162e-09, -2.927955e-09, -3.106139e-09, 
    -3.261135e-09, -3.506368e-09, -3.758853e-09, -4.056717e-09, -4.657815e-09,
  -2.890452e-09, -2.656953e-09, -2.478553e-09, -2.362084e-09, -2.317977e-09, 
    -2.338234e-09, -2.464677e-09, -2.622941e-09, -2.803813e-09, -2.99307e-09, 
    -3.17699e-09, -3.431176e-09, -3.715368e-09, -3.995389e-09, -4.512101e-09,
  -2.713904e-09, -2.525791e-09, -2.366854e-09, -2.249318e-09, -2.233969e-09, 
    -2.288995e-09, -2.421793e-09, -2.550942e-09, -2.705247e-09, 
    -2.911602e-09, -3.10447e-09, -3.365988e-09, -3.67726e-09, -3.996647e-09, 
    -4.412012e-09,
  -2.584668e-09, -2.400709e-09, -2.285663e-09, -2.213733e-09, -2.165093e-09, 
    -2.192817e-09, -2.356837e-09, -2.463386e-09, -2.641578e-09, 
    -2.898201e-09, -3.068729e-09, -3.296469e-09, -3.619269e-09, 
    -4.004702e-09, -4.432069e-09,
  -2.46192e-09, -2.330591e-09, -2.219606e-09, -2.16155e-09, -2.177356e-09, 
    -2.212611e-09, -2.323345e-09, -2.477395e-09, -2.666134e-09, -2.87327e-09, 
    -3.068258e-09, -3.412971e-09, -3.727005e-09, -4.060272e-09, -4.448584e-09,
  -1.042821e-08, -1.017612e-08, -9.874756e-09, -9.633676e-09, -9.485309e-09, 
    -9.51574e-09, -9.601519e-09, -9.743732e-09, -9.759258e-09, -9.792791e-09, 
    -9.832904e-09, -9.940833e-09, -1.012815e-08, -1.061764e-08, -1.140042e-08,
  -9.844381e-09, -9.619699e-09, -9.336069e-09, -9.017541e-09, -8.781863e-09, 
    -8.671167e-09, -8.612954e-09, -8.611197e-09, -8.608815e-09, 
    -8.674362e-09, -8.798803e-09, -8.952466e-09, -9.132176e-09, -9.39465e-09, 
    -9.824406e-09,
  -9.499789e-09, -9.324149e-09, -9.107688e-09, -8.749852e-09, -8.414492e-09, 
    -8.147823e-09, -7.999459e-09, -7.866818e-09, -7.740392e-09, 
    -7.722272e-09, -7.872137e-09, -8.100655e-09, -8.348836e-09, 
    -8.562391e-09, -8.871531e-09,
  -8.972187e-09, -8.818827e-09, -8.63972e-09, -8.336947e-09, -7.978348e-09, 
    -7.602512e-09, -7.385029e-09, -7.198397e-09, -7.052347e-09, 
    -6.957385e-09, -6.993845e-09, -7.176406e-09, -7.462746e-09, 
    -7.732064e-09, -7.995816e-09,
  -8.531625e-09, -8.451279e-09, -8.278219e-09, -8.050764e-09, -7.721627e-09, 
    -7.337306e-09, -7.017468e-09, -6.78494e-09, -6.638115e-09, -6.533748e-09, 
    -6.526242e-09, -6.533815e-09, -6.700537e-09, -6.963006e-09, -7.190234e-09,
  -7.905722e-09, -7.898434e-09, -7.788444e-09, -7.661825e-09, -7.373118e-09, 
    -7.074597e-09, -6.723847e-09, -6.457401e-09, -6.301305e-09, 
    -6.207853e-09, -6.144588e-09, -6.114072e-09, -6.139049e-09, -6.26658e-09, 
    -6.481311e-09,
  -7.359251e-09, -7.435762e-09, -7.366783e-09, -7.307643e-09, -7.091688e-09, 
    -6.860799e-09, -6.572781e-09, -6.296606e-09, -6.064977e-09, 
    -5.925046e-09, -5.83224e-09, -5.714541e-09, -5.67608e-09, -5.640746e-09, 
    -5.722884e-09,
  -6.558604e-09, -6.782691e-09, -6.860974e-09, -6.835932e-09, -6.752539e-09, 
    -6.558908e-09, -6.382662e-09, -6.125844e-09, -5.887757e-09, 
    -5.650206e-09, -5.532059e-09, -5.385388e-09, -5.268587e-09, 
    -5.215039e-09, -5.182487e-09,
  -5.763774e-09, -5.97363e-09, -6.272667e-09, -6.438079e-09, -6.445405e-09, 
    -6.272961e-09, -6.102193e-09, -5.85511e-09, -5.606998e-09, -5.318587e-09, 
    -5.066032e-09, -4.904357e-09, -4.789784e-09, -4.723364e-09, -4.740897e-09,
  -5.00632e-09, -5.291537e-09, -5.555908e-09, -5.886478e-09, -5.932917e-09, 
    -6.039238e-09, -5.978147e-09, -5.732258e-09, -5.43415e-09, -5.103307e-09, 
    -4.789166e-09, -4.551953e-09, -4.458014e-09, -4.402321e-09, -4.407878e-09,
  -1.373805e-08, -1.400086e-08, -1.399263e-08, -1.504785e-08, -1.555283e-08, 
    -1.597079e-08, -1.556463e-08, -1.919447e-08, -1.911531e-08, 
    -1.603786e-08, -1.856179e-08, -2.269934e-08, -2.191153e-08, 
    -2.167342e-08, -2.174452e-08,
  -1.283299e-08, -1.32916e-08, -1.33933e-08, -1.35991e-08, -1.427243e-08, 
    -1.520395e-08, -1.530796e-08, -1.666684e-08, -1.922738e-08, 
    -1.788751e-08, -1.732568e-08, -1.97642e-08, -2.16909e-08, -2.219621e-08, 
    -2.197418e-08,
  -1.2198e-08, -1.22411e-08, -1.262093e-08, -1.265482e-08, -1.318009e-08, 
    -1.374308e-08, -1.470921e-08, -1.505475e-08, -1.732985e-08, -1.89055e-08, 
    -1.775962e-08, -1.824685e-08, -1.943208e-08, -2.15957e-08, -2.172252e-08,
  -1.177894e-08, -1.176077e-08, -1.176517e-08, -1.186781e-08, -1.206757e-08, 
    -1.273193e-08, -1.329528e-08, -1.413497e-08, -1.490474e-08, 
    -1.745461e-08, -1.818809e-08, -1.779664e-08, -1.805865e-08, 
    -1.949612e-08, -2.099807e-08,
  -1.066863e-08, -1.104189e-08, -1.116825e-08, -1.126593e-08, -1.130685e-08, 
    -1.156717e-08, -1.233921e-08, -1.285039e-08, -1.373002e-08, 
    -1.485294e-08, -1.697451e-08, -1.786878e-08, -1.767231e-08, 
    -1.807934e-08, -1.946188e-08,
  -9.671902e-09, -9.83768e-09, -1.024325e-08, -1.058165e-08, -1.075193e-08, 
    -1.081968e-08, -1.117524e-08, -1.195821e-08, -1.245207e-08, 
    -1.353327e-08, -1.481707e-08, -1.663653e-08, -1.729831e-08, 
    -1.738955e-08, -1.80015e-08,
  -8.657175e-09, -8.868164e-09, -9.088732e-09, -9.613739e-09, -9.987045e-09, 
    -1.026773e-08, -1.038381e-08, -1.089965e-08, -1.162941e-08, 
    -1.223467e-08, -1.321742e-08, -1.485378e-08, -1.632353e-08, 
    -1.687284e-08, -1.709182e-08,
  -7.436807e-09, -7.939682e-09, -8.154441e-09, -8.488247e-09, -8.957236e-09, 
    -9.319685e-09, -9.718715e-09, -9.95713e-09, -1.063352e-08, -1.126443e-08, 
    -1.207172e-08, -1.293566e-08, -1.4584e-08, -1.597596e-08, -1.658085e-08,
  -5.972303e-09, -6.453139e-09, -7.098709e-09, -7.452015e-09, -7.930748e-09, 
    -8.424001e-09, -8.805556e-09, -9.216712e-09, -9.584941e-09, 
    -1.035744e-08, -1.097753e-08, -1.197186e-08, -1.277243e-08, 
    -1.435327e-08, -1.554113e-08,
  -4.733839e-09, -5.115039e-09, -5.61437e-09, -6.168252e-09, -6.617511e-09, 
    -7.303025e-09, -7.897156e-09, -8.373316e-09, -8.727684e-09, 
    -9.255061e-09, -1.002197e-08, -1.076884e-08, -1.168303e-08, 
    -1.257522e-08, -1.39716e-08,
  -1.120914e-08, -1.28334e-08, -1.354407e-08, -1.41218e-08, -1.424786e-08, 
    -1.51542e-08, -1.676491e-08, -1.782924e-08, -1.729297e-08, -1.724944e-08, 
    -1.892041e-08, -2.121993e-08, -2.173718e-08, -2.155921e-08, -2.087739e-08,
  -1.045249e-08, -1.156884e-08, -1.297037e-08, -1.37495e-08, -1.420686e-08, 
    -1.463828e-08, -1.528104e-08, -1.780685e-08, -1.799933e-08, 
    -1.745064e-08, -1.760405e-08, -1.988639e-08, -2.109578e-08, 
    -2.137876e-08, -2.067191e-08,
  -1.027326e-08, -1.02539e-08, -1.171053e-08, -1.299692e-08, -1.361291e-08, 
    -1.43664e-08, -1.478407e-08, -1.604206e-08, -1.806619e-08, -1.815714e-08, 
    -1.744366e-08, -1.881888e-08, -2.006141e-08, -2.077124e-08, -2.054152e-08,
  -9.795201e-09, -1.009979e-08, -1.037172e-08, -1.199315e-08, -1.291234e-08, 
    -1.381911e-08, -1.433105e-08, -1.493694e-08, -1.69168e-08, -1.823014e-08, 
    -1.792511e-08, -1.814971e-08, -1.934121e-08, -2.002792e-08, -2.022124e-08,
  -9.445934e-09, -9.817188e-09, -1.008969e-08, -1.074971e-08, -1.221494e-08, 
    -1.296205e-08, -1.404751e-08, -1.436867e-08, -1.534744e-08, -1.76852e-08, 
    -1.828381e-08, -1.807041e-08, -1.887311e-08, -1.935868e-08, -1.972905e-08,
  -9.109857e-09, -9.42457e-09, -9.813262e-09, -1.007488e-08, -1.121717e-08, 
    -1.22935e-08, -1.312828e-08, -1.396674e-08, -1.444255e-08, -1.59672e-08, 
    -1.808936e-08, -1.839952e-08, -1.863522e-08, -1.892409e-08, -1.922561e-08,
  -8.949198e-09, -9.218923e-09, -9.435788e-09, -9.804596e-09, -1.023715e-08, 
    -1.150778e-08, -1.243443e-08, -1.344479e-08, -1.387699e-08, 
    -1.455905e-08, -1.666761e-08, -1.812601e-08, -1.883284e-08, 
    -1.871033e-08, -1.876718e-08,
  -9.044182e-09, -9.067923e-09, -9.269543e-09, -9.493163e-09, -9.740405e-09, 
    -1.041558e-08, -1.167882e-08, -1.253448e-08, -1.374881e-08, 
    -1.382196e-08, -1.509031e-08, -1.715778e-08, -1.863388e-08, 
    -1.891519e-08, -1.864311e-08,
  -9.311012e-09, -9.262702e-09, -9.240058e-09, -9.412154e-09, -9.56913e-09, 
    -9.756395e-09, -1.05531e-08, -1.174059e-08, -1.264633e-08, -1.382813e-08, 
    -1.394793e-08, -1.558798e-08, -1.781922e-08, -1.876664e-08, -1.875416e-08,
  -9.305502e-09, -9.402821e-09, -9.505516e-09, -9.458121e-09, -9.527794e-09, 
    -9.63904e-09, -9.858336e-09, -1.071405e-08, -1.181932e-08, -1.283229e-08, 
    -1.383265e-08, -1.426665e-08, -1.621199e-08, -1.826938e-08, -1.879733e-08,
  -1.520524e-08, -1.530426e-08, -1.585239e-08, -1.582349e-08, -1.504698e-08, 
    -1.443458e-08, -1.40671e-08, -1.396349e-08, -1.352629e-08, -1.287107e-08, 
    -1.286362e-08, -1.332604e-08, -1.618852e-08, -1.884835e-08, -1.98772e-08,
  -1.592348e-08, -1.596392e-08, -1.588907e-08, -1.529364e-08, -1.449866e-08, 
    -1.445002e-08, -1.361004e-08, -1.296767e-08, -1.280097e-08, 
    -1.237811e-08, -1.24258e-08, -1.278366e-08, -1.463281e-08, -1.786222e-08, 
    -1.980064e-08,
  -1.625183e-08, -1.604377e-08, -1.560572e-08, -1.490833e-08, -1.436519e-08, 
    -1.402414e-08, -1.291759e-08, -1.231782e-08, -1.229114e-08, 
    -1.195224e-08, -1.192322e-08, -1.245384e-08, -1.346117e-08, 
    -1.689909e-08, -1.915061e-08,
  -1.517483e-08, -1.520195e-08, -1.481748e-08, -1.430056e-08, -1.375132e-08, 
    -1.29573e-08, -1.231535e-08, -1.202425e-08, -1.188302e-08, -1.188449e-08, 
    -1.178006e-08, -1.219259e-08, -1.303597e-08, -1.564541e-08, -1.847909e-08,
  -1.421686e-08, -1.413618e-08, -1.390207e-08, -1.348516e-08, -1.307098e-08, 
    -1.235164e-08, -1.202724e-08, -1.190566e-08, -1.174309e-08, 
    -1.159557e-08, -1.163828e-08, -1.182594e-08, -1.279323e-08, 
    -1.430303e-08, -1.754447e-08,
  -1.37714e-08, -1.360528e-08, -1.329374e-08, -1.297564e-08, -1.256823e-08, 
    -1.20427e-08, -1.185814e-08, -1.1838e-08, -1.16244e-08, -1.155114e-08, 
    -1.160408e-08, -1.158351e-08, -1.24223e-08, -1.339163e-08, -1.631472e-08,
  -1.332133e-08, -1.31676e-08, -1.308496e-08, -1.277693e-08, -1.236024e-08, 
    -1.199148e-08, -1.172938e-08, -1.167541e-08, -1.144412e-08, 
    -1.131899e-08, -1.141678e-08, -1.138425e-08, -1.208267e-08, 
    -1.291787e-08, -1.494673e-08,
  -1.255839e-08, -1.261538e-08, -1.255177e-08, -1.239351e-08, -1.219531e-08, 
    -1.197574e-08, -1.168579e-08, -1.161244e-08, -1.146815e-08, 
    -1.117854e-08, -1.115125e-08, -1.11862e-08, -1.185623e-08, -1.25652e-08, 
    -1.3863e-08,
  -1.141918e-08, -1.154781e-08, -1.171995e-08, -1.182477e-08, -1.194764e-08, 
    -1.18454e-08, -1.151039e-08, -1.137942e-08, -1.131757e-08, -1.114009e-08, 
    -1.091762e-08, -1.094485e-08, -1.141048e-08, -1.226297e-08, -1.325494e-08,
  -1.024748e-08, -1.060141e-08, -1.079701e-08, -1.114223e-08, -1.135074e-08, 
    -1.159336e-08, -1.153821e-08, -1.129139e-08, -1.112687e-08, 
    -1.105742e-08, -1.08244e-08, -1.075571e-08, -1.103277e-08, -1.182871e-08, 
    -1.288425e-08,
  -1.617395e-08, -1.662803e-08, -1.695638e-08, -1.721133e-08, -1.74496e-08, 
    -1.731667e-08, -1.741112e-08, -1.855245e-08, -1.930849e-08, 
    -2.017685e-08, -2.061849e-08, -2.085058e-08, -2.088207e-08, 
    -2.013308e-08, -1.937378e-08,
  -1.608415e-08, -1.636126e-08, -1.65393e-08, -1.694931e-08, -1.738394e-08, 
    -1.737873e-08, -1.78974e-08, -1.845014e-08, -1.884111e-08, -1.933543e-08, 
    -1.915043e-08, -1.914511e-08, -1.886593e-08, -1.829918e-08, -1.76583e-08,
  -1.564479e-08, -1.595193e-08, -1.631039e-08, -1.664023e-08, -1.703353e-08, 
    -1.748995e-08, -1.798916e-08, -1.820148e-08, -1.828692e-08, -1.81996e-08, 
    -1.822719e-08, -1.774403e-08, -1.73341e-08, -1.708096e-08, -1.677466e-08,
  -1.546858e-08, -1.548456e-08, -1.584052e-08, -1.627407e-08, -1.657064e-08, 
    -1.707233e-08, -1.760635e-08, -1.781366e-08, -1.777673e-08, 
    -1.786792e-08, -1.771317e-08, -1.744781e-08, -1.672911e-08, 
    -1.650933e-08, -1.624852e-08,
  -1.55054e-08, -1.53199e-08, -1.548324e-08, -1.573202e-08, -1.616964e-08, 
    -1.66218e-08, -1.699993e-08, -1.732205e-08, -1.749627e-08, -1.749429e-08, 
    -1.744513e-08, -1.706545e-08, -1.634412e-08, -1.582407e-08, -1.558093e-08,
  -1.520221e-08, -1.544248e-08, -1.557769e-08, -1.561016e-08, -1.588276e-08, 
    -1.632568e-08, -1.671735e-08, -1.707172e-08, -1.717339e-08, 
    -1.732784e-08, -1.727139e-08, -1.700506e-08, -1.638323e-08, 
    -1.581146e-08, -1.553508e-08,
  -1.399575e-08, -1.482061e-08, -1.531628e-08, -1.557021e-08, -1.568145e-08, 
    -1.581695e-08, -1.611553e-08, -1.645235e-08, -1.691704e-08, 
    -1.720438e-08, -1.730528e-08, -1.71513e-08, -1.657825e-08, -1.591075e-08, 
    -1.551972e-08,
  -1.267754e-08, -1.345972e-08, -1.426308e-08, -1.508448e-08, -1.562052e-08, 
    -1.591535e-08, -1.591999e-08, -1.599785e-08, -1.632049e-08, 
    -1.669026e-08, -1.705729e-08, -1.699505e-08, -1.668986e-08, 
    -1.606317e-08, -1.563837e-08,
  -1.25455e-08, -1.238254e-08, -1.278311e-08, -1.359793e-08, -1.461533e-08, 
    -1.540077e-08, -1.579564e-08, -1.592946e-08, -1.602018e-08, 
    -1.626119e-08, -1.674469e-08, -1.697178e-08, -1.682329e-08, 
    -1.636662e-08, -1.587373e-08,
  -1.271092e-08, -1.256735e-08, -1.221389e-08, -1.229774e-08, -1.284616e-08, 
    -1.394898e-08, -1.484852e-08, -1.541578e-08, -1.571607e-08, -1.5987e-08, 
    -1.625511e-08, -1.658679e-08, -1.678319e-08, -1.649495e-08, -1.617144e-08,
  -1.300613e-08, -1.293336e-08, -1.291123e-08, -1.278977e-08, -1.29959e-08, 
    -1.342984e-08, -1.396807e-08, -1.44475e-08, -1.478592e-08, -1.483894e-08, 
    -1.491468e-08, -1.513656e-08, -1.54865e-08, -1.621001e-08, -1.677267e-08,
  -1.227083e-08, -1.2305e-08, -1.225e-08, -1.214846e-08, -1.213971e-08, 
    -1.227088e-08, -1.245412e-08, -1.276933e-08, -1.309321e-08, 
    -1.349962e-08, -1.391105e-08, -1.427901e-08, -1.450678e-08, 
    -1.502561e-08, -1.580646e-08,
  -1.17967e-08, -1.186261e-08, -1.186505e-08, -1.178863e-08, -1.175677e-08, 
    -1.179316e-08, -1.185736e-08, -1.189152e-08, -1.205203e-08, 
    -1.234956e-08, -1.278613e-08, -1.326658e-08, -1.36408e-08, -1.396367e-08, 
    -1.464123e-08,
  -1.123293e-08, -1.127066e-08, -1.139468e-08, -1.144578e-08, -1.14368e-08, 
    -1.147797e-08, -1.153192e-08, -1.150601e-08, -1.153218e-08, 
    -1.167207e-08, -1.190707e-08, -1.234864e-08, -1.275038e-08, 
    -1.309412e-08, -1.358713e-08,
  -1.068187e-08, -1.075626e-08, -1.087801e-08, -1.09998e-08, -1.105634e-08, 
    -1.109824e-08, -1.119222e-08, -1.119719e-08, -1.119615e-08, 
    -1.126048e-08, -1.141029e-08, -1.16432e-08, -1.205869e-08, -1.234621e-08, 
    -1.273488e-08,
  -9.98382e-09, -1.014081e-08, -1.027556e-08, -1.051513e-08, -1.063018e-08, 
    -1.071238e-08, -1.083129e-08, -1.089662e-08, -1.090182e-08, 
    -1.094513e-08, -1.10667e-08, -1.121116e-08, -1.157782e-08, -1.186411e-08, 
    -1.208643e-08,
  -9.321544e-09, -9.52177e-09, -9.652326e-09, -9.867893e-09, -1.017378e-08, 
    -1.033218e-08, -1.04984e-08, -1.061638e-08, -1.066302e-08, -1.066807e-08, 
    -1.073799e-08, -1.085618e-08, -1.108387e-08, -1.153418e-08, -1.174001e-08,
  -8.806776e-09, -8.969729e-09, -9.123642e-09, -9.238435e-09, -9.511544e-09, 
    -9.806347e-09, -1.002147e-08, -1.025124e-08, -1.039286e-08, 
    -1.047124e-08, -1.054103e-08, -1.061574e-08, -1.071645e-08, -1.11347e-08, 
    -1.145481e-08,
  -8.397611e-09, -8.533318e-09, -8.742718e-09, -8.930717e-09, -9.102407e-09, 
    -9.289276e-09, -9.468352e-09, -9.712713e-09, -9.931882e-09, -1.01309e-08, 
    -1.027019e-08, -1.04761e-08, -1.058918e-08, -1.091061e-08, -1.124765e-08,
  -7.916182e-09, -8.15106e-09, -8.338991e-09, -8.60847e-09, -8.861292e-09, 
    -9.052659e-09, -9.084799e-09, -9.26739e-09, -9.532096e-09, -9.73376e-09, 
    -9.935348e-09, -1.014774e-08, -1.037478e-08, -1.072615e-08, -1.104958e-08,
  -1.406925e-08, -1.315869e-08, -1.167955e-08, -1.047697e-08, -9.967856e-09, 
    -1.066459e-08, -1.241893e-08, -1.332526e-08, -1.38044e-08, -1.527268e-08, 
    -1.609514e-08, -1.680699e-08, -1.746738e-08, -1.806925e-08, -1.883521e-08,
  -1.404038e-08, -1.405102e-08, -1.341229e-08, -1.277259e-08, -1.236931e-08, 
    -1.296399e-08, -1.33341e-08, -1.376539e-08, -1.406292e-08, -1.453718e-08, 
    -1.461154e-08, -1.522164e-08, -1.597384e-08, -1.678727e-08, -1.75142e-08,
  -1.325895e-08, -1.463106e-08, -1.512143e-08, -1.478052e-08, -1.465847e-08, 
    -1.415688e-08, -1.403285e-08, -1.399385e-08, -1.400868e-08, 
    -1.379569e-08, -1.366613e-08, -1.384453e-08, -1.424192e-08, 
    -1.469589e-08, -1.537003e-08,
  -1.148538e-08, -1.214474e-08, -1.310629e-08, -1.346524e-08, -1.333914e-08, 
    -1.328679e-08, -1.323882e-08, -1.319465e-08, -1.313608e-08, -1.3014e-08, 
    -1.301503e-08, -1.304149e-08, -1.322941e-08, -1.347311e-08, -1.374389e-08,
  -1.050853e-08, -1.086199e-08, -1.13096e-08, -1.173056e-08, -1.184982e-08, 
    -1.19784e-08, -1.208594e-08, -1.220259e-08, -1.226575e-08, -1.22434e-08, 
    -1.235377e-08, -1.250484e-08, -1.275754e-08, -1.303704e-08, -1.330345e-08,
  -9.716703e-09, -9.864094e-09, -1.013714e-08, -1.046806e-08, -1.07491e-08, 
    -1.089652e-08, -1.106453e-08, -1.11869e-08, -1.126281e-08, -1.130554e-08, 
    -1.140114e-08, -1.152518e-08, -1.169187e-08, -1.195689e-08, -1.225472e-08,
  -9.212627e-09, -9.292727e-09, -9.397607e-09, -9.601854e-09, -9.924023e-09, 
    -1.017239e-08, -1.03448e-08, -1.047258e-08, -1.061148e-08, -1.07736e-08, 
    -1.090222e-08, -1.103362e-08, -1.114613e-08, -1.127662e-08, -1.146853e-08,
  -8.935364e-09, -9.038363e-09, -9.096228e-09, -9.184107e-09, -9.374302e-09, 
    -9.664544e-09, -9.858866e-09, -1.00072e-08, -1.019222e-08, -1.040683e-08, 
    -1.058826e-08, -1.077637e-08, -1.094903e-08, -1.102799e-08, -1.110616e-08,
  -8.570981e-09, -8.692212e-09, -8.773896e-09, -8.889755e-09, -9.028456e-09, 
    -9.228872e-09, -9.401159e-09, -9.598833e-09, -9.783308e-09, 
    -1.002298e-08, -1.021435e-08, -1.042046e-08, -1.068251e-08, 
    -1.092465e-08, -1.104345e-08,
  -7.709578e-09, -8.179151e-09, -8.360965e-09, -8.505755e-09, -8.628916e-09, 
    -8.978479e-09, -9.16864e-09, -9.459291e-09, -9.687169e-09, -9.798139e-09, 
    -9.844448e-09, -9.968816e-09, -1.016479e-08, -1.050577e-08, -1.075143e-08,
  -1.837232e-08, -1.861519e-08, -1.881903e-08, -1.87351e-08, -1.841164e-08, 
    -1.689689e-08, -1.55302e-08, -1.588462e-08, -1.710766e-08, -1.741335e-08, 
    -1.801917e-08, -1.905254e-08, -2.004142e-08, -2.046678e-08, -2.059348e-08,
  -1.497256e-08, -1.530572e-08, -1.553533e-08, -1.571362e-08, -1.5732e-08, 
    -1.474592e-08, -1.420599e-08, -1.486721e-08, -1.592549e-08, 
    -1.680506e-08, -1.781958e-08, -1.807941e-08, -1.863272e-08, 
    -1.926234e-08, -1.973555e-08,
  -1.220477e-08, -1.244337e-08, -1.297328e-08, -1.363788e-08, -1.397875e-08, 
    -1.4367e-08, -1.43467e-08, -1.491737e-08, -1.558807e-08, -1.685417e-08, 
    -1.782283e-08, -1.804769e-08, -1.817812e-08, -1.820242e-08, -1.836794e-08,
  -9.630881e-09, -9.826335e-09, -1.039786e-08, -1.16375e-08, -1.276832e-08, 
    -1.343489e-08, -1.41451e-08, -1.477257e-08, -1.553911e-08, -1.654337e-08, 
    -1.715693e-08, -1.746224e-08, -1.731925e-08, -1.683562e-08, -1.666617e-08,
  -8.106075e-09, -8.24108e-09, -8.535739e-09, -9.086789e-09, -9.742664e-09, 
    -1.060482e-08, -1.151569e-08, -1.225621e-08, -1.279252e-08, 
    -1.384105e-08, -1.474485e-08, -1.541403e-08, -1.55733e-08, -1.512723e-08, 
    -1.554844e-08,
  -7.413692e-09, -7.484415e-09, -7.619596e-09, -7.87181e-09, -8.155212e-09, 
    -8.475905e-09, -8.842707e-09, -9.19864e-09, -9.664778e-09, -1.000823e-08, 
    -1.033799e-08, -1.085605e-08, -1.162423e-08, -1.23612e-08, -1.295928e-08,
  -7.050634e-09, -7.135903e-09, -7.167118e-09, -7.032198e-09, -7.007213e-09, 
    -7.096183e-09, -7.113409e-09, -7.061006e-09, -6.963574e-09, 
    -7.153774e-09, -7.739803e-09, -8.365551e-09, -9.106846e-09, 
    -9.875756e-09, -1.080086e-08,
  -6.490732e-09, -6.655808e-09, -6.699971e-09, -6.615328e-09, -6.463638e-09, 
    -6.415944e-09, -6.327321e-09, -6.308183e-09, -6.452417e-09, 
    -6.606185e-09, -6.995224e-09, -7.524829e-09, -8.205935e-09, 
    -8.919909e-09, -9.426966e-09,
  -5.771105e-09, -5.822863e-09, -5.89708e-09, -5.975573e-09, -6.037434e-09, 
    -6.076719e-09, -6.171689e-09, -6.183994e-09, -6.48227e-09, -6.879536e-09, 
    -7.208603e-09, -7.603626e-09, -8.038688e-09, -8.338846e-09, -8.598383e-09,
  -4.937264e-09, -5.038311e-09, -5.136176e-09, -5.288624e-09, -5.43742e-09, 
    -5.602485e-09, -5.970691e-09, -6.186102e-09, -6.437441e-09, 
    -6.932559e-09, -7.247862e-09, -7.397796e-09, -7.604902e-09, 
    -7.863838e-09, -8.134112e-09,
  -2.370796e-08, -2.430793e-08, -2.465707e-08, -2.50418e-08, -2.543917e-08, 
    -2.563613e-08, -2.589764e-08, -2.644337e-08, -2.703631e-08, 
    -2.769428e-08, -2.802509e-08, -2.818415e-08, -2.828889e-08, 
    -2.829958e-08, -2.828841e-08,
  -2.078919e-08, -2.161526e-08, -2.224058e-08, -2.279068e-08, -2.334807e-08, 
    -2.363011e-08, -2.39109e-08, -2.433287e-08, -2.475509e-08, -2.522401e-08, 
    -2.551342e-08, -2.577578e-08, -2.601188e-08, -2.625459e-08, -2.64165e-08,
  -1.669215e-08, -1.76504e-08, -1.863588e-08, -1.960079e-08, -2.023784e-08, 
    -2.07594e-08, -2.118097e-08, -2.163598e-08, -2.199284e-08, -2.239636e-08, 
    -2.266469e-08, -2.292231e-08, -2.315637e-08, -2.344178e-08, -2.367913e-08,
  -1.307978e-08, -1.367493e-08, -1.457958e-08, -1.565022e-08, -1.649055e-08, 
    -1.723025e-08, -1.799288e-08, -1.863488e-08, -1.921831e-08, 
    -1.963745e-08, -1.998303e-08, -2.02271e-08, -2.038641e-08, -2.05433e-08, 
    -2.06059e-08,
  -9.594711e-09, -1.049313e-08, -1.154261e-08, -1.252035e-08, -1.316903e-08, 
    -1.37459e-08, -1.446781e-08, -1.527125e-08, -1.593946e-08, -1.655324e-08, 
    -1.691311e-08, -1.716127e-08, -1.729126e-08, -1.733459e-08, -1.724119e-08,
  -6.19504e-09, -7.081129e-09, -8.12759e-09, -9.255372e-09, -1.024799e-08, 
    -1.101634e-08, -1.174852e-08, -1.243172e-08, -1.308697e-08, 
    -1.356337e-08, -1.395327e-08, -1.416009e-08, -1.423272e-08, 
    -1.421977e-08, -1.407387e-08,
  -4.713134e-09, -5.100304e-09, -5.828528e-09, -6.511395e-09, -7.169712e-09, 
    -8.016646e-09, -8.878401e-09, -9.686999e-09, -1.034361e-08, 
    -1.078189e-08, -1.099644e-08, -1.114387e-08, -1.120728e-08, 
    -1.120763e-08, -1.12029e-08,
  -5.055166e-09, -5.028908e-09, -5.21472e-09, -5.388087e-09, -5.701344e-09, 
    -6.356391e-09, -7.107133e-09, -7.728952e-09, -8.211979e-09, -8.4605e-09, 
    -8.528226e-09, -8.558705e-09, -8.574512e-09, -8.570452e-09, -8.603413e-09,
  -5.150859e-09, -5.234239e-09, -5.341783e-09, -5.353869e-09, -5.54406e-09, 
    -5.971339e-09, -6.583933e-09, -6.926898e-09, -6.940962e-09, 
    -6.936882e-09, -6.804771e-09, -6.745401e-09, -6.707082e-09, -6.69535e-09, 
    -6.641725e-09,
  -4.053197e-09, -4.322569e-09, -4.446878e-09, -4.557003e-09, -4.833827e-09, 
    -5.509254e-09, -6.033611e-09, -6.200217e-09, -5.514751e-09, 
    -5.359574e-09, -5.424711e-09, -5.748459e-09, -6.023531e-09, 
    -6.165572e-09, -6.259798e-09,
  -2.219186e-08, -2.213906e-08, -2.246284e-08, -2.309137e-08, -2.358706e-08, 
    -2.384765e-08, -2.396549e-08, -2.412896e-08, -2.429252e-08, 
    -2.452721e-08, -2.480704e-08, -2.500688e-08, -2.525882e-08, -2.55933e-08, 
    -2.586702e-08,
  -2.202216e-08, -2.236838e-08, -2.230479e-08, -2.241107e-08, -2.285929e-08, 
    -2.350541e-08, -2.388331e-08, -2.407057e-08, -2.424147e-08, 
    -2.426609e-08, -2.43731e-08, -2.473169e-08, -2.506552e-08, -2.536241e-08, 
    -2.552351e-08,
  -2.215637e-08, -2.218252e-08, -2.253941e-08, -2.250196e-08, -2.247624e-08, 
    -2.26355e-08, -2.314041e-08, -2.37043e-08, -2.397285e-08, -2.429833e-08, 
    -2.437412e-08, -2.448824e-08, -2.472839e-08, -2.516232e-08, -2.550067e-08,
  -1.982968e-08, -2.137894e-08, -2.213465e-08, -2.252132e-08, -2.273437e-08, 
    -2.279141e-08, -2.264137e-08, -2.283891e-08, -2.344739e-08, 
    -2.389663e-08, -2.428401e-08, -2.447018e-08, -2.462905e-08, 
    -2.490577e-08, -2.537576e-08,
  -1.787803e-08, -1.928826e-08, -2.077643e-08, -2.207567e-08, -2.223746e-08, 
    -2.267596e-08, -2.308463e-08, -2.319501e-08, -2.321767e-08, 
    -2.351074e-08, -2.393244e-08, -2.443112e-08, -2.482853e-08, 
    -2.509019e-08, -2.536414e-08,
  -1.207548e-08, -1.585216e-08, -1.800995e-08, -1.96632e-08, -2.147338e-08, 
    -2.211631e-08, -2.220916e-08, -2.25511e-08, -2.314061e-08, -2.367225e-08, 
    -2.408669e-08, -2.426449e-08, -2.451171e-08, -2.481999e-08, -2.508268e-08,
  -7.419628e-09, -1.009671e-08, -1.337418e-08, -1.615475e-08, -1.802061e-08, 
    -1.977925e-08, -2.147467e-08, -2.196506e-08, -2.185585e-08, 
    -2.199521e-08, -2.275226e-08, -2.355941e-08, -2.430696e-08, 
    -2.474954e-08, -2.49486e-08,
  -7.038195e-09, -7.710339e-09, -9.026025e-09, -1.13116e-08, -1.394049e-08, 
    -1.641919e-08, -1.800144e-08, -1.974734e-08, -2.113703e-08, 
    -2.172091e-08, -2.146023e-08, -2.190058e-08, -2.239996e-08, 
    -2.306759e-08, -2.381713e-08,
  -5.896995e-09, -6.896761e-09, -7.411129e-09, -8.29332e-09, -9.767571e-09, 
    -1.197109e-08, -1.452448e-08, -1.661964e-08, -1.805845e-08, -1.97283e-08, 
    -2.072206e-08, -2.073148e-08, -2.091787e-08, -2.123385e-08, -2.161656e-08,
  -3.600049e-09, -4.659249e-09, -5.56079e-09, -6.403658e-09, -7.033523e-09, 
    -8.504341e-09, -1.067275e-08, -1.27523e-08, -1.430321e-08, -1.610438e-08, 
    -1.769383e-08, -1.901982e-08, -1.945801e-08, -1.91508e-08, -1.940223e-08,
  -1.686735e-08, -1.808865e-08, -2.000484e-08, -2.132634e-08, -2.248634e-08, 
    -2.337912e-08, -2.483608e-08, -2.569589e-08, -2.566798e-08, 
    -2.562831e-08, -2.52837e-08, -2.530187e-08, -2.557194e-08, -2.566629e-08, 
    -2.537691e-08,
  -1.720174e-08, -1.723912e-08, -1.809075e-08, -1.939223e-08, -2.07983e-08, 
    -2.22796e-08, -2.340288e-08, -2.479939e-08, -2.547853e-08, -2.552651e-08, 
    -2.537043e-08, -2.529228e-08, -2.54034e-08, -2.563357e-08, -2.559902e-08,
  -1.965472e-08, -1.792171e-08, -1.749344e-08, -1.812293e-08, -1.907169e-08, 
    -2.036922e-08, -2.17564e-08, -2.318771e-08, -2.457462e-08, -2.53441e-08, 
    -2.55285e-08, -2.52149e-08, -2.513911e-08, -2.536922e-08, -2.558459e-08,
  -1.875761e-08, -1.97026e-08, -1.870415e-08, -1.781247e-08, -1.807378e-08, 
    -1.886859e-08, -1.992692e-08, -2.120349e-08, -2.277451e-08, -2.42379e-08, 
    -2.517031e-08, -2.557857e-08, -2.513688e-08, -2.491673e-08, -2.514149e-08,
  -1.521409e-08, -1.821136e-08, -1.985672e-08, -1.99358e-08, -1.849812e-08, 
    -1.823059e-08, -1.883391e-08, -1.964951e-08, -2.073973e-08, -2.23413e-08, 
    -2.371308e-08, -2.497718e-08, -2.54365e-08, -2.518737e-08, -2.488706e-08,
  -8.898237e-09, -1.354735e-08, -1.690969e-08, -1.887925e-08, -2.009713e-08, 
    -1.928692e-08, -1.859792e-08, -1.886283e-08, -1.943651e-08, 
    -2.036752e-08, -2.174267e-08, -2.318416e-08, -2.438718e-08, 
    -2.517048e-08, -2.525672e-08,
  -6.758194e-09, -8.076955e-09, -1.185974e-08, -1.568378e-08, -1.837615e-08, 
    -2.005623e-08, -2.037546e-08, -1.921966e-08, -1.892742e-08, 
    -1.931553e-08, -2.003788e-08, -2.117903e-08, -2.256048e-08, 
    -2.375906e-08, -2.474504e-08,
  -5.817594e-09, -6.572728e-09, -7.558993e-09, -1.00951e-08, -1.417457e-08, 
    -1.746065e-08, -1.924906e-08, -2.064012e-08, -2.029855e-08, 
    -1.933305e-08, -1.919456e-08, -1.972048e-08, -2.06286e-08, -2.186021e-08, 
    -2.316495e-08,
  -4.42272e-09, -5.189522e-09, -6.06513e-09, -6.970754e-09, -8.71295e-09, 
    -1.255874e-08, -1.620585e-08, -1.834489e-08, -1.987769e-08, 
    -2.088125e-08, -2.017013e-08, -1.933985e-08, -1.953465e-08, 
    -2.012442e-08, -2.10407e-08,
  -3.422735e-09, -3.84616e-09, -4.474091e-09, -5.320877e-09, -5.818795e-09, 
    -7.390236e-09, -1.078739e-08, -1.471724e-08, -1.715603e-08, 
    -1.872344e-08, -2.048677e-08, -2.094985e-08, -2.01225e-08, -1.951356e-08, 
    -1.982636e-08,
  -1.597545e-08, -1.660189e-08, -1.787586e-08, -1.939187e-08, -2.128796e-08, 
    -2.362704e-08, -2.489861e-08, -2.513696e-08, -2.486692e-08, 
    -2.486384e-08, -2.519119e-08, -2.567557e-08, -2.59633e-08, -2.621836e-08, 
    -2.643872e-08,
  -1.653301e-08, -1.618798e-08, -1.662519e-08, -1.747524e-08, -1.884025e-08, 
    -2.059442e-08, -2.310108e-08, -2.463748e-08, -2.5284e-08, -2.53338e-08, 
    -2.497574e-08, -2.524554e-08, -2.559109e-08, -2.610955e-08, -2.639823e-08,
  -1.687903e-08, -1.705441e-08, -1.661536e-08, -1.665236e-08, -1.72706e-08, 
    -1.825781e-08, -1.97971e-08, -2.220965e-08, -2.431627e-08, -2.529284e-08, 
    -2.549255e-08, -2.51785e-08, -2.515189e-08, -2.544441e-08, -2.595589e-08,
  -1.569282e-08, -1.65217e-08, -1.714874e-08, -1.723649e-08, -1.690449e-08, 
    -1.721833e-08, -1.789585e-08, -1.905764e-08, -2.107123e-08, 
    -2.361038e-08, -2.513097e-08, -2.567854e-08, -2.552662e-08, 
    -2.526862e-08, -2.534314e-08,
  -1.433643e-08, -1.528549e-08, -1.603473e-08, -1.684692e-08, -1.745786e-08, 
    -1.730894e-08, -1.737688e-08, -1.779136e-08, -1.865334e-08, 
    -2.009226e-08, -2.255897e-08, -2.467074e-08, -2.559437e-08, 
    -2.570467e-08, -2.552302e-08,
  -1.253376e-08, -1.363852e-08, -1.494083e-08, -1.568671e-08, -1.641819e-08, 
    -1.718302e-08, -1.761978e-08, -1.762892e-08, -1.780047e-08, 
    -1.843654e-08, -1.949608e-08, -2.134388e-08, -2.384716e-08, 
    -2.520619e-08, -2.573049e-08,
  -1.088224e-08, -1.178995e-08, -1.29151e-08, -1.434496e-08, -1.567826e-08, 
    -1.625649e-08, -1.687582e-08, -1.746496e-08, -1.786398e-08, 
    -1.794818e-08, -1.833548e-08, -1.915217e-08, -2.04371e-08, -2.252734e-08, 
    -2.44502e-08,
  -8.325299e-09, -9.764106e-09, -1.08061e-08, -1.189148e-08, -1.33612e-08, 
    -1.518242e-08, -1.625404e-08, -1.663796e-08, -1.714449e-08, 
    -1.767815e-08, -1.808224e-08, -1.827112e-08, -1.889791e-08, 
    -1.985759e-08, -2.13281e-08,
  -5.795375e-09, -6.778223e-09, -8.083862e-09, -9.425157e-09, -1.07241e-08, 
    -1.218395e-08, -1.425133e-08, -1.578282e-08, -1.636719e-08, 
    -1.689797e-08, -1.735624e-08, -1.789874e-08, -1.827713e-08, 
    -1.867197e-08, -1.944884e-08,
  -4.232913e-09, -4.764576e-09, -5.461403e-09, -6.517942e-09, -7.62008e-09, 
    -9.226431e-09, -1.120178e-08, -1.320711e-08, -1.478835e-08, 
    -1.608266e-08, -1.669689e-08, -1.710789e-08, -1.755197e-08, 
    -1.802929e-08, -1.841728e-08,
  -1.86443e-08, -1.957849e-08, -2.040281e-08, -2.133816e-08, -2.214328e-08, 
    -2.29852e-08, -2.36087e-08, -2.419773e-08, -2.452046e-08, -2.485933e-08, 
    -2.510846e-08, -2.505192e-08, -2.484576e-08, -2.44725e-08, -2.423248e-08,
  -1.632713e-08, -1.756316e-08, -1.864333e-08, -1.960367e-08, -2.064145e-08, 
    -2.159897e-08, -2.252446e-08, -2.338215e-08, -2.409981e-08, 
    -2.439772e-08, -2.475219e-08, -2.497982e-08, -2.506135e-08, 
    -2.482251e-08, -2.452526e-08,
  -1.382092e-08, -1.499038e-08, -1.637988e-08, -1.755739e-08, -1.862259e-08, 
    -1.972635e-08, -2.087304e-08, -2.191702e-08, -2.296943e-08, 
    -2.384509e-08, -2.440688e-08, -2.469002e-08, -2.491809e-08, 
    -2.502142e-08, -2.481573e-08,
  -1.149023e-08, -1.241269e-08, -1.36099e-08, -1.502447e-08, -1.635619e-08, 
    -1.758689e-08, -1.87506e-08, -2.002507e-08, -2.124132e-08, -2.24767e-08, 
    -2.353731e-08, -2.437292e-08, -2.478357e-08, -2.496788e-08, -2.503888e-08,
  -9.577478e-09, -1.032902e-08, -1.119084e-08, -1.234857e-08, -1.369234e-08, 
    -1.507062e-08, -1.645572e-08, -1.770829e-08, -1.904091e-08, 
    -2.042225e-08, -2.181022e-08, -2.313631e-08, -2.41529e-08, -2.491315e-08, 
    -2.520386e-08,
  -8.148679e-09, -8.713441e-09, -9.412068e-09, -1.021554e-08, -1.129326e-08, 
    -1.25107e-08, -1.386296e-08, -1.528781e-08, -1.666408e-08, -1.802399e-08, 
    -1.941826e-08, -2.094713e-08, -2.244425e-08, -2.374777e-08, -2.480777e-08,
  -7.075744e-09, -7.602767e-09, -8.134757e-09, -8.723152e-09, -9.473959e-09, 
    -1.043533e-08, -1.154749e-08, -1.283236e-08, -1.418679e-08, 
    -1.563733e-08, -1.706715e-08, -1.84605e-08, -1.996056e-08, -2.161005e-08, 
    -2.312106e-08,
  -5.986037e-09, -6.717448e-09, -7.239537e-09, -7.673272e-09, -8.205858e-09, 
    -8.89249e-09, -9.736067e-09, -1.075478e-08, -1.192994e-08, -1.320679e-08, 
    -1.462756e-08, -1.610869e-08, -1.754185e-08, -1.897881e-08, -2.057344e-08,
  -4.724009e-09, -5.419542e-09, -6.205707e-09, -6.798087e-09, -7.266753e-09, 
    -7.809722e-09, -8.550693e-09, -9.303343e-09, -1.013499e-08, 
    -1.115933e-08, -1.233569e-08, -1.368259e-08, -1.51676e-08, -1.665675e-08, 
    -1.808429e-08,
  -3.624492e-09, -3.998553e-09, -4.596772e-09, -5.460357e-09, -6.106907e-09, 
    -6.817149e-09, -7.575361e-09, -8.354691e-09, -9.025567e-09, 
    -9.752923e-09, -1.058233e-08, -1.161531e-08, -1.282795e-08, 
    -1.421317e-08, -1.567077e-08,
  -2.213919e-08, -2.231249e-08, -2.252489e-08, -2.262022e-08, -2.271754e-08, 
    -2.298004e-08, -2.301018e-08, -2.301584e-08, -2.323631e-08, 
    -2.335166e-08, -2.328965e-08, -2.329685e-08, -2.332986e-08, 
    -2.345072e-08, -2.333529e-08,
  -2.094094e-08, -2.128557e-08, -2.162477e-08, -2.202889e-08, -2.24412e-08, 
    -2.26501e-08, -2.293267e-08, -2.312206e-08, -2.304146e-08, -2.325975e-08, 
    -2.342018e-08, -2.355452e-08, -2.362187e-08, -2.364788e-08, -2.379302e-08,
  -1.946947e-08, -1.999152e-08, -2.040491e-08, -2.074738e-08, -2.121422e-08, 
    -2.175273e-08, -2.226054e-08, -2.270039e-08, -2.302023e-08, 
    -2.311624e-08, -2.318477e-08, -2.332567e-08, -2.349806e-08, 
    -2.363412e-08, -2.381852e-08,
  -1.805288e-08, -1.860249e-08, -1.905633e-08, -1.951983e-08, -1.995641e-08, 
    -2.037252e-08, -2.085338e-08, -2.139006e-08, -2.206726e-08, 
    -2.261048e-08, -2.306987e-08, -2.31195e-08, -2.326042e-08, -2.338933e-08, 
    -2.34703e-08,
  -1.613772e-08, -1.67613e-08, -1.738518e-08, -1.802346e-08, -1.857913e-08, 
    -1.910582e-08, -1.958614e-08, -2.002809e-08, -2.054509e-08, 
    -2.119215e-08, -2.198434e-08, -2.267196e-08, -2.297562e-08, 
    -2.316936e-08, -2.326513e-08,
  -1.325224e-08, -1.419333e-08, -1.522827e-08, -1.616178e-08, -1.693702e-08, 
    -1.751517e-08, -1.807631e-08, -1.86607e-08, -1.919462e-08, -1.970681e-08, 
    -2.033267e-08, -2.111615e-08, -2.198035e-08, -2.260413e-08, -2.290458e-08,
  -1.089152e-08, -1.134237e-08, -1.203353e-08, -1.30052e-08, -1.419806e-08, 
    -1.546294e-08, -1.637199e-08, -1.702785e-08, -1.761271e-08, 
    -1.816917e-08, -1.878391e-08, -1.9431e-08, -2.020262e-08, -2.115106e-08, 
    -2.196154e-08,
  -8.253984e-09, -9.143344e-09, -9.741851e-09, -1.026646e-08, -1.092093e-08, 
    -1.201687e-08, -1.323595e-08, -1.456864e-08, -1.565248e-08, 
    -1.648926e-08, -1.712849e-08, -1.771591e-08, -1.836908e-08, 
    -1.920323e-08, -2.015037e-08,
  -5.556041e-09, -6.28591e-09, -7.096732e-09, -7.911415e-09, -8.594723e-09, 
    -9.276923e-09, -1.0251e-08, -1.120987e-08, -1.231558e-08, -1.371531e-08, 
    -1.490405e-08, -1.594235e-08, -1.659577e-08, -1.7249e-08, -1.804264e-08,
  -3.952304e-09, -4.173696e-09, -4.604727e-09, -5.21315e-09, -5.733634e-09, 
    -6.781058e-09, -7.838956e-09, -8.923353e-09, -9.619448e-09, 
    -1.062269e-08, -1.168198e-08, -1.299609e-08, -1.429026e-08, 
    -1.543021e-08, -1.618089e-08,
  -1.819312e-08, -1.539094e-08, -1.386102e-08, -1.315978e-08, -1.32201e-08, 
    -1.382327e-08, -1.447231e-08, -1.518845e-08, -1.564357e-08, 
    -1.617048e-08, -1.674467e-08, -1.745519e-08, -1.82247e-08, -1.87172e-08, 
    -1.895381e-08,
  -2.360158e-08, -2.053804e-08, -1.690718e-08, -1.466565e-08, -1.39219e-08, 
    -1.383393e-08, -1.420786e-08, -1.463612e-08, -1.517877e-08, 
    -1.573041e-08, -1.642264e-08, -1.713114e-08, -1.785434e-08, 
    -1.856815e-08, -1.899094e-08,
  -2.329781e-08, -2.401729e-08, -2.31408e-08, -1.933704e-08, -1.583905e-08, 
    -1.443647e-08, -1.428879e-08, -1.46865e-08, -1.502678e-08, -1.52644e-08, 
    -1.576455e-08, -1.653039e-08, -1.740951e-08, -1.82814e-08, -1.891893e-08,
  -2.00025e-08, -2.160575e-08, -2.288768e-08, -2.377111e-08, -2.193002e-08, 
    -1.814895e-08, -1.561437e-08, -1.480873e-08, -1.492357e-08, 
    -1.539328e-08, -1.565001e-08, -1.602489e-08, -1.676285e-08, 
    -1.772273e-08, -1.868987e-08,
  -1.731908e-08, -1.838402e-08, -1.979821e-08, -2.151825e-08, -2.281975e-08, 
    -2.313388e-08, -2.040793e-08, -1.763049e-08, -1.590088e-08, 
    -1.536778e-08, -1.560931e-08, -1.595069e-08, -1.642731e-08, 
    -1.712836e-08, -1.8022e-08,
  -1.639338e-08, -1.670538e-08, -1.711716e-08, -1.821327e-08, -1.996283e-08, 
    -2.161516e-08, -2.269613e-08, -2.223142e-08, -1.955126e-08, 
    -1.763531e-08, -1.647919e-08, -1.610209e-08, -1.622575e-08, 
    -1.673173e-08, -1.743275e-08,
  -1.505245e-08, -1.559376e-08, -1.603497e-08, -1.66182e-08, -1.735498e-08, 
    -1.864732e-08, -2.032362e-08, -2.176533e-08, -2.241513e-08, 
    -2.122855e-08, -1.920933e-08, -1.786674e-08, -1.711012e-08, 
    -1.686775e-08, -1.710245e-08,
  -1.32476e-08, -1.356957e-08, -1.425383e-08, -1.500396e-08, -1.582026e-08, 
    -1.656847e-08, -1.763991e-08, -1.915126e-08, -2.072728e-08, 
    -2.195714e-08, -2.201885e-08, -2.064667e-08, -1.91264e-08, -1.816923e-08, 
    -1.775447e-08,
  -1.024009e-08, -1.056118e-08, -1.156151e-08, -1.248374e-08, -1.35002e-08, 
    -1.460105e-08, -1.567207e-08, -1.673931e-08, -1.789611e-08, 
    -1.956316e-08, -2.090408e-08, -2.182106e-08, -2.142033e-08, 
    -2.016118e-08, -1.920699e-08,
  -9.078252e-09, -9.121676e-09, -9.109825e-09, -9.457964e-09, -1.005858e-08, 
    -1.136593e-08, -1.301262e-08, -1.463006e-08, -1.581083e-08, 
    -1.707311e-08, -1.835187e-08, -1.979769e-08, -2.113619e-08, 
    -2.152727e-08, -2.079379e-08,
  -1.413734e-08, -1.387654e-08, -1.40152e-08, -1.437324e-08, -1.467901e-08, 
    -1.492202e-08, -1.531599e-08, -1.565461e-08, -1.579595e-08, 
    -1.593657e-08, -1.62153e-08, -1.662944e-08, -1.713897e-08, -1.789642e-08, 
    -1.824683e-08,
  -1.488478e-08, -1.458336e-08, -1.42904e-08, -1.393465e-08, -1.391871e-08, 
    -1.418364e-08, -1.454036e-08, -1.491728e-08, -1.533282e-08, 
    -1.555351e-08, -1.567293e-08, -1.577743e-08, -1.586901e-08, -1.63089e-08, 
    -1.68233e-08,
  -1.581087e-08, -1.576384e-08, -1.552738e-08, -1.514003e-08, -1.453512e-08, 
    -1.385205e-08, -1.368571e-08, -1.382668e-08, -1.414657e-08, 
    -1.459251e-08, -1.508863e-08, -1.542858e-08, -1.562262e-08, 
    -1.562008e-08, -1.589425e-08,
  -1.689694e-08, -1.680875e-08, -1.697719e-08, -1.692732e-08, -1.671902e-08, 
    -1.609935e-08, -1.504823e-08, -1.402964e-08, -1.355745e-08, 
    -1.345814e-08, -1.365607e-08, -1.40362e-08, -1.449208e-08, -1.484004e-08, 
    -1.51827e-08,
  -1.728388e-08, -1.713234e-08, -1.715473e-08, -1.732984e-08, -1.745272e-08, 
    -1.759069e-08, -1.738282e-08, -1.67758e-08, -1.555017e-08, -1.430383e-08, 
    -1.35908e-08, -1.326533e-08, -1.332569e-08, -1.353475e-08, -1.390769e-08,
  -1.789567e-08, -1.773535e-08, -1.765432e-08, -1.759479e-08, -1.768923e-08, 
    -1.776533e-08, -1.803524e-08, -1.80142e-08, -1.796194e-08, -1.709341e-08, 
    -1.575648e-08, -1.465692e-08, -1.37801e-08, -1.33497e-08, -1.316454e-08,
  -1.799824e-08, -1.808793e-08, -1.811476e-08, -1.808019e-08, -1.8092e-08, 
    -1.806038e-08, -1.818981e-08, -1.820893e-08, -1.834628e-08, 
    -1.844176e-08, -1.818039e-08, -1.717672e-08, -1.59541e-08, -1.497373e-08, 
    -1.423711e-08,
  -1.742317e-08, -1.76966e-08, -1.796003e-08, -1.816383e-08, -1.825609e-08, 
    -1.832664e-08, -1.83537e-08, -1.843401e-08, -1.852059e-08, -1.862643e-08, 
    -1.87373e-08, -1.878618e-08, -1.82223e-08, -1.718431e-08, -1.610479e-08,
  -1.590485e-08, -1.611329e-08, -1.673869e-08, -1.734507e-08, -1.779493e-08, 
    -1.803224e-08, -1.826603e-08, -1.838719e-08, -1.851019e-08, 
    -1.864939e-08, -1.877199e-08, -1.898565e-08, -1.912218e-08, -1.89992e-08, 
    -1.82406e-08,
  -1.358429e-08, -1.355171e-08, -1.384023e-08, -1.44672e-08, -1.524451e-08, 
    -1.601354e-08, -1.672748e-08, -1.720034e-08, -1.755719e-08, 
    -1.797334e-08, -1.836748e-08, -1.875641e-08, -1.913046e-08, 
    -1.947713e-08, -1.965318e-08,
  -1.381734e-08, -1.407483e-08, -1.421526e-08, -1.44721e-08, -1.498751e-08, 
    -1.602884e-08, -1.819145e-08, -1.961385e-08, -2.034942e-08, 
    -2.085381e-08, -2.12819e-08, -2.126827e-08, -2.142857e-08, -2.137993e-08, 
    -2.11867e-08,
  -1.306706e-08, -1.358403e-08, -1.400704e-08, -1.419179e-08, -1.447022e-08, 
    -1.491936e-08, -1.559637e-08, -1.713368e-08, -1.837835e-08, 
    -1.939923e-08, -1.999274e-08, -2.05773e-08, -2.091411e-08, -2.128666e-08, 
    -2.15316e-08,
  -1.248009e-08, -1.281504e-08, -1.34283e-08, -1.388968e-08, -1.411359e-08, 
    -1.442827e-08, -1.479103e-08, -1.531508e-08, -1.640313e-08, 
    -1.748862e-08, -1.855296e-08, -1.921227e-08, -1.967277e-08, 
    -2.019555e-08, -2.068933e-08,
  -1.21449e-08, -1.228926e-08, -1.257332e-08, -1.314438e-08, -1.36776e-08, 
    -1.40645e-08, -1.437581e-08, -1.474257e-08, -1.520961e-08, -1.594719e-08, 
    -1.667167e-08, -1.757309e-08, -1.835976e-08, -1.888075e-08, -1.942553e-08,
  -1.21513e-08, -1.2091e-08, -1.216652e-08, -1.235949e-08, -1.28078e-08, 
    -1.339693e-08, -1.393677e-08, -1.437351e-08, -1.472288e-08, 
    -1.521556e-08, -1.574986e-08, -1.628046e-08, -1.689057e-08, 
    -1.761737e-08, -1.819781e-08,
  -1.259517e-08, -1.209049e-08, -1.194926e-08, -1.199738e-08, -1.213169e-08, 
    -1.248555e-08, -1.301051e-08, -1.367086e-08, -1.424352e-08, 
    -1.471252e-08, -1.515483e-08, -1.558884e-08, -1.60613e-08, -1.644145e-08, 
    -1.697619e-08,
  -1.286266e-08, -1.260435e-08, -1.209047e-08, -1.190506e-08, -1.184908e-08, 
    -1.19498e-08, -1.222108e-08, -1.264195e-08, -1.327838e-08, -1.391985e-08, 
    -1.451888e-08, -1.501603e-08, -1.540666e-08, -1.586677e-08, -1.617755e-08,
  -1.27994e-08, -1.275384e-08, -1.252807e-08, -1.225669e-08, -1.198024e-08, 
    -1.184784e-08, -1.188389e-08, -1.208166e-08, -1.243242e-08, 
    -1.292659e-08, -1.351249e-08, -1.41157e-08, -1.470522e-08, -1.513673e-08, 
    -1.556142e-08,
  -1.263821e-08, -1.264985e-08, -1.25711e-08, -1.242718e-08, -1.236334e-08, 
    -1.217665e-08, -1.1975e-08, -1.188931e-08, -1.202567e-08, -1.230554e-08, 
    -1.270373e-08, -1.316667e-08, -1.368808e-08, -1.42231e-08, -1.469808e-08,
  -1.162651e-08, -1.249331e-08, -1.262993e-08, -1.250071e-08, -1.221321e-08, 
    -1.234857e-08, -1.236285e-08, -1.229464e-08, -1.217132e-08, 
    -1.216383e-08, -1.229449e-08, -1.255457e-08, -1.291463e-08, 
    -1.332068e-08, -1.375688e-08,
  -1.77685e-08, -1.835576e-08, -1.910957e-08, -2.028632e-08, -2.080961e-08, 
    -2.124385e-08, -2.172169e-08, -2.236803e-08, -2.396909e-08, 
    -2.529123e-08, -2.633632e-08, -2.625666e-08, -2.580859e-08, 
    -2.498232e-08, -2.418019e-08,
  -1.638979e-08, -1.699833e-08, -1.76104e-08, -1.829337e-08, -1.91597e-08, 
    -1.978788e-08, -2.040403e-08, -2.109265e-08, -2.180133e-08, -2.29708e-08, 
    -2.448601e-08, -2.552594e-08, -2.58031e-08, -2.572696e-08, -2.545631e-08,
  -1.49137e-08, -1.550652e-08, -1.612186e-08, -1.671608e-08, -1.738497e-08, 
    -1.813678e-08, -1.873511e-08, -1.93947e-08, -2.008103e-08, -2.078486e-08, 
    -2.185036e-08, -2.312072e-08, -2.426547e-08, -2.487e-08, -2.513759e-08,
  -1.372402e-08, -1.413721e-08, -1.460287e-08, -1.521349e-08, -1.577204e-08, 
    -1.641918e-08, -1.709844e-08, -1.766282e-08, -1.826957e-08, 
    -1.893157e-08, -1.966624e-08, -2.066593e-08, -2.171392e-08, 
    -2.274984e-08, -2.360546e-08,
  -1.279004e-08, -1.315455e-08, -1.3524e-08, -1.389471e-08, -1.43807e-08, 
    -1.489505e-08, -1.547455e-08, -1.608566e-08, -1.65727e-08, -1.714414e-08, 
    -1.768041e-08, -1.837222e-08, -1.928455e-08, -2.023384e-08, -2.116139e-08,
  -1.205197e-08, -1.223835e-08, -1.251247e-08, -1.286686e-08, -1.325155e-08, 
    -1.364096e-08, -1.410536e-08, -1.461345e-08, -1.513719e-08, 
    -1.555569e-08, -1.603918e-08, -1.64724e-08, -1.708138e-08, -1.781264e-08, 
    -1.871484e-08,
  -1.133123e-08, -1.154867e-08, -1.171901e-08, -1.193918e-08, -1.221308e-08, 
    -1.263101e-08, -1.302103e-08, -1.340412e-08, -1.384782e-08, 
    -1.428906e-08, -1.466846e-08, -1.501457e-08, -1.53879e-08, -1.585743e-08, 
    -1.645023e-08,
  -1.05042e-08, -1.077751e-08, -1.100622e-08, -1.119492e-08, -1.140732e-08, 
    -1.164298e-08, -1.203474e-08, -1.239907e-08, -1.277881e-08, 
    -1.317334e-08, -1.357748e-08, -1.391803e-08, -1.420053e-08, 
    -1.449071e-08, -1.481002e-08,
  -9.535567e-09, -9.845692e-09, -1.010386e-08, -1.038747e-08, -1.068016e-08, 
    -1.094401e-08, -1.120172e-08, -1.150707e-08, -1.180677e-08, 
    -1.214537e-08, -1.2508e-08, -1.287583e-08, -1.32202e-08, -1.351337e-08, 
    -1.380251e-08,
  -8.240439e-09, -8.68391e-09, -9.026847e-09, -9.317986e-09, -9.594198e-09, 
    -9.988306e-09, -1.045345e-08, -1.078342e-08, -1.10867e-08, -1.134758e-08, 
    -1.164234e-08, -1.192341e-08, -1.222123e-08, -1.250996e-08, -1.279417e-08,
  -1.920345e-08, -1.955272e-08, -2.014206e-08, -2.072404e-08, -2.128711e-08, 
    -2.197804e-08, -2.236707e-08, -2.226636e-08, -2.22921e-08, -2.278436e-08, 
    -2.443137e-08, -2.574669e-08, -2.629001e-08, -2.600265e-08, -2.567413e-08,
  -1.880411e-08, -1.938577e-08, -1.973081e-08, -2.032094e-08, -2.11245e-08, 
    -2.158804e-08, -2.222224e-08, -2.260257e-08, -2.257183e-08, 
    -2.266473e-08, -2.328271e-08, -2.467465e-08, -2.57366e-08, -2.613799e-08, 
    -2.598151e-08,
  -1.835802e-08, -1.868134e-08, -1.919111e-08, -1.958952e-08, -2.031596e-08, 
    -2.124131e-08, -2.179872e-08, -2.22747e-08, -2.259722e-08, -2.271255e-08, 
    -2.296689e-08, -2.359577e-08, -2.466438e-08, -2.555939e-08, -2.596349e-08,
  -1.782452e-08, -1.816232e-08, -1.852666e-08, -1.910056e-08, -1.964918e-08, 
    -2.038854e-08, -2.131425e-08, -2.200926e-08, -2.249909e-08, -2.27226e-08, 
    -2.287673e-08, -2.317765e-08, -2.378288e-08, -2.475694e-08, -2.551609e-08,
  -1.695069e-08, -1.760981e-08, -1.795981e-08, -1.836929e-08, -1.896419e-08, 
    -1.96628e-08, -2.042603e-08, -2.129678e-08, -2.207659e-08, -2.264781e-08, 
    -2.28277e-08, -2.294431e-08, -2.320658e-08, -2.396821e-08, -2.482431e-08,
  -1.649274e-08, -1.677093e-08, -1.735385e-08, -1.765047e-08, -1.80754e-08, 
    -1.872897e-08, -1.947461e-08, -2.032035e-08, -2.119729e-08, 
    -2.201107e-08, -2.261132e-08, -2.290447e-08, -2.29642e-08, -2.329699e-08, 
    -2.411098e-08,
  -1.621535e-08, -1.639832e-08, -1.656671e-08, -1.705286e-08, -1.735626e-08, 
    -1.778547e-08, -1.845611e-08, -1.911832e-08, -1.999621e-08, 
    -2.090182e-08, -2.1709e-08, -2.232925e-08, -2.273351e-08, -2.295618e-08, 
    -2.331139e-08,
  -1.538676e-08, -1.592773e-08, -1.62689e-08, -1.648363e-08, -1.673802e-08, 
    -1.70373e-08, -1.750636e-08, -1.807123e-08, -1.86691e-08, -1.951436e-08, 
    -2.046345e-08, -2.128775e-08, -2.198961e-08, -2.254278e-08, -2.286701e-08,
  -1.389556e-08, -1.480051e-08, -1.554657e-08, -1.610701e-08, -1.653541e-08, 
    -1.672867e-08, -1.687698e-08, -1.716314e-08, -1.751407e-08, 
    -1.801825e-08, -1.879398e-08, -1.97852e-08, -2.066745e-08, -2.15844e-08, 
    -2.221775e-08,
  -1.196346e-08, -1.294637e-08, -1.400651e-08, -1.488593e-08, -1.56071e-08, 
    -1.626711e-08, -1.672825e-08, -1.699719e-08, -1.704143e-08, 
    -1.718353e-08, -1.744118e-08, -1.809734e-08, -1.898629e-08, 
    -2.002644e-08, -2.109644e-08,
  -1.294271e-08, -1.338228e-08, -1.379401e-08, -1.420459e-08, -1.457892e-08, 
    -1.501359e-08, -1.546347e-08, -1.576834e-08, -1.593747e-08, 
    -1.591037e-08, -1.583096e-08, -1.581181e-08, -1.609964e-08, 
    -1.641042e-08, -1.653958e-08,
  -1.253907e-08, -1.294984e-08, -1.338575e-08, -1.369632e-08, -1.408413e-08, 
    -1.450056e-08, -1.514311e-08, -1.567424e-08, -1.605788e-08, 
    -1.619265e-08, -1.630776e-08, -1.634084e-08, -1.64936e-08, -1.677898e-08, 
    -1.703035e-08,
  -1.229206e-08, -1.265869e-08, -1.300531e-08, -1.338007e-08, -1.359617e-08, 
    -1.402326e-08, -1.461074e-08, -1.53781e-08, -1.595264e-08, -1.623562e-08, 
    -1.634066e-08, -1.657099e-08, -1.686751e-08, -1.71123e-08, -1.736934e-08,
  -1.192258e-08, -1.238067e-08, -1.275452e-08, -1.311233e-08, -1.33732e-08, 
    -1.362914e-08, -1.413078e-08, -1.485613e-08, -1.563431e-08, 
    -1.619014e-08, -1.640192e-08, -1.65727e-08, -1.698426e-08, -1.741625e-08, 
    -1.773755e-08,
  -1.150131e-08, -1.203308e-08, -1.256297e-08, -1.293414e-08, -1.321069e-08, 
    -1.342752e-08, -1.378381e-08, -1.434657e-08, -1.504751e-08, 
    -1.578085e-08, -1.634841e-08, -1.664386e-08, -1.691182e-08, 
    -1.739626e-08, -1.794278e-08,
  -1.080427e-08, -1.142783e-08, -1.214109e-08, -1.276422e-08, -1.313446e-08, 
    -1.340278e-08, -1.362922e-08, -1.410681e-08, -1.465849e-08, 
    -1.532871e-08, -1.597976e-08, -1.652345e-08, -1.690652e-08, 
    -1.719396e-08, -1.774364e-08,
  -1.022041e-08, -1.082072e-08, -1.148106e-08, -1.231903e-08, -1.296588e-08, 
    -1.339434e-08, -1.369666e-08, -1.394339e-08, -1.448125e-08, -1.50671e-08, 
    -1.570873e-08, -1.62542e-08, -1.673341e-08, -1.703385e-08, -1.744404e-08,
  -9.423699e-09, -1.00783e-08, -1.066151e-08, -1.15384e-08, -1.243302e-08, 
    -1.319885e-08, -1.377722e-08, -1.424973e-08, -1.448073e-08, 
    -1.501226e-08, -1.56297e-08, -1.615207e-08, -1.660056e-08, -1.682083e-08, 
    -1.706837e-08,
  -8.607066e-09, -9.195639e-09, -9.929431e-09, -1.070541e-08, -1.170622e-08, 
    -1.248894e-08, -1.332975e-08, -1.409588e-08, -1.483701e-08, 
    -1.508381e-08, -1.559609e-08, -1.614351e-08, -1.659456e-08, 
    -1.688284e-08, -1.697452e-08,
  -7.833058e-09, -8.457744e-09, -9.092458e-09, -9.909079e-09, -1.084999e-08, 
    -1.207269e-08, -1.273949e-08, -1.361431e-08, -1.463107e-08, -1.54588e-08, 
    -1.590078e-08, -1.622374e-08, -1.669636e-08, -1.69008e-08, -1.710733e-08,
  -2.100267e-08, -2.086071e-08, -2.080557e-08, -2.08517e-08, -2.07338e-08, 
    -2.044624e-08, -2.032855e-08, -2.020948e-08, -2.020198e-08, 
    -2.025951e-08, -2.01406e-08, -1.996463e-08, -1.959065e-08, -1.947708e-08, 
    -1.947826e-08,
  -2.088958e-08, -2.053576e-08, -2.002062e-08, -1.93285e-08, -1.849295e-08, 
    -1.775344e-08, -1.737406e-08, -1.732273e-08, -1.745872e-08, 
    -1.788881e-08, -1.83189e-08, -1.851753e-08, -1.847417e-08, -1.839274e-08, 
    -1.841298e-08,
  -1.964633e-08, -1.866431e-08, -1.788508e-08, -1.702029e-08, -1.595579e-08, 
    -1.493466e-08, -1.44199e-08, -1.426937e-08, -1.447469e-08, -1.502076e-08, 
    -1.574288e-08, -1.650623e-08, -1.704543e-08, -1.729367e-08, -1.744641e-08,
  -1.646279e-08, -1.514445e-08, -1.447173e-08, -1.369615e-08, -1.259542e-08, 
    -1.188537e-08, -1.154313e-08, -1.146196e-08, -1.164659e-08, 
    -1.206447e-08, -1.280229e-08, -1.379392e-08, -1.4833e-08, -1.571842e-08, 
    -1.632662e-08,
  -1.282738e-08, -1.172349e-08, -1.098218e-08, -1.047493e-08, -9.596979e-09, 
    -9.370067e-09, -9.504287e-09, -9.611715e-09, -9.725722e-09, 
    -9.973097e-09, -1.047851e-08, -1.13293e-08, -1.246167e-08, -1.358361e-08, 
    -1.465382e-08,
  -1.041573e-08, -9.45608e-09, -8.539226e-09, -7.512285e-09, -7.042456e-09, 
    -7.043018e-09, -7.528915e-09, -7.923057e-09, -8.185842e-09, 
    -8.522774e-09, -8.958207e-09, -9.646358e-09, -1.067241e-08, 
    -1.191104e-08, -1.308441e-08,
  -8.126738e-09, -7.743233e-09, -6.958926e-09, -5.444832e-09, -4.83808e-09, 
    -5.235021e-09, -5.789303e-09, -6.33415e-09, -6.675931e-09, -7.088748e-09, 
    -7.584132e-09, -8.229319e-09, -9.100718e-09, -1.028566e-08, -1.157873e-08,
  -6.01203e-09, -5.978227e-09, -5.927643e-09, -5.000723e-09, -3.760667e-09, 
    -3.91536e-09, -4.582135e-09, -5.346398e-09, -5.738418e-09, -5.922855e-09, 
    -6.269423e-09, -6.886529e-09, -7.758561e-09, -8.895224e-09, -1.016381e-08,
  -5.450977e-09, -4.833574e-09, -4.920748e-09, -5.316882e-09, -4.760585e-09, 
    -3.694058e-09, -3.760193e-09, -4.485042e-09, -5.272156e-09, -5.44585e-09, 
    -5.399534e-09, -5.711108e-09, -6.255825e-09, -7.336356e-09, -8.74382e-09,
  -6.423988e-09, -5.780484e-09, -5.297561e-09, -5.63271e-09, -5.807844e-09, 
    -5.083388e-09, -4.697859e-09, -4.616807e-09, -5.063781e-09, 
    -5.390482e-09, -5.422503e-09, -5.281876e-09, -5.424978e-09, 
    -6.010988e-09, -7.206919e-09,
  -2.083133e-08, -2.120341e-08, -2.15767e-08, -2.186346e-08, -2.205852e-08, 
    -2.213476e-08, -2.224502e-08, -2.238696e-08, -2.254203e-08, 
    -2.273511e-08, -2.29336e-08, -2.316976e-08, -2.329234e-08, -2.346009e-08, 
    -2.352475e-08,
  -2.077318e-08, -2.089105e-08, -2.116904e-08, -2.151016e-08, -2.173542e-08, 
    -2.1888e-08, -2.192104e-08, -2.196897e-08, -2.199208e-08, -2.207756e-08, 
    -2.223933e-08, -2.246491e-08, -2.271378e-08, -2.293485e-08, -2.308727e-08,
  -2.038557e-08, -2.050443e-08, -2.060373e-08, -2.08975e-08, -2.11709e-08, 
    -2.135966e-08, -2.144675e-08, -2.145619e-08, -2.143122e-08, -2.14444e-08, 
    -2.154858e-08, -2.168415e-08, -2.18876e-08, -2.203897e-08, -2.207604e-08,
  -1.979809e-08, -1.98985e-08, -2.001975e-08, -2.02789e-08, -2.045551e-08, 
    -2.064962e-08, -2.078501e-08, -2.083602e-08, -2.088866e-08, 
    -2.090955e-08, -2.095403e-08, -2.100966e-08, -2.105272e-08, 
    -2.106091e-08, -2.108465e-08,
  -1.937411e-08, -1.936404e-08, -1.941831e-08, -1.968782e-08, -1.984964e-08, 
    -1.99536e-08, -2.004791e-08, -2.00644e-08, -2.018658e-08, -2.023074e-08, 
    -2.022721e-08, -2.013972e-08, -2.003337e-08, -1.987001e-08, -1.978684e-08,
  -1.94188e-08, -1.927356e-08, -1.930187e-08, -1.926139e-08, -1.930129e-08, 
    -1.929354e-08, -1.933958e-08, -1.936273e-08, -1.941831e-08, 
    -1.945025e-08, -1.949102e-08, -1.948939e-08, -1.949267e-08, 
    -1.951303e-08, -1.953183e-08,
  -1.966781e-08, -1.962022e-08, -1.960848e-08, -1.94483e-08, -1.928944e-08, 
    -1.924313e-08, -1.913268e-08, -1.911241e-08, -1.909032e-08, 
    -1.915533e-08, -1.919182e-08, -1.921137e-08, -1.922058e-08, 
    -1.929136e-08, -1.940856e-08,
  -1.922101e-08, -1.946086e-08, -1.961448e-08, -1.955218e-08, -1.940761e-08, 
    -1.942222e-08, -1.929909e-08, -1.928436e-08, -1.940244e-08, 
    -1.954913e-08, -1.957389e-08, -1.955026e-08, -1.947663e-08, 
    -1.938274e-08, -1.930564e-08,
  -1.829935e-08, -1.858421e-08, -1.878079e-08, -1.897947e-08, -1.911177e-08, 
    -1.919551e-08, -1.932086e-08, -1.941416e-08, -1.960655e-08, 
    -1.975376e-08, -1.965519e-08, -1.949896e-08, -1.928255e-08, 
    -1.909046e-08, -1.888041e-08,
  -1.635975e-08, -1.682102e-08, -1.71338e-08, -1.741584e-08, -1.7523e-08, 
    -1.764651e-08, -1.806002e-08, -1.846249e-08, -1.872391e-08, 
    -1.897892e-08, -1.887757e-08, -1.867759e-08, -1.84377e-08, -1.817339e-08, 
    -1.795485e-08,
  -1.458592e-08, -1.525771e-08, -1.597019e-08, -1.650339e-08, -1.698456e-08, 
    -1.743752e-08, -1.794306e-08, -1.837262e-08, -1.875675e-08, 
    -1.917332e-08, -1.969313e-08, -2.025344e-08, -2.0818e-08, -2.130649e-08, 
    -2.174314e-08,
  -1.45283e-08, -1.513545e-08, -1.585153e-08, -1.652229e-08, -1.716765e-08, 
    -1.763834e-08, -1.805145e-08, -1.849141e-08, -1.892155e-08, 
    -1.933279e-08, -1.974808e-08, -2.018412e-08, -2.064402e-08, -2.10774e-08, 
    -2.153402e-08,
  -1.440683e-08, -1.507757e-08, -1.575596e-08, -1.639032e-08, -1.710813e-08, 
    -1.771549e-08, -1.818242e-08, -1.863607e-08, -1.906373e-08, 
    -1.944639e-08, -1.982495e-08, -2.020398e-08, -2.058838e-08, 
    -2.098849e-08, -2.137431e-08,
  -1.427059e-08, -1.481282e-08, -1.557784e-08, -1.633929e-08, -1.708276e-08, 
    -1.774935e-08, -1.824925e-08, -1.871008e-08, -1.914471e-08, 
    -1.959491e-08, -1.996201e-08, -2.029705e-08, -2.060242e-08, 
    -2.096595e-08, -2.127594e-08,
  -1.445456e-08, -1.469571e-08, -1.516149e-08, -1.596991e-08, -1.68422e-08, 
    -1.769943e-08, -1.831652e-08, -1.880992e-08, -1.919341e-08, 
    -1.959025e-08, -1.997111e-08, -2.031957e-08, -2.064239e-08, 
    -2.097899e-08, -2.127253e-08,
  -1.432081e-08, -1.473123e-08, -1.5086e-08, -1.559546e-08, -1.636013e-08, 
    -1.721154e-08, -1.798754e-08, -1.861635e-08, -1.90316e-08, -1.933835e-08, 
    -1.967672e-08, -1.997471e-08, -2.027659e-08, -2.059519e-08, -2.09346e-08,
  -1.371601e-08, -1.451147e-08, -1.478123e-08, -1.526676e-08, -1.580474e-08, 
    -1.654005e-08, -1.730326e-08, -1.804585e-08, -1.86811e-08, -1.904421e-08, 
    -1.926284e-08, -1.946949e-08, -1.971503e-08, -2.000391e-08, -2.03432e-08,
  -1.334787e-08, -1.404986e-08, -1.448755e-08, -1.487061e-08, -1.528265e-08, 
    -1.586292e-08, -1.656253e-08, -1.735403e-08, -1.805614e-08, 
    -1.855314e-08, -1.878989e-08, -1.89447e-08, -1.911387e-08, -1.93382e-08, 
    -1.962729e-08,
  -1.292117e-08, -1.342146e-08, -1.399384e-08, -1.433355e-08, -1.470101e-08, 
    -1.499716e-08, -1.558457e-08, -1.635069e-08, -1.71144e-08, -1.771363e-08, 
    -1.789556e-08, -1.807027e-08, -1.821108e-08, -1.846454e-08, -1.877508e-08,
  -1.289819e-08, -1.28933e-08, -1.339544e-08, -1.37691e-08, -1.395357e-08, 
    -1.429819e-08, -1.467988e-08, -1.53449e-08, -1.595891e-08, -1.644834e-08, 
    -1.678008e-08, -1.699959e-08, -1.721088e-08, -1.74259e-08, -1.771951e-08,
  -7.083037e-09, -7.093123e-09, -7.042374e-09, -6.940126e-09, -6.825275e-09, 
    -6.747977e-09, -6.686662e-09, -6.651911e-09, -6.603784e-09, 
    -6.556167e-09, -6.522902e-09, -6.577884e-09, -6.798096e-09, 
    -7.089081e-09, -7.498107e-09,
  -7.155899e-09, -7.114735e-09, -7.072577e-09, -6.997774e-09, -6.929418e-09, 
    -6.888766e-09, -6.847707e-09, -6.783128e-09, -6.729974e-09, 
    -6.654299e-09, -6.601268e-09, -6.538094e-09, -6.620366e-09, 
    -6.832323e-09, -7.143281e-09,
  -7.381508e-09, -7.236726e-09, -7.166325e-09, -7.087158e-09, -7.048358e-09, 
    -7.071057e-09, -7.056294e-09, -7.034113e-09, -6.954886e-09, 
    -6.859099e-09, -6.771504e-09, -6.676564e-09, -6.650477e-09, 
    -6.770176e-09, -6.962346e-09,
  -7.66146e-09, -7.430998e-09, -7.274714e-09, -7.177249e-09, -7.118572e-09, 
    -7.168333e-09, -7.235359e-09, -7.225684e-09, -7.249057e-09, 
    -7.152078e-09, -7.086391e-09, -7.006017e-09, -6.918841e-09, 
    -6.901466e-09, -6.98122e-09,
  -7.967187e-09, -7.721317e-09, -7.479833e-09, -7.356645e-09, -7.216705e-09, 
    -7.192033e-09, -7.286302e-09, -7.334161e-09, -7.394072e-09, 
    -7.401113e-09, -7.386275e-09, -7.362502e-09, -7.26941e-09, -7.208234e-09, 
    -7.161608e-09,
  -8.249319e-09, -8.016997e-09, -7.780713e-09, -7.616029e-09, -7.462349e-09, 
    -7.38248e-09, -7.433507e-09, -7.504712e-09, -7.540796e-09, -7.585331e-09, 
    -7.592645e-09, -7.624317e-09, -7.635504e-09, -7.582398e-09, -7.507521e-09,
  -8.405901e-09, -8.24404e-09, -8.024985e-09, -7.809581e-09, -7.670538e-09, 
    -7.529475e-09, -7.524563e-09, -7.571633e-09, -7.604738e-09, 
    -7.678426e-09, -7.771511e-09, -7.854704e-09, -7.909782e-09, 
    -7.903957e-09, -7.855915e-09,
  -8.498554e-09, -8.401056e-09, -8.217155e-09, -8.013372e-09, -7.84211e-09, 
    -7.808174e-09, -7.72788e-09, -7.703343e-09, -7.677523e-09, -7.753667e-09, 
    -7.900659e-09, -8.045053e-09, -8.198049e-09, -8.26229e-09, -8.242138e-09,
  -8.362704e-09, -8.258657e-09, -8.177084e-09, -8.057833e-09, -7.956837e-09, 
    -7.931845e-09, -7.92109e-09, -7.900902e-09, -7.86342e-09, -7.916004e-09, 
    -8.114475e-09, -8.297238e-09, -8.450616e-09, -8.57029e-09, -8.549565e-09,
  -8.365715e-09, -8.184403e-09, -8.075453e-09, -8.058053e-09, -8.048915e-09, 
    -8.109634e-09, -8.068392e-09, -8.085174e-09, -8.081504e-09, 
    -8.200468e-09, -8.377709e-09, -8.584999e-09, -8.712893e-09, 
    -8.860554e-09, -8.914803e-09,
  -1.566623e-08, -1.603258e-08, -1.574581e-08, -1.576167e-08, -1.563449e-08, 
    -1.51927e-08, -1.452899e-08, -1.395803e-08, -1.347743e-08, -1.321821e-08, 
    -1.306285e-08, -1.298076e-08, -1.296448e-08, -1.293804e-08, -1.288925e-08,
  -1.357864e-08, -1.36572e-08, -1.357808e-08, -1.377792e-08, -1.369375e-08, 
    -1.343006e-08, -1.310794e-08, -1.282177e-08, -1.258393e-08, 
    -1.239157e-08, -1.223753e-08, -1.215234e-08, -1.207887e-08, 
    -1.207035e-08, -1.202403e-08,
  -1.19551e-08, -1.190829e-08, -1.18778e-08, -1.191913e-08, -1.184487e-08, 
    -1.172791e-08, -1.162037e-08, -1.150699e-08, -1.141484e-08, -1.13256e-08, 
    -1.121226e-08, -1.111905e-08, -1.108362e-08, -1.113237e-08, -1.116474e-08,
  -1.049766e-08, -1.044524e-08, -1.04175e-08, -1.037984e-08, -1.031237e-08, 
    -1.023832e-08, -1.018962e-08, -1.018003e-08, -1.017354e-08, 
    -1.018542e-08, -1.01709e-08, -1.013979e-08, -1.00803e-08, -1.00772e-08, 
    -1.013749e-08,
  -9.173289e-09, -9.149273e-09, -9.142249e-09, -9.155907e-09, -9.166574e-09, 
    -9.182881e-09, -9.163613e-09, -9.149681e-09, -9.182691e-09, 
    -9.243148e-09, -9.309169e-09, -9.336647e-09, -9.313053e-09, 
    -9.278072e-09, -9.278521e-09,
  -7.922845e-09, -7.973484e-09, -7.998829e-09, -8.071916e-09, -8.135892e-09, 
    -8.228332e-09, -8.275967e-09, -8.297121e-09, -8.316363e-09, -8.39903e-09, 
    -8.515061e-09, -8.613782e-09, -8.662945e-09, -8.692258e-09, -8.684264e-09,
  -6.957433e-09, -7.067266e-09, -7.119879e-09, -7.165644e-09, -7.288097e-09, 
    -7.394138e-09, -7.504764e-09, -7.590208e-09, -7.637376e-09, 
    -7.712329e-09, -7.821505e-09, -7.933992e-09, -8.024662e-09, 
    -8.100327e-09, -8.161027e-09,
  -6.161848e-09, -6.279019e-09, -6.408444e-09, -6.455484e-09, -6.536836e-09, 
    -6.68781e-09, -6.825915e-09, -6.965647e-09, -7.049509e-09, -7.148243e-09, 
    -7.277407e-09, -7.397373e-09, -7.49042e-09, -7.571177e-09, -7.664809e-09,
  -5.540432e-09, -5.66062e-09, -5.798862e-09, -5.913588e-09, -6.000162e-09, 
    -6.108356e-09, -6.269748e-09, -6.413371e-09, -6.551484e-09, 
    -6.666997e-09, -6.82464e-09, -7.001543e-09, -7.11736e-09, -7.223957e-09, 
    -7.334633e-09,
  -4.928312e-09, -5.120294e-09, -5.212411e-09, -5.332709e-09, -5.319951e-09, 
    -5.479141e-09, -5.749533e-09, -5.940512e-09, -6.065903e-09, 
    -6.251632e-09, -6.37542e-09, -6.55867e-09, -6.685356e-09, -6.800651e-09, 
    -6.938293e-09,
  -2.316246e-08, -2.319987e-08, -2.310366e-08, -2.291599e-08, -2.292402e-08, 
    -2.312987e-08, -2.330613e-08, -2.337294e-08, -2.338555e-08, 
    -2.315814e-08, -2.275749e-08, -2.22996e-08, -2.188042e-08, -2.153383e-08, 
    -2.13042e-08,
  -2.28103e-08, -2.256072e-08, -2.250902e-08, -2.240321e-08, -2.228255e-08, 
    -2.217681e-08, -2.20249e-08, -2.190442e-08, -2.170311e-08, -2.145342e-08, 
    -2.119624e-08, -2.090409e-08, -2.061384e-08, -2.029897e-08, -2.002653e-08,
  -2.21664e-08, -2.20971e-08, -2.205424e-08, -2.190306e-08, -2.170705e-08, 
    -2.152238e-08, -2.13631e-08, -2.114204e-08, -2.086032e-08, -2.055501e-08, 
    -2.025536e-08, -1.995032e-08, -1.966271e-08, -1.933397e-08, -1.902641e-08,
  -2.111981e-08, -2.121575e-08, -2.120272e-08, -2.114394e-08, -2.100427e-08, 
    -2.085624e-08, -2.066322e-08, -2.038505e-08, -2.006295e-08, 
    -1.968123e-08, -1.92595e-08, -1.876154e-08, -1.829338e-08, -1.781076e-08, 
    -1.734482e-08,
  -1.960386e-08, -1.96085e-08, -1.962123e-08, -1.953265e-08, -1.947855e-08, 
    -1.933582e-08, -1.910167e-08, -1.877483e-08, -1.837529e-08, 
    -1.790506e-08, -1.736718e-08, -1.680172e-08, -1.622134e-08, 
    -1.562324e-08, -1.511289e-08,
  -1.781177e-08, -1.783464e-08, -1.77903e-08, -1.770582e-08, -1.755417e-08, 
    -1.742633e-08, -1.721497e-08, -1.683388e-08, -1.634893e-08, 
    -1.577902e-08, -1.519261e-08, -1.465043e-08, -1.410624e-08, 
    -1.357568e-08, -1.307128e-08,
  -1.531813e-08, -1.54777e-08, -1.556384e-08, -1.549409e-08, -1.538406e-08, 
    -1.518866e-08, -1.497059e-08, -1.458274e-08, -1.411249e-08, 
    -1.355582e-08, -1.30424e-08, -1.254102e-08, -1.209799e-08, -1.165015e-08, 
    -1.121387e-08,
  -1.240157e-08, -1.277639e-08, -1.299525e-08, -1.304731e-08, -1.29708e-08, 
    -1.280888e-08, -1.255432e-08, -1.217707e-08, -1.172813e-08, 
    -1.128584e-08, -1.087361e-08, -1.050019e-08, -1.015839e-08, 
    -9.837336e-09, -9.51436e-09,
  -9.493809e-09, -9.775698e-09, -1.000118e-08, -1.009642e-08, -1.017208e-08, 
    -1.015027e-08, -1.003676e-08, -9.742395e-09, -9.443057e-09, -9.16018e-09, 
    -8.899508e-09, -8.680882e-09, -8.447277e-09, -8.239911e-09, -8.028856e-09,
  -7.119429e-09, -7.272619e-09, -7.350414e-09, -7.407938e-09, -7.422219e-09, 
    -7.570856e-09, -7.791955e-09, -7.801601e-09, -7.57352e-09, -7.43859e-09, 
    -7.305018e-09, -7.188488e-09, -7.066791e-09, -6.967272e-09, -6.873263e-09,
  -2.519996e-08, -2.502859e-08, -2.48313e-08, -2.482497e-08, -2.477638e-08, 
    -2.45641e-08, -2.43218e-08, -2.409752e-08, -2.399517e-08, -2.392853e-08, 
    -2.395992e-08, -2.395516e-08, -2.396291e-08, -2.387425e-08, -2.373956e-08,
  -2.487038e-08, -2.484368e-08, -2.476343e-08, -2.467206e-08, -2.451917e-08, 
    -2.441524e-08, -2.416078e-08, -2.399558e-08, -2.388425e-08, 
    -2.372516e-08, -2.36629e-08, -2.354953e-08, -2.346851e-08, -2.339801e-08, 
    -2.32958e-08,
  -2.47512e-08, -2.485571e-08, -2.489983e-08, -2.485161e-08, -2.457416e-08, 
    -2.437406e-08, -2.406324e-08, -2.390983e-08, -2.376812e-08, 
    -2.363418e-08, -2.354325e-08, -2.340314e-08, -2.331902e-08, 
    -2.325864e-08, -2.317569e-08,
  -2.464948e-08, -2.459002e-08, -2.454377e-08, -2.469481e-08, -2.464288e-08, 
    -2.448628e-08, -2.4205e-08, -2.39751e-08, -2.377871e-08, -2.36215e-08, 
    -2.344753e-08, -2.334706e-08, -2.316947e-08, -2.301602e-08, -2.283057e-08,
  -2.423744e-08, -2.46901e-08, -2.466728e-08, -2.446e-08, -2.433892e-08, 
    -2.419417e-08, -2.403131e-08, -2.373755e-08, -2.365572e-08, 
    -2.346706e-08, -2.343107e-08, -2.333173e-08, -2.322308e-08, -2.30813e-08, 
    -2.280048e-08,
  -2.432777e-08, -2.404024e-08, -2.44379e-08, -2.470616e-08, -2.449133e-08, 
    -2.431596e-08, -2.413346e-08, -2.387721e-08, -2.371609e-08, 
    -2.353897e-08, -2.346159e-08, -2.338812e-08, -2.330548e-08, 
    -2.307623e-08, -2.264637e-08,
  -2.42686e-08, -2.399385e-08, -2.391036e-08, -2.420714e-08, -2.434387e-08, 
    -2.432861e-08, -2.416319e-08, -2.396555e-08, -2.376597e-08, 
    -2.356249e-08, -2.339316e-08, -2.317033e-08, -2.281257e-08, 
    -2.226297e-08, -2.156802e-08,
  -2.305886e-08, -2.31398e-08, -2.326669e-08, -2.339607e-08, -2.355713e-08, 
    -2.382247e-08, -2.3763e-08, -2.359837e-08, -2.335981e-08, -2.311926e-08, 
    -2.281703e-08, -2.229499e-08, -2.159494e-08, -2.080142e-08, -2.004871e-08,
  -2.152746e-08, -2.164079e-08, -2.205918e-08, -2.205045e-08, -2.22496e-08, 
    -2.235175e-08, -2.249183e-08, -2.236317e-08, -2.201975e-08, 
    -2.183283e-08, -2.144758e-08, -2.084225e-08, -2.011412e-08, 
    -1.944948e-08, -1.881453e-08,
  -2.079921e-08, -2.056324e-08, -2.089628e-08, -2.088802e-08, -2.075942e-08, 
    -2.090952e-08, -2.109609e-08, -2.126478e-08, -2.086453e-08, -2.0672e-08, 
    -2.021054e-08, -1.970852e-08, -1.918641e-08, -1.854582e-08, -1.799367e-08,
  -2.082703e-08, -2.151856e-08, -2.179066e-08, -2.228352e-08, -2.285399e-08, 
    -2.333504e-08, -2.367962e-08, -2.380769e-08, -2.393453e-08, 
    -2.425038e-08, -2.459484e-08, -2.493612e-08, -2.513214e-08, -2.54362e-08, 
    -2.557128e-08,
  -2.062697e-08, -2.144639e-08, -2.190238e-08, -2.215005e-08, -2.264713e-08, 
    -2.342124e-08, -2.383139e-08, -2.394679e-08, -2.40781e-08, -2.433205e-08, 
    -2.459267e-08, -2.492254e-08, -2.519086e-08, -2.533799e-08, -2.547469e-08,
  -2.011619e-08, -2.109591e-08, -2.167033e-08, -2.219786e-08, -2.248438e-08, 
    -2.312126e-08, -2.376483e-08, -2.406145e-08, -2.421817e-08, 
    -2.433311e-08, -2.458235e-08, -2.495672e-08, -2.526745e-08, 
    -2.541297e-08, -2.539179e-08,
  -1.981422e-08, -2.076013e-08, -2.135339e-08, -2.199662e-08, -2.23115e-08, 
    -2.291211e-08, -2.354909e-08, -2.401572e-08, -2.422735e-08, 
    -2.442192e-08, -2.452401e-08, -2.480568e-08, -2.515503e-08, 
    -2.524641e-08, -2.530119e-08,
  -1.937817e-08, -2.034694e-08, -2.097288e-08, -2.16304e-08, -2.227469e-08, 
    -2.272059e-08, -2.352836e-08, -2.411807e-08, -2.434676e-08, -2.4535e-08, 
    -2.467242e-08, -2.480721e-08, -2.507826e-08, -2.511106e-08, -2.512045e-08,
  -1.876342e-08, -1.974504e-08, -2.052181e-08, -2.118051e-08, -2.185594e-08, 
    -2.262375e-08, -2.314192e-08, -2.402681e-08, -2.455757e-08, 
    -2.461171e-08, -2.471407e-08, -2.487972e-08, -2.501301e-08, 
    -2.513575e-08, -2.508013e-08,
  -1.755849e-08, -1.891768e-08, -1.990366e-08, -2.080296e-08, -2.148039e-08, 
    -2.23554e-08, -2.310237e-08, -2.354323e-08, -2.432428e-08, -2.483222e-08, 
    -2.49515e-08, -2.501206e-08, -2.512594e-08, -2.528982e-08, -2.531942e-08,
  -1.595239e-08, -1.767783e-08, -1.892055e-08, -2.024427e-08, -2.098972e-08, 
    -2.183787e-08, -2.283477e-08, -2.372644e-08, -2.415018e-08, 
    -2.457021e-08, -2.498145e-08, -2.518579e-08, -2.527769e-08, 
    -2.528091e-08, -2.544796e-08,
  -1.420167e-08, -1.613e-08, -1.813297e-08, -1.935997e-08, -2.059187e-08, 
    -2.114826e-08, -2.208273e-08, -2.300954e-08, -2.407277e-08, 
    -2.443522e-08, -2.465428e-08, -2.509413e-08, -2.54732e-08, -2.560398e-08, 
    -2.566438e-08,
  -1.228417e-08, -1.444372e-08, -1.668159e-08, -1.833982e-08, -1.953643e-08, 
    -2.084009e-08, -2.151159e-08, -2.22594e-08, -2.311822e-08, -2.387779e-08, 
    -2.427278e-08, -2.437409e-08, -2.475021e-08, -2.501368e-08, -2.516289e-08,
  -1.707718e-08, -1.747105e-08, -1.780662e-08, -1.803582e-08, -1.819667e-08, 
    -1.849939e-08, -1.904392e-08, -1.975914e-08, -2.03561e-08, -2.089002e-08, 
    -2.128581e-08, -2.171855e-08, -2.203929e-08, -2.223326e-08, -2.22753e-08,
  -1.638878e-08, -1.683971e-08, -1.741115e-08, -1.781831e-08, -1.812231e-08, 
    -1.829846e-08, -1.869862e-08, -1.936692e-08, -2.00993e-08, -2.080005e-08, 
    -2.131238e-08, -2.181603e-08, -2.201882e-08, -2.226861e-08, -2.242574e-08,
  -1.57945e-08, -1.611197e-08, -1.668897e-08, -1.722717e-08, -1.767289e-08, 
    -1.794661e-08, -1.829986e-08, -1.884014e-08, -1.95336e-08, -2.031297e-08, 
    -2.094566e-08, -2.157929e-08, -2.192431e-08, -2.220809e-08, -2.238821e-08,
  -1.527069e-08, -1.559769e-08, -1.600085e-08, -1.655928e-08, -1.707059e-08, 
    -1.744733e-08, -1.780673e-08, -1.833809e-08, -1.898931e-08, 
    -1.974377e-08, -2.047832e-08, -2.117845e-08, -2.165193e-08, 
    -2.216844e-08, -2.239075e-08,
  -1.451431e-08, -1.509479e-08, -1.544413e-08, -1.590472e-08, -1.63897e-08, 
    -1.693243e-08, -1.725794e-08, -1.777729e-08, -1.840163e-08, 
    -1.911524e-08, -1.994948e-08, -2.068533e-08, -2.133727e-08, 
    -2.192151e-08, -2.238189e-08,
  -1.356961e-08, -1.419826e-08, -1.486301e-08, -1.532315e-08, -1.579332e-08, 
    -1.632001e-08, -1.670437e-08, -1.718648e-08, -1.785034e-08, 
    -1.855136e-08, -1.932154e-08, -2.015369e-08, -2.088269e-08, 
    -2.160581e-08, -2.21684e-08,
  -1.252109e-08, -1.321696e-08, -1.383188e-08, -1.451029e-08, -1.514885e-08, 
    -1.572863e-08, -1.614568e-08, -1.653538e-08, -1.715229e-08, 
    -1.794365e-08, -1.876547e-08, -1.959193e-08, -2.040031e-08, 
    -2.117612e-08, -2.182886e-08,
  -1.123314e-08, -1.2075e-08, -1.274189e-08, -1.353834e-08, -1.428935e-08, 
    -1.505608e-08, -1.562391e-08, -1.604086e-08, -1.654953e-08, 
    -1.724869e-08, -1.810661e-08, -1.896981e-08, -1.984541e-08, 
    -2.071149e-08, -2.140009e-08,
  -9.803882e-09, -1.065526e-08, -1.160703e-08, -1.245324e-08, -1.337436e-08, 
    -1.412277e-08, -1.474772e-08, -1.53042e-08, -1.588683e-08, -1.664326e-08, 
    -1.746578e-08, -1.828598e-08, -1.913439e-08, -2.003564e-08, -2.091677e-08,
  -8.865171e-09, -9.549598e-09, -1.033021e-08, -1.135835e-08, -1.239035e-08, 
    -1.351307e-08, -1.394938e-08, -1.456059e-08, -1.513956e-08, 
    -1.588836e-08, -1.683294e-08, -1.770291e-08, -1.846656e-08, 
    -1.922319e-08, -2.00953e-08,
  -2.12744e-08, -2.095584e-08, -2.054446e-08, -2.018984e-08, -1.973594e-08, 
    -1.932163e-08, -1.89547e-08, -1.871832e-08, -1.857772e-08, -1.852238e-08, 
    -1.850139e-08, -1.847955e-08, -1.859525e-08, -1.875434e-08, -1.901062e-08,
  -2.068737e-08, -2.036721e-08, -1.977608e-08, -1.931978e-08, -1.881428e-08, 
    -1.837996e-08, -1.802271e-08, -1.776232e-08, -1.756602e-08, 
    -1.755595e-08, -1.75992e-08, -1.76145e-08, -1.76787e-08, -1.789043e-08, 
    -1.814968e-08,
  -2.040785e-08, -1.990089e-08, -1.937745e-08, -1.886932e-08, -1.843827e-08, 
    -1.808349e-08, -1.770369e-08, -1.742225e-08, -1.716987e-08, 
    -1.712348e-08, -1.713697e-08, -1.717438e-08, -1.725814e-08, 
    -1.744879e-08, -1.769074e-08,
  -1.964356e-08, -1.910209e-08, -1.853555e-08, -1.802948e-08, -1.75806e-08, 
    -1.721924e-08, -1.692813e-08, -1.670328e-08, -1.652564e-08, 
    -1.643037e-08, -1.647835e-08, -1.658488e-08, -1.675916e-08, 
    -1.702998e-08, -1.733044e-08,
  -1.8838e-08, -1.835085e-08, -1.78331e-08, -1.740962e-08, -1.701716e-08, 
    -1.671231e-08, -1.644849e-08, -1.618178e-08, -1.595457e-08, 
    -1.581094e-08, -1.581345e-08, -1.592631e-08, -1.613875e-08, 
    -1.645062e-08, -1.688401e-08,
  -1.817834e-08, -1.768321e-08, -1.728273e-08, -1.685796e-08, -1.639068e-08, 
    -1.606296e-08, -1.576079e-08, -1.550023e-08, -1.53011e-08, -1.515586e-08, 
    -1.511366e-08, -1.521241e-08, -1.542281e-08, -1.569305e-08, -1.6159e-08,
  -1.741209e-08, -1.710353e-08, -1.675925e-08, -1.633615e-08, -1.586217e-08, 
    -1.546668e-08, -1.517655e-08, -1.493297e-08, -1.473132e-08, 
    -1.460616e-08, -1.455304e-08, -1.463204e-08, -1.480214e-08, 
    -1.506148e-08, -1.542279e-08,
  -1.664074e-08, -1.637694e-08, -1.606728e-08, -1.563248e-08, -1.507003e-08, 
    -1.469369e-08, -1.442236e-08, -1.421455e-08, -1.406664e-08, 
    -1.396888e-08, -1.391337e-08, -1.396555e-08, -1.414525e-08, 
    -1.438544e-08, -1.472557e-08,
  -1.559625e-08, -1.543172e-08, -1.508236e-08, -1.46594e-08, -1.416978e-08, 
    -1.379838e-08, -1.352884e-08, -1.33361e-08, -1.321327e-08, -1.313744e-08, 
    -1.310251e-08, -1.314036e-08, -1.330052e-08, -1.355439e-08, -1.387306e-08,
  -1.44448e-08, -1.42324e-08, -1.406569e-08, -1.35379e-08, -1.315364e-08, 
    -1.267682e-08, -1.253477e-08, -1.232814e-08, -1.217264e-08, 
    -1.208918e-08, -1.208385e-08, -1.216834e-08, -1.232854e-08, 
    -1.259327e-08, -1.292402e-08,
  -2.653931e-08, -2.697931e-08, -2.747473e-08, -2.792034e-08, -2.815835e-08, 
    -2.83489e-08, -2.856291e-08, -2.863218e-08, -2.857531e-08, -2.830311e-08, 
    -2.784899e-08, -2.75404e-08, -2.711988e-08, -2.627175e-08, -2.48588e-08,
  -2.738253e-08, -2.754519e-08, -2.770159e-08, -2.79468e-08, -2.80641e-08, 
    -2.816641e-08, -2.840787e-08, -2.872915e-08, -2.865783e-08, 
    -2.786435e-08, -2.692162e-08, -2.614862e-08, -2.540482e-08, 
    -2.433192e-08, -2.305847e-08,
  -2.787297e-08, -2.78328e-08, -2.78341e-08, -2.792986e-08, -2.789697e-08, 
    -2.803471e-08, -2.810007e-08, -2.804083e-08, -2.738655e-08, -2.65585e-08, 
    -2.545054e-08, -2.468037e-08, -2.421968e-08, -2.336258e-08, -2.240191e-08,
  -2.827712e-08, -2.803883e-08, -2.793903e-08, -2.799788e-08, -2.808461e-08, 
    -2.804031e-08, -2.782728e-08, -2.749996e-08, -2.692163e-08, 
    -2.601159e-08, -2.507187e-08, -2.420942e-08, -2.34598e-08, -2.246587e-08, 
    -2.155448e-08,
  -2.828332e-08, -2.811141e-08, -2.810844e-08, -2.800752e-08, -2.793785e-08, 
    -2.751046e-08, -2.723859e-08, -2.680945e-08, -2.638898e-08, 
    -2.560545e-08, -2.437067e-08, -2.330834e-08, -2.232605e-08, 
    -2.123647e-08, -2.023212e-08,
  -2.776636e-08, -2.765379e-08, -2.788423e-08, -2.782354e-08, -2.752918e-08, 
    -2.715642e-08, -2.686102e-08, -2.66253e-08, -2.610408e-08, -2.505695e-08, 
    -2.379904e-08, -2.261954e-08, -2.146636e-08, -2.03621e-08, -1.935679e-08,
  -2.716927e-08, -2.713384e-08, -2.762229e-08, -2.795079e-08, -2.73841e-08, 
    -2.669624e-08, -2.64059e-08, -2.621399e-08, -2.55734e-08, -2.450432e-08, 
    -2.326164e-08, -2.214421e-08, -2.08222e-08, -1.977624e-08, -1.882919e-08,
  -2.669667e-08, -2.671621e-08, -2.723068e-08, -2.766878e-08, -2.726037e-08, 
    -2.646762e-08, -2.593302e-08, -2.545988e-08, -2.474935e-08, 
    -2.387998e-08, -2.273911e-08, -2.146634e-08, -2.031198e-08, 
    -1.932789e-08, -1.850448e-08,
  -2.548176e-08, -2.573931e-08, -2.635528e-08, -2.646465e-08, -2.620554e-08, 
    -2.546271e-08, -2.469631e-08, -2.403332e-08, -2.372763e-08, 
    -2.307922e-08, -2.201834e-08, -2.115475e-08, -2.013198e-08, 
    -1.910766e-08, -1.832078e-08,
  -2.402264e-08, -2.392778e-08, -2.48734e-08, -2.553282e-08, -2.526679e-08, 
    -2.412738e-08, -2.338727e-08, -2.293235e-08, -2.277608e-08, 
    -2.212093e-08, -2.132954e-08, -2.060628e-08, -1.950854e-08, 
    -1.864878e-08, -1.780586e-08,
  -2.769162e-08, -2.778599e-08, -2.812362e-08, -2.79592e-08, -2.782172e-08, 
    -2.756978e-08, -2.762595e-08, -2.790305e-08, -2.826271e-08, 
    -2.913685e-08, -3.009037e-08, -3.034038e-08, -3.021456e-08, 
    -3.042554e-08, -3.121357e-08,
  -2.871297e-08, -2.761128e-08, -2.718839e-08, -2.750409e-08, -2.792445e-08, 
    -2.829566e-08, -2.852634e-08, -2.875781e-08, -2.909777e-08, 
    -2.981409e-08, -3.027194e-08, -3.036941e-08, -3.051264e-08, 
    -3.051789e-08, -3.094094e-08,
  -3.068221e-08, -2.929063e-08, -2.800453e-08, -2.720642e-08, -2.713709e-08, 
    -2.722668e-08, -2.760304e-08, -2.814569e-08, -2.881432e-08, 
    -2.983683e-08, -3.001064e-08, -3.048484e-08, -3.027467e-08, 
    -3.005268e-08, -2.996104e-08,
  -3.054968e-08, -3.072576e-08, -3.03318e-08, -2.917715e-08, -2.819074e-08, 
    -2.770748e-08, -2.769908e-08, -2.786445e-08, -2.844942e-08, 
    -2.895086e-08, -2.936452e-08, -3.006611e-08, -2.979023e-08, 
    -2.973202e-08, -2.960073e-08,
  -2.975854e-08, -3.034009e-08, -3.12577e-08, -3.167472e-08, -3.070841e-08, 
    -2.968927e-08, -2.90666e-08, -2.875877e-08, -2.885777e-08, -2.891124e-08, 
    -2.926804e-08, -2.950425e-08, -2.943215e-08, -2.947266e-08, -2.975467e-08,
  -2.715473e-08, -2.859126e-08, -2.948935e-08, -3.034587e-08, -3.065638e-08, 
    -3.049538e-08, -3.029571e-08, -3.016888e-08, -2.979259e-08, 
    -2.972278e-08, -2.951491e-08, -2.98615e-08, -2.967049e-08, -2.984282e-08, 
    -3.00368e-08,
  -2.480911e-08, -2.620709e-08, -2.745345e-08, -2.871412e-08, -2.918048e-08, 
    -2.920777e-08, -2.923603e-08, -2.937056e-08, -2.931692e-08, 
    -2.908208e-08, -2.917728e-08, -2.90634e-08, -2.861157e-08, -2.854753e-08, 
    -2.799286e-08,
  -2.196995e-08, -2.359556e-08, -2.479621e-08, -2.619035e-08, -2.733076e-08, 
    -2.814895e-08, -2.837267e-08, -2.843148e-08, -2.827936e-08, 
    -2.809182e-08, -2.785121e-08, -2.75071e-08, -2.709021e-08, -2.669817e-08, 
    -2.620868e-08,
  -2.01714e-08, -2.105314e-08, -2.217819e-08, -2.325028e-08, -2.444822e-08, 
    -2.573393e-08, -2.685086e-08, -2.763569e-08, -2.786312e-08, 
    -2.777493e-08, -2.744529e-08, -2.695433e-08, -2.605502e-08, 
    -2.553562e-08, -2.614217e-08,
  -1.837866e-08, -1.948611e-08, -2.029126e-08, -2.095717e-08, -2.168882e-08, 
    -2.261375e-08, -2.372841e-08, -2.469773e-08, -2.515409e-08, 
    -2.522534e-08, -2.52718e-08, -2.503222e-08, -2.456745e-08, -2.510449e-08, 
    -2.630523e-08,
  -2.319143e-08, -2.409437e-08, -2.453476e-08, -2.467648e-08, -2.494216e-08, 
    -2.526369e-08, -2.541931e-08, -2.55419e-08, -2.552604e-08, -2.565407e-08, 
    -2.561396e-08, -2.557817e-08, -2.558707e-08, -2.562106e-08, -2.564666e-08,
  -2.1691e-08, -2.259863e-08, -2.324845e-08, -2.380706e-08, -2.411486e-08, 
    -2.444583e-08, -2.474625e-08, -2.494065e-08, -2.511488e-08, 
    -2.521606e-08, -2.544128e-08, -2.553915e-08, -2.556524e-08, 
    -2.563853e-08, -2.570543e-08,
  -2.040797e-08, -2.117664e-08, -2.176403e-08, -2.236542e-08, -2.284087e-08, 
    -2.326883e-08, -2.365262e-08, -2.40463e-08, -2.443917e-08, -2.478933e-08, 
    -2.512944e-08, -2.543168e-08, -2.567551e-08, -2.58232e-08, -2.596174e-08,
  -1.930046e-08, -1.99896e-08, -2.058517e-08, -2.111647e-08, -2.154747e-08, 
    -2.196134e-08, -2.239207e-08, -2.277488e-08, -2.31434e-08, -2.346796e-08, 
    -2.380994e-08, -2.41334e-08, -2.443306e-08, -2.469363e-08, -2.493268e-08,
  -1.81685e-08, -1.889295e-08, -1.944722e-08, -2.016188e-08, -2.067185e-08, 
    -2.109091e-08, -2.148753e-08, -2.190775e-08, -2.220052e-08, 
    -2.252464e-08, -2.272312e-08, -2.294365e-08, -2.314459e-08, 
    -2.332028e-08, -2.366866e-08,
  -1.697516e-08, -1.754105e-08, -1.8122e-08, -1.873877e-08, -1.938763e-08, 
    -2.000784e-08, -2.054034e-08, -2.099364e-08, -2.136091e-08, 
    -2.169487e-08, -2.203654e-08, -2.233798e-08, -2.268619e-08, 
    -2.307269e-08, -2.350365e-08,
  -1.608675e-08, -1.658293e-08, -1.698883e-08, -1.752653e-08, -1.798151e-08, 
    -1.850041e-08, -1.902212e-08, -1.953603e-08, -1.997152e-08, 
    -2.036064e-08, -2.068863e-08, -2.102223e-08, -2.133148e-08, 
    -2.173631e-08, -2.21343e-08,
  -1.49891e-08, -1.549841e-08, -1.605977e-08, -1.652366e-08, -1.691599e-08, 
    -1.730977e-08, -1.766156e-08, -1.805928e-08, -1.845758e-08, 
    -1.887277e-08, -1.92781e-08, -1.969552e-08, -2.008857e-08, -2.043049e-08, 
    -2.070739e-08,
  -1.397002e-08, -1.436417e-08, -1.488849e-08, -1.537512e-08, -1.588906e-08, 
    -1.627094e-08, -1.657963e-08, -1.691426e-08, -1.717565e-08, -1.74995e-08, 
    -1.783417e-08, -1.816648e-08, -1.853242e-08, -1.87744e-08, -1.900779e-08,
  -1.285931e-08, -1.332236e-08, -1.377462e-08, -1.420524e-08, -1.459601e-08, 
    -1.510965e-08, -1.551766e-08, -1.590741e-08, -1.615469e-08, -1.64579e-08, 
    -1.675786e-08, -1.701977e-08, -1.728322e-08, -1.742263e-08, -1.758861e-08,
  -2.840888e-08, -2.824467e-08, -2.804074e-08, -2.788715e-08, -2.765823e-08, 
    -2.750015e-08, -2.740019e-08, -2.720411e-08, -2.714925e-08, 
    -2.702943e-08, -2.69626e-08, -2.679973e-08, -2.666423e-08, -2.647952e-08, 
    -2.629688e-08,
  -2.781928e-08, -2.821071e-08, -2.832856e-08, -2.837501e-08, -2.834099e-08, 
    -2.825965e-08, -2.823366e-08, -2.808972e-08, -2.80289e-08, -2.786547e-08, 
    -2.77872e-08, -2.770996e-08, -2.75954e-08, -2.747442e-08, -2.728902e-08,
  -2.572157e-08, -2.636067e-08, -2.69632e-08, -2.741077e-08, -2.770823e-08, 
    -2.788318e-08, -2.797927e-08, -2.800105e-08, -2.797499e-08, 
    -2.792856e-08, -2.788645e-08, -2.787061e-08, -2.782104e-08, 
    -2.778724e-08, -2.769117e-08,
  -2.34969e-08, -2.379071e-08, -2.408452e-08, -2.447064e-08, -2.477327e-08, 
    -2.49622e-08, -2.512825e-08, -2.523881e-08, -2.525942e-08, -2.524096e-08, 
    -2.516654e-08, -2.50726e-08, -2.491793e-08, -2.47505e-08, -2.453597e-08,
  -2.209515e-08, -2.223855e-08, -2.222747e-08, -2.232037e-08, -2.238096e-08, 
    -2.233591e-08, -2.23199e-08, -2.225999e-08, -2.221591e-08, -2.208582e-08, 
    -2.195114e-08, -2.176908e-08, -2.155122e-08, -2.133285e-08, -2.109684e-08,
  -2.100908e-08, -2.095631e-08, -2.089473e-08, -2.075824e-08, -2.069493e-08, 
    -2.056401e-08, -2.046488e-08, -2.036564e-08, -2.028321e-08, 
    -2.019335e-08, -2.008662e-08, -2.001149e-08, -1.989927e-08, 
    -1.978156e-08, -1.96786e-08,
  -1.970709e-08, -1.963065e-08, -1.941129e-08, -1.931334e-08, -1.919902e-08, 
    -1.893244e-08, -1.892394e-08, -1.885724e-08, -1.88989e-08, -1.891672e-08, 
    -1.896535e-08, -1.898794e-08, -1.901068e-08, -1.902661e-08, -1.904109e-08,
  -1.98543e-08, -1.964025e-08, -1.945022e-08, -1.932824e-08, -1.910688e-08, 
    -1.893432e-08, -1.882345e-08, -1.879233e-08, -1.882377e-08, -1.88916e-08, 
    -1.893759e-08, -1.895699e-08, -1.892435e-08, -1.885048e-08, -1.876034e-08,
  -1.967317e-08, -1.955287e-08, -1.938452e-08, -1.924759e-08, -1.913469e-08, 
    -1.894842e-08, -1.882705e-08, -1.8757e-08, -1.871523e-08, -1.86831e-08, 
    -1.857889e-08, -1.842513e-08, -1.821355e-08, -1.797968e-08, -1.769611e-08,
  -1.854883e-08, -1.868058e-08, -1.873408e-08, -1.862035e-08, -1.83591e-08, 
    -1.805654e-08, -1.822635e-08, -1.80842e-08, -1.791808e-08, -1.765227e-08, 
    -1.726107e-08, -1.681796e-08, -1.633302e-08, -1.581656e-08, -1.529473e-08,
  -2.84617e-08, -2.778992e-08, -2.821044e-08, -2.806285e-08, -2.774432e-08, 
    -2.75569e-08, -2.752838e-08, -2.750019e-08, -2.745008e-08, -2.735634e-08, 
    -2.731458e-08, -2.732043e-08, -2.727065e-08, -2.716679e-08, -2.701903e-08,
  -2.818222e-08, -2.761067e-08, -2.781368e-08, -2.766633e-08, -2.75875e-08, 
    -2.742165e-08, -2.744739e-08, -2.743141e-08, -2.742402e-08, -2.74215e-08, 
    -2.745963e-08, -2.744656e-08, -2.746213e-08, -2.741668e-08, -2.741678e-08,
  -2.81583e-08, -2.769868e-08, -2.778395e-08, -2.775572e-08, -2.774721e-08, 
    -2.776788e-08, -2.779204e-08, -2.775088e-08, -2.772922e-08, 
    -2.771376e-08, -2.770574e-08, -2.769907e-08, -2.770454e-08, 
    -2.771521e-08, -2.772437e-08,
  -2.810023e-08, -2.797024e-08, -2.80848e-08, -2.826667e-08, -2.82969e-08, 
    -2.82885e-08, -2.822326e-08, -2.816131e-08, -2.810405e-08, -2.803794e-08, 
    -2.79199e-08, -2.773017e-08, -2.748933e-08, -2.722726e-08, -2.697932e-08,
  -2.845514e-08, -2.868037e-08, -2.832178e-08, -2.801765e-08, -2.784788e-08, 
    -2.775316e-08, -2.756039e-08, -2.732885e-08, -2.707161e-08, 
    -2.672255e-08, -2.634202e-08, -2.592692e-08, -2.551985e-08, 
    -2.507904e-08, -2.466248e-08,
  -2.862656e-08, -2.86379e-08, -2.829084e-08, -2.775399e-08, -2.734265e-08, 
    -2.697695e-08, -2.642474e-08, -2.583548e-08, -2.51589e-08, -2.450854e-08, 
    -2.388635e-08, -2.333415e-08, -2.285657e-08, -2.248492e-08, -2.222092e-08,
  -2.782773e-08, -2.775215e-08, -2.700684e-08, -2.6523e-08, -2.579058e-08, 
    -2.504639e-08, -2.428119e-08, -2.360457e-08, -2.298119e-08, 
    -2.244782e-08, -2.206837e-08, -2.183439e-08, -2.173259e-08, -2.17851e-08, 
    -2.192797e-08,
  -2.597976e-08, -2.562434e-08, -2.497662e-08, -2.440401e-08, -2.367288e-08, 
    -2.3064e-08, -2.259636e-08, -2.223394e-08, -2.203878e-08, -2.200511e-08, 
    -2.209767e-08, -2.228063e-08, -2.250445e-08, -2.266424e-08, -2.271012e-08,
  -2.389801e-08, -2.35799e-08, -2.31679e-08, -2.270708e-08, -2.239996e-08, 
    -2.21303e-08, -2.20306e-08, -2.203832e-08, -2.214024e-08, -2.227387e-08, 
    -2.234175e-08, -2.236645e-08, -2.231377e-08, -2.214478e-08, -2.176139e-08,
  -2.261156e-08, -2.25585e-08, -2.230655e-08, -2.215081e-08, -2.196371e-08, 
    -2.172327e-08, -2.197546e-08, -2.211975e-08, -2.206345e-08, 
    -2.188576e-08, -2.16603e-08, -2.130536e-08, -2.064509e-08, -1.967536e-08, 
    -1.852872e-08,
  -2.732809e-08, -2.685312e-08, -2.707593e-08, -2.72769e-08, -2.70267e-08, 
    -2.678931e-08, -2.640284e-08, -2.610981e-08, -2.58752e-08, -2.570485e-08, 
    -2.543361e-08, -2.505809e-08, -2.468155e-08, -2.452239e-08, -2.447686e-08,
  -2.66445e-08, -2.628437e-08, -2.657529e-08, -2.673193e-08, -2.640055e-08, 
    -2.591569e-08, -2.559335e-08, -2.557904e-08, -2.551954e-08, 
    -2.530893e-08, -2.511569e-08, -2.497002e-08, -2.493365e-08, 
    -2.486863e-08, -2.488238e-08,
  -2.563448e-08, -2.568935e-08, -2.533987e-08, -2.533315e-08, -2.541712e-08, 
    -2.529748e-08, -2.515415e-08, -2.508231e-08, -2.519071e-08, 
    -2.523049e-08, -2.527705e-08, -2.5351e-08, -2.543569e-08, -2.554494e-08, 
    -2.562707e-08,
  -2.474222e-08, -2.507913e-08, -2.513342e-08, -2.494523e-08, -2.516725e-08, 
    -2.514154e-08, -2.514824e-08, -2.516617e-08, -2.53532e-08, -2.55888e-08, 
    -2.578228e-08, -2.591569e-08, -2.605635e-08, -2.615342e-08, -2.621974e-08,
  -2.498914e-08, -2.489227e-08, -2.457695e-08, -2.472547e-08, -2.523007e-08, 
    -2.551476e-08, -2.585177e-08, -2.600383e-08, -2.630578e-08, 
    -2.661499e-08, -2.682218e-08, -2.693462e-08, -2.692621e-08, 
    -2.683289e-08, -2.665566e-08,
  -2.443632e-08, -2.552202e-08, -2.563601e-08, -2.500673e-08, -2.504975e-08, 
    -2.546982e-08, -2.594123e-08, -2.640588e-08, -2.671974e-08, 
    -2.686385e-08, -2.691999e-08, -2.68604e-08, -2.671344e-08, -2.65117e-08, 
    -2.62789e-08,
  -2.45757e-08, -2.528155e-08, -2.586787e-08, -2.627428e-08, -2.644003e-08, 
    -2.661109e-08, -2.6832e-08, -2.693177e-08, -2.694418e-08, -2.687108e-08, 
    -2.667298e-08, -2.635583e-08, -2.595443e-08, -2.55187e-08, -2.515569e-08,
  -2.553625e-08, -2.558583e-08, -2.555615e-08, -2.641392e-08, -2.696513e-08, 
    -2.705578e-08, -2.686879e-08, -2.677475e-08, -2.649781e-08, 
    -2.607013e-08, -2.551581e-08, -2.499324e-08, -2.457873e-08, 
    -2.424932e-08, -2.388898e-08,
  -2.611823e-08, -2.641446e-08, -2.644193e-08, -2.612363e-08, -2.611759e-08, 
    -2.594048e-08, -2.580175e-08, -2.563877e-08, -2.519083e-08, 
    -2.468435e-08, -2.421513e-08, -2.390843e-08, -2.359107e-08, 
    -2.312724e-08, -2.25506e-08,
  -2.590361e-08, -2.642536e-08, -2.676368e-08, -2.685791e-08, -2.723072e-08, 
    -2.693321e-08, -2.530296e-08, -2.450527e-08, -2.408212e-08, 
    -2.362576e-08, -2.330417e-08, -2.285329e-08, -2.23084e-08, -2.145757e-08, 
    -2.03466e-08,
  -1.673437e-08, -1.7519e-08, -1.834952e-08, -1.902179e-08, -1.955569e-08, 
    -2.03754e-08, -2.1179e-08, -2.224892e-08, -2.287812e-08, -2.341464e-08, 
    -2.408211e-08, -2.450245e-08, -2.475198e-08, -2.459725e-08, -2.473729e-08,
  -1.728203e-08, -1.802199e-08, -1.894336e-08, -1.95198e-08, -2.004213e-08, 
    -2.085038e-08, -2.160707e-08, -2.254824e-08, -2.340518e-08, 
    -2.397306e-08, -2.446721e-08, -2.480339e-08, -2.48708e-08, -2.456165e-08, 
    -2.434995e-08,
  -1.787984e-08, -1.860853e-08, -1.952164e-08, -2.013134e-08, -2.070256e-08, 
    -2.138627e-08, -2.20179e-08, -2.285955e-08, -2.36382e-08, -2.408115e-08, 
    -2.434974e-08, -2.454323e-08, -2.462844e-08, -2.452991e-08, -2.41833e-08,
  -1.877491e-08, -1.949578e-08, -2.034522e-08, -2.08728e-08, -2.131166e-08, 
    -2.190979e-08, -2.25662e-08, -2.318798e-08, -2.369704e-08, -2.407551e-08, 
    -2.423939e-08, -2.435451e-08, -2.449345e-08, -2.458579e-08, -2.45363e-08,
  -1.939011e-08, -2.024961e-08, -2.133251e-08, -2.177508e-08, -2.210688e-08, 
    -2.264996e-08, -2.299631e-08, -2.343283e-08, -2.382271e-08, 
    -2.415108e-08, -2.436893e-08, -2.459079e-08, -2.490787e-08, -2.52061e-08, 
    -2.547809e-08,
  -1.978238e-08, -2.091341e-08, -2.172897e-08, -2.217319e-08, -2.236367e-08, 
    -2.293945e-08, -2.364598e-08, -2.401579e-08, -2.44453e-08, -2.486705e-08, 
    -2.525931e-08, -2.546861e-08, -2.572968e-08, -2.600135e-08, -2.60395e-08,
  -2.030655e-08, -2.127701e-08, -2.228305e-08, -2.252276e-08, -2.28772e-08, 
    -2.330197e-08, -2.385959e-08, -2.44931e-08, -2.515979e-08, -2.584814e-08, 
    -2.616042e-08, -2.610873e-08, -2.610634e-08, -2.625054e-08, -2.611811e-08,
  -2.049057e-08, -2.073742e-08, -2.170053e-08, -2.301195e-08, -2.330964e-08, 
    -2.39556e-08, -2.469367e-08, -2.554527e-08, -2.601846e-08, -2.637355e-08, 
    -2.666657e-08, -2.689308e-08, -2.675901e-08, -2.654106e-08, -2.626561e-08,
  -1.983831e-08, -2.07221e-08, -2.125582e-08, -2.238279e-08, -2.357e-08, 
    -2.419575e-08, -2.501199e-08, -2.556786e-08, -2.639521e-08, -2.67812e-08, 
    -2.713463e-08, -2.710391e-08, -2.691703e-08, -2.662927e-08, -2.635962e-08,
  -1.972268e-08, -2.064127e-08, -2.275466e-08, -2.364982e-08, -2.510793e-08, 
    -2.633714e-08, -2.475787e-08, -2.516899e-08, -2.610635e-08, 
    -2.700844e-08, -2.715559e-08, -2.719464e-08, -2.695676e-08, 
    -2.680468e-08, -2.659099e-08,
  -9.48911e-09, -9.571104e-09, -9.545241e-09, -9.562558e-09, -9.587533e-09, 
    -9.689845e-09, -9.731908e-09, -9.722017e-09, -9.763687e-09, 
    -9.954455e-09, -1.014527e-08, -1.034861e-08, -1.068342e-08, 
    -1.098174e-08, -1.139558e-08,
  -9.776025e-09, -9.663306e-09, -9.661706e-09, -9.660658e-09, -9.766978e-09, 
    -9.924831e-09, -1.000401e-08, -1.000746e-08, -9.901312e-09, 
    -9.897144e-09, -1.004921e-08, -1.020497e-08, -1.046894e-08, 
    -1.076112e-08, -1.113415e-08,
  -1.013263e-08, -9.921814e-09, -9.835568e-09, -9.864979e-09, -9.919771e-09, 
    -1.005961e-08, -1.016841e-08, -1.022153e-08, -1.018136e-08, 
    -1.006538e-08, -1.009722e-08, -1.02354e-08, -1.044877e-08, -1.066657e-08, 
    -1.093903e-08,
  -1.032519e-08, -1.022319e-08, -1.003606e-08, -1.004248e-08, -1.009099e-08, 
    -1.023002e-08, -1.041644e-08, -1.051161e-08, -1.051143e-08, 
    -1.047871e-08, -1.044106e-08, -1.043472e-08, -1.056636e-08, 
    -1.080363e-08, -1.10632e-08,
  -1.080908e-08, -1.055636e-08, -1.032126e-08, -1.024495e-08, -1.019126e-08, 
    -1.022396e-08, -1.031825e-08, -1.0468e-08, -1.05585e-08, -1.058835e-08, 
    -1.057152e-08, -1.060446e-08, -1.065037e-08, -1.094494e-08, -1.118257e-08,
  -1.078562e-08, -1.08037e-08, -1.071784e-08, -1.056834e-08, -1.04527e-08, 
    -1.046329e-08, -1.048798e-08, -1.042856e-08, -1.044034e-08, 
    -1.044576e-08, -1.048778e-08, -1.05525e-08, -1.077044e-08, -1.099726e-08, 
    -1.139634e-08,
  -1.119116e-08, -1.113528e-08, -1.095113e-08, -1.09573e-08, -1.076902e-08, 
    -1.061555e-08, -1.060656e-08, -1.060482e-08, -1.064243e-08, 
    -1.062604e-08, -1.062064e-08, -1.066908e-08, -1.076113e-08, 
    -1.097682e-08, -1.142951e-08,
  -1.250302e-08, -1.215201e-08, -1.179824e-08, -1.175984e-08, -1.156723e-08, 
    -1.130035e-08, -1.122258e-08, -1.110696e-08, -1.106024e-08, 
    -1.109975e-08, -1.117354e-08, -1.125542e-08, -1.12708e-08, -1.145831e-08, 
    -1.183168e-08,
  -1.328896e-08, -1.325329e-08, -1.351623e-08, -1.317544e-08, -1.270502e-08, 
    -1.239742e-08, -1.271263e-08, -1.294427e-08, -1.309601e-08, 
    -1.304126e-08, -1.300307e-08, -1.298418e-08, -1.294461e-08, 
    -1.291094e-08, -1.316679e-08,
  -1.351555e-08, -1.423761e-08, -1.48482e-08, -1.51069e-08, -1.480234e-08, 
    -1.452218e-08, -1.33399e-08, -1.3387e-08, -1.369877e-08, -1.421548e-08, 
    -1.470541e-08, -1.517022e-08, -1.546452e-08, -1.558283e-08, -1.56905e-08,
  -1.124874e-08, -1.133999e-08, -1.142735e-08, -1.142223e-08, -1.139741e-08, 
    -1.130856e-08, -1.126665e-08, -1.125429e-08, -1.131051e-08, -1.13993e-08, 
    -1.15277e-08, -1.16663e-08, -1.18289e-08, -1.195838e-08, -1.208073e-08,
  -1.096044e-08, -1.108887e-08, -1.104497e-08, -1.098038e-08, -1.094872e-08, 
    -1.088971e-08, -1.088237e-08, -1.091417e-08, -1.097028e-08, 
    -1.102503e-08, -1.10848e-08, -1.114458e-08, -1.119619e-08, -1.122747e-08, 
    -1.123753e-08,
  -1.071201e-08, -1.074344e-08, -1.069215e-08, -1.061327e-08, -1.057873e-08, 
    -1.052871e-08, -1.052781e-08, -1.054517e-08, -1.057903e-08, 
    -1.061536e-08, -1.064558e-08, -1.06599e-08, -1.065549e-08, -1.062002e-08, 
    -1.057351e-08,
  -1.047083e-08, -1.052205e-08, -1.048132e-08, -1.04192e-08, -1.036802e-08, 
    -1.031176e-08, -1.030159e-08, -1.02894e-08, -1.029614e-08, -1.028903e-08, 
    -1.030334e-08, -1.029253e-08, -1.026252e-08, -1.021381e-08, -1.013792e-08,
  -1.005326e-08, -1.010347e-08, -1.010139e-08, -1.006727e-08, -1.00325e-08, 
    -1.000282e-08, -9.982177e-09, -9.986502e-09, -9.992236e-09, 
    -1.000136e-08, -1.000331e-08, -1.000707e-08, -9.991822e-09, 
    -9.973303e-09, -9.908399e-09,
  -9.828188e-09, -9.852655e-09, -9.868683e-09, -9.856294e-09, -9.801919e-09, 
    -9.806421e-09, -9.840542e-09, -9.890114e-09, -9.93634e-09, -9.940091e-09, 
    -9.938337e-09, -9.943864e-09, -9.942402e-09, -9.933387e-09, -9.907488e-09,
  -9.546385e-09, -9.594037e-09, -9.600584e-09, -9.642721e-09, -9.637238e-09, 
    -9.733832e-09, -9.852243e-09, -9.954078e-09, -9.969887e-09, 
    -9.958537e-09, -9.925574e-09, -9.923824e-09, -9.94248e-09, -9.935194e-09, 
    -9.934372e-09,
  -9.378581e-09, -9.441399e-09, -9.461449e-09, -9.550226e-09, -9.671026e-09, 
    -9.820444e-09, -9.919724e-09, -9.996857e-09, -1.000398e-08, 
    -9.980092e-09, -9.961337e-09, -9.98081e-09, -9.984847e-09, -1.002727e-08, 
    -1.000509e-08,
  -9.180667e-09, -9.247485e-09, -9.348513e-09, -9.487104e-09, -9.660755e-09, 
    -9.825097e-09, -9.913235e-09, -1.002025e-08, -1.011475e-08, 
    -1.024589e-08, -1.03755e-08, -1.053596e-08, -1.066035e-08, -1.073003e-08, 
    -1.074122e-08,
  -8.889332e-09, -9.114117e-09, -9.243295e-09, -9.524139e-09, -9.728792e-09, 
    -1.020189e-08, -1.01622e-08, -1.027647e-08, -1.044004e-08, -1.057408e-08, 
    -1.074147e-08, -1.094969e-08, -1.126018e-08, -1.158978e-08, -1.188856e-08,
  -1.702127e-08, -1.672818e-08, -1.661357e-08, -1.653824e-08, -1.642541e-08, 
    -1.60966e-08, -1.576549e-08, -1.537817e-08, -1.502653e-08, -1.474899e-08, 
    -1.455346e-08, -1.445383e-08, -1.441604e-08, -1.442536e-08, -1.446031e-08,
  -1.677632e-08, -1.657978e-08, -1.635954e-08, -1.630615e-08, -1.604052e-08, 
    -1.564648e-08, -1.52004e-08, -1.478349e-08, -1.442447e-08, -1.411408e-08, 
    -1.392106e-08, -1.381557e-08, -1.379839e-08, -1.382617e-08, -1.389239e-08,
  -1.661149e-08, -1.638929e-08, -1.620085e-08, -1.61173e-08, -1.587171e-08, 
    -1.537609e-08, -1.487258e-08, -1.4452e-08, -1.40531e-08, -1.375255e-08, 
    -1.350021e-08, -1.335584e-08, -1.326878e-08, -1.323185e-08, -1.324084e-08,
  -1.627993e-08, -1.610303e-08, -1.590672e-08, -1.576807e-08, -1.548845e-08, 
    -1.499544e-08, -1.454213e-08, -1.414176e-08, -1.381861e-08, 
    -1.349368e-08, -1.325112e-08, -1.308831e-08, -1.298711e-08, 
    -1.293538e-08, -1.2886e-08,
  -1.557791e-08, -1.542887e-08, -1.519172e-08, -1.50161e-08, -1.467277e-08, 
    -1.427804e-08, -1.389109e-08, -1.355161e-08, -1.32739e-08, -1.301498e-08, 
    -1.282784e-08, -1.270255e-08, -1.26336e-08, -1.259466e-08, -1.256763e-08,
  -1.492007e-08, -1.480222e-08, -1.46453e-08, -1.440667e-08, -1.400638e-08, 
    -1.366751e-08, -1.333713e-08, -1.30428e-08, -1.278647e-08, -1.258216e-08, 
    -1.242962e-08, -1.233681e-08, -1.230381e-08, -1.228372e-08, -1.227277e-08,
  -1.412877e-08, -1.400516e-08, -1.384935e-08, -1.363684e-08, -1.329105e-08, 
    -1.294853e-08, -1.269847e-08, -1.245205e-08, -1.224929e-08, 
    -1.210496e-08, -1.197544e-08, -1.191555e-08, -1.19073e-08, -1.191168e-08, 
    -1.193102e-08,
  -1.331891e-08, -1.317748e-08, -1.306104e-08, -1.293352e-08, -1.268083e-08, 
    -1.240547e-08, -1.219915e-08, -1.2013e-08, -1.185844e-08, -1.172542e-08, 
    -1.163627e-08, -1.158017e-08, -1.15902e-08, -1.16206e-08, -1.16722e-08,
  -1.247625e-08, -1.240611e-08, -1.234021e-08, -1.222605e-08, -1.206002e-08, 
    -1.186489e-08, -1.166496e-08, -1.153703e-08, -1.141304e-08, 
    -1.133892e-08, -1.129009e-08, -1.124373e-08, -1.124099e-08, 
    -1.128574e-08, -1.135941e-08,
  -1.153651e-08, -1.148677e-08, -1.154494e-08, -1.151062e-08, -1.141312e-08, 
    -1.131049e-08, -1.115573e-08, -1.099486e-08, -1.096648e-08, 
    -1.092467e-08, -1.091204e-08, -1.08961e-08, -1.088148e-08, -1.092673e-08, 
    -1.098796e-08,
  -2.026734e-08, -2.050359e-08, -2.07233e-08, -2.09228e-08, -2.11068e-08, 
    -2.131721e-08, -2.145937e-08, -2.163038e-08, -2.172156e-08, 
    -2.171927e-08, -2.164457e-08, -2.148371e-08, -2.121164e-08, 
    -2.108174e-08, -2.097736e-08,
  -1.894484e-08, -1.935621e-08, -1.976649e-08, -2.006022e-08, -2.026025e-08, 
    -2.047689e-08, -2.065647e-08, -2.084671e-08, -2.09104e-08, -2.093112e-08, 
    -2.080538e-08, -2.062636e-08, -2.034746e-08, -2.022512e-08, -2.011413e-08,
  -1.77989e-08, -1.81902e-08, -1.866161e-08, -1.897681e-08, -1.927436e-08, 
    -1.951669e-08, -1.976477e-08, -1.999225e-08, -2.008836e-08, 
    -2.014192e-08, -2.006826e-08, -1.990734e-08, -1.971187e-08, 
    -1.956988e-08, -1.944046e-08,
  -1.635784e-08, -1.688367e-08, -1.735959e-08, -1.776181e-08, -1.804788e-08, 
    -1.827539e-08, -1.848056e-08, -1.865452e-08, -1.877079e-08, 
    -1.887037e-08, -1.884589e-08, -1.876162e-08, -1.859637e-08, 
    -1.847149e-08, -1.835273e-08,
  -1.477164e-08, -1.531772e-08, -1.585309e-08, -1.628069e-08, -1.662982e-08, 
    -1.693246e-08, -1.713809e-08, -1.733937e-08, -1.746425e-08, 
    -1.756941e-08, -1.756862e-08, -1.753378e-08, -1.742347e-08, 
    -1.728444e-08, -1.720361e-08,
  -1.323171e-08, -1.373745e-08, -1.426632e-08, -1.471569e-08, -1.507837e-08, 
    -1.541872e-08, -1.566012e-08, -1.585647e-08, -1.595373e-08, 
    -1.603187e-08, -1.604063e-08, -1.604061e-08, -1.595921e-08, 
    -1.585976e-08, -1.577878e-08,
  -1.171959e-08, -1.22785e-08, -1.267339e-08, -1.314288e-08, -1.347266e-08, 
    -1.379727e-08, -1.406973e-08, -1.425441e-08, -1.437528e-08, 
    -1.444982e-08, -1.450778e-08, -1.451905e-08, -1.44743e-08, -1.443096e-08, 
    -1.437781e-08,
  -1.023243e-08, -1.066438e-08, -1.106435e-08, -1.14343e-08, -1.178657e-08, 
    -1.210558e-08, -1.237682e-08, -1.257758e-08, -1.272735e-08, 
    -1.285261e-08, -1.294928e-08, -1.299115e-08, -1.299342e-08, 
    -1.297942e-08, -1.295636e-08,
  -8.908398e-09, -9.107032e-09, -9.487057e-09, -9.866886e-09, -1.015363e-08, 
    -1.044918e-08, -1.069098e-08, -1.090025e-08, -1.107009e-08, -1.12124e-08, 
    -1.135007e-08, -1.144271e-08, -1.148208e-08, -1.153589e-08, -1.15706e-08,
  -7.700442e-09, -7.944756e-09, -8.135094e-09, -8.426428e-09, -8.707728e-09, 
    -9.001584e-09, -9.149465e-09, -9.333821e-09, -9.505322e-09, 
    -9.633801e-09, -9.749857e-09, -9.871963e-09, -9.963286e-09, 
    -1.004957e-08, -1.013835e-08 ;

 sftlf =
  0.1986115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9611561, 0.1583273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7949425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7552791, 0.2484612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.9872221, 0.4156101, 0.04560489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.8345782, 0.2958934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.7792858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9990003, 0.3505592, 0.06537855, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.8140894, 0.2409153, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.9453563, 0.02902743, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  1.522432, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  122.465, 2.830728, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  113.0215, 29.31339, 0.004701966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  140.0874, 33.71546, 1.141547, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  141.9684, 87.21121, 14.52402, 0.1304746, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  165.7051, 185.2302, 111.1391, 5.227489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  172.6293, 232.1111, 238.8028, 89.74486, 0.6524738, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  149.5705, 217.5222, 183.4477, 142.7244, 6.651272, 0.2006134, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  253.9191, 270.7406, 160.8987, 135.4378, 83.93595, 3.422685, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  248.2018, 381.5977, 396.3867, 296.0411, 147.8827, 85.51294, 0.2661929, 0, 
    0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
