netcdf ocean_static.hfgeou {
dimensions:
	time = UNLIMITED ; // (1 currently)
	yh = 10 ;
	xh = 15 ;
	xq = 15 ;
	yq = 10 ;
variables:
	float hfgeou(yh, xh) ;
		hfgeou:_FillValue = 1.e+20f ;
		hfgeou:missing_value = 1.e+20f ;
		hfgeou:units = "W m-2" ;
		hfgeou:long_name = "Upward geothermal heat flux at sea floor" ;
		hfgeou:cell_methods = "area:mean yh:mean xh:mean time: point" ;
		hfgeou:standard_name = "upward_geothermal_heat_flux_at_sea_floor" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
	double xh(xh) ;
		xh:units = "degrees_east" ;
		xh:long_name = "h point nominal longitude" ;
		xh:axis = "X" ;
	double xq(xq) ;
		xq:units = "degrees_east" ;
		xq:long_name = "q point nominal longitude" ;
		xq:axis = "X" ;
	double yh(yh) ;
		yh:units = "degrees_north" ;
		yh:long_name = "h point nominal latitude" ;
		yh:axis = "Y" ;
	double yq(yq) ;
		yq:units = "degrees_north" ;
		yq:long_name = "q point nominal latitude" ;
		yq:axis = "Y" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:43:25 2025: ncks -d xh,532,546 -d yh,526,535 -d xq,532,546 -d yq,526,535 /work/Carolyn.Whitlock/scratch//00010101.ocean_static.nc -O /work/Carolyn.Whitlock/scratch/ocean_subset/raw//00010101.ocean_static.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 hfgeou =
  0.07096534, 0.07089603, 0.07082672, 0.0707574, 0.07068809, 0.07061878, 
    0.07054947, 0.07048015, 0.07044549, 0.07044549, 0.07044549, 0.07044549, 
    0.07044549, 0.07044549, 0.07044549,
  0.07095248, 0.07085741, 0.07076235, 0.07066729, 0.07057223, 0.07047717, 
    0.0703821, 0.07028704, 0.07023951, 0.07023951, 0.07023951, 0.07023951, 
    0.07023951, 0.07023951, 0.07023951,
  0.07093959, 0.07081874, 0.07069791, 0.07057708, 0.07045624, 0.0703354, 
    0.07021457, 0.07009373, 0.07003331, 0.07003331, 0.07003331, 0.07003331, 
    0.07003331, 0.07003331, 0.07003331,
  0.07092668, 0.07078005, 0.0706334, 0.07048677, 0.07034013, 0.07019349, 
    0.07004685, 0.06990021, 0.06982689, 0.06982689, 0.06982689, 0.06982689, 
    0.06982689, 0.06982689, 0.06982689,
  0.07091377, 0.0707413, 0.07056884, 0.07039636, 0.0702239, 0.07005143, 
    0.06987897, 0.0697065, 0.06962027, 0.06962027, 0.06962027, 0.06962027, 
    0.06962027, 0.06962027, 0.06962027,
  0.07090084, 0.07070252, 0.0705042, 0.07030588, 0.07010756, 0.06990923, 
    0.06971091, 0.06951259, 0.06941342, 0.06941342, 0.06941342, 0.06941342, 
    0.06941342, 0.06941342, 0.06941342,
  0.07061216, 0.07041199, 0.07021181, 0.07001164, 0.06981146, 0.06961128, 
    0.06941111, 0.06921093, 0.06912883, 0.0691648, 0.06920077, 0.06923673, 
    0.0692727, 0.06930867, 0.06934464,
  0.07001173, 0.06983684, 0.06966195, 0.06948706, 0.06931216, 0.06913728, 
    0.06896238, 0.06878749, 0.06875634, 0.06886895, 0.06898155, 0.06909415, 
    0.06920676, 0.06931936, 0.06943196,
  0.06940359, 0.06925463, 0.06910566, 0.0689567, 0.06880774, 0.06865878, 
    0.06850982, 0.06836086, 0.0683815, 0.06857174, 0.06876198, 0.06895223, 
    0.06914247, 0.0693327, 0.06952295,
  0.06879488, 0.06867187, 0.06854886, 0.06842586, 0.06830285, 0.06817984, 
    0.06805684, 0.06793383, 0.0680063, 0.06827425, 0.0685422, 0.06881016, 
    0.06907811, 0.06934606, 0.06961402 ;

 time = 0 ;

 xh = -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375 ;

 xq = -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, -165, 
    -164.75, -164.5, -164.25, -164, -163.75, -163.5 ;

 yh = -14.3476556382336, -14.1053228834302, -13.862732304759, 
    -13.6198879813569, -13.3767940148509, -13.1334545290505, 
    -12.889873669635, -12.6460556038367, -12.4020045201193, -12.1577246278516 ;

 yq = -14.4687240631789, -14.2265217428746, -13.9840595676627, 
    -13.7413416053212, -13.4983719462701, -13.2551547032665, 
    -13.011694011094, -12.7679940262485, -12.5240589266184, -12.279892911161 ;
}
