netcdf \00010101.atmos_daily.tile1.ps {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float ps(time, grid_yt, grid_xt) ;
		ps:_FillValue = 1.e+20f ;
		ps:missing_value = 1.e+20f ;
		ps:units = "Pa" ;
		ps:long_name = "Surface Air Pressure" ;
		ps:cell_methods = "time: mean" ;
		ps:cell_measures = "area: area" ;
		ps:time_avg_info = "average_T1,average_T2,average_DT" ;
		ps:standard_name = "surface_air_pressure" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:53:52 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile1.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile1.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.1986115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9611561, 0.1583273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7949425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7552791, 0.2484612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.9872221, 0.4156101, 0.04560489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.8345782, 0.2958934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.7792858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9990003, 0.3505592, 0.06537855, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.8140894, 0.2409153, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.9453563, 0.02902743, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 ps =
  101882.4, 101966.1, 101989.7, 101996.6, 101986.1, 101968.2, 101943.2, 
    101913.1, 101864.9, 101812.7, 101752.6, 101683.9, 101601.9, 101517.6, 
    101425.3,
  100465.8, 101929.3, 101998, 102012.4, 102022.6, 102020.9, 102005.2, 
    101980.3, 101946, 101899.7, 101845.2, 101787.1, 101718.5, 101641, 101555.1,
  100568.7, 101604.9, 102001, 102024.1, 102037.4, 102046.7, 102045.4, 
    102034.9, 102004, 101964, 101915.8, 101863.5, 101803.8, 101735, 101661.2,
  100216.1, 101540.5, 101970, 102020.1, 102045, 102068.2, 102075.8, 102069.6, 
    102053.6, 102026.3, 101981.7, 101932.9, 101880.2, 101817.5, 101751.9,
  100139.1, 100848.8, 101784.1, 101999.9, 102037, 102068.1, 102086.2, 
    102088.4, 102080.1, 102063.1, 102034.1, 101989.5, 101941.4, 101889.2, 
    101829.8,
  99821.64, 99668.84, 100608.7, 101907.1, 102015.9, 102050.9, 102084.9, 
    102099.4, 102102.4, 102095.5, 102069, 102032.9, 101989.6, 101940, 101887.9,
  99676.62, 99087.6, 99089.15, 100891.8, 101983.6, 102037.5, 102069.2, 
    102098.3, 102104.6, 102100.8, 102084.5, 102057.3, 102022.4, 101981.1, 
    101934.2,
  99838.28, 99200.09, 99668.33, 100225.1, 101866.2, 102001, 102045.6, 
    102079.9, 102089.7, 102093.7, 102081.7, 102061.3, 102030.4, 101992.9, 
    101952.6,
  98560.73, 98498.51, 99841.91, 100263.3, 100924.7, 101927.3, 102006, 
    102037.9, 102056.9, 102067.2, 102059.2, 102047.4, 102025.9, 102001, 
    101973.1,
  98497.87, 97137.93, 97077.64, 98313.65, 100062.5, 100899.4, 101968.9, 
    102021.1, 102016.4, 102041, 102031.1, 102030.4, 102011.3, 101993.2, 
    101974.9,
  100935.8, 101054.8, 101124.5, 101162.2, 101195.8, 101218.9, 101237.8, 
    101247.6, 101247.6, 101236.2, 101208.9, 101172.3, 101124.9, 101070.4, 
    101011.8,
  99596.44, 101042, 101160.4, 101204.3, 101253.5, 101294, 101326, 101347.9, 
    101358.5, 101357.7, 101348.5, 101326.5, 101292.2, 101247.5, 101192.9,
  99749.81, 100776, 101201.4, 101251.4, 101304.1, 101351.7, 101392.4, 
    101424.9, 101448.9, 101464.1, 101464.1, 101454.3, 101430.5, 101399.2, 
    101358.8,
  99455.93, 100738.8, 101199.7, 101279.6, 101338.6, 101396.7, 101448.7, 
    101490.4, 101525.9, 101551.5, 101564.1, 101566.6, 101556.2, 101533.8, 
    101503.9,
  99422.81, 100108.2, 101045.8, 101296.2, 101366, 101423.3, 101484.3, 
    101536.4, 101581.1, 101617.9, 101642.5, 101654.3, 101654.7, 101644.4, 
    101625.9,
  99146.71, 98999.48, 99925.27, 101225.3, 101375.7, 101445.8, 101512, 
    101573.5, 101629.3, 101672.3, 101704.6, 101727.5, 101739.3, 101735.9, 
    101725.6,
  99040.81, 98467.48, 98493.64, 100251.9, 101361.6, 101452.4, 101524.4, 
    101597.2, 101659.3, 101710.4, 101752.9, 101779.7, 101797.7, 101806.7, 
    101808.9,
  99246.14, 98579.99, 99081.82, 99658.66, 101268.4, 101445, 101529.8, 
    101610.2, 101680.4, 101741.2, 101787, 101823.2, 101847, 101866.2, 101873.4,
  98086.02, 97933.85, 99223.7, 99701.17, 100383.2, 101385.9, 101531.6, 
    101607.8, 101684.9, 101761.2, 101809.2, 101850.6, 101873.4, 101900.1, 
    101914.8,
  98102.59, 96710.05, 96595.82, 97770.69, 99548.92, 100352, 101505.2, 
    101626.3, 101678.1, 101768.2, 101812.4, 101861.9, 101890.2, 101921.8, 
    101943.1,
  100310.9, 100283, 100292, 100305, 100307.9, 100311.1, 100297, 100262, 
    100237, 100233.1, 100252.8, 100275.9, 100304.3, 100333.9, 100361.2,
  98965.8, 100294.4, 100339.2, 100339.3, 100358.5, 100371.9, 100375.8, 
    100375.7, 100376, 100386.5, 100404.4, 100431.8, 100463.1, 100496.3, 
    100537.4,
  99105.68, 100070.9, 100407.9, 100401.4, 100415.8, 100430.4, 100461.9, 
    100486.9, 100502.9, 100523.3, 100549.2, 100580.8, 100620, 100664.5, 
    100711.8,
  98888.26, 100066, 100456.1, 100456.2, 100459.9, 100485.1, 100520, 100553.9, 
    100592.3, 100625.8, 100662.8, 100705.3, 100750.3, 100802.9, 100860.5,
  98889.95, 99523.93, 100361.7, 100520.4, 100518.3, 100542.7, 100589.9, 
    100653.6, 100710.9, 100752, 100789.7, 100836.7, 100888.6, 100945.9, 101005,
  98570.38, 98421.54, 99273.23, 100490.3, 100568.1, 100582.4, 100631, 
    100706.1, 100781.5, 100855.1, 100910.4, 100964.4, 101017.1, 101073.6, 
    101131.8,
  98505.52, 97902.43, 97867.3, 99550.12, 100589.8, 100638.7, 100688.5, 
    100755.9, 100835.6, 100915, 100987.2, 101051.4, 101112.7, 101177.3, 
    101239.6,
  98716.48, 97998.17, 98456.09, 98957.97, 100524.3, 100660.8, 100730.3, 
    100799.2, 100881, 100958.6, 101041.8, 101112.5, 101185.6, 101256.4, 
    101322.4,
  97630.82, 97410.23, 98638.87, 99015.49, 99659.86, 100620.6, 100749.7, 
    100831.4, 100920.6, 101003.6, 101090, 101166.3, 101243, 101313.8, 101384.6,
  97702.09, 96265.67, 96113.66, 97201.76, 98872.55, 99670.64, 100736.7, 
    100861.1, 100946.5, 101040.1, 101126.7, 101206.1, 101285.1, 101357.7, 
    101430.1,
  101211.2, 101278.8, 101287.8, 101286.2, 101273.3, 101252.2, 101223.8, 
    101194, 101156.4, 101113.1, 101066.1, 101015.6, 100957.7, 100898.2, 100841,
  99796.11, 101219.9, 101284.9, 101284.3, 101279.6, 101260.2, 101241, 
    101213.2, 101180.5, 101144.8, 101105.9, 101062.9, 101018, 100974.4, 
    100918.4,
  99881.77, 100897.4, 101265.3, 101269.7, 101270.4, 101259.2, 101242.4, 
    101218.5, 101191.9, 101158.4, 101126.6, 101091.2, 101054.3, 101014.1, 
    100973.6,
  99528.44, 100809.4, 101216.6, 101246.2, 101239, 101231.9, 101219.8, 
    101205.3, 101183, 101157, 101128.3, 101102.5, 101073, 101039.9, 101005.3,
  99424.82, 100133.7, 101015.1, 101197.5, 101204.3, 101196.6, 101187.1, 
    101173.1, 101156.4, 101140.1, 101118.2, 101087.8, 101058.1, 101031.8, 
    101010.6,
  99073, 98928.88, 99828.12, 101085.5, 101154.6, 101150.9, 101144.8, 
    101135.9, 101123.7, 101110.4, 101090.7, 101071.7, 101050.2, 101030.4, 
    101019,
  98937.3, 98338.16, 98307.78, 100067.9, 101096.8, 101097.1, 101092.4, 
    101090.5, 101080.3, 101073, 101062.2, 101051.4, 101037.3, 101031.5, 
    101038.3,
  99153.7, 98453.15, 98877.36, 99384.76, 100975.1, 101064.4, 101045.8, 
    101038.5, 101032.4, 101034.7, 101030, 101040.1, 101047.3, 101057.5, 
    101067.8,
  97884.74, 97781.73, 99082.42, 99424.7, 100026.4, 100980.3, 101010.2, 
    100991.2, 100990.6, 100998.7, 101015.3, 101030.3, 101050.1, 101071.3, 
    101093.4,
  97904.62, 96493.01, 96376.22, 97543.76, 99211.4, 99984.95, 100967.4, 
    100963.5, 100931.6, 100951, 100968.6, 101007.4, 101055.5, 101102.2, 101138,
  100181.9, 100266.8, 100337.7, 100417.2, 100520.1, 100627.2, 100744.4, 
    100862.6, 100983.1, 101096.6, 101203.8, 101302.3, 101392.4, 101472.2, 
    101546.9,
  98865.98, 100268.6, 100384.8, 100443.2, 100531.8, 100627.4, 100733.4, 
    100844.9, 100961.4, 101077.7, 101189.5, 101291.9, 101386, 101471.7, 
    101551.9,
  99025.93, 100016.6, 100407, 100463.9, 100547.6, 100630.5, 100725.3, 100830, 
    100941.1, 101058.2, 101173, 101277.1, 101373, 101460.6, 101545.4,
  98748.55, 99990.51, 100417.3, 100489, 100560.7, 100638, 100724.7, 100822.6, 
    100927.5, 101039.5, 101152.1, 101255.6, 101355.8, 101443.1, 101525,
  98766.08, 99410.33, 100293, 100515.1, 100578.2, 100650.4, 100725.3, 
    100812.5, 100911.7, 101018.2, 101131, 101233.1, 101334.1, 101424, 101508.2,
  98513.76, 98334.88, 99200.98, 100466.9, 100598.7, 100656.2, 100726.2, 
    100803.8, 100895.8, 100999.4, 101109.2, 101208.6, 101309.7, 101398.8, 
    101479.8,
  98465.81, 97858.16, 97835.98, 99531.05, 100603.1, 100663.3, 100720.7, 
    100789.4, 100873.9, 100970.6, 101081.4, 101182.2, 101284.6, 101374.4, 
    101456.8,
  98718.73, 98033.41, 98464.03, 98966.79, 100533.1, 100666.5, 100718.2, 
    100777.2, 100852.4, 100949.1, 101055.6, 101156.5, 101261.8, 101353.1, 
    101438.8,
  97590.43, 97443.36, 98702.65, 99074.04, 99696.5, 100644.1, 100721.7, 
    100759.1, 100832.6, 100923, 101033.6, 101136.6, 101245.4, 101338.9, 
    101428.8,
  97650.98, 96250.57, 96112.52, 97250.56, 98934.46, 99697.33, 100735.6, 
    100763.7, 100810.5, 100914.1, 101019.8, 101120.5, 101232.3, 101337, 101436,
  100789.5, 100759.2, 100720.2, 100648.3, 100580.4, 100500.3, 100425.6, 
    100345, 100276.8, 100229.5, 100209.8, 100201.3, 100211.1, 100232.6, 
    100270.9,
  99424.1, 100727.5, 100750.3, 100693.6, 100652.4, 100579.3, 100487.9, 
    100402.4, 100347.7, 100321.8, 100306.8, 100297.7, 100307, 100332.4, 
    100379.4,
  99538.45, 100461.8, 100786.4, 100729.3, 100677.5, 100612, 100550.2, 
    100502.7, 100469.6, 100440.8, 100420.4, 100415, 100431.9, 100457.3, 
    100505.3,
  99270.72, 100440.7, 100787.8, 100754.5, 100712.2, 100655.6, 100608.9, 
    100570.7, 100537.2, 100513.1, 100509.4, 100518.5, 100545, 100570.2, 
    100615.2,
  99254.88, 99841.81, 100641.3, 100780.4, 100744.5, 100706.1, 100670.3, 
    100634.2, 100611.6, 100615.5, 100626.9, 100629.6, 100655.3, 100686.9, 
    100735.7,
  98956.76, 98718.43, 99529.77, 100724.9, 100757.8, 100716, 100696.8, 100700, 
    100709.9, 100699.5, 100697, 100713, 100744.3, 100787.3, 100846.5,
  98858.95, 98202.2, 98113.76, 99786.04, 100784.2, 100771.3, 100761, 
    100761.8, 100752.5, 100751.6, 100765.1, 100786.9, 100825.4, 100879.4, 
    100939.2,
  99086.14, 98354.51, 98724.63, 99197.71, 100718, 100791.9, 100766.3, 
    100766.5, 100781.1, 100793.6, 100813.5, 100845.5, 100895.4, 100957.6, 
    101022,
  97915.05, 97732.18, 98954.39, 99284.12, 99868.78, 100771.3, 100776.5, 
    100782.9, 100809.3, 100830.5, 100863.9, 100916.2, 100969.9, 101030.1, 
    101098.7,
  97896.9, 96476.48, 96312.8, 97425.59, 99082.88, 99839.77, 100828.4, 
    100835.6, 100851.9, 100894.6, 100933.3, 100987.1, 101034, 101097.9, 
    101177.4,
  101785.2, 101819.5, 101813.6, 101802.3, 101800.3, 101786.6, 101766.8, 
    101741.3, 101713.1, 101676.3, 101634.9, 101594.9, 101555.7, 101517, 
    101474.6,
  100393.3, 101786, 101828, 101811.5, 101807.7, 101803.9, 101785.8, 101762.8, 
    101738.2, 101711.7, 101682.1, 101647, 101607.2, 101567.3, 101526,
  100496.6, 101480.6, 101829.2, 101822.4, 101825.4, 101828.5, 101829.9, 
    101817.5, 101798.5, 101772.5, 101745.3, 101711.1, 101675.9, 101636.8, 
    101596.6,
  100178.8, 101411.8, 101786.7, 101802.8, 101800.2, 101808.1, 101811.4, 
    101810.5, 101803.2, 101786.6, 101768.7, 101745, 101712.6, 101675.9, 
    101638.9,
  100109.7, 100763.3, 101614.5, 101777.7, 101774.9, 101786.8, 101815.1, 
    101821.4, 101822.3, 101812.7, 101795.9, 101771.4, 101749.9, 101725.9, 
    101698.8,
  99798.7, 99592.72, 100457, 101673.2, 101751.2, 101759.9, 101785.9, 
    101792.9, 101797, 101791.6, 101790.5, 101786.7, 101778.7, 101759.2, 
    101730.2,
  99638.5, 98980.45, 98931.09, 100668.3, 101722.1, 101746.6, 101772.7, 
    101786.5, 101797.1, 101802, 101800.6, 101793.4, 101778.3, 101763.8, 
    101752.3,
  99876.38, 99150.66, 99568.69, 100072.1, 101665.4, 101751.6, 101760.7, 
    101771.5, 101776.9, 101788.7, 101792.3, 101790.3, 101786.4, 101791.2, 
    101802,
  98637.04, 98472.87, 99755.23, 100093.6, 100732.2, 101690.6, 101757.9, 
    101778.6, 101795.6, 101801.9, 101799.9, 101804.1, 101810.5, 101825.4, 
    101821.8,
  98565.93, 97141.2, 97046.69, 98225.32, 99968.08, 100739.5, 101764.5, 
    101768.4, 101753, 101752.4, 101764.1, 101792.4, 101804.6, 101793.8, 
    101779.2,
  101690.9, 101780.5, 101826.1, 101851.5, 101879.8, 101903.1, 101923.6, 
    101938.6, 101950.6, 101959.2, 101962.8, 101963.8, 101962.1, 101957.5, 
    101950.4,
  100326.6, 101757.7, 101842.3, 101880.8, 101919.4, 101955.8, 101986.2, 
    102008.4, 102027, 102039.9, 102051.6, 102059.9, 102064.6, 102065.6, 
    102063.1,
  100441.8, 101459.8, 101851.1, 101897.8, 101936.9, 101981.4, 102017.9, 
    102047.7, 102077, 102098.6, 102119, 102131.2, 102142.5, 102149, 102152.4,
  100116.6, 101398.7, 101824.9, 101894.5, 101936.6, 101989.5, 102038, 
    102076.2, 102113.5, 102140.4, 102164.5, 102184.8, 102200.9, 102209.3, 
    102216,
  100053.6, 100749.1, 101653.5, 101878.1, 101928.4, 101979.9, 102031.3, 
    102072.8, 102115.5, 102153.9, 102187, 102213.6, 102234.9, 102250.9, 
    102261.8,
  99720.36, 99568.2, 100486.7, 101788.6, 101904.2, 101959.9, 102017, 
    102066.6, 102114.2, 102155.7, 102193, 102226.6, 102253.9, 102276.6, 
    102293.6,
  99594.22, 98984.47, 98979.16, 100768.9, 101860.2, 101922.5, 101978.4, 
    102028.9, 102074.6, 102124, 102168.8, 102210.1, 102245.8, 102278.6, 
    102306.6,
  99794.8, 99115.96, 99583.86, 100120.7, 101746.3, 101878.3, 101932.3, 
    101995.3, 102042.3, 102087.2, 102129.1, 102169, 102209, 102240.7, 102270.5,
  98539.2, 98421.62, 99763.16, 100156.5, 100820.7, 101801.5, 101874.9, 
    101910.5, 101959.8, 101996.4, 102040.8, 102078.5, 102119.2, 102158.4, 
    102198.3,
  98501.47, 97072.26, 96978.02, 98218.07, 99987.36, 100755.6, 101844.7, 
    101862.5, 101897.7, 101929.9, 101961.9, 102007.9, 102053.1, 102099, 
    102140.9,
  101036.9, 101146.7, 101209.5, 101258.4, 101315.2, 101369.5, 101414.8, 
    101459.3, 101502.1, 101541.9, 101575.5, 101607.4, 101633.8, 101659.3, 
    101681.7,
  99696.16, 101115.9, 101220.9, 101275.8, 101333.2, 101395, 101451.6, 
    101506.5, 101556.7, 101602.3, 101644.5, 101686.8, 101724.3, 101761, 
    101792.2,
  99800.02, 100805, 101209.1, 101282.9, 101340.4, 101411.2, 101473.5, 
    101535.3, 101590.7, 101643.8, 101693.6, 101741.8, 101787.6, 101831.2, 
    101871.7,
  99495.55, 100773.7, 101173.3, 101254, 101311.8, 101397.1, 101468.3, 
    101539.2, 101598.7, 101658.7, 101717.3, 101776.9, 101832.1, 101883.8, 
    101931.9,
  99431.09, 100121.3, 101016, 101250.9, 101297.4, 101376.9, 101457.8, 101530, 
    101589.6, 101652.1, 101717.2, 101784.2, 101847.7, 101906.6, 101962.2,
  99136.84, 98968.46, 99854.28, 101137.9, 101269.9, 101345.8, 101432.8, 
    101524.4, 101588.8, 101642.3, 101707.2, 101784.5, 101850.2, 101913.5, 
    101976.6,
  99037.59, 98410.8, 98404.25, 100144.4, 101262.1, 101330.7, 101415.1, 
    101500.5, 101575.5, 101638.3, 101699.4, 101767.8, 101834.8, 101903, 
    101968.7,
  99247.12, 98534.61, 99002.16, 99520.79, 101137.6, 101304.5, 101389.8, 
    101476, 101558.9, 101626.9, 101689.4, 101750.8, 101821.2, 101890, 101955.5,
  98059.49, 97895.41, 99181.83, 99579.02, 100246.3, 101244.8, 101357.9, 
    101425.4, 101513.9, 101591.1, 101668, 101736.3, 101803.2, 101866.8, 
    101933.5,
  98106.77, 96666.9, 96549.33, 97708.91, 99442.6, 100211.4, 101315.7, 101397, 
    101473.5, 101573.4, 101643.2, 101718.1, 101791.7, 101853.5, 101916.2,
  100293.8, 100349.3, 100381.5, 100392.8, 100421.5, 100448.7, 100476.7, 
    100513.9, 100563.3, 100612.8, 100658.8, 100711.7, 100767.2, 100823.2, 
    100864.4,
  98974.43, 100334.6, 100420.8, 100445.6, 100465.4, 100489.5, 100510.8, 
    100531.9, 100569, 100618, 100673.5, 100738.5, 100800.4, 100872.7, 100935.5,
  99140.17, 100089.6, 100441.3, 100465.2, 100473.2, 100486.9, 100495, 
    100511.7, 100541.3, 100590.2, 100648.9, 100719.6, 100805.2, 100895.6, 
    100976.3,
  98904.23, 100089.5, 100457.4, 100491.9, 100487.8, 100489.4, 100482.9, 
    100473.9, 100496.6, 100540.7, 100604.3, 100675.5, 100770.1, 100882.8, 
    100996.6,
  98901.19, 99515.52, 100326.8, 100513.5, 100512.7, 100501.7, 100482.3, 
    100461.4, 100455.2, 100468.8, 100530.7, 100629.1, 100734.7, 100850, 
    100979.4,
  98688.46, 98453.62, 99242.84, 100454.6, 100535.2, 100524.4, 100515.5, 
    100496.6, 100485.9, 100490.5, 100530, 100606.6, 100708.6, 100843.2, 
    100990.1,
  98658.94, 97983.16, 97888.27, 99506.09, 100533.1, 100549.4, 100541.1, 
    100539.9, 100537.6, 100554.4, 100604.5, 100672, 100762, 100873.3, 101019.5,
  98942.45, 98183.9, 98537.97, 98969.8, 100479.6, 100568.8, 100572.5, 
    100581.1, 100594.2, 100615.8, 100653.8, 100718.1, 100816.4, 100931, 
    101055.8,
  97838.04, 97604.81, 98809.97, 99113.16, 99668.48, 100559.9, 100612.8, 
    100627.8, 100647.7, 100672.5, 100710.5, 100779, 100862.4, 100961.4, 101084,
  97925.06, 96446.71, 96270.01, 97348.2, 98976.48, 99691.33, 100665.6, 
    100704.9, 100727.6, 100762.9, 100793.8, 100842, 100922.4, 101018.9, 
    101117.8,
  100251, 100299.1, 100324.8, 100354.1, 100384.5, 100403.6, 100403.1, 
    100392.7, 100376.9, 100362.1, 100341.9, 100323.3, 100300.8, 100280.3, 
    100261.3,
  98907.34, 100231.5, 100336.6, 100362.8, 100399.9, 100423.1, 100445.5, 
    100445.1, 100438.6, 100424.3, 100408.4, 100387, 100363.3, 100339.6, 
    100320.2,
  99109.13, 100020.7, 100381.5, 100401.7, 100420.6, 100444.8, 100462.1, 
    100482.8, 100484.3, 100484.6, 100468.2, 100448.4, 100420.1, 100388.9, 
    100359.9,
  98879.3, 100055.7, 100418.8, 100457.1, 100473.9, 100490.9, 100516.5, 
    100533.9, 100544.6, 100546, 100532.5, 100507, 100471.4, 100426.1, 100389.6,
  98895.63, 99512.16, 100329.8, 100520.4, 100537.9, 100550, 100564.4, 100588, 
    100598.9, 100611.5, 100600.4, 100571, 100531.4, 100480.1, 100433.8,
  98652.02, 98453.64, 99271.28, 100478.5, 100573.4, 100594.8, 100613.6, 
    100640.3, 100657.4, 100670.4, 100663.7, 100642.5, 100603.2, 100548.8, 
    100499.1,
  98600.28, 97955.77, 97894.66, 99554.01, 100586.6, 100624.9, 100644.7, 
    100672.7, 100699.3, 100717.7, 100720.6, 100710.9, 100684, 100643.5, 
    100603.5,
  98860.6, 98125.68, 98519.48, 98977.43, 100516.6, 100631.2, 100665.8, 
    100700.7, 100726.8, 100755.1, 100768.5, 100765.8, 100756, 100728.4, 
    100705.3,
  97748.83, 97559.7, 98773.42, 99075.35, 99664.49, 100598.4, 100672.3, 
    100700.9, 100739.4, 100771.8, 100794.4, 100805.3, 100811.2, 100805.5, 
    100801.5,
  97818.34, 96362.56, 96198.84, 97297.84, 98942.75, 99664.78, 100675.8, 
    100709.5, 100737.6, 100778.4, 100810.5, 100837.8, 100852, 100868.1, 
    100878.3,
  100225.7, 100318.1, 100396.3, 100447, 100499, 100550.4, 100604.1, 100668.5, 
    100741.9, 100816.5, 100899.8, 100975, 101040.2, 101094.8, 101140,
  98949.41, 100332.1, 100463.2, 100526.4, 100582, 100633.9, 100690.9, 
    100753.7, 100822.1, 100892.6, 100971.5, 101044.7, 101113.5, 101179.2, 
    101233.5,
  99157.72, 100116.9, 100515.7, 100582.4, 100641.2, 100698.6, 100760.7, 
    100824.3, 100891.9, 100962.4, 101044.1, 101117.7, 101187.3, 101252.1, 
    101312.9,
  98916.23, 100118.5, 100544.9, 100627.7, 100692.7, 100751.7, 100820.1, 
    100889.6, 100961.1, 101033.1, 101112.2, 101181.5, 101247.9, 101318.4, 
    101379.1,
  98926.95, 99554.81, 100425.3, 100647, 100723.4, 100786.9, 100864, 100938.8, 
    101016.2, 101090.9, 101170.7, 101239, 101307.9, 101375.1, 101436.5,
  98676.92, 98487.05, 99348.5, 100584.3, 100733.6, 100803.4, 100890.5, 
    100974.1, 101062.5, 101140.2, 101220, 101291.8, 101359.3, 101424.8, 
    101486.1,
  98625.39, 97982.98, 97963.9, 99633.72, 100715.2, 100809.4, 100906.9, 
    100996.1, 101091.1, 101174.5, 101259.2, 101330.2, 101400.2, 101465, 
    101528.3,
  98872.01, 98144.68, 98567.48, 99054.62, 100617.1, 100793.1, 100907.9, 
    101003.1, 101106.5, 101195.4, 101283.6, 101357.4, 101430.7, 101497.8, 
    101566.4,
  97744.06, 97563.3, 98789.82, 99112.95, 99754.38, 100740.1, 100913, 
    101005.8, 101111.7, 101204.3, 101293.6, 101369.4, 101446, 101517.5, 
    101591.3,
  97804.95, 96362.73, 96218.12, 97330.27, 99007.09, 99746.4, 100885.5, 
    101006.5, 101103.1, 101205.1, 101294.5, 101374.3, 101451.3, 101528.2, 
    101607.5,
  100539.8, 100614.4, 100715.4, 100819.4, 100911.9, 101002.6, 101086.1, 
    101162.3, 101235.3, 101300.7, 101361.4, 101418, 101466.9, 101509.2, 
    101546.4,
  99206.26, 100569.8, 100701.3, 100800, 100897.2, 100998.6, 101098.9, 
    101193.1, 101287.9, 101377.7, 101461.6, 101536.5, 101600.8, 101660.6, 
    101713.9,
  99357.24, 100310.9, 100704.7, 100802.1, 100904.8, 101009.8, 101120.5, 
    101223.9, 101322.6, 101412.9, 101502.4, 101582.6, 101655.1, 101721.6, 
    101780.5,
  99052.56, 100264.9, 100687.9, 100796.2, 100905.5, 101014, 101131.5, 
    101242.9, 101353.3, 101458.4, 101558.6, 101649.7, 101734.2, 101812.5, 
    101881.9,
  99050.88, 99684.34, 100546.5, 100791, 100905.4, 101016.9, 101138.5, 
    101255.4, 101375, 101483.1, 101587.9, 101685.1, 101775.7, 101860.4, 
    101936.4,
  98775.74, 98597.3, 99458.92, 100715.1, 100893.1, 101009.6, 101137.3, 
    101259.9, 101387.8, 101507.6, 101618.9, 101721.2, 101817.2, 101908.2, 
    101991.9,
  98725.3, 98090.45, 98079.2, 99762.21, 100866.9, 100997.2, 101135.6, 
    101264.5, 101398.5, 101520.3, 101628.4, 101731.5, 101829.8, 101923.9, 
    102011.4,
  98958.04, 98248.39, 98687.58, 99186.72, 100767, 100970.6, 101125, 101260.9, 
    101395.5, 101522.5, 101631.6, 101734.6, 101836, 101931.8, 102024,
  97827.54, 97674.33, 98918, 99259.7, 99906.57, 100908.7, 101115.6, 101251.6, 
    101382.4, 101509.4, 101619, 101724.5, 101827.1, 101924.3, 102017.8,
  97880.41, 96475.66, 96330.07, 97480.12, 99172.15, 99903.2, 101076.4, 
    101236.4, 101351.5, 101486.9, 101600.7, 101710.1, 101815.9, 101914.1, 
    102010.8,
  100733.9, 100796, 100870.2, 100943.1, 101013.5, 101085.9, 101162.1, 
    101229.5, 101294.4, 101354.7, 101407.9, 101455.5, 101498.9, 101540.1, 
    101574.4,
  99402.88, 100772.7, 100869.2, 100939.9, 101025.8, 101111.9, 101198.3, 
    101277.6, 101356.8, 101425.3, 101492.3, 101552.3, 101604.1, 101653.9, 
    101695,
  99525.73, 100490.7, 100877.2, 100951.3, 101034.9, 101129.4, 101225.6, 
    101318, 101403.2, 101483.3, 101560.7, 101625.7, 101686.5, 101743.9, 
    101793.9,
  99222.71, 100447.3, 100863.5, 100942.1, 101040, 101139.6, 101240.8, 
    101343.7, 101438.2, 101528.4, 101611.1, 101688.2, 101761.1, 101827.2, 
    101891.4,
  99214.92, 99860.23, 100726.7, 100937.5, 101034.4, 101141.2, 101247.3, 
    101358.1, 101461.1, 101561.6, 101651.1, 101736.9, 101817.2, 101890, 
    101962.8,
  98950.94, 98778.73, 99632.32, 100881.3, 101024.9, 101133.6, 101246.4, 
    101364.3, 101474.5, 101583.4, 101681, 101774.3, 101862.1, 101940.8, 
    102019.4,
  98888.45, 98282.43, 98261.52, 99930.28, 101014.9, 101123.1, 101245.4, 
    101368.9, 101481.4, 101599.6, 101701.5, 101799.8, 101892.3, 101976.3, 
    102055,
  99144.48, 98440.98, 98877.5, 99366.59, 100929.1, 101110.8, 101241.7, 
    101371.6, 101486, 101609.1, 101715.7, 101816.4, 101911.7, 101996, 102078.2,
  98005.38, 97858.65, 99112.08, 99460.69, 100072.6, 101075, 101250.2, 
    101381.4, 101490.3, 101614.9, 101723.6, 101823.7, 101918.8, 102006.3, 
    102088.9,
  98068.23, 96654.88, 96515.1, 97651.12, 99354.06, 100097.3, 101220.4, 
    101388.1, 101487.7, 101613.8, 101723, 101821.8, 101916.8, 102004.7, 
    102088.8,
  100395.6, 100497.3, 100559.3, 100629.8, 100698.3, 100774.1, 100842.9, 
    100909.1, 100971.3, 101031.2, 101090.6, 101151.6, 101212.3, 101267.9, 
    101312,
  99095.07, 100480.4, 100576.3, 100653.8, 100738.1, 100823.3, 100902.6, 
    100978.6, 101049.8, 101123.3, 101193.7, 101260.1, 101319.3, 101368.3, 
    101412.8,
  99256.92, 100230.1, 100611, 100681.9, 100769.8, 100859.9, 100951, 101039.3, 
    101119.1, 101198.6, 101275.3, 101347.4, 101416.6, 101478.8, 101533.4,
  98997.23, 100208.9, 100623, 100698, 100798.7, 100894.2, 100991.3, 101092, 
    101182.3, 101274.9, 101358.3, 101434.7, 101506.5, 101571.1, 101627.5,
  99013.84, 99642.27, 100507, 100719.3, 100819.1, 100922.1, 101023.8, 
    101133.9, 101232.8, 101333.9, 101424.3, 101506.2, 101585, 101654.1, 
    101717.4,
  98772.27, 98587.61, 99439.12, 100682.9, 100834.3, 100936.4, 101047.7, 
    101163.6, 101271.1, 101380, 101475.4, 101561.1, 101641.5, 101712.2, 
    101776.4,
  98738.17, 98109.79, 98085.64, 99760.37, 100846.2, 100953.3, 101073, 
    101191.6, 101299.1, 101409.1, 101506.1, 101593.4, 101677.7, 101752.3, 
    101821.6,
  99002.67, 98285.96, 98725.33, 99215.84, 100788.1, 100958.8, 101090.2, 
    101213.9, 101320.2, 101430.3, 101526.4, 101613.6, 101698.8, 101775.8, 
    101847.9,
  97889.56, 97723.02, 98972.52, 99315.82, 99956.26, 100933.8, 101114.4, 
    101238.4, 101336.2, 101445.1, 101539.3, 101627.2, 101713, 101791.3, 
    101867.2,
  97959.65, 96537.91, 96396.23, 97529.3, 99224.9, 99966.47, 101093.1, 
    101255.9, 101342.5, 101455.1, 101550, 101636.8, 101722.1, 101802.2, 
    101877.6,
  100375.9, 100381.3, 100376.1, 100385.3, 100398.5, 100403.6, 100405.6, 
    100403.6, 100402.4, 100395.2, 100381.8, 100364.2, 100352, 100350.5, 
    100368.9,
  99046.17, 100406.3, 100432.4, 100428.5, 100445.1, 100463.9, 100479.2, 
    100491.3, 100501, 100510.4, 100516.5, 100520.5, 100526.7, 100538.7, 100555,
  99138.77, 100101.3, 100450.2, 100459.1, 100479.1, 100502.1, 100532.9, 
    100565.9, 100600.9, 100630.6, 100650.9, 100668, 100685.4, 100708.9, 
    100739.9,
  98870.55, 100056.2, 100441.1, 100469.4, 100511.4, 100548.3, 100587.8, 
    100631.9, 100673.1, 100711.3, 100750.8, 100787.1, 100821.7, 100859.5, 
    100895.6,
  98885.55, 99494.87, 100339.8, 100520.9, 100554.3, 100595.8, 100640.6, 
    100696.1, 100750.9, 100805.2, 100856.8, 100902.5, 100947.5, 100994, 
    101043.2,
  98644.88, 98449.34, 99271.78, 100485.8, 100584.5, 100633.8, 100697.6, 
    100765.6, 100828.3, 100889.8, 100951.9, 101010.7, 101068.4, 101123.8, 
    101178.6,
  98616.48, 97979.16, 97935.97, 99586.59, 100623.3, 100692.8, 100762.7, 
    100840.5, 100909.9, 100982.2, 101050.6, 101113.7, 101173.7, 101232.1, 
    101289.4,
  98888.8, 98168.5, 98582.2, 99063.13, 100588.3, 100731.2, 100810, 100902, 
    100982, 101058.2, 101132, 101198.4, 101263, 101324.7, 101387.4,
  97775.49, 97618.98, 98835.22, 99168.74, 99772.3, 100729.8, 100859.5, 
    100959.9, 101042.1, 101118.6, 101195.8, 101264.4, 101332.9, 101398.3, 
    101462.9,
  97847.28, 96433.11, 96276.38, 97391.62, 99057.68, 99790.51, 100864.9, 
    101000.6, 101075, 101160.3, 101241.9, 101314.6, 101384.4, 101450.4, 
    101516.5,
  101247.8, 101256, 101268.5, 101282.1, 101301.1, 101314.6, 101341.2, 
    101366.5, 101387.6, 101408.5, 101428.1, 101439.9, 101449.5, 101448.7, 
    101447,
  99810.23, 101203.6, 101243.6, 101254.7, 101263, 101266.9, 101283.2, 
    101290.6, 101327.2, 101357.4, 101389.9, 101412.7, 101428.5, 101437.4, 
    101434.2,
  99907.43, 100898.1, 101182, 101164.4, 101172.8, 101194.8, 101222.2, 
    101253.2, 101270.4, 101298.2, 101325.1, 101355.9, 101386.5, 101413.6, 
    101429.5,
  99464.29, 100706.8, 101069.3, 101071, 101059.7, 101075.9, 101066.7, 
    101059.8, 101043.4, 101066.8, 101106.9, 101162.3, 101204.7, 101250.5, 
    101300.9,
  99340.58, 100006.6, 100801.9, 100918.2, 100877.4, 100906.3, 100923.7, 
    100940.6, 100936.2, 100960.6, 101008.6, 101081.3, 101147.1, 101206.2, 
    101259.3,
  98964.48, 98784, 99597.14, 100776.2, 100825.5, 100841, 100871.7, 100902.3, 
    100932.2, 100983, 101047.3, 101117.8, 101179.3, 101237.3, 101293.2,
  98787.09, 98165.78, 98123.28, 99776.52, 100775.5, 100801.9, 100849.1, 
    100915, 100975.3, 101037.2, 101107.5, 101182.5, 101252.1, 101318, 101378.9,
  98998.81, 98281.93, 98683.82, 99165.8, 100687.9, 100793.9, 100864.8, 
    100947.2, 101019.4, 101090, 101169.1, 101244.5, 101313.9, 101382.8, 
    101445.2,
  97855.27, 97685.8, 98910.45, 99238.84, 99830.59, 100760.9, 100881.8, 
    100974.1, 101061.9, 101138.6, 101220.8, 101296.8, 101368.2, 101436.4, 
    101498.3,
  97912.59, 96486.04, 96341.58, 97451.05, 99113.46, 99839.77, 100877.9, 
    101001, 101085.8, 101168.9, 101250.8, 101323.9, 101394.3, 101461, 101526.1,
  101383.5, 101460.7, 101506.8, 101547.5, 101578.4, 101602.6, 101621.6, 
    101637.2, 101655.7, 101667.9, 101677.1, 101683.8, 101688.2, 101691.4, 
    101701,
  99933.9, 101360.7, 101432, 101469.3, 101498.4, 101522.2, 101543.9, 
    101564.1, 101578.1, 101596, 101608.1, 101617, 101624.6, 101636.1, 101645.1,
  99960.62, 100957.8, 101336.7, 101387.7, 101422.8, 101441.3, 101446.5, 
    101453.7, 101454.7, 101467.2, 101482.8, 101501.5, 101517.9, 101535.4, 
    101553,
  99587.73, 100858.3, 101240.1, 101280.2, 101296.5, 101335.5, 101348.5, 
    101374.5, 101401.6, 101418, 101414.9, 101419.6, 101424.2, 101420, 101417.9,
  99430.59, 100159.7, 101036.4, 101248.3, 101244, 101272.8, 101282.2, 
    101298.2, 101281.8, 101268, 101255.6, 101267.8, 101281, 101303.3, 101319,
  99049.43, 98895.07, 99771.81, 101041.5, 101132.5, 101156, 101178.9, 
    101182.2, 101159.2, 101149.7, 101160.8, 101199, 101230, 101259.8, 101288.9,
  98916.85, 98299.8, 98284.13, 99994.47, 101017, 101030.9, 101048.6, 101065, 
    101083.8, 101106.3, 101143.4, 101191.5, 101245.1, 101297.7, 101346.5,
  99065.92, 98365.99, 98818.55, 99299.55, 100831.2, 100914, 100955.5, 
    101020.8, 101072.8, 101119.5, 101175.5, 101227.6, 101282.5, 101337, 
    101391.2,
  97879.77, 97728.44, 98971.42, 99319.73, 99893.94, 100837.1, 100906.8, 
    100990.9, 101059.8, 101114.8, 101176.5, 101234.3, 101299.6, 101364.2, 
    101429.2,
  97924.21, 96494.09, 96347.41, 97482.62, 99159.12, 99865.29, 100871.5, 
    100959.7, 101041.2, 101110.2, 101182.9, 101250.9, 101320.6, 101388.5, 
    101456.6,
  101045.8, 101079.4, 101086.9, 101111.3, 101148.7, 101183.7, 101209.2, 
    101228.9, 101233, 101250.9, 101273.6, 101309.9, 101355.8, 101453.4, 
    101547.4,
  99610.4, 101005.2, 101053.6, 101055.5, 101062, 101074.5, 101093, 101107.6, 
    101124.7, 101141.8, 101151.3, 101193.3, 101249.2, 101349.7, 101457.6,
  99626.84, 100609.6, 100946.7, 100977.3, 101021.1, 101048.4, 101054.7, 
    101069.2, 101062, 101061.7, 101065.8, 101116.4, 101167.7, 101255.4, 
    101342.7,
  99236.55, 100444.3, 100824.2, 100862, 100900.7, 100954.1, 100979, 100984.1, 
    100986.3, 100979.2, 101008.8, 101070.5, 101130, 101203.7, 101286,
  99165.58, 99780.59, 100596.4, 100765.2, 100801.6, 100854.5, 100916.7, 
    100928.6, 100941.5, 100968.4, 101005, 101054, 101108.3, 101163.5, 101230.4,
  98885.66, 98667.55, 99479.93, 100663.9, 100753.8, 100768, 100818.3, 
    100864.9, 100913.5, 100971.7, 101027.1, 101082, 101137.5, 101196.9, 
    101251.8,
  98798.84, 98138.9, 98073.69, 99710.55, 100727.5, 100767.2, 100810.7, 
    100875.4, 100932, 100981.7, 101041.6, 101101.4, 101161.8, 101223.1, 
    101282.2,
  99033.75, 98308.46, 98694.85, 99149.89, 100665.8, 100754.7, 100805.3, 
    100855.9, 100919.6, 100986.1, 101061.2, 101129.2, 101197.6, 101261, 
    101322.7,
  97870.11, 97712.05, 98936.57, 99256.62, 99821.14, 100733, 100812.8, 
    100873.7, 100937.6, 101000.8, 101071.9, 101138.6, 101208, 101277.9, 
    101342.3,
  97925.01, 96480.61, 96325.88, 97441.57, 99086.58, 99805.13, 100814.8, 
    100876.3, 100931, 101000.7, 101071.6, 101141.7, 101215.4, 101281, 101350.7,
  101073, 101116.4, 101118.5, 101106.8, 101094.4, 101071.4, 101039.3, 
    101008.5, 100969, 100936.1, 100900.6, 100848.3, 100771.8, 100690, 100612.1,
  99734.25, 101110.4, 101145.9, 101129.4, 101113.4, 101091.1, 101061.4, 
    101030.7, 100992.4, 100955.8, 100913, 100867.6, 100802.1, 100722.9, 
    100635.3,
  99850.96, 100821.2, 101159.1, 101142.1, 101128.6, 101108.1, 101072.5, 
    101034.3, 100993.1, 100957.1, 100919.6, 100882.3, 100831, 100770.6, 
    100716.1,
  99556.12, 100774.5, 101142.7, 101153.6, 101127.6, 101100.6, 101067.2, 
    101031.5, 100991.7, 100953.7, 100905.9, 100860.1, 100818.6, 100779, 
    100743.2,
  99501.08, 100147.6, 100977.7, 101143.9, 101119.2, 101089.4, 101055.5, 
    101015.6, 100968.6, 100918.8, 100876.3, 100840, 100807.4, 100782.5, 
    100751.3,
  99193.95, 99006.03, 99858.81, 101063.3, 101103.4, 101065.4, 101033.4, 
    100997.9, 100945.7, 100901.9, 100860.5, 100818.6, 100780.5, 100757.1, 
    100736.6,
  99056.94, 98425.04, 98370.4, 100080.4, 101069.9, 101044.2, 101009.1, 
    100980.9, 100942.5, 100903.8, 100861.5, 100822.5, 100792.1, 100765.8, 
    100749.4,
  99251.8, 98550.63, 98944.96, 99437.21, 100974.9, 101025, 101000.2, 
    100976.3, 100949.1, 100919.2, 100893.2, 100869.7, 100848.1, 100829.2, 
    100817.4,
  98026.01, 97892.91, 99146.26, 99466.78, 100067.4, 100965.8, 100983, 
    100958.7, 100939.8, 100923.3, 100904.2, 100891.1, 100884.1, 100883.3, 
    100884.9,
  98021.89, 96596.91, 96486.34, 97628.06, 99280.23, 100014.3, 100971.1, 
    100957, 100927.5, 100925.5, 100922.6, 100927.9, 100926.1, 100939.5, 
    100950.4,
  100898.8, 100957.1, 100968.4, 100953.2, 100937.8, 100915.9, 100887.6, 
    100858, 100822.3, 100782.3, 100744.7, 100708.8, 100670.5, 100633.9, 
    100596.6,
  99593.05, 100954.3, 101017.6, 101022.9, 101018.9, 101006.7, 100986.5, 
    100961.3, 100932.4, 100905.2, 100873.1, 100841.8, 100809.3, 100775.1, 
    100739.9,
  99736.16, 100698.5, 101060.5, 101075.1, 101076.9, 101074.2, 101064.1, 
    101048.3, 101026.3, 101000.5, 100972.6, 100945.6, 100917.8, 100886, 
    100856.5,
  99444.88, 100668.3, 101066.4, 101111.7, 101118.6, 101124.9, 101125.3, 
    101120, 101106.6, 101089.4, 101068.8, 101043.2, 101021.8, 100995.8, 
    100965.9,
  99407.97, 100057, 100925.8, 101124.1, 101145.6, 101156.5, 101168.4, 
    101170.8, 101166, 101156.5, 101140.2, 101127.9, 101105.1, 101078.4, 
    101045.7,
  99095.3, 98921.44, 99800.76, 101051.7, 101148.8, 101169.7, 101186.4, 
    101200.4, 101203.4, 101201.3, 101194.6, 101181.8, 101165.1, 101143.3, 
    101115.7,
  98978.15, 98362.9, 98343.2, 100067.5, 101125.2, 101167.3, 101188.3, 
    101207.2, 101217, 101223.3, 101221.4, 101215.2, 101204.1, 101185.9, 101160,
  99157.18, 98478.03, 98922.52, 99438.59, 101019.8, 101141.9, 101173.6, 
    101193.6, 101208.7, 101218.1, 101223.7, 101224.9, 101220.2, 101211.6, 
    101194.9,
  97939.84, 97817.04, 99104.66, 99463.51, 100112.7, 101080.9, 101147.5, 
    101168.3, 101184.6, 101199, 101204.7, 101214.1, 101214.8, 101215.6, 
    101207.4,
  97912.76, 96516.4, 96403.83, 97602.59, 99301.8, 100081.2, 101112.8, 
    101139.4, 101142.1, 101168.7, 101175.4, 101189.5, 101194.3, 101204.7, 
    101209.4,
  100880.4, 101003.5, 101085.8, 101159.6, 101238.4, 101301.1, 101363.4, 
    101398.4, 101426.1, 101437.2, 101439.8, 101423.5, 101399, 101367.2, 
    101322.4,
  99482.95, 100904.8, 101017.5, 101086.4, 101162.8, 101230.2, 101291.1, 
    101344.1, 101387.2, 101417.6, 101432.6, 101438.7, 101431.1, 101409.8, 
    101380.3,
  99539.08, 100561.7, 100976.1, 101045.4, 101113, 101174.4, 101227, 101276.7, 
    101327.4, 101366.6, 101397.8, 101416.3, 101426.4, 101426.4, 101413.6,
  99191.74, 100456.1, 100903.2, 100994.6, 101065.6, 101137, 101199.7, 
    101249.4, 101292.2, 101327.9, 101362.7, 101392.9, 101419.1, 101426.2, 
    101427.8,
  99115.5, 99793.56, 100707.1, 100944.6, 101020.8, 101090.8, 101167.4, 
    101225.9, 101275, 101314.8, 101347.9, 101372.8, 101395.5, 101415.1, 
    101424.7,
  98787.51, 98632.99, 99524.5, 100819.5, 100966, 101041.9, 101120.8, 
    101192.5, 101251.4, 101304.7, 101347.5, 101383.5, 101409.6, 101429.1, 
    101442,
  98669.98, 98069.37, 98075.2, 99798.17, 100903.8, 100992.4, 101073.8, 
    101151.9, 101216.9, 101275.6, 101326.3, 101373, 101412.3, 101445.4, 
    101468.1,
  98849.42, 98174, 98635.55, 99166.78, 100759.6, 100937.4, 101021.5, 
    101102.5, 101180.5, 101244.2, 101299.7, 101351.9, 101396, 101441, 101474.8,
  97657.3, 97537.54, 98808.49, 99182.13, 99846.57, 100856.8, 100986.8, 
    101056, 101138.2, 101210.5, 101271.1, 101329.2, 101379.6, 101428.5, 
    101468.6,
  97657.96, 96278.23, 96161.46, 97339.98, 99027.72, 99814.74, 100930.5, 
    101016.7, 101087.6, 101174.4, 101239.2, 101304.4, 101360.4, 101417.8, 
    101465.8,
  101030.8, 101122.4, 101196.4, 101271.5, 101348, 101424, 101498.3, 101574.3, 
    101653.3, 101716, 101772.3, 101809.4, 101843.6, 101863.3, 101876.5,
  99522.12, 100906.8, 100982.3, 101023.7, 101129.8, 101212.9, 101302.2, 
    101387.9, 101462.6, 101538.2, 101606.6, 101665.5, 101719.8, 101766.9, 
    101810.3,
  99482.53, 100493.6, 100887.9, 100927.1, 100997.5, 101067.2, 101139, 
    101209.3, 101289, 101370.4, 101452.9, 101527.5, 101593.9, 101655, 101716,
  99092.67, 100310.9, 100757.4, 100828.6, 100902.7, 100975.3, 101049.7, 
    101114.6, 101174.8, 101233.3, 101304.2, 101379.5, 101449.6, 101510.6, 
    101565.6,
  98998.35, 99667.25, 100546.7, 100766.2, 100849.2, 100920, 101012.1, 
    101087.8, 101152.7, 101210.4, 101261.2, 101311.4, 101362.2, 101411.2, 
    101460.2,
  98712.11, 98525.48, 99373.04, 100622.4, 100769, 100854.7, 100955, 101048.3, 
    101138.2, 101210.2, 101272.9, 101334.3, 101387.3, 101436.5, 101478.2,
  98616.99, 97945.85, 97890.94, 99591.24, 100679.9, 100785.1, 100894.8, 
    100996.7, 101100.2, 101187.1, 101263.7, 101337, 101400.2, 101460.4, 
    101511.5,
  98745.66, 98063.6, 98442.32, 98948.58, 100519.4, 100701, 100823.3, 
    100932.1, 101052, 101154.8, 101247.4, 101333.1, 101409, 101481.1, 101542.9,
  97564.03, 97424.42, 98614.12, 98957.27, 99603.93, 100593.5, 100770.6, 
    100870.6, 100997.2, 101109.1, 101212.3, 101310, 101397.3, 101481.9, 
    101554.4,
  97596.28, 96140.39, 95997.88, 97127.56, 98827.92, 99548.39, 100695.2, 
    100817.3, 100936.6, 101064.8, 101177.4, 101284.2, 101380, 101471.8, 101554,
  101542.6, 101544.5, 101529.1, 101521.7, 101507.1, 101494.6, 101481.3, 
    101476.9, 101489.9, 101509.5, 101527.4, 101531, 101526.6, 101513.5, 
    101493.6,
  100078.6, 101400.9, 101390.7, 101350.1, 101321.1, 101309.7, 101304.9, 
    101304.7, 101307.8, 101315.1, 101328.2, 101343.9, 101361.4, 101367.9, 
    101377.1,
  99996.41, 100959.2, 101247.2, 101195.6, 101161.1, 101135.1, 101128.9, 
    101130.7, 101145.6, 101171.9, 101210.2, 101238.1, 101254.4, 101268.8, 
    101280.9,
  99583.9, 100776.1, 101077.7, 101015.4, 100947.3, 100898.4, 100877, 
    100872.8, 100894.8, 100927.1, 100956.7, 100995.9, 101028.9, 101056.9, 
    101088.5,
  99414.19, 99997.31, 100767.8, 100863.8, 100778, 100712.9, 100683.6, 
    100676.3, 100701.9, 100727, 100776.7, 100838.5, 100853.5, 100881, 100924.2,
  99032.68, 98791.07, 99582.55, 100684.6, 100645.5, 100534.4, 100473.7, 
    100475.2, 100509.8, 100573.3, 100641, 100695.2, 100738.5, 100753.5, 
    100799.2,
  98870.36, 98152.27, 98005.98, 99629.62, 100508.2, 100405.3, 100264.3, 
    100208.1, 100216.1, 100308, 100378.5, 100458.9, 100583.8, 100658.5, 
    100762.1,
  99083.06, 98248.56, 98507.23, 98932.72, 100339.7, 100320.3, 100177.3, 
    100079.2, 100044.9, 100081.6, 100164.9, 100309, 100463.2, 100598.8, 
    100707.4,
  97866.61, 97603.55, 98697.93, 98918.71, 99400.71, 100219.1, 100175.4, 
    100086.8, 100047.3, 100056.9, 100145.2, 100286.3, 100436.5, 100588.1, 
    100724.8,
  97843.43, 96341.86, 96097.12, 97100.65, 98641.33, 99279.23, 100157.5, 
    100122, 100073.1, 100095.9, 100182.6, 100310, 100445.7, 100590.7, 100730.8,
  101689.7, 101691, 101647.1, 101614.8, 101570.7, 101517.7, 101473.7, 
    101426.3, 101382.8, 101347.4, 101317.2, 101290.9, 101275.6, 101270.9, 
    101268,
  100272.2, 101636.6, 101616.6, 101583.5, 101531.8, 101475.7, 101423.8, 
    101362.9, 101307.2, 101248.3, 101198.7, 101156.5, 101123.6, 101092.2, 
    101080,
  100334.7, 101291.6, 101589.8, 101544.2, 101490.6, 101430.8, 101361.1, 
    101283.9, 101199.9, 101120, 101049.6, 100980.3, 100928.5, 100904.4, 
    100913.4,
  99997.46, 101209.3, 101543, 101519.8, 101454.8, 101384.4, 101298.6, 101205, 
    101097.4, 100987.4, 100862.2, 100756.5, 100683.7, 100624.4, 100566.8,
  99930.05, 100560.9, 101351.2, 101487.9, 101412.8, 101338, 101243.9, 
    101130.8, 100987.4, 100831.8, 100663.8, 100542.7, 100413.3, 100344.4, 
    100330.4,
  99610.66, 99379.88, 100208.9, 101392.9, 101386.6, 101300.7, 101196.4, 
    101067.1, 100892.8, 100712, 100493.7, 100296.2, 100095.9, 100009.2, 
    99947.78,
  99481.6, 98786.71, 98690.44, 100390.2, 101352, 101276, 101161.2, 101021.6, 
    100830.7, 100620.1, 100343.8, 99997.64, 99727.81, 99626.8, 99544.51,
  99681.93, 98920.37, 99280.71, 99751.67, 101263, 101257.8, 101147.6, 
    101005.3, 100815.3, 100593.1, 100288.5, 99869.84, 99503.92, 99301.7, 
    99214.64,
  98428.52, 98268.85, 99503.65, 99798.88, 100356.1, 101215.2, 101147.6, 
    101003.9, 100822.5, 100619.4, 100337.9, 99991.5, 99633.4, 99364.51, 
    99218.02,
  98363.49, 96908.81, 96775.34, 97933.96, 99556.85, 100278.5, 101147.2, 
    101045.9, 100857, 100670.9, 100418.7, 100131.2, 99822.9, 99556.52, 
    99388.32,
  101548.3, 101594.8, 101594.9, 101575.1, 101557.1, 101524.5, 101481.2, 
    101428.4, 101364.5, 101293.1, 101215, 101133.5, 101045.8, 100955.5, 
    100858.3,
  100140.6, 101558.1, 101595.8, 101586.8, 101568.5, 101544.2, 101508.1, 
    101459.2, 101399.9, 101329.4, 101250.4, 101163.3, 101070, 100971.2, 
    100865.7,
  100233.6, 101234.1, 101590.4, 101589.9, 101571.8, 101551.7, 101520.2, 
    101476, 101420.4, 101352.7, 101275.8, 101187, 101092.2, 100982.9, 100867.2,
  99899.77, 101164.5, 101546.5, 101583.2, 101570.4, 101552.2, 101525.9, 
    101488.7, 101438.2, 101371.2, 101297.5, 101209.3, 101112, 100996.2, 
    100864.5,
  99847.27, 100518.6, 101373.5, 101560.4, 101560.4, 101544.2, 101523.8, 
    101491, 101445.1, 101385.9, 101315.1, 101228.3, 101129.4, 101005, 100857.9,
  99533.41, 99333.83, 100227, 101466.1, 101539.1, 101531, 101518.8, 101492, 
    101448, 101394.4, 101328.7, 101246.8, 101148, 101020.6, 100869.7,
  99395.57, 98742.24, 98712.29, 100460.3, 101500.4, 101512.6, 101497.5, 
    101480.4, 101444, 101396.3, 101336.2, 101260.7, 101168.8, 101042.5, 
    100891.4,
  99585.23, 98866.84, 99292.75, 99805.88, 101397.4, 101483.8, 101476.7, 
    101458.9, 101429.6, 101391.4, 101338.9, 101272.6, 101188.9, 101078.7, 
    100936.5,
  98331.58, 98206.2, 99494.3, 99832.88, 100476.9, 101423.2, 101455.3, 
    101432.8, 101412.4, 101380.4, 101334.4, 101276.1, 101204.8, 101111.5, 
    100988,
  98292.94, 96854.16, 96747.09, 97964.87, 99664.22, 100427.1, 101424.2, 
    101431.4, 101391.5, 101368.5, 101323.4, 101278.9, 101219.9, 101146.4, 
    101046.1,
  101494.1, 101589.5, 101639.4, 101677, 101715.4, 101743.3, 101761.1, 
    101774.6, 101781.8, 101787, 101785, 101781.2, 101785.7, 101800, 101806.1,
  100120.8, 101554.6, 101639.6, 101680.2, 101724.9, 101761.9, 101785.5, 
    101798.8, 101806.1, 101811.4, 101802.9, 101795.3, 101797.5, 101804.4, 
    101813.6,
  100211.4, 101234.1, 101635.7, 101683.8, 101721.8, 101764.1, 101795.1, 
    101818.6, 101831.3, 101845, 101844.4, 101837.8, 101827, 101815.1, 101808.8,
  99880.98, 101165.4, 101591.7, 101663.6, 101701.2, 101745.7, 101787.2, 
    101815.4, 101838, 101848, 101851.9, 101859.8, 101854, 101845.2, 101834.9,
  99810.3, 100502.7, 101404.5, 101627.8, 101678.6, 101719.5, 101762.1, 
    101795.3, 101821.2, 101843.3, 101859, 101868.7, 101867.7, 101868.6, 
    101858.8,
  99488.17, 99318.63, 100226.1, 101511.5, 101627.6, 101681.3, 101726.5, 
    101765.2, 101796.8, 101822.3, 101842.4, 101858.8, 101868.8, 101871.5, 
    101870.2,
  99357.06, 98732.92, 98728.77, 100487.6, 101568.5, 101628.8, 101676.9, 
    101718.7, 101754.1, 101784.1, 101810.8, 101832.6, 101848.7, 101864, 
    101867.4,
  99541.47, 98843.86, 99298.86, 99824.25, 101433.2, 101564.5, 101612.8, 
    101659.6, 101699.7, 101734.7, 101767, 101797.9, 101821, 101839.6, 101851.4,
  98290.52, 98177.59, 99477.54, 99840.7, 100501.7, 101479.9, 101554.7, 
    101596, 101638.1, 101680.4, 101714, 101748.9, 101778, 101806.4, 101824.2,
  98261.39, 96839.39, 96733.22, 97956.59, 99654.62, 100435.6, 101490.1, 
    101535.9, 101561.1, 101608.9, 101649.5, 101690.5, 101726.2, 101755, 
    101783.8,
  100928.4, 101031.1, 101086, 101135.7, 101206.5, 101266.9, 101333.3, 
    101395.4, 101464.8, 101528.6, 101589.3, 101646.7, 101696.9, 101744.9, 
    101789.3,
  99581.08, 100997.9, 101101, 101153.6, 101222.3, 101287.9, 101357.4, 
    101423.9, 101497.2, 101566.4, 101625.5, 101685.1, 101739.4, 101790.5, 
    101839.1,
  99697.18, 100702.8, 101102.1, 101156.1, 101221.9, 101292.4, 101364.3, 
    101430.8, 101508.4, 101579.2, 101641.9, 101708.3, 101764.5, 101817.1, 
    101870,
  99392.07, 100648.9, 101079.2, 101149.3, 101210.3, 101276.2, 101356.1, 
    101428.6, 101506.1, 101581, 101647, 101712, 101770.6, 101827.8, 101879.8,
  99360.92, 100015.6, 100915.7, 101131.7, 101197.3, 101253.4, 101332.4, 
    101407.8, 101487, 101565.4, 101635.2, 101700.8, 101762.5, 101820.1, 
    101879.5,
  99059.62, 98878.95, 99763.51, 101036.1, 101168.9, 101228.3, 101301.6, 
    101379.6, 101458.4, 101536, 101608.7, 101677.4, 101739.4, 101799.2, 
    101853.8,
  98958.12, 98326.57, 98320.53, 100033.6, 101128.2, 101194.8, 101266.4, 
    101339.1, 101420.1, 101496.3, 101567.6, 101639.5, 101702.9, 101765.2, 
    101825.2,
  99165.02, 98455.73, 98903.77, 99407.1, 101006.1, 101153.8, 101226.4, 
    101297.5, 101372.9, 101448.3, 101517.6, 101586.7, 101652.1, 101716, 
    101779.1,
  97967.33, 97818.13, 99093.56, 99453.65, 100099.4, 101084.4, 101190.3, 
    101248.8, 101319.6, 101390.8, 101458.4, 101523.8, 101590, 101655.6, 101717,
  97975.63, 96543.12, 96414.42, 97583.27, 99272.8, 100049.8, 101138.6, 
    101212.1, 101266.2, 101331.6, 101396.3, 101461.1, 101517.8, 101582.3, 
    101649.4,
  100173, 100234.3, 100277, 100313.7, 100355.6, 100401.5, 100457.9, 100519.1, 
    100585.6, 100655.3, 100725.4, 100796.5, 100868, 100941.1, 101013.2,
  98865.02, 100219.9, 100320.9, 100367.1, 100422.2, 100475, 100535.8, 
    100602.1, 100668.6, 100734.1, 100797.7, 100865.4, 100926.1, 100994.9, 
    101059.7,
  99019.13, 99978.36, 100356.1, 100410.4, 100467.3, 100520.8, 100586.8, 
    100652.5, 100716.4, 100780.4, 100842, 100907.5, 100963.9, 101029.5, 
    101087.2,
  98754.55, 99957.24, 100374.6, 100446.8, 100508.8, 100561.6, 100630, 
    100694.6, 100757, 100813.4, 100870, 100926.8, 100979.6, 101035.6, 101088.7,
  98769.72, 99392.18, 100247.7, 100470, 100536.9, 100591.9, 100655.3, 100720, 
    100778.4, 100832.5, 100885.6, 100934.5, 100980.6, 101025.9, 101067.2,
  98516.98, 98323.78, 99164.05, 100414.9, 100552.4, 100610.2, 100673, 
    100734.7, 100794.3, 100843.1, 100890.5, 100933.6, 100967.8, 100997.6, 
    101023.8,
  98456.23, 97827.7, 97785.59, 99461.59, 100547.8, 100618.9, 100677, 
    100735.5, 100795.7, 100843.8, 100887.6, 100919.4, 100945.3, 100958.3, 
    100968.8,
  98705.91, 97983.52, 98396.88, 98884.59, 100460.2, 100615.5, 100677, 
    100731.8, 100790.3, 100835.6, 100872.8, 100896.8, 100914.2, 100915.2, 
    100915.3,
  97572.5, 97392.52, 98626.04, 98968.98, 99591.25, 100567.7, 100674.6, 
    100715.1, 100776.4, 100818, 100850.5, 100870.4, 100882.1, 100878.8, 
    100869.1,
  97636.66, 96195.31, 96031.48, 97153.99, 98829.55, 99587.41, 100667.5, 
    100713.8, 100744.6, 100793.6, 100816.3, 100834.2, 100842.8, 100839.4, 
    100828.9,
  101190.6, 101157.5, 101090.6, 101014.2, 100953.6, 100875.5, 100798.4, 
    100738.6, 100683.8, 100624.9, 100548.2, 100473, 100409.8, 100364.3, 
    100325.2,
  99737.02, 101088.5, 101076.7, 101006.3, 100958.8, 100895.7, 100839.2, 
    100767.7, 100691.8, 100623.6, 100572.4, 100526.6, 100486.8, 100450.1, 
    100414.8,
  99760, 100734.1, 101044.1, 100972.9, 100938.1, 100885.1, 100830.1, 100772, 
    100720.7, 100673.3, 100631.7, 100595.9, 100563, 100527.7, 100490.4,
  99400.24, 100628.4, 100979.7, 100944.3, 100910, 100869.5, 100831.2, 100787, 
    100743.8, 100705.5, 100671.5, 100643.1, 100619.2, 100587.6, 100551.6,
  99306.41, 99971.63, 100797.5, 100920, 100881, 100851.4, 100821.2, 100789.1, 
    100757.6, 100731.5, 100710.4, 100690, 100667.8, 100640.4, 100607,
  98968.09, 98800.42, 99640.76, 100839.9, 100861.5, 100835.4, 100817.1, 
    100800.1, 100778.5, 100763.6, 100745.8, 100730.8, 100712.5, 100690.1, 
    100659.5,
  98816.81, 98213.18, 98168.11, 99839.01, 100835.6, 100827.8, 100805.6, 
    100797.2, 100785.6, 100778.8, 100768.6, 100757.7, 100744.2, 100728.3, 
    100706.2,
  99041.54, 98313.12, 98719.26, 99215.18, 100742, 100808.8, 100796.7, 
    100790.8, 100787.7, 100786.5, 100779.8, 100770.9, 100763.2, 100751.4, 
    100736.4,
  97868.59, 97690.28, 98921.38, 99274.91, 99850.05, 100747.6, 100772.3, 
    100762.6, 100770.8, 100779.1, 100780.7, 100782.4, 100773.4, 100773.3, 
    100764.1,
  97901.68, 96462.89, 96302, 97415.02, 99065.31, 99794.59, 100769.6, 
    100772.4, 100753.4, 100773.6, 100775.5, 100784.2, 100785.3, 100788.3, 
    100793.2,
  101514.1, 101597.5, 101621.2, 101627.1, 101647.9, 101647.3, 101643.3, 
    101636.5, 101621.9, 101603.5, 101577.2, 101545.8, 101508.5, 101470.2, 
    101424.2,
  100138.9, 101561.6, 101634.1, 101637.5, 101666, 101664.1, 101659.7, 
    101656.1, 101645.9, 101634.6, 101612.1, 101587.8, 101554.1, 101516.3, 
    101475.1,
  100216.4, 101247.8, 101619.4, 101639.4, 101657.4, 101666.4, 101672.8, 
    101673, 101665.5, 101653.8, 101635.2, 101616.8, 101589.4, 101557.7, 
    101518.7,
  99874.88, 101165.9, 101581.2, 101637.8, 101654.1, 101668, 101668.3, 
    101666.2, 101666.2, 101663.3, 101646.9, 101628.8, 101605.6, 101577.2, 
    101541,
  99800.54, 100507.6, 101407.4, 101604.7, 101635.4, 101650.5, 101662, 
    101660.8, 101661.7, 101657.4, 101645.4, 101630.1, 101608.2, 101581.5, 
    101552.6,
  99461.91, 99312.27, 100236.5, 101519.4, 101602.1, 101615, 101631.8, 
    101640.6, 101638.3, 101635.8, 101629.9, 101617.1, 101597.4, 101574.6, 
    101547.4,
  99304, 98717.9, 98702.51, 100476.5, 101545.7, 101583.8, 101593, 101598.5, 
    101604, 101607.3, 101595.3, 101585.1, 101565.8, 101542.4, 101515.5,
  99490.59, 98819.26, 99263.42, 99806.59, 101418, 101526, 101545.3, 101555.9, 
    101558.9, 101558.3, 101548.2, 101536.6, 101519.7, 101502.2, 101484.2,
  98238.55, 98136.42, 99452.11, 99828.82, 100478.7, 101445.3, 101498.5, 
    101499.3, 101506.8, 101504.5, 101493.3, 101484, 101466.1, 101448.2, 
    101424.2,
  98202.16, 96812.06, 96714.95, 97924.23, 99635.98, 100436.2, 101450.3, 
    101462.5, 101440.8, 101441.6, 101428.7, 101418.4, 101396.6, 101380, 
    101364.9,
  100940.4, 101052.9, 101126.9, 101210.3, 101301.9, 101379.9, 101456.7, 
    101527.4, 101596.9, 101661, 101719, 101769.9, 101814.8, 101855.8, 101889,
  99571.16, 100999.6, 101118.1, 101200.1, 101290.1, 101380.3, 101459.8, 
    101533.9, 101606.6, 101672.9, 101732.9, 101793.7, 101843.8, 101887.2, 
    101928,
  99650.09, 100676.8, 101094.5, 101181.9, 101266.9, 101361, 101446.6, 101523, 
    101596.2, 101665.9, 101729, 101791.1, 101846.7, 101896, 101939.2,
  99309.8, 100589.8, 101049.1, 101151.4, 101240.3, 101334.4, 101424.6, 
    101505.6, 101580.3, 101648.8, 101714.7, 101778.8, 101837.6, 101891.8, 
    101936.9,
  99237.08, 99915.45, 100854, 101107.5, 101198.8, 101291.4, 101385.8, 
    101473.5, 101546.5, 101620.4, 101685.9, 101751.4, 101810.9, 101869.9, 
    101919,
  98908.3, 98752.48, 99663.29, 100989.3, 101151.5, 101244.3, 101337.7, 
    101431.7, 101508.1, 101581.9, 101646.6, 101713.6, 101774.7, 101836.7, 
    101890.4,
  98789.54, 98190.2, 98207.3, 99952.88, 101089.2, 101194.2, 101285.2, 
    101379.6, 101460.1, 101530.4, 101597.1, 101659.4, 101720, 101780.4, 101839,
  98983.88, 98307.59, 98776.89, 99318.76, 100946.4, 101129.8, 101225.9, 
    101316.5, 101403.4, 101476.8, 101539.9, 101600.1, 101655.9, 101713.4, 
    101769.5,
  97789.06, 97659.7, 98955.41, 99349.55, 100029.1, 101053.1, 101181, 
    101257.8, 101340.6, 101413.9, 101473.7, 101531.2, 101584.2, 101636.2, 
    101689.5,
  97807.69, 96404.14, 96292.53, 97474.15, 99195.78, 100000.6, 101130.2, 
    101209.4, 101274.2, 101347.7, 101400.8, 101448.6, 101491.5, 101538.7, 
    101591,
  100790.1, 100799.9, 100805.1, 100797.1, 100818.1, 100823.9, 100838.9, 
    100857.8, 100889.3, 100928.7, 100976.3, 101028.6, 101078.6, 101118.4, 
    101163.5,
  99342.13, 100693.9, 100755.3, 100752.2, 100782.4, 100803.1, 100826.6, 
    100853.6, 100885, 100928.5, 100975.7, 101030.9, 101092.7, 101133.4, 
    101166.2,
  99349.83, 100331.7, 100708.3, 100720.5, 100751.3, 100793.6, 100833, 
    100867.2, 100903.8, 100946.6, 100992.2, 101041.7, 101092.3, 101132.2, 
    101165.9,
  98980.73, 100212.1, 100624.2, 100665, 100707.9, 100756.8, 100812.2, 
    100858.8, 100903.4, 100940.6, 100984.5, 101033.1, 101076.5, 101109.8, 
    101143.2,
  98894.05, 99539.59, 100417.8, 100611.4, 100663.4, 100710.9, 100784.8, 
    100850.9, 100905.5, 100950, 100989.9, 101024.3, 101061.2, 101096.3, 
    101142.7,
  98578.47, 98385.03, 99245.33, 100491.3, 100607.1, 100656.9, 100734.2, 
    100802.7, 100872.7, 100929.4, 100973.3, 101012.3, 101047.9, 101093.4, 
    101139.8,
  98473.59, 97830.62, 97800.74, 99481.56, 100542, 100596.1, 100679, 100768.8, 
    100849.5, 100918.1, 100964.9, 101008.2, 101044.3, 101084.7, 101128.6,
  98688.3, 97943.45, 98350.02, 98849.85, 100420, 100537.3, 100624.2, 
    100721.8, 100809.7, 100892, 100950.1, 100997.8, 101034.4, 101075.9, 
    101120.5,
  97533.53, 97355.86, 98586.5, 98921.98, 99507.77, 100462.4, 100592.5, 
    100691.4, 100785.3, 100869.9, 100937.1, 100985.7, 101026.2, 101067.3, 
    101121,
  97580.52, 96165.22, 95999.34, 97111.06, 98785.54, 99494.42, 100563.9, 
    100667.9, 100753.9, 100847.2, 100916.2, 100971.9, 101017.5, 101059.8, 
    101123.4,
  100800.9, 100810.8, 100802.3, 100794.5, 100780.6, 100760.5, 100746.5, 
    100724.9, 100709.5, 100683.5, 100658.9, 100637.4, 100630.5, 100637.1, 
    100669,
  99340.11, 100692.4, 100719.6, 100702, 100700.6, 100685.4, 100677.8, 
    100660.3, 100646.1, 100626.6, 100615.7, 100593.4, 100588.5, 100596.7, 
    100594.6,
  99338.75, 100308.2, 100641.3, 100632.5, 100628.6, 100619.9, 100615.6, 
    100602.2, 100584.7, 100557.8, 100527.5, 100502.9, 100493.3, 100486.4, 
    100537,
  98937.48, 100175.8, 100548.6, 100552, 100529.3, 100530.8, 100524.2, 
    100523.4, 100528.5, 100528.4, 100525.8, 100519.3, 100516.4, 100547.8, 
    100620.6,
  98844, 99473.16, 100294.5, 100458.3, 100444.5, 100441.8, 100455.5, 
    100464.7, 100467.8, 100479.2, 100474.8, 100453.4, 100453.5, 100504.4, 
    100582.1,
  98427.24, 98268.98, 99101.6, 100310.2, 100354, 100363.8, 100381.6, 
    100400.9, 100426.2, 100448.8, 100464.1, 100479.1, 100500.4, 100576.3, 
    100679,
  98240.91, 97669.28, 97569.67, 99259.18, 100265.9, 100289.2, 100321.8, 
    100367.2, 100404.7, 100446.7, 100485.7, 100526.5, 100569.9, 100629.9, 
    100699.7,
  98423.48, 97741.23, 98130.12, 98624.52, 100150.2, 100234.4, 100256.5, 
    100318.2, 100373, 100429.9, 100484, 100538.3, 100592.2, 100672, 100764.7,
  97307.93, 97118.74, 98327.74, 98668.77, 99259.6, 100186.6, 100248, 
    100296.7, 100367.4, 100437.6, 100508.1, 100580.3, 100645.8, 100729.4, 
    100803.5,
  97423.24, 95937.34, 95781.44, 96885.27, 98546.23, 99245.15, 100235.8, 
    100284.2, 100349.9, 100440.1, 100512.7, 100597.9, 100675, 100764.7, 
    100853.5,
  100977.5, 100997.6, 100983.5, 100966.7, 100953, 100923.3, 100901, 100878.2, 
    100860.9, 100842.1, 100812.4, 100772.9, 100729.3, 100688.2, 100655.6,
  99577.43, 100925.7, 100927.6, 100885.4, 100870.1, 100841.6, 100827.5, 
    100801.5, 100780.2, 100760.6, 100740.6, 100710.6, 100670.9, 100619.5, 
    100561.6,
  99631.55, 100573.8, 100888.1, 100871.7, 100849.8, 100812.6, 100797.2, 
    100769, 100749.5, 100726.4, 100693.1, 100640.7, 100587.4, 100524.8, 
    100461.3,
  99288.27, 100481.8, 100829, 100812.9, 100794.3, 100783.1, 100744.3, 
    100702.9, 100667.5, 100637.8, 100612, 100585.1, 100531.4, 100442.3, 
    100352.6,
  99227, 99831.5, 100649.9, 100798.7, 100768.2, 100734.8, 100692.5, 100656.5, 
    100616.2, 100582.4, 100535.6, 100483.6, 100415.9, 100351.4, 100310.7,
  98920.28, 98668.51, 99509.72, 100683.7, 100693.9, 100652.7, 100604.4, 
    100552.5, 100482.7, 100438.1, 100409.4, 100391.3, 100362.2, 100319.2, 
    100281.6,
  98783.49, 98092.03, 97989.75, 99658.36, 100611.1, 100560.6, 100512, 
    100470.8, 100411.4, 100371.5, 100336, 100316, 100288.7, 100258.3, 100240.6,
  98980.27, 98222, 98549.73, 98999.49, 100502.6, 100541.1, 100475.6, 
    100437.2, 100385.9, 100350.4, 100324.9, 100321.7, 100320.1, 100321.2, 
    100323.6,
  97772.9, 97585.36, 98776.23, 99081.71, 99634.21, 100492.1, 100478.4, 
    100436.3, 100401.3, 100387.4, 100378.9, 100383.4, 100389.7, 100404.7, 
    100427,
  97780.59, 96312.81, 96147.62, 97244.79, 98869.13, 99590.44, 100513.6, 
    100491.3, 100428.8, 100435.6, 100429.1, 100447.2, 100468.2, 100501.9, 
    100532.2,
  101495.5, 101549.1, 101566.3, 101562.1, 101564.9, 101553.3, 101542.6, 
    101528.5, 101508.4, 101482.8, 101453.8, 101423, 101388.9, 101351.2, 
    101314.4,
  100120, 101526.9, 101584.1, 101586.7, 101597.5, 101591.5, 101582.4, 
    101567.8, 101551.3, 101528.7, 101504, 101476, 101442.7, 101407, 101368.6,
  100244.1, 101231.6, 101597.1, 101604.5, 101612.6, 101606.3, 101604.4, 
    101589.9, 101576.6, 101556.9, 101536, 101512.2, 101483.2, 101451, 101413.3,
  99930.84, 101178.3, 101572.2, 101602.2, 101606.3, 101614.2, 101611.5, 
    101602.1, 101591.4, 101576.4, 101556.3, 101533.6, 101508.1, 101477, 
    101439.9,
  99880.05, 100543.1, 101395.8, 101588.2, 101600.5, 101604.8, 101606.9, 
    101602.9, 101593.6, 101577, 101559.5, 101536.4, 101512.4, 101480.5, 
    101444.3,
  99567.73, 99385.09, 100265.6, 101502.9, 101578.7, 101585.6, 101588.9, 
    101590.5, 101579, 101562.2, 101540.9, 101516.7, 101490.4, 101457.4, 
    101417.5,
  99437.71, 98796.09, 98759.04, 100506.2, 101543.3, 101563.7, 101563.3, 
    101561.5, 101548.2, 101529.6, 101507.3, 101480.4, 101450.5, 101414.2, 
    101377.4,
  99635.18, 98928.7, 99352.73, 99867.48, 101446, 101532.6, 101535.2, 
    101529.7, 101510, 101489.9, 101461.4, 101427.7, 101389.8, 101355.1, 101319,
  98382.93, 98257.85, 99530.83, 99878.48, 100509.6, 101460.4, 101500.6, 
    101481.5, 101463.9, 101438.2, 101400.8, 101365.7, 101327.7, 101292.4, 
    101253.6,
  98344.02, 96926.55, 96831.22, 98020.73, 99706.13, 100464.3, 101443.4, 
    101451.2, 101402, 101380.1, 101336.9, 101307.2, 101258.1, 101212.8, 
    101175.3,
  100908.5, 100971.9, 100987.2, 100982, 100982.3, 100979.6, 100978.4, 
    100975.7, 100973.4, 100971.7, 100969.4, 100970.9, 100973.3, 100983.2, 
    100998.8,
  99643.1, 101031, 101089.6, 101095.8, 101102.2, 101107.2, 101110.2, 
    101110.7, 101116.3, 101113.8, 101114, 101111.7, 101115.8, 101120.9, 
    101131.2,
  99826.16, 100802, 101154.8, 101176, 101186, 101197.6, 101206.5, 101212.1, 
    101216.9, 101221.1, 101226.3, 101227.9, 101238, 101240.7, 101248.5,
  99557.12, 100795.4, 101195.2, 101237.1, 101249.2, 101270.1, 101283, 
    101295.6, 101303.3, 101310.1, 101314.8, 101320.9, 101325.9, 101331.4, 
    101338.5,
  99537.76, 100189.9, 101054.4, 101261.5, 101284.5, 101307.2, 101326.5, 
    101346.8, 101357.1, 101366.8, 101373.9, 101381.3, 101389.6, 101397.5, 
    101404.6,
  99247.45, 99060.65, 99941.51, 101198.8, 101300.9, 101329.2, 101350.9, 
    101375.8, 101385.7, 101397.6, 101405.3, 101415.2, 101422.5, 101428.3, 
    101434.2,
  99137.45, 98506.91, 98484.66, 100219, 101282.7, 101325.4, 101349.5, 
    101373.8, 101391.5, 101403.5, 101410.7, 101419.7, 101426.1, 101435.4, 
    101437.1,
  99337.92, 98644.52, 99079.77, 99590.31, 101186.7, 101304.9, 101335.9, 
    101358.5, 101376.2, 101388.9, 101394.6, 101401.5, 101406.4, 101410.9, 
    101411.5,
  98094.42, 97981.76, 99279.75, 99636.48, 100280.8, 101249, 101311.2, 
    101329.7, 101344.7, 101355.8, 101359.7, 101366.3, 101367.5, 101372.8, 
    101370.9,
  98083.59, 96668.59, 96555.68, 97769.47, 99462.55, 100242.6, 101283.1, 
    101305.4, 101300.6, 101308.5, 101306.9, 101311.2, 101312.1, 101315, 
    101305.8,
  100587.9, 100602.5, 100590.7, 100577.2, 100571.4, 100562, 100551.4, 
    100536.8, 100516.6, 100495, 100474.1, 100454.9, 100441.3, 100429.7, 
    100421.2,
  99197.08, 100564.7, 100604.5, 100599.7, 100601.3, 100595.6, 100587.3, 
    100577, 100567.4, 100557.5, 100549.9, 100541.6, 100533.4, 100527.9, 100528,
  99266.62, 100248, 100598.2, 100594.6, 100600.6, 100601.6, 100604, 100607, 
    100607.9, 100608.5, 100608, 100608.1, 100614.7, 100623.4, 100636,
  98966.88, 100185.3, 100589.1, 100612.4, 100622.3, 100630.4, 100638.6, 
    100646.2, 100651, 100656.2, 100662.8, 100671.6, 100684.6, 100697.6, 
    100712.6,
  98925.12, 99563.8, 100425.2, 100615.1, 100625.9, 100635.1, 100650.9, 
    100667.6, 100679.5, 100693.8, 100704.1, 100713.2, 100727.6, 100744.1, 
    100769.2,
  98635.74, 98444.91, 99300.74, 100547.3, 100629.4, 100641.9, 100661.9, 
    100686.1, 100702.7, 100713, 100722.4, 100732.5, 100746, 100765.4, 100777.1,
  98532.02, 97900.81, 97845.89, 99546.51, 100609.5, 100638.1, 100653.8, 
    100683, 100705, 100716, 100720.5, 100725.1, 100729.4, 100742.8, 100751,
  98763.98, 98044.19, 98430.89, 98919.87, 100500.5, 100613.4, 100641.1, 
    100667.6, 100686.7, 100699.5, 100698.8, 100697.3, 100689.6, 100698.4, 
    100719.7,
  97580.24, 97406.14, 98639.09, 98973.65, 99576.56, 100538.9, 100621, 
    100643.4, 100659.8, 100675.4, 100663.9, 100658.8, 100642.7, 100658.8, 
    100675,
  97626.57, 96165.7, 96009.48, 97111.59, 98771.17, 99525.98, 100587.1, 
    100623.8, 100627.2, 100654.8, 100627.9, 100609.8, 100592.8, 100590.8, 
    100601.7,
  101532.4, 101522.5, 101470, 101417.7, 101388.2, 101356.9, 101330.6, 
    101310.8, 101286.7, 101261.7, 101232, 101197.8, 101162.8, 101130.9, 
    101095.5,
  100044, 101444.3, 101462.6, 101400, 101372.5, 101330.1, 101296.7, 101266, 
    101237.7, 101209.2, 101183.1, 101155.4, 101123.8, 101087.8, 101055.6,
  100108.5, 101093.6, 101427.2, 101373.7, 101345.2, 101302.3, 101265.9, 
    101232.3, 101204.7, 101180.6, 101152, 101121.4, 101089.5, 101056.6, 
    101019.5,
  99740.58, 100984.1, 101364.1, 101340.6, 101306.5, 101266.2, 101227.6, 
    101193.3, 101161.2, 101130.3, 101098.4, 101066.9, 101036.9, 101008.3, 
    100975.5,
  99631.45, 100289.7, 101141.5, 101291.8, 101263.1, 101226.6, 101188.3, 
    101145.3, 101111.1, 101074.3, 101048.1, 101019.5, 100992.2, 100963.5, 
    100932.8,
  99281.86, 99098.61, 99960.16, 101177.9, 101216.6, 101176.3, 101142.8, 
    101106, 101064, 101035.4, 101001.9, 100966.7, 100935, 100908.4, 100883.4,
  99115.92, 98501.87, 98444.95, 100162.8, 101162.5, 101145.3, 101105.9, 
    101073.7, 101034.3, 100998.2, 100963.8, 100924, 100899.9, 100871.1, 
    100833.8,
  99299.84, 98597.45, 99007.63, 99505.23, 101054.5, 101110.7, 101077.4, 
    101046.5, 101007.1, 100968.4, 100936.2, 100900.4, 100865.1, 100830.2, 
    100794.6,
  98068, 97934.26, 99198.57, 99535.66, 100133.9, 101039.6, 101046.4, 
    101009.8, 100972.2, 100943.4, 100909, 100883.7, 100841.4, 100812, 100777.4,
  98042.62, 96621.16, 96499.4, 97658.79, 99315.28, 100074.5, 101013.1, 
    100996.5, 100934.3, 100915, 100876.7, 100848.8, 100816.5, 100785.4, 
    100753.7,
  101830.8, 101886.4, 101889, 101880, 101896.7, 101893.4, 101912.4, 101918.4, 
    101920.7, 101916.4, 101907.6, 101897.5, 101885.7, 101863.3, 101837.3,
  100419.7, 101829.4, 101871.4, 101858, 101888.1, 101882.4, 101893.9, 
    101895.5, 101897.3, 101892.8, 101882, 101871.3, 101855.4, 101836.8, 
    101809.1,
  100512.4, 101509.4, 101855.6, 101851, 101860.8, 101854.5, 101863.5, 
    101862.8, 101870, 101863.4, 101850.3, 101840.2, 101821.1, 101795.9, 
    101761.9,
  100161.5, 101432.5, 101813.5, 101836.4, 101831.1, 101830.4, 101837.2, 
    101836.4, 101837.2, 101829.9, 101821.5, 101803.2, 101777.3, 101748.8, 
    101711,
  100084.7, 100773.5, 101627.3, 101801.3, 101795.7, 101801, 101801.5, 
    101797.1, 101799, 101786.9, 101774.7, 101754, 101730.7, 101694.7, 101648.6,
  99748.94, 99578.77, 100474.4, 101709.1, 101771.2, 101762.9, 101760.6, 
    101757.5, 101750.1, 101742.3, 101728.1, 101704.9, 101673.3, 101636.4, 
    101591.6,
  99589.7, 98963.92, 98929.8, 100697, 101727.9, 101732.8, 101720.8, 101714.6, 
    101701.6, 101691.6, 101673.2, 101649.4, 101619.2, 101575.5, 101522.1,
  99760.64, 99067.1, 99500.24, 100019.3, 101615, 101692, 101678.5, 101672.5, 
    101652.8, 101642.2, 101616.1, 101585.9, 101547.1, 101507.8, 101459.3,
  98469.16, 98364.9, 99664.02, 100031.5, 100658.5, 101605.3, 101645.6, 
    101627, 101607.9, 101588.2, 101552.3, 101522.6, 101486.2, 101448, 101395.3,
  98416.8, 97015.72, 96911.69, 98121.3, 99823.76, 100616.9, 101602.5, 
    101603.8, 101558.4, 101540.5, 101497.6, 101467.2, 101423.8, 101387.1, 
    101337,
  101758.2, 101847.9, 101872.9, 101892, 101923.6, 101935, 101954, 101961.6, 
    101965.7, 101964.7, 101955.6, 101942.2, 101919.8, 101890.5, 101857.1,
  100405.8, 101826.5, 101890.5, 101914.3, 101946.7, 101966.3, 101985.7, 
    101999.1, 102012.6, 102017.6, 102019.1, 102009.5, 101996, 101969.4, 
    101937.6,
  100502.2, 101515.7, 101889.3, 101923.7, 101954.4, 101982.6, 102001.6, 
    102018.2, 102037, 102041.3, 102050.1, 102050.4, 102036.4, 102018.9, 
    101989.2,
  100168.5, 101447.7, 101860.2, 101915.2, 101951.1, 101983.6, 102008.4, 
    102028.6, 102045, 102057.8, 102062.6, 102063, 102059.6, 102044.6, 102021.7,
  100095.2, 100789.2, 101669.1, 101887.1, 101924.7, 101968.6, 101995.4, 
    102022.4, 102037.5, 102050.7, 102060.7, 102061.8, 102060.2, 102045.4, 
    102026.9,
  99752.6, 99591.6, 100502.2, 101781.1, 101888, 101936.6, 101971, 102001, 
    102013.9, 102030.7, 102034.7, 102039.2, 102038.7, 102029, 102009.6,
  99599.1, 98979.8, 98976.18, 100751.1, 101830.1, 101890.3, 101926.3, 101960, 
    101979.6, 101998.2, 102003.6, 102012.7, 102010.3, 101997.6, 101979.8,
  99758.62, 99076.57, 99528.44, 100068, 101695.1, 101822.9, 101875, 101907.9, 
    101931.5, 101951.8, 101960.2, 101965.1, 101957.2, 101951.9, 101935.1,
  98473.18, 98380.57, 99696.09, 100071.2, 100734.4, 101724.8, 101803.2, 
    101845.3, 101869.7, 101893.4, 101899, 101910.6, 101905.1, 101902.1, 
    101886.2,
  98431.27, 97025.8, 96921.5, 98153.23, 99893.06, 100688.2, 101735.7, 
    101783.6, 101793.2, 101824, 101827.8, 101841.1, 101837, 101839.4, 101829.3,
  101674, 101787.3, 101827.4, 101858.3, 101898.3, 101924, 101940.5, 101954.8, 
    101954.3, 101953.9, 101940.5, 101922.9, 101904.3, 101874.9, 101850.3,
  100310.5, 101750.1, 101832.6, 101879.5, 101924.9, 101958.9, 101980.7, 
    101999.2, 102012.3, 102017.5, 102020, 102009.3, 101993.9, 101969.2, 
    101947.1,
  100393.8, 101428.7, 101817.7, 101872.7, 101920.4, 101965.3, 101994.2, 
    102022.9, 102047.1, 102062.3, 102072.2, 102077.8, 102076, 102067.3, 
    102051.4,
  100054.5, 101345.7, 101780.2, 101853.4, 101905.5, 101960.8, 101994.7, 
    102030.7, 102059, 102086.2, 102101, 102115.3, 102121.7, 102119.8, 102112.7,
  99979.63, 100677.8, 101581.8, 101815.1, 101867, 101929.4, 101972, 102015.2, 
    102056.2, 102088, 102109.3, 102131, 102145.7, 102152, 102154.1,
  99633.62, 99481.77, 100407, 101701, 101821.5, 101882.4, 101937.9, 101976.4, 
    102013.5, 102050.1, 102083.8, 102115.1, 102130.6, 102147, 102155.3,
  99485.43, 98881.35, 98887.88, 100664.2, 101760.6, 101825.5, 101883.5, 
    101935.2, 101971, 102011.5, 102038, 102072.5, 102096.9, 102118.2, 102131.2,
  99655.28, 98981.5, 99454.5, 99995.16, 101622.6, 101761, 101816.6, 101875, 
    101915.7, 101957.1, 101984.1, 102018.5, 102039.5, 102063.6, 102079.5,
  98403.75, 98297.07, 99622.66, 100002.6, 100674, 101672.4, 101759.3, 
    101810.6, 101855.8, 101895.2, 101923.8, 101950.9, 101969.8, 101994.3, 
    102010.2,
  98373.82, 96973.38, 96876.5, 98093.63, 99845.85, 100631.4, 101702.6, 
    101751, 101787.4, 101823.7, 101853.3, 101875.8, 101897.3, 101917, 101934.8,
  101788.3, 101928.9, 101988.1, 102047.7, 102090.1, 102117, 102130.4, 
    102134.9, 102129.8, 102120.5, 102109.8, 102097.4, 102080.1, 102051.2, 
    102019,
  100398.6, 101855.9, 101959.3, 102030.6, 102084.1, 102122, 102145.2, 
    102162.2, 102167.8, 102163.6, 102156, 102143, 102129.3, 102109.1, 102081.6,
  100453.6, 101504.4, 101916.7, 101992.1, 102052.6, 102102.4, 102138.9, 
    102167.5, 102185.6, 102195.8, 102197.8, 102197, 102187.7, 102172.4, 
    102149.9,
  100102.9, 101410.8, 101855.5, 101951, 102017.8, 102076.2, 102119.9, 
    102154.2, 102182.2, 102203.1, 102216.5, 102219.6, 102217.7, 102211.8, 
    102198.6,
  100023.9, 100733.5, 101645.1, 101889.4, 101958.4, 102026.1, 102077.7, 
    102124.6, 102158.7, 102189.3, 102213.3, 102228.8, 102237.8, 102241.9, 
    102235.9,
  99682.37, 99536.16, 100462.5, 101763.9, 101895.3, 101966, 102021.9, 102070, 
    102112.6, 102150.2, 102178.1, 102202.3, 102218.5, 102231.7, 102235.6,
  99547.26, 98936.38, 98949.48, 100719.7, 101820.2, 101889.2, 101951.3, 
    102005.2, 102049.4, 102090.6, 102122.1, 102151.8, 102173.2, 102191.4, 
    102202.9,
  99726.94, 99040.27, 99509.9, 100048.6, 101672.8, 101807.8, 101868.9, 
    101921.9, 101967.3, 102011.6, 102047.1, 102079.4, 102102, 102125.4, 
    102140.7,
  98477.45, 98373.73, 99687.46, 100051.1, 100726.9, 101712.7, 101794.6, 
    101839.9, 101882, 101919.8, 101949.9, 101979, 102003.4, 102025.5, 102044.7,
  98452.9, 97044.98, 96934.5, 98163.91, 99888.38, 100662.6, 101721.4, 
    101764.7, 101798.2, 101830.8, 101859.4, 101883.1, 101906.9, 101925.7, 
    101945.5,
  101738.6, 101870.4, 101937, 102002.3, 102056.3, 102101.3, 102141.4, 
    102173.1, 102204.3, 102222, 102234.9, 102275.9, 102306.7, 102329.1, 
    102357.9,
  100358.1, 101802.6, 101911.7, 101983.1, 102047, 102093.9, 102133.2, 102171, 
    102199.2, 102215.7, 102230.2, 102250.5, 102289.9, 102324.2, 102337.4,
  100425.8, 101463.7, 101876.8, 101947.2, 102014.6, 102070.5, 102118.1, 
    102158.8, 102192.5, 102217.6, 102237, 102244.3, 102261, 102282.8, 102303.2,
  100086.7, 101375.4, 101816, 101904.8, 101972.4, 102038.4, 102086.8, 
    102129.6, 102166.3, 102195.1, 102215, 102228.2, 102240, 102249.8, 102255.3,
  100009.7, 100706.8, 101610.7, 101850.8, 101914.1, 101984.1, 102044.7, 
    102092.2, 102130.4, 102163.7, 102187.7, 102206.3, 102217.4, 102224.6, 
    102231.3,
  99683.87, 99520.51, 100431.8, 101729.2, 101856.2, 101919.5, 101980.4, 
    102033.4, 102076, 102110.6, 102137.1, 102159.6, 102175.4, 102189, 102199,
  99552.57, 98931.44, 98933.89, 100691.4, 101790.2, 101855.4, 101911.5, 
    101965.4, 102004.9, 102046, 102072.6, 102095.7, 102112.1, 102130.1, 
    102142.2,
  99736.09, 99041.87, 99502.04, 100028.2, 101644.2, 101780.2, 101834.2, 
    101886.3, 101925.6, 101962.1, 101988.4, 102016.3, 102036.1, 102052.3, 
    102065.2,
  98497.88, 98381.93, 99688.11, 100049, 100711, 101689.4, 101767.7, 101806.2, 
    101843.7, 101875.6, 101903.7, 101925.9, 101945.7, 101962.8, 101975,
  98481.69, 97062.7, 96950.84, 98169.44, 99879.38, 100644.1, 101696.4, 
    101730.7, 101759.1, 101786.1, 101810.5, 101830.4, 101848.6, 101862.4, 
    101868.8,
  101643.7, 101784.2, 101851.5, 101920.5, 101979.1, 102026.6, 102074.7, 
    102110.8, 102146.8, 102173.2, 102199.3, 102233.9, 102262.8, 102278.6, 
    102292.1,
  100279.3, 101720.1, 101832.1, 101904.9, 101967.9, 102012.1, 102057.9, 
    102099.8, 102134, 102169.6, 102190.4, 102230.9, 102259.4, 102291.2, 
    102297.3,
  100345.9, 101383.1, 101794.2, 101864, 101930.9, 101980.4, 102021.3, 
    102058.3, 102089.9, 102128, 102160.5, 102201.5, 102233.5, 102266.2, 
    102285.5,
  100012, 101301.4, 101741.6, 101825.1, 101884.3, 101944.2, 101985.8, 
    102020.7, 102049, 102078.2, 102107.7, 102135.7, 102170.7, 102198, 102232.6,
  99935.82, 100629.9, 101539.9, 101774, 101834.5, 101886.8, 101932, 101964.2, 
    101991, 102014.3, 102036.3, 102059.3, 102079.3, 102104.3, 102134.3,
  99606.07, 99449.63, 100369.4, 101658.7, 101780.5, 101832.6, 101873.5, 
    101901.8, 101922.8, 101939.3, 101952.1, 101963, 101974.8, 101994.1, 
    102025.7,
  99475.03, 98862.66, 98863.3, 100630.7, 101718.2, 101776.9, 101812.6, 
    101836.5, 101847.4, 101858, 101860.6, 101859, 101856.5, 101863, 101886.3,
  99673.49, 98973.48, 99427.09, 99959.5, 101576.8, 101709.5, 101744.7, 
    101766.8, 101772.2, 101774.1, 101767.6, 101758, 101744.1, 101739.8, 
    101751.4,
  98444.98, 98312.92, 99616.81, 99979.3, 100637.9, 101615.6, 101683.1, 
    101694.7, 101698.3, 101694.3, 101682.8, 101667.6, 101647.6, 101632.1, 
    101629.7,
  98437.47, 97008.69, 96885.38, 98089.1, 99808.04, 100585.9, 101616.1, 
    101630.1, 101614.8, 101607.3, 101596.1, 101581.3, 101569.5, 101557.7, 
    101555.4,
  101462.6, 101592.5, 101655.9, 101721, 101773.3, 101825.1, 101875.7, 
    101931.8, 101991.4, 102055.3, 102118.5, 102178.1, 102233.9, 102282.9, 
    102328.2,
  100101.8, 101538.2, 101633.5, 101689, 101738.2, 101787.3, 101834.6, 
    101887.8, 101945.1, 102010, 102075, 102139.5, 102202, 102261.8, 102316.6,
  100177.3, 101206.8, 101606.5, 101659, 101700, 101743.3, 101783.6, 101832.9, 
    101887.9, 101950.3, 102016.1, 102084.1, 102150.9, 102215.9, 102275.9,
  99855.16, 101132.7, 101556.4, 101622.5, 101659.9, 101698.3, 101734.5, 
    101775.1, 101822.6, 101880.1, 101944.3, 102013.1, 102084.4, 102153.9, 
    102220.2,
  99787.01, 100474.5, 101363.8, 101582.8, 101620.2, 101651.4, 101683.6, 
    101717, 101757.9, 101808.8, 101865.6, 101932.6, 102005.6, 102080.6, 
    102153.4,
  99468.77, 99302.73, 100201.8, 101469.7, 101573.5, 101604.1, 101633.5, 
    101664.6, 101693.6, 101736, 101786.2, 101848.8, 101920.4, 101999, 102077.4,
  99338.35, 98724.23, 98714.21, 100449.6, 101516.4, 101555.5, 101580, 
    101608.5, 101635.4, 101667.7, 101710.9, 101767.6, 101834.7, 101912.1, 
    101989.4,
  99530, 98838.24, 99281.68, 99791.48, 101378.9, 101493.1, 101525, 101552.3, 
    101579.8, 101608.8, 101639.8, 101691.4, 101751.1, 101823.4, 101898.5,
  98298.08, 98187.44, 99477.16, 99818.53, 100451.1, 101408.1, 101467.5, 
    101485.6, 101514.7, 101543.1, 101574.9, 101619.7, 101673.1, 101740.3, 
    101804.5,
  98281.32, 96873.06, 96760.61, 97966.15, 99646.37, 100397.5, 101411.8, 
    101437, 101440.1, 101467.9, 101493.7, 101532.8, 101582.6, 101640.4, 
    101702.7,
  101254.4, 101363.2, 101427, 101487.3, 101556.9, 101611.9, 101669, 101727.7, 
    101784.6, 101846.1, 101907.2, 101968.5, 102024.9, 102083.8, 102139,
  99888.37, 101313.8, 101422.8, 101477.2, 101545.6, 101601.2, 101659.3, 
    101713.7, 101770.9, 101834.1, 101898.8, 101960.7, 102020.3, 102080.1, 
    102132.1,
  99983.21, 100981.4, 101393.5, 101449.9, 101511.4, 101573.9, 101632.4, 
    101688.4, 101745, 101803, 101867.1, 101930, 101989.1, 102050.8, 102111.1,
  99654.22, 100911.7, 101348.1, 101422.1, 101478.5, 101536.4, 101595.1, 
    101646.2, 101703.6, 101760.2, 101821.9, 101884.9, 101946.6, 102009.7, 
    102069,
  99594.58, 100257.1, 101151.5, 101375.7, 101432.5, 101487.5, 101544, 
    101595.9, 101648.7, 101704.1, 101758.9, 101818.3, 101879.9, 101943.7, 
    102006.1,
  99275.9, 99098.66, 99992.62, 101266.1, 101381.4, 101432.7, 101484.3, 
    101533.2, 101582, 101632.9, 101687, 101742.5, 101802, 101863.4, 101929.6,
  99145.7, 98530.84, 98505.62, 100246.7, 101314, 101369.6, 101415.7, 
    101458.7, 101502.9, 101546.8, 101593.4, 101644.9, 101701.8, 101765.3, 
    101832.8,
  99339.9, 98643.86, 99069.95, 99584.13, 101176.6, 101296.2, 101339.1, 
    101376.4, 101413.3, 101450.8, 101491.5, 101538.8, 101591.6, 101654.3, 
    101721.5,
  98122.58, 97988.51, 99256.91, 99601.66, 100242.7, 101196.9, 101260.8, 
    101280.3, 101311.9, 101344.7, 101377.7, 101423.9, 101470.5, 101529.8, 
    101591.8,
  98106.8, 96699.97, 96570.79, 97750.95, 99419.65, 100165, 101176.7, 
    101204.5, 101197.3, 101227.9, 101253.1, 101293.2, 101339.1, 101395, 
    101451.8,
  101246.9, 101353.6, 101407.6, 101457.8, 101491.5, 101518.2, 101534.3, 
    101544.6, 101566.5, 101590.3, 101605.3, 101624.5, 101633.6, 101643.1, 
    101664.5,
  99859.59, 101294.9, 101388.4, 101434.5, 101471.4, 101499.5, 101523.9, 
    101540.2, 101550.2, 101567.7, 101580.2, 101593.9, 101610.5, 101621.7, 
    101632.6,
  99933.52, 100948.3, 101350.4, 101394.8, 101428.4, 101452.6, 101471.9, 
    101489, 101501.4, 101518.9, 101531.3, 101543.5, 101551.8, 101558.3, 
    101573.3,
  99605.07, 100866.3, 101294.9, 101359, 101390.1, 101413.1, 101430.4, 
    101440.5, 101446, 101449, 101452, 101457, 101464.8, 101473.8, 101477.1,
  99531.23, 100202.3, 101087, 101305.1, 101339.2, 101352.8, 101364.5, 
    101365.1, 101367.1, 101368.2, 101370.4, 101374.7, 101379.6, 101378.9, 
    101374.5,
  99209.8, 99037.6, 99941.59, 101189.9, 101277.8, 101288.7, 101292.5, 
    101294.5, 101289.4, 101284.5, 101280.9, 101281.2, 101281.1, 101276.5, 
    101264.8,
  99062.88, 98447.85, 98425.87, 100170.6, 101200.4, 101226, 101222.7, 
    101220.3, 101210.2, 101201.4, 101194.2, 101191.2, 101186, 101178.1, 
    101156.4,
  99253.19, 98560.59, 98982.03, 99491.48, 101065, 101154.4, 101154, 101143.9, 
    101128.2, 101116.5, 101103.1, 101099.3, 101092, 101085.4, 101059.3,
  98024.45, 97897.18, 99163.62, 99500.08, 100121.7, 101061.5, 101087.6, 
    101065.9, 101049.8, 101034.7, 101017.1, 101011, 100998.5, 100992.7, 
    100968.4,
  98000.95, 96594.99, 96470.31, 97649.9, 99309.73, 100057.9, 101025.7, 
    101018.6, 100970.9, 100953.2, 100926.1, 100912.3, 100903, 100900.1, 
    100884.9,
  101543.5, 101628, 101673.1, 101690.8, 101704.8, 101708.9, 101712.9, 
    101711.4, 101720.2, 101724.9, 101729.1, 101731.5, 101737, 101736.8, 
    101730.1,
  100144, 101566.1, 101640.2, 101661.7, 101673.6, 101671.4, 101666.4, 
    101659.3, 101657.6, 101650.8, 101647.7, 101654.5, 101653.5, 101648.8, 
    101642.3,
  100193.2, 101211.6, 101594.4, 101623.9, 101638.9, 101643.2, 101639.8, 
    101634.2, 101628.3, 101622, 101614.9, 101607.9, 101596.7, 101582.4, 
    101565.1,
  99839.51, 101121.3, 101537.3, 101585.1, 101596.5, 101606.6, 101606.3, 
    101603.5, 101594.3, 101587.4, 101579.3, 101565.7, 101548.8, 101527.1, 
    101498,
  99743.79, 100431.9, 101310, 101519.2, 101542.4, 101551.6, 101559.1, 
    101555.3, 101553.8, 101545.5, 101532.6, 101517.9, 101495.8, 101470.7, 
    101430.5,
  99401.91, 99244.78, 100143.8, 101388.4, 101474.1, 101482.4, 101493.5, 
    101495.8, 101493.9, 101488.2, 101478.6, 101462.4, 101438.9, 101412, 101371,
  99238.93, 98628.6, 98603.34, 100352.9, 101391.5, 101423, 101428.8, 
    101432.9, 101428.3, 101425.3, 101411.6, 101396.4, 101374.9, 101347.6, 
    101314.1,
  99412.91, 98726.86, 99151.23, 99667.84, 101253.4, 101353.1, 101360.5, 
    101363.3, 101356.7, 101351.4, 101338.1, 101323.5, 101303.7, 101283.5, 
    101252.5,
  98160.27, 98047.53, 99326.9, 99673.78, 100304.7, 101255.2, 101298.4, 
    101291.2, 101285.5, 101276.1, 101258.6, 101241, 101218, 101195.6, 101177,
  98119.99, 96731.16, 96617.45, 97815.2, 99493.2, 100258.9, 101239.9, 
    101244.1, 101212.1, 101198.1, 101175.5, 101154.8, 101136.2, 101117.9, 
    101114.2,
  101472.1, 101612, 101674.1, 101738.2, 101804.6, 101869.3, 101943, 102004.1, 
    102070.9, 102130.7, 102186.1, 102234.2, 102281.6, 102320.1, 102358.7,
  100096, 101535.5, 101628, 101688.7, 101746.6, 101800.1, 101863.6, 101923.9, 
    101983.8, 102039.3, 102091.5, 102136.6, 102177.8, 102215.4, 102252.1,
  100151.8, 101192.5, 101594.5, 101652.9, 101702.8, 101754.4, 101800.1, 
    101847.6, 101895.8, 101944.9, 101989.2, 102030.2, 102067.4, 102101, 
    102133.4,
  99806.24, 101098.5, 101534.8, 101609.6, 101652.9, 101700.8, 101743.4, 
    101781.8, 101820, 101857.9, 101893.8, 101926.9, 101957.9, 101986.4, 102013,
  99726.72, 100423.6, 101331.4, 101559.7, 101608.9, 101647, 101685.7, 
    101712.9, 101741.8, 101769, 101794.8, 101821.7, 101847.4, 101872.4, 
    101895.8,
  99377.52, 99234.81, 100160.6, 101440.3, 101555.3, 101592.9, 101625, 
    101648.9, 101669.7, 101690.2, 101706.2, 101725.5, 101743.9, 101764.2, 
    101783.8,
  99225.53, 98636.62, 98643.32, 100415, 101484.6, 101540.4, 101565.5, 
    101585.4, 101596.2, 101609.7, 101618.2, 101628.3, 101638.6, 101652.5, 
    101666.4,
  99386.31, 98738.91, 99191.33, 99739.16, 101344.9, 101468.7, 101498.5, 
    101514.3, 101521, 101525.1, 101523.4, 101524.9, 101524.8, 101529.2, 
    101532.3,
  98127.57, 98051.56, 99370.57, 99748.93, 100405.9, 101378.1, 101438.7, 
    101445.5, 101446.2, 101442.3, 101432.9, 101425.9, 101415.2, 101407.9, 
    101403.4,
  98072.86, 96716.12, 96632.54, 97861.53, 99584.23, 100367.6, 101380.1, 
    101399.5, 101374.6, 101366.1, 101345, 101326.7, 101305.4, 101286.8, 
    101268.2,
  101239, 101398.7, 101488.6, 101581.7, 101662.6, 101739.5, 101817.3, 
    101894.7, 101970.5, 102047.4, 102122.7, 102197.3, 102269.1, 102339, 
    102409.1,
  99871.35, 101324, 101447.6, 101531.3, 101620.3, 101698.6, 101773.5, 
    101849.5, 101922.2, 101993.5, 102062.3, 102132.5, 102201.2, 102273.9, 
    102344.2,
  99928.53, 100976.4, 101413.1, 101496.9, 101578.4, 101657.2, 101730.2, 
    101801.5, 101870, 101938.5, 102003, 102069.1, 102134.2, 102198.8, 102264.1,
  99591.97, 100884.2, 101347.5, 101446.1, 101524.3, 101603.2, 101680.8, 
    101745.9, 101810.8, 101870.4, 101929.3, 101987.1, 102046.6, 102109.3, 
    102172.5,
  99523.78, 100218.4, 101139.7, 101398.6, 101477.6, 101550.6, 101623.8, 
    101688.8, 101749.1, 101804, 101854.8, 101903.9, 101954.4, 102007.8, 
    102066.1,
  99187.31, 99046.87, 99964.64, 101265.5, 101415.2, 101491.9, 101562.7, 
    101625.3, 101680.4, 101730.2, 101775.3, 101817.9, 101860.3, 101905.1, 
    101954.1,
  99050.5, 98466.25, 98491.22, 100240.6, 101348, 101428.5, 101500.3, 101559, 
    101610, 101655.2, 101690.5, 101726, 101757.9, 101794.3, 101836,
  99221.59, 98564.92, 99041.22, 99585.45, 101199.6, 101360.7, 101431.6, 
    101493.4, 101538, 101578.3, 101606, 101631.3, 101652.5, 101678.8, 101709.6,
  97990.95, 97898.55, 99207.43, 99611.23, 100276, 101266.9, 101367.7, 
    101423.1, 101470.8, 101504, 101524.4, 101537.5, 101545.9, 101557.8, 
    101573.4,
  97962.3, 96598.29, 96492.84, 97699.42, 99446.93, 100245.2, 101311.4, 
    101359.6, 101398.5, 101427.4, 101443.9, 101445.5, 101441.6, 101436.7, 
    101433.5,
  101237, 101367.6, 101459.5, 101548.4, 101629, 101703.5, 101774.8, 101847.3, 
    101920, 101998.2, 102072.3, 102148.5, 102223.5, 102303.4, 102380.8,
  99855.6, 101300, 101438.3, 101515, 101597.2, 101667.7, 101736.9, 101805.9, 
    101875.1, 101953.3, 102030.6, 102111.3, 102188.4, 102272.4, 102354,
  99931.37, 100959.6, 101397.5, 101481.4, 101558.2, 101634.9, 101703.2, 
    101772.2, 101840.8, 101917.2, 101995.8, 102074, 102153.5, 102243, 102321.6,
  99596.88, 100875.4, 101339.5, 101441.2, 101513.6, 101585.6, 101655.7, 
    101722, 101790.4, 101861.6, 101941, 102022.7, 102103.3, 102189.8, 102272.4,
  99528.62, 100218.4, 101136.6, 101395.8, 101472.3, 101539.9, 101606.6, 
    101671.6, 101736.4, 101805.2, 101880, 101962.1, 102043.5, 102132.8, 
    102219.1,
  99200.57, 99064.31, 99975.38, 101274.6, 101419.5, 101485.9, 101548.3, 
    101606.8, 101667.3, 101735.6, 101807, 101886.6, 101971.8, 102058.2, 
    102144.8,
  99062.44, 98489.62, 98505.81, 100258, 101361.9, 101435.5, 101491.7, 
    101545.6, 101597.5, 101658.2, 101723.2, 101803.2, 101886.7, 101977.4, 
    102064.4,
  99251.56, 98591.71, 99061.96, 99609.28, 101219.5, 101377.6, 101431.4, 
    101478.3, 101522.1, 101575.9, 101632.9, 101707.8, 101789.2, 101882, 
    101972.9,
  98046.15, 97927.52, 99224.88, 99626.02, 100302.4, 101300, 101386.7, 
    101420.2, 101455.8, 101495, 101542.2, 101608.4, 101687.1, 101775.2, 
    101868.4,
  98056.95, 96649.05, 96534.73, 97734.36, 99479.41, 100272.1, 101344.4, 
    101380.8, 101392.7, 101421.5, 101456.8, 101506.7, 101576.9, 101659.9, 
    101753,
  101386.5, 101495.9, 101557.9, 101623.8, 101700.4, 101771.6, 101846.9, 
    101910.1, 101975.6, 102048.6, 102119.4, 102189, 102249.2, 102311.4, 
    102360.8,
  99990.05, 101429.4, 101542.6, 101606, 101679.8, 101748.7, 101818.4, 
    101888.8, 101958.5, 102036.7, 102114.2, 102190.3, 102260.5, 102326.7, 
    102381.2,
  100081.7, 101094.2, 101504.1, 101567.4, 101631.6, 101714.9, 101790.5, 
    101859.7, 101933.2, 102011.3, 102092.1, 102172.6, 102246.7, 102320.9, 
    102386.4,
  99755.37, 101010.1, 101452.1, 101534.2, 101594.9, 101667.4, 101746.8, 
    101821.8, 101898.1, 101976.7, 102058.7, 102144.1, 102220.7, 102297.9, 
    102368.7,
  99693.75, 100361, 101253.8, 101487.4, 101553.9, 101620.2, 101704, 101779.6, 
    101853.9, 101935.7, 102018.6, 102106, 102188.2, 102267.8, 102344.8,
  99377.39, 99215.66, 100109.3, 101371.7, 101506.9, 101570.9, 101650.2, 
    101729.1, 101807.1, 101886.6, 101971.6, 102059.1, 102141.4, 102227.3, 
    102302.2,
  99244.62, 98645.8, 98633.68, 100364.3, 101447, 101522.5, 101596, 101675.2, 
    101751.2, 101830.4, 101912.5, 102002.2, 102087.1, 102176.5, 102258.2,
  99424.22, 98757.78, 99200.3, 99728.02, 101313.7, 101467.3, 101536.6, 
    101609.3, 101685.4, 101765, 101846.1, 101934.7, 102022.4, 102111.8, 
    102196.8,
  98206.47, 98095.1, 99371.14, 99746.09, 100409.4, 101399.2, 101498.2, 
    101552.7, 101625.4, 101695.7, 101773.5, 101857.6, 101948.5, 102038, 
    102129.3,
  98189.02, 96797.6, 96674.02, 97860.77, 99583.93, 100358.9, 101455.6, 
    101511.5, 101562.6, 101630.6, 101700.4, 101777.9, 101865.9, 101955.4, 
    102045.8,
  101569.2, 101686.5, 101759.7, 101825.8, 101886.6, 101949.9, 102002.7, 
    102064.5, 102109.6, 102177.2, 102219.1, 102259.7, 102298.2, 102333.1, 
    102361.7,
  100175.4, 101600.1, 101708.1, 101772.7, 101847.3, 101906.4, 101971.2, 
    102040.5, 102101.8, 102167.6, 102231.2, 102285.6, 102330.1, 102374.3, 
    102409.6,
  100204, 101236.4, 101646.8, 101724.9, 101790.6, 101877.4, 101945.2, 
    102016.3, 102079.6, 102153.3, 102213.3, 102273.5, 102324.7, 102375.6, 
    102419.6,
  99872.62, 101150.6, 101578.9, 101668.8, 101734.8, 101811.1, 101891.4, 
    101973.2, 102048.5, 102128.1, 102197.7, 102266, 102322.7, 102377.6, 
    102423.7,
  99798.54, 100476.3, 101368.5, 101613.3, 101688.4, 101765.6, 101851.3, 
    101922.4, 102002.7, 102082, 102160.7, 102231.7, 102293.8, 102354.2, 102405,
  99453.39, 99308.96, 100204.1, 101483.6, 101626.2, 101699.6, 101786.9, 
    101880.6, 101958.2, 102040, 102117.5, 102195, 102260.3, 102324.4, 102378.6,
  99315.55, 98725.09, 98728.21, 100469.9, 101563.9, 101647.8, 101725.2, 
    101815.3, 101895.2, 101987.4, 102061.1, 102143.5, 102211.9, 102278.5, 
    102338.7,
  99502.3, 98830.54, 99291.3, 99826.91, 101422.5, 101584.4, 101661, 101754.8, 
    101835.8, 101926.4, 102003.1, 102083.8, 102156.5, 102224.1, 102286.1,
  98278.46, 98166.67, 99439.69, 99836.3, 100499.2, 101505.8, 101618.3, 
    101687.2, 101773.3, 101859.8, 101939, 102018, 102092.9, 102164.5, 102227.4,
  98257.97, 96881.16, 96763.38, 97953.77, 99680.3, 100457.1, 101566.2, 
    101641.2, 101710.4, 101793.1, 101868.6, 101947, 102021.9, 102091.9, 
    102156.9,
  101344.3, 101486.3, 101580, 101680, 101770.6, 101859.6, 101935.5, 102014.7, 
    102090.6, 102163.3, 102230.9, 102293.9, 102349.5, 102401.7, 102443.7,
  99969.75, 101411.4, 101543.8, 101628.8, 101730.3, 101823.3, 101909.4, 
    101993.4, 102072.8, 102146.6, 102218.1, 102286.2, 102347.7, 102406.1, 
    102458.4,
  100021.1, 101052.9, 101491.4, 101580.9, 101678, 101780.2, 101869.6, 
    101950.7, 102032.9, 102109.8, 102180.6, 102251, 102317.4, 102382, 102441.6,
  99690.63, 100959.9, 101419.2, 101539, 101625, 101717.2, 101822.1, 101908.6, 
    101988.3, 102069.6, 102144, 102217.1, 102285.9, 102353.4, 102416.5,
  99613.86, 100290.6, 101210.5, 101466.4, 101567, 101659.7, 101761.1, 
    101860.1, 101938.4, 102016.3, 102086.3, 102158.8, 102228.2, 102298, 102364,
  99292.72, 99146.41, 100047.7, 101351.5, 101516.3, 101602.3, 101698.7, 
    101798, 101880.9, 101962.9, 102033.2, 102105, 102171.4, 102242.6, 102309.9,
  99174.99, 98575.67, 98585.56, 100335.2, 101441.4, 101549.8, 101638, 
    101737.1, 101819.7, 101901, 101963.8, 102033.6, 102093.9, 102163.9, 
    102233.2,
  99378.06, 98691.38, 99162.48, 99699.83, 101312.8, 101490.4, 101576.6, 
    101671.1, 101758.5, 101840.3, 101906.2, 101965.8, 102021, 102080.9, 
    102148.5,
  98162.84, 98039.34, 99318.98, 99722.62, 100391.2, 101410.2, 101532.3, 
    101610, 101694.8, 101775.8, 101841.6, 101892.3, 101942.8, 101990.5, 
    102053.7,
  98154.13, 96756.97, 96639.62, 97846.05, 99572.97, 100356.8, 101474.2, 
    101557.8, 101637.5, 101713.4, 101783.6, 101834, 101870.9, 101909.1, 101957,
  101285.3, 101444.3, 101546.8, 101649.6, 101735.7, 101805.1, 101871.1, 
    101938.1, 102001.4, 102067.2, 102134.8, 102204.6, 102275.6, 102348.2, 
    102422.4,
  99906, 101358.2, 101495.4, 101589, 101682.6, 101764, 101825.5, 101884.6, 
    101941.1, 102008, 102075.1, 102147, 102224.2, 102302.2, 102384.3,
  99964.64, 100995.6, 101437.9, 101542.4, 101629.3, 101715.9, 101781.5, 
    101840.2, 101896.3, 101954.7, 102021.7, 102091.7, 102167.8, 102247.7, 
    102344.9,
  99618.12, 100895.3, 101363.3, 101482.4, 101578, 101659.4, 101740.4, 
    101795.7, 101848.7, 101899.6, 101962.1, 102031.4, 102116.4, 102194.2, 
    102306.1,
  99552.45, 100225.4, 101146.3, 101410.7, 101521.1, 101607, 101693.3, 
    101754.9, 101806, 101857.3, 101914.7, 101982.8, 102058.2, 102146.2, 
    102247.8,
  99226.52, 99082.16, 99985.91, 101293.8, 101454.7, 101551.5, 101637.8, 
    101713.1, 101765.2, 101815.1, 101865.5, 101930.8, 102004.9, 102096, 
    102189.5,
  99108.05, 98515.28, 98524.83, 100271.6, 101382.1, 101494, 101585.6, 
    101668.8, 101728, 101779, 101828.3, 101882.3, 101957.2, 102042.4, 102141.1,
  99307.61, 98629.54, 99099.09, 99640.55, 101251.8, 101432.7, 101525, 
    101616.6, 101686, 101740.6, 101790.4, 101843.7, 101909.5, 101985.6, 
    102087.3,
  98108.02, 97983.05, 99261.31, 99666.23, 100335.8, 101353.1, 101486.3, 
    101562, 101641.5, 101701.8, 101750.8, 101802.2, 101866.4, 101952.3, 
    102031.1,
  98121.07, 96721.96, 96599.94, 97794.27, 99530.41, 100314.4, 101432.1, 
    101519.4, 101593.5, 101661.3, 101714.4, 101770.7, 101829.2, 101909.6, 
    101991.9,
  101299.5, 101453.4, 101544, 101622, 101688.9, 101740.2, 101794, 101854.5, 
    101927.2, 101998.4, 102061.7, 102120.1, 102183.7, 102235.6, 102288.7,
  99932.4, 101374.3, 101496.2, 101569.1, 101639.3, 101701.3, 101754.4, 
    101810, 101883.2, 101960.3, 102035.9, 102108.4, 102178.3, 102244.5, 102313,
  99986.2, 101022.1, 101451.6, 101529.4, 101595, 101653.3, 101698.5, 
    101757.8, 101831.5, 101931.2, 102012.9, 102083.9, 102168.6, 102242.9, 
    102317.9,
  99649.62, 100924.2, 101382, 101481, 101547, 101607, 101655.4, 101707.2, 
    101772.2, 101871, 101964, 102045.6, 102128.4, 102217.1, 102304.3,
  99574.85, 100261.6, 101170, 101423.8, 101499.2, 101560.2, 101615.8, 
    101659.1, 101719.8, 101809.5, 101924.5, 102012.4, 102103.4, 102187.7, 
    102278.7,
  99256.17, 99100.77, 100012.5, 101298.5, 101446.8, 101515.1, 101577, 
    101623.4, 101677.8, 101754.8, 101861.3, 101957.3, 102053.7, 102140.4, 
    102235.4,
  99128.51, 98530.27, 98537.27, 100280.6, 101379.1, 101465.3, 101534.6, 
    101595.4, 101642.7, 101707.1, 101797.5, 101891.6, 101987.1, 102088.1, 
    102170.2,
  99328.66, 98648.2, 99106.84, 99634.73, 101239.9, 101408.9, 101485.7, 
    101559.5, 101615.2, 101675.9, 101740.9, 101840, 101908.6, 102013.4, 
    102094.6,
  98131.07, 97991.02, 99266.77, 99670.25, 100317, 101326.7, 101445.5, 
    101517.5, 101585.9, 101649.1, 101698.9, 101779.5, 101846.2, 101945.8, 
    102019.7,
  98162.12, 96734.76, 96592.84, 97767.91, 99503.84, 100285.1, 101402.9, 
    101484.5, 101554.1, 101620.9, 101668.9, 101737.8, 101803.9, 101870, 
    101960.5,
  101313.5, 101425.8, 101493.4, 101552.9, 101597.7, 101628.4, 101669, 
    101736.5, 101815.8, 101867.1, 101933.8, 102001.1, 102089.7, 102149.7, 
    102207.5,
  99928.02, 101331.6, 101418.9, 101483.9, 101543.9, 101600.3, 101656.6, 
    101722.3, 101792.4, 101842.9, 101905.3, 101967.5, 102048.7, 102115.8, 
    102183.4,
  99975.92, 100974.7, 101377.1, 101440.5, 101510.7, 101573.1, 101633.2, 
    101699.9, 101765.8, 101811.4, 101870.9, 101907.9, 102000.6, 102071.8, 
    102131.9,
  99624.46, 100871.8, 101297.7, 101373.6, 101455.7, 101524.5, 101605, 
    101674.4, 101747.4, 101798.8, 101857.1, 101895.4, 101970.5, 102041.2, 
    102106,
  99550.81, 100211.1, 101091.8, 101322.3, 101403, 101475, 101565.8, 101638.4, 
    101715.5, 101777.9, 101836.3, 101877.5, 101943.5, 102009.3, 102076.9,
  99229.14, 99050.1, 99935.76, 101200.2, 101346.9, 101421.4, 101516.3, 
    101601.6, 101686.5, 101757.9, 101817.8, 101871.4, 101928.8, 101997.9, 
    102058.1,
  99103.24, 98488.3, 98469.53, 100182, 101279.9, 101370, 101459.7, 101552.1, 
    101640.6, 101725.5, 101793.1, 101848.3, 101910.6, 101969.1, 102038.9,
  99312.44, 98606.12, 99045.92, 99551.37, 101144.9, 101316, 101408, 101498.6, 
    101592.1, 101682.3, 101757.4, 101827.8, 101881.3, 101949.9, 102016.9,
  98120.48, 97969.94, 99228.25, 99586.51, 100229.2, 101220, 101365.7, 
    101441.9, 101533.6, 101635, 101711.7, 101790.5, 101858.9, 101918.4, 
    101980.6,
  98135.73, 96712.68, 96561.03, 97704.29, 99436.77, 100195.7, 101318, 
    101399.1, 101480.9, 101577.7, 101665.3, 101748.4, 101817.9, 101885, 
    101946.8,
  100956.8, 101040.7, 101107.6, 101189.8, 101268, 101357.6, 101448.3, 
    101540.6, 101631.4, 101702.2, 101768.4, 101828.5, 101910.9, 101970.4, 
    102014,
  99574.62, 100978.6, 101075.2, 101153.8, 101240, 101339.3, 101423.6, 
    101517.8, 101603.6, 101675.3, 101756.8, 101826.8, 101892.3, 101948.8, 
    101995.8,
  99649.95, 100643.1, 101046.9, 101121.2, 101206.8, 101302.7, 101399.2, 
    101493.1, 101582.1, 101661.4, 101733.3, 101804, 101870.5, 101930.4, 
    101989.2,
  99328.45, 100564.8, 100998, 101079.6, 101177.9, 101261.2, 101367.5, 
    101466.6, 101552.1, 101632.9, 101714, 101783.6, 101854.8, 101911, 101978.4,
  99268.05, 99922.52, 100805.1, 101049.8, 101132.3, 101229.9, 101335.6, 
    101434.1, 101523.4, 101607.6, 101680.2, 101757.4, 101821.8, 101888.8, 
    101953,
  98978.04, 98795.01, 99661.5, 100936.6, 101091.5, 101189.2, 101294, 
    101401.9, 101493.2, 101579.4, 101653.5, 101730, 101789.8, 101860.4, 
    101925.8,
  98870.12, 98245.65, 98227.48, 99933.5, 101033.8, 101147.5, 101252.3, 
    101366.4, 101458.8, 101548.4, 101623.4, 101698.7, 101762, 101822.5, 
    101893.7,
  99082.59, 98372.27, 98801.38, 99307.3, 100903.7, 101094.6, 101210.1, 
    101320, 101424.7, 101520.8, 101595.3, 101667, 101735.2, 101790.7, 101855.9,
  97891.61, 97748.84, 99000.07, 99342.55, 99992.72, 101001.4, 101173.5, 
    101271.5, 101386.5, 101482.5, 101564.2, 101637.9, 101702.9, 101761.5, 
    101818.1,
  97896.37, 96487.7, 96334.57, 97481.78, 99206.71, 99970.41, 101130.1, 
    101233.1, 101338, 101445.2, 101531.8, 101606.2, 101670.7, 101735.3, 
    101788.4,
  100566.9, 100631.5, 100697.7, 100768.3, 100852.3, 100941.4, 101034.5, 
    101136.4, 101235, 101332, 101425.3, 101505.1, 101582.3, 101661, 101736.9,
  99207.01, 100584.4, 100706.6, 100779.3, 100873.5, 100971.8, 101065.3, 
    101162.1, 101255.9, 101348.9, 101444.6, 101531.8, 101613, 101695.2, 
    101771.5,
  99329, 100288.3, 100689.7, 100770.8, 100860.7, 100957.8, 101060.8, 
    101164.4, 101264.4, 101360.7, 101456.4, 101546, 101627.9, 101715.2, 
    101799.7,
  99023.66, 100239, 100658.9, 100759.2, 100857.8, 100956.4, 101063.8, 
    101171.4, 101269.5, 101365.9, 101460.2, 101548.7, 101636.2, 101721.4, 
    101807.1,
  98994.23, 99625.77, 100492.9, 100737.2, 100833.1, 100939.5, 101047, 
    101158.3, 101263.1, 101361.3, 101455, 101544.8, 101630, 101715.9, 101805.8,
  98710.99, 98531.29, 99378.61, 100650.2, 100807.7, 100914.7, 101031.7, 
    101144.4, 101250.2, 101350.8, 101441.4, 101529.9, 101618.9, 101705.6, 
    101797.1,
  98620.41, 97995.77, 97973.96, 99672.99, 100765.4, 100882.7, 101000.7, 
    101116.8, 101226.5, 101330.9, 101420.1, 101510.6, 101596.6, 101685, 
    101779.3,
  98849.97, 98129.29, 98565.33, 99073.64, 100653.8, 100842.6, 100972.2, 
    101084.1, 101199.4, 101306.4, 101396.6, 101485.6, 101571.5, 101662.1, 
    101753.2,
  97684.08, 97530.66, 98772.38, 99136.3, 99787.54, 100768.2, 100944.7, 
    101053.3, 101166.8, 101276.7, 101368.3, 101457, 101541.4, 101629.6, 
    101719.1,
  97717.88, 96312.39, 96167.19, 97305.62, 99002.52, 99760.98, 100907.8, 
    101034.2, 101128.5, 101246.8, 101337.6, 101426.5, 101508.3, 101597.4, 
    101678.2,
  100797.8, 100782.9, 100768.9, 100777.2, 100807.6, 100833.8, 100855.7, 
    100888.7, 100926.9, 100977, 101027.4, 101088.4, 101151.7, 101225.5, 101302,
  99367.98, 100719.8, 100740.4, 100766.9, 100801, 100850, 100895.8, 100950, 
    101000.5, 101060.4, 101123.5, 101194.7, 101264, 101341.4, 101414.1,
  99452.51, 100387.2, 100737.8, 100775.2, 100810.6, 100870.6, 100929.2, 
    100996.1, 101054.5, 101120.8, 101182, 101252.7, 101321.9, 101400.2, 
    101474.5,
  99120.32, 100302.2, 100691.1, 100753.2, 100803.5, 100875.3, 100947.5, 
    101023.4, 101096.4, 101171.6, 101241.5, 101318.7, 101392.9, 101470.4, 
    101546.1,
  99066.86, 99679.5, 100511, 100732.3, 100795.1, 100872.9, 100954.4, 
    101039.5, 101117.5, 101207.2, 101281.6, 101361.9, 101436.4, 101515.2, 
    101592.7,
  98780.36, 98560.77, 99396.77, 100645.9, 100779.7, 100858.1, 100955, 
    101047.2, 101131.8, 101230.2, 101313, 101397.5, 101477.5, 101557.4, 
    101638.7,
  98682.38, 98011.48, 97970.04, 99670.29, 100740.5, 100831.3, 100934.6, 
    101039.3, 101133, 101238.3, 101325.3, 101410.5, 101496.1, 101575.2, 
    101659.7,
  98916.91, 98157.3, 98560.7, 99057.58, 100625.7, 100782.1, 100887.9, 
    101007.8, 101107.4, 101224.3, 101316.6, 101411.6, 101498.4, 101582.2, 
    101664.6,
  97748.88, 97574.31, 98778.08, 99113.21, 99731.79, 100698.1, 100852.7, 
    100979.1, 101078.2, 101198.2, 101298.8, 101394, 101483.8, 101570.8, 
    101656.4,
  97782.58, 96380.23, 96194.2, 97305.51, 98980.15, 99715.07, 100811.8, 
    100956.6, 101047.4, 101169.4, 101270.6, 101371.3, 101462.7, 101553.5, 
    101642.5,
  101427.5, 101442.4, 101435.7, 101426.5, 101423.8, 101425.7, 101422.8, 
    101416.7, 101397.4, 101381.1, 101367.8, 101377.4, 101403.8, 101432.6, 
    101425.8,
  99989.88, 101347.1, 101375.7, 101369.4, 101362.3, 101360.1, 101358.6, 
    101354.9, 101348, 101348.5, 101348, 101353.8, 101365.8, 101415.5, 101456.6,
  100012, 100980.2, 101309.3, 101291, 101300.7, 101312.3, 101327.7, 101344.5, 
    101350.2, 101353.9, 101355.2, 101357.3, 101412.5, 101504.3, 101567.6,
  99616.88, 100837.9, 101196.1, 101233.5, 101253.6, 101292.5, 101316.8, 
    101337.6, 101353.4, 101368.3, 101391.4, 101420.8, 101501.8, 101575.2, 
    101632.7,
  99488.84, 100134.6, 100973.2, 101180.8, 101209.4, 101250.1, 101294.7, 
    101349.4, 101375.8, 101409.2, 101444.6, 101496.3, 101576.2, 101660.2, 
    101743.9,
  99121.03, 98941.34, 99821.14, 101029.9, 101148.5, 101215.6, 101279.1, 
    101336.9, 101381.9, 101433.5, 101478.7, 101529.9, 101611.2, 101673.9, 
    101753,
  98958.23, 98329.74, 98296.35, 100001.3, 101048.9, 101128.2, 101216.6, 
    101294.7, 101361.5, 101427.5, 101484, 101538.8, 101609.2, 101681.8, 
    101760.1,
  99131.88, 98409.19, 98810.67, 99307.59, 100891.1, 101045.7, 101156.4, 
    101248.8, 101331.6, 101418.4, 101485.5, 101552, 101622.2, 101696.5, 
    101771.1,
  97928.8, 97780.97, 98993.53, 99320.31, 99931.92, 100920.7, 101090.6, 
    101195.9, 101293.4, 101389.9, 101471.4, 101547.8, 101622.2, 101698.8, 
    101776.5,
  97904.06, 96491.38, 96346.55, 97484.83, 99165.43, 99896.53, 101017.8, 
    101154.4, 101251.1, 101357.9, 101448.4, 101532.6, 101615.4, 101693.4, 
    101769.7,
  101333.5, 101412.6, 101450.4, 101487.8, 101525.9, 101554.1, 101583.4, 
    101595.7, 101595, 101548.5, 101489, 101410.4, 101440.1, 101566.4, 101745.3,
  99897.56, 101298.6, 101367.4, 101406.3, 101449.1, 101488.1, 101523.2, 
    101539.5, 101529.2, 101493.6, 101433.6, 101354.7, 101364.4, 101508.8, 
    101676,
  99909.1, 100903.6, 101282.2, 101323.2, 101369.1, 101416.3, 101456.5, 
    101505.1, 101529.8, 101528, 101492.1, 101454.6, 101483.2, 101578.1, 
    101686.4,
  99528.41, 100778.1, 101181.1, 101255.4, 101304, 101353.3, 101400.8, 
    101446.8, 101474.2, 101510.4, 101525.1, 101521.6, 101562.8, 101630, 
    101704.7,
  99410.61, 100085, 100966.4, 101198.3, 101262.5, 101318.2, 101376.4, 
    101430.4, 101479.4, 101517.4, 101557.1, 101590.2, 101632, 101678.8, 
    101753.3,
  99065.95, 98895.98, 99790.74, 101050.5, 101202, 101271.2, 101338.6, 
    101399.7, 101459.4, 101508.4, 101562.7, 101613, 101664, 101723.2, 101784.2,
  98900.51, 98291.24, 98288.54, 100020.6, 101108.1, 101206.5, 101290.4, 
    101363.1, 101433.1, 101489.4, 101551, 101611.8, 101680.5, 101728.9, 
    101788.2,
  99063.2, 98372.15, 98802.59, 99335.73, 100944, 101124.4, 101226.2, 
    101309.6, 101394.9, 101460.5, 101520.1, 101577.8, 101642, 101710.9, 101774,
  97849.95, 97717.8, 98973.09, 99324.22, 99988.68, 101018.2, 101175.8, 
    101252.7, 101347.6, 101426.2, 101491.6, 101557.3, 101620.1, 101684.6, 
    101749.3,
  97814.99, 96448.71, 96302.34, 97489.5, 99166.4, 99942.67, 101105.9, 
    101208.7, 101293.8, 101381.4, 101449.4, 101510.4, 101575, 101642, 101709.3,
  100761.5, 100852.5, 100907.3, 100954.3, 100996.7, 101036.8, 101068, 
    101099.1, 101130.4, 101152.6, 101163.1, 101158, 101144.9, 101129.4, 
    101117.6,
  99385, 100782.5, 100880.5, 100929.2, 100981.8, 101026.4, 101063.4, 
    101105.1, 101134.2, 101154, 101168.6, 101176.2, 101178.5, 101185.2, 
    101192.1,
  99452.49, 100447.3, 100846.6, 100911, 100969, 101022.3, 101071.2, 101113.4, 
    101156.9, 101182.9, 101203.1, 101223.5, 101241.8, 101256.5, 101274.1,
  99107.92, 100353.5, 100776.6, 100873.6, 100934.7, 101002.7, 101060.6, 
    101115.7, 101160.7, 101189.9, 101221.6, 101248.4, 101272.9, 101300.8, 
    101329.9,
  99030.96, 99691.48, 100574.9, 100823.3, 100902.3, 100976.6, 101047, 
    101106.4, 101164, 101202.7, 101242, 101274.4, 101312, 101340.6, 101377,
  98719.17, 98547.62, 99425.47, 100697.3, 100855.8, 100936.2, 101020.1, 
    101089, 101151.2, 101198.6, 101244.5, 101286.7, 101320, 101364, 101399.9,
  98602.54, 97988.98, 97981.18, 99695.04, 100790.5, 100893.2, 100986.7, 
    101064.4, 101136.6, 101192.6, 101238.9, 101282.3, 101328.6, 101374, 
    101417.2,
  98848.09, 98111.22, 98557.42, 99067.45, 100652.7, 100839.6, 100938.7, 
    101024.5, 101105.5, 101173.6, 101225.5, 101275.5, 101322.9, 101371.3, 
    101419.5,
  97690.44, 97507.22, 98768.23, 99125.37, 99762.76, 100764.7, 100914.5, 
    100988.1, 101074.6, 101148.6, 101207.6, 101259, 101314.7, 101362.1, 
    101413.9,
  97724.73, 96290.24, 96158.61, 97325.52, 98999.62, 99728.46, 100861.9, 
    100951.4, 101035.2, 101114.4, 101181.2, 101239.6, 101292.8, 101347.8, 
    101397.3,
  100628.6, 100603.1, 100571.4, 100528.4, 100496.1, 100463.9, 100433.6, 
    100403, 100386, 100368.8, 100359.6, 100348.6, 100339.3, 100341.2, 100358.5,
  99214.95, 100527, 100561, 100527.6, 100509.7, 100489.8, 100475.6, 100465.2, 
    100461.1, 100456, 100453.7, 100447, 100451.3, 100466.1, 100479.8,
  99265.35, 100205, 100537.6, 100515.5, 100507.4, 100498.1, 100496.2, 100500, 
    100507.4, 100515.9, 100522.4, 100529.8, 100539.7, 100553.6, 100567.4,
  98914.06, 100110.1, 100489.4, 100491.5, 100488.2, 100494.9, 100511, 
    100523.2, 100546.2, 100563.1, 100580.5, 100598.9, 100618.8, 100637.6, 
    100661.8,
  98836.27, 99466.98, 100291, 100462, 100477.5, 100482.6, 100507.4, 100532.8, 
    100563.2, 100588.6, 100616.3, 100646.6, 100677.2, 100709.1, 100743.8,
  98529.83, 98336.38, 99168.44, 100362, 100450.2, 100465.7, 100496.9, 
    100533.2, 100574.4, 100614.6, 100652, 100689.9, 100730.2, 100771.5, 
    100814.2,
  98418.12, 97788.84, 97731.59, 99390.98, 100416.5, 100445.3, 100476.4, 
    100529.6, 100576.8, 100628.9, 100672.7, 100718.6, 100767.5, 100815, 
    100867.3,
  98661.7, 97913.84, 98296.41, 98768.21, 100294.2, 100412.2, 100456.4, 
    100516.4, 100573.2, 100632, 100686.5, 100739.7, 100789.1, 100846.8, 
    100907.7,
  97510.04, 97317.98, 98527.79, 98832.96, 99408.15, 100329, 100424.7, 
    100491.6, 100553.4, 100623.5, 100684.3, 100749.6, 100805.6, 100869.9, 
    100929.9,
  97570.66, 96120.73, 95945.18, 97038.68, 98667.17, 99364.6, 100395.4, 
    100478.2, 100528.9, 100607.1, 100672.6, 100744.3, 100807.5, 100876.5, 
    100946.3,
  101706, 101685.4, 101623.4, 101542.8, 101460.8, 101377.4, 101286.6, 
    101199.5, 101110.4, 101016.9, 100925.9, 100838.7, 100753.1, 100671.1, 
    100596.6,
  100289, 101618.6, 101612, 101534.3, 101460, 101382.3, 101300, 101216.7, 
    101131.2, 101044.8, 100960.3, 100879.5, 100796.8, 100714.9, 100646.8,
  100344.3, 101296.5, 101591.9, 101524.4, 101455.9, 101382, 101308.4, 
    101232.5, 101157.7, 101080.5, 101004.4, 100924.2, 100851.4, 100782, 
    100718.8,
  99995.53, 101211.2, 101553, 101496.9, 101434.7, 101368.4, 101298.2, 
    101226.9, 101156.4, 101079, 101005.2, 100932.4, 100861.9, 100791.7, 
    100720.5,
  99908.48, 100537.6, 101333.6, 101472.3, 101409.8, 101339.2, 101274.9, 
    101207.7, 101139.7, 101068.8, 100997.9, 100925.2, 100849.2, 100784.5, 
    100719,
  99541.19, 99343.76, 100174.3, 101362.7, 101378.8, 101314.8, 101245.5, 
    101178, 101110.8, 101037.6, 100962.4, 100892.2, 100826.6, 100760, 100696.4,
  99366.14, 98720.73, 98646.03, 100349.2, 101329.1, 101270.3, 101205.9, 
    101135.9, 101068.8, 100996.8, 100931.7, 100865.3, 100795.3, 100740.7, 
    100693.5,
  99514.36, 98794.23, 99183.65, 99688.52, 101212.5, 101242.3, 101169, 
    101100.9, 101030, 100954.5, 100886.4, 100821.8, 100766.6, 100716, 100673.8,
  98245.91, 98114.35, 99371.1, 99699.02, 100272.9, 101142.1, 101123.8, 
    101053, 100979.5, 100913.9, 100839.9, 100775.5, 100734.6, 100693.1, 
    100670.8,
  98186.17, 96775.65, 96642.84, 97803.93, 99447.42, 100188.8, 101080.3, 
    101033.8, 100933.5, 100875.8, 100802.5, 100751.6, 100711.5, 100690, 
    100673.5,
  102223, 102286.5, 102277.2, 102263.9, 102232.7, 102196, 102151.8, 102116.4, 
    102096.9, 102060.3, 102013.2, 101953.3, 101883.7, 101808.8, 101734.3,
  100819.8, 102224.7, 102271, 102266.3, 102246.8, 102216.4, 102181.2, 
    102150.1, 102124.4, 102091.4, 102053.2, 101999, 101932.6, 101855.9, 101780,
  100883.5, 101892.9, 102248.4, 102258.8, 102250.4, 102236.4, 102203.4, 
    102171.8, 102150.4, 102118.6, 102083.9, 102035.6, 101976.3, 101904.4, 
    101829.1,
  100524.6, 101800.2, 102198.6, 102235.3, 102234.4, 102226.8, 102208.5, 
    102188, 102167.2, 102136.8, 102099.6, 102057.7, 102003.6, 101935.4, 
    101862.7,
  100443.4, 101124.7, 101993.3, 102193.5, 102206.6, 102202.6, 102194.8, 
    102183.5, 102168.6, 102140.8, 102108.2, 102066.8, 102017.9, 101956.7, 
    101889,
  100098, 99920.6, 100823.4, 102071.3, 102159.4, 102160, 102164.4, 102161.6, 
    102148.8, 102124.7, 102095, 102055.7, 102010.7, 101955.7, 101894.5,
  99945.66, 99302.34, 99282.66, 101043.7, 102092.1, 102126.1, 102127.2, 
    102123.5, 102114.2, 102096.3, 102072.5, 102039.6, 101998.4, 101952, 
    101897.2,
  100115.8, 99409.09, 99841.46, 100368.6, 101964.3, 102064.8, 102077.7, 
    102079.9, 102067.3, 102056, 102034.4, 102001.7, 101966.4, 101924.1, 
    101876.8,
  98844.68, 98733.01, 100021.2, 100367.5, 101015, 101977.9, 102032.3, 
    102028.7, 102025.8, 102015.7, 101992.9, 101968.6, 101938.3, 101903.4, 
    101861.3,
  98776.19, 97351.61, 97256.07, 98475.48, 100178.4, 100950.8, 101969.7, 
    101997.3, 101975.3, 101975.4, 101948.9, 101926.4, 101893, 101861.1, 
    101826.2,
  102165.7, 102257.9, 102296.6, 102328, 102351.2, 102380.7, 102413.7, 
    102450.6, 102478, 102510.7, 102511.9, 102506.5, 102504.5, 102499.2, 
    102482.2,
  100753.4, 102177, 102246.2, 102283, 102315.5, 102350.1, 102386.5, 102426.7, 
    102459.1, 102487.3, 102500.7, 102509.9, 102498.2, 102486, 102472.7,
  100805.7, 101830.9, 102213.2, 102251.4, 102283.2, 102319.3, 102351.5, 
    102396.5, 102430.9, 102469.4, 102490.2, 102499.8, 102500.1, 102489.1, 
    102474.7,
  100450.9, 101731.6, 102145, 102205.7, 102235.7, 102274.6, 102310.1, 
    102356.8, 102391.3, 102425, 102456.8, 102473, 102482.6, 102483.9, 102472.6,
  100375.6, 101059.4, 101942.3, 102159.7, 102194, 102225.2, 102261.2, 
    102300.4, 102338.5, 102374.4, 102406.8, 102432.6, 102448.2, 102455.1, 
    102459.5,
  100034.6, 99861.8, 100767.1, 102032, 102139.3, 102173.9, 102207.7, 
    102244.6, 102277.8, 102310.3, 102341.5, 102365.8, 102386, 102402.5, 
    102413.6,
  99891.63, 99253.58, 99243.03, 101003.5, 102071.3, 102120.8, 102149.6, 
    102181.7, 102216.5, 102249.2, 102275.7, 102299.5, 102322.6, 102342.5, 
    102357.9,
  100067.6, 99356.77, 99799.1, 100321.6, 101928.1, 102047.4, 102086.6, 
    102115.1, 102144.8, 102172.5, 102192.2, 102216.9, 102239.4, 102263.5, 
    102281.1,
  98806.04, 98690.21, 99982.8, 100324.2, 100976.6, 101947.6, 102015.3, 
    102041.3, 102067.4, 102091.5, 102108.4, 102133.1, 102154.6, 102180.3, 
    102199.8,
  98764.74, 97330.6, 97221.94, 98438.98, 100138.3, 100904.9, 101942.2, 
    101981.2, 101978, 102004.6, 102017.1, 102036.9, 102057.5, 102082.6, 102109,
  101920.3, 102024.6, 102076.9, 102143.1, 102196.6, 102257.1, 102313.2, 
    102365.2, 102410.3, 102456.7, 102503.1, 102544.1, 102581.8, 102631.6, 
    102691.1,
  100508.8, 101933.7, 102022.1, 102085.6, 102143.1, 102196.2, 102246.3, 
    102298.2, 102341.9, 102384.5, 102422, 102462.7, 102504.7, 102546.3, 
    102599.8,
  100561.5, 101578, 101967.9, 102024.1, 102077.5, 102132.7, 102181.5, 102231, 
    102276.1, 102321.2, 102360.6, 102396.4, 102430.1, 102465.1, 102510.8,
  100206.9, 101472.1, 101893.8, 101961.1, 102004.2, 102054.7, 102105, 
    102154.8, 102199.2, 102245, 102288, 102329.1, 102369.1, 102407.5, 102447,
  100133.9, 100801.7, 101683.1, 101897.3, 101942.7, 101984.1, 102027.7, 
    102074.4, 102118.1, 102163.6, 102208.5, 102251.3, 102292.8, 102333.9, 
    102379.1,
  99794.96, 99613.88, 100502.7, 101764.8, 101867.5, 101908.6, 101948.1, 
    101990.4, 102029.7, 102068.5, 102109.6, 102151.2, 102198.6, 102250.1, 
    102297.7,
  99658.85, 99017.77, 98990.46, 100734.5, 101791.6, 101837.1, 101865.6, 
    101896.4, 101930.9, 101964.8, 101999.1, 102037.3, 102074.4, 102109.2, 
    102156.7,
  99836.88, 99126.37, 99550.59, 100058.3, 101641.2, 101752.2, 101779, 
    101804.1, 101822.9, 101844.4, 101862.8, 101883.9, 101903.7, 101960.5, 
    102021.2,
  98585.36, 98459.8, 99735.76, 100065.1, 100703.1, 101655.6, 101705.1, 
    101708.4, 101714.2, 101725.1, 101730.4, 101735.4, 101768.9, 101814.8, 
    101871,
  98554.34, 97113.16, 96994.58, 98194.63, 99857.03, 100610.4, 101622.2, 
    101634.2, 101599.8, 101597.8, 101567.5, 101557.6, 101587.2, 101632.9, 
    101683.8,
  101614.8, 101709.8, 101759.7, 101807, 101851.1, 101895.9, 101939.8, 101980, 
    102016, 102051.5, 102094.3, 102141.8, 102211, 102278.5, 102347.6,
  100226.3, 101643, 101725.2, 101768.3, 101805.1, 101840.6, 101874.1, 
    101906.2, 101932.4, 101964.7, 101997.8, 102041.5, 102086.7, 102143.6, 
    102219.6,
  100298.4, 101303.9, 101683.5, 101720.2, 101752, 101781.4, 101804.8, 
    101825.4, 101839.8, 101856.5, 101879.1, 101915.6, 101957.7, 102017.1, 
    102100.7,
  99963.57, 101222.6, 101627.9, 101674.8, 101693.1, 101711.2, 101727.3, 
    101739.6, 101739.6, 101743.7, 101756.4, 101760.5, 101793.1, 101858.9, 
    101925,
  99909.15, 100568.9, 101428.6, 101628.7, 101644.9, 101650, 101653, 101649.8, 
    101634.2, 101618.5, 101604.2, 101588.4, 101627, 101668.5, 101715.7,
  99596.15, 99411.55, 100287.6, 101519, 101594.9, 101592.1, 101581, 101563.2, 
    101529, 101488.5, 101451.2, 101407.7, 101430.9, 101411.1, 101427.5,
  99483.37, 98839.57, 98787.7, 100517.7, 101540.9, 101542.1, 101516, 
    101476.2, 101423.9, 101358.3, 101289.9, 101227.6, 101179.4, 101134.8, 
    101138.4,
  99691.73, 98971.65, 99376.96, 99867.24, 101416.1, 101485, 101455.2, 
    101396.8, 101320.2, 101233.3, 101128.1, 101036, 100929.5, 100860.5, 
    100868.8,
  98470.81, 98329.78, 99586.92, 99893.59, 100501, 101408.3, 101403.4, 
    101323.7, 101233.2, 101121.8, 100987.2, 100831.6, 100671.9, 100589.8, 
    100615.7,
  98460.96, 97020.92, 96894.86, 98060.36, 99703.88, 100424.6, 101353.5, 
    101290.2, 101152.9, 101021.2, 100850.3, 100641.1, 100430.6, 100353, 
    100390.5,
  101479.1, 101505.5, 101497.9, 101486.7, 101479, 101467.3, 101460.8, 
    101441.7, 101418.5, 101385.2, 101344.3, 101289.7, 101230.5, 101165.5, 
    101127.4,
  100091.8, 101468.6, 101517.6, 101513.3, 101511.7, 101499.1, 101482.2, 
    101459, 101429.3, 101375.5, 101312.3, 101226.8, 101143.7, 101083.5, 
    100989.5,
  100198.5, 101186.4, 101539.2, 101536.5, 101530.7, 101522.4, 101498.8, 
    101467.1, 101421.1, 101347.8, 101262.8, 101152.6, 101065.9, 100947.1, 
    100849.1,
  99912.34, 101146.9, 101532.5, 101555.4, 101548, 101541.8, 101511.3, 
    101476.7, 101416.8, 101327.2, 101224.5, 101089.5, 100972.2, 100796.6, 
    100706.2,
  99897.53, 100539.2, 101376, 101568.1, 101566, 101554.2, 101523.4, 101477.3, 
    101409, 101306.2, 101188.1, 101042.1, 100875.3, 100678.1, 100590.4,
  99608.65, 99427.12, 100286.6, 101510.2, 101583, 101563.8, 101537, 101484.3, 
    101411.2, 101301.7, 101170.4, 101013.2, 100805.7, 100620.6, 100535.2,
  99526.66, 98899.05, 98835.01, 100549.3, 101584.8, 101578.4, 101547.3, 
    101490.1, 101415.4, 101309, 101175.2, 101014.6, 100804.3, 100631.2, 
    100538.1,
  99778.01, 99052.33, 99459.43, 99944.05, 101494.3, 101577.7, 101557.6, 
    101504.1, 101426, 101329.3, 101199.5, 101043, 100845.3, 100683.6, 100581.7,
  98578.48, 98424.62, 99705.67, 100015, 100619.2, 101539.7, 101563.7, 
    101511.2, 101442.2, 101356.6, 101237.6, 101097.2, 100917.2, 100774.6, 
    100671.1,
  98591.92, 97135.9, 97001.38, 98184.46, 99858.84, 100584.3, 101567.1, 
    101536.3, 101454.4, 101385.8, 101282.9, 101164.3, 101010.1, 100879, 
    100786.5,
  102071, 102049.3, 101989.6, 101904.5, 101857.2, 101811.7, 101757.6, 
    101705.8, 101649.8, 101598.2, 101546.3, 101495.2, 101438, 101381.5, 
    101325.4,
  100604.1, 101966.7, 101974.2, 101903.1, 101858.1, 101811, 101761.3, 
    101719.6, 101672.9, 101629.7, 101581, 101534.9, 101480.1, 101429.8, 
    101374.8,
  100629.4, 101621.4, 101954.9, 101898.3, 101862.7, 101820.9, 101776.7, 
    101734.1, 101688.1, 101647, 101604.5, 101561, 101516.9, 101470.8, 101422.9,
  100302.9, 101537.8, 101909.6, 101889.8, 101867.1, 101835.8, 101799.7, 
    101765.1, 101725.9, 101689.5, 101653, 101614.2, 101567.9, 101523.9, 
    101475.9,
  100244.9, 100876.7, 101726.2, 101889, 101876.3, 101854.2, 101825.9, 
    101795.9, 101768.4, 101735.5, 101701.7, 101666.8, 101623.6, 101579.4, 
    101538.3,
  99923.91, 99736.34, 100602.8, 101821.8, 101888.7, 101874.9, 101858, 101838, 
    101817.3, 101790.4, 101758.2, 101728.4, 101690.4, 101646.9, 101605.6,
  99806.34, 99192.12, 99132.93, 100850, 101889.6, 101908.4, 101891.9, 101879, 
    101858.6, 101838.1, 101813.7, 101787.8, 101755.3, 101715.5, 101673.1,
  100045.9, 99335.1, 99739.62, 100230.3, 101795.8, 101907.9, 101924.6, 
    101922, 101904.2, 101889.4, 101869.5, 101844, 101815.9, 101778.6, 101736.1,
  98837.95, 98697.66, 99971.16, 100294.2, 100915.3, 101874.2, 101942, 
    101933.5, 101931.6, 101917.8, 101895.5, 101879.2, 101851.1, 101816.4, 
    101774.8,
  98856.68, 97398.12, 97262.1, 98424.65, 100120.7, 100870.5, 101936.6, 
    101949.2, 101931.6, 101933.2, 101913.5, 101896.1, 101867, 101837.6, 101800,
  102204.5, 102264.3, 102288.9, 102291.4, 102311.7, 102321.3, 102319.2, 
    102298.8, 102271.2, 102235.2, 102188.5, 102136.1, 102076.6, 102011.4, 
    101943.1,
  100766.9, 102201.3, 102264.7, 102297, 102316.2, 102331.4, 102330.1, 
    102322.9, 102304.1, 102277.4, 102241.4, 102200.7, 102150, 102093.4, 
    102031.7,
  100851.1, 101854.1, 102219.8, 102258.6, 102288.5, 102310.3, 102317.6, 
    102321.2, 102314.3, 102298.3, 102272.9, 102241.2, 102199.9, 102150.2, 
    102097.2,
  100472.4, 101744.7, 102162.8, 102214.5, 102242.6, 102266.7, 102286.8, 
    102297.8, 102300, 102293.6, 102281.9, 102256.5, 102228.1, 102187, 102139.9,
  100416.9, 101086.9, 101961.8, 102170, 102194.3, 102217.7, 102237.8, 102261, 
    102267.7, 102269.8, 102266.4, 102255.9, 102239.7, 102209.5, 102168.9,
  100072.7, 99912.41, 100801.3, 102055.8, 102154.2, 102171.6, 102196.2, 
    102212.7, 102223.2, 102235.5, 102239.2, 102234, 102222.9, 102203.7, 
    102170.4,
  99956.16, 99339.79, 99288.98, 101042.2, 102086.9, 102119.2, 102142.6, 
    102158.4, 102177.3, 102185.1, 102191.8, 102193.3, 102194, 102177.9, 
    102155.2,
  100169.9, 99466.13, 99881.84, 100384.3, 101966.2, 102078.2, 102094.7, 
    102112.3, 102124, 102141.4, 102148.8, 102153.6, 102150.6, 102143.6, 
    102135.5,
  98957.85, 98828.98, 100109, 100442.1, 101071.6, 102029, 102088.9, 102092, 
    102094.5, 102104.1, 102097.5, 102104.2, 102105.4, 102105.2, 102102.9,
  98933.36, 97507.35, 97384.16, 98573.66, 100274.4, 101035.1, 102088.2, 
    102111.3, 102087.4, 102094.2, 102080.7, 102085.8, 102083.7, 102091.4, 
    102095.8,
  101591.1, 101686.8, 101773.9, 101856.4, 101933.7, 101996.3, 102053.2, 
    102107.1, 102154, 102189.7, 102221.1, 102237.7, 102239.5, 102234.1, 
    102224.1,
  100204, 101632.6, 101747.8, 101829.7, 101913.7, 101989.9, 102055, 102111.1, 
    102160.4, 102200.3, 102233, 102251, 102265.8, 102269.5, 102267,
  100307.6, 101325.5, 101726.4, 101802.7, 101885.1, 101961.2, 102034.4, 
    102094.1, 102151, 102199.7, 102238.8, 102267.1, 102288.9, 102301.7, 
    102304.1,
  99984.82, 101263, 101687.5, 101775.2, 101847.9, 101928.1, 102008.6, 
    102075.4, 102131.6, 102182.3, 102226.2, 102263.9, 102295.7, 102320.4, 
    102334.8,
  99946.63, 100631.9, 101516.3, 101745.7, 101810.5, 101884.9, 101967.4, 
    102040.6, 102099.8, 102152.7, 102200.5, 102245.1, 102280.3, 102312.8, 
    102338.9,
  99636.55, 99491.65, 100381.9, 101659.7, 101775.4, 101838.9, 101910.7, 
    101993.8, 102057.1, 102113.5, 102160.1, 102203.2, 102246.8, 102288, 102324,
  99541.73, 98937.84, 98920.33, 100662.4, 101742.3, 101803.6, 101863.2, 
    101930.3, 101992.3, 102044.8, 102099.1, 102140, 102184.5, 102231.7, 
    102281.6,
  99772.95, 99078.75, 99528.68, 100039.7, 101634.3, 101764.7, 101816.4, 
    101875.3, 101930.8, 101976.2, 102014.3, 102051.1, 102088.3, 102137.8, 
    102193,
  98577.91, 98438.52, 99741.21, 100106.2, 100752.3, 101716.8, 101797.2, 
    101827.3, 101874.1, 101901.6, 101922.5, 101945.5, 101984.6, 102042.4, 
    102112.7,
  98575.96, 97158.2, 97033.7, 98207.21, 99932.15, 100699.8, 101787.4, 
    101808.2, 101830.1, 101855.4, 101849.4, 101851.7, 101857, 101907.8, 
    102004.8,
  101012.1, 101087.6, 101148.6, 101196.7, 101246.3, 101301.3, 101358.9, 
    101420.8, 101470.8, 101522.7, 101572.4, 101617.1, 101655.8, 101724.2, 
    101773.7,
  99666.02, 101077.9, 101181.6, 101229.5, 101279, 101333.9, 101391.4, 
    101454.2, 101501.6, 101546.7, 101577.6, 101612.9, 101660.7, 101689.1, 
    101739.5,
  99810.08, 100812.2, 101202.6, 101257.4, 101307.9, 101361.3, 101413, 
    101472.8, 101513.2, 101552.1, 101577.9, 101602.1, 101625.6, 101651.4, 
    101734.7,
  99546.38, 100782.8, 101202.7, 101276.6, 101323.1, 101373.7, 101426.6, 
    101482, 101521.9, 101554.3, 101568.8, 101576.8, 101576.4, 101628.2, 
    101723.9,
  99530.27, 100194.3, 101064, 101283.3, 101332.6, 101380.2, 101432.1, 101481, 
    101522.7, 101551, 101553, 101546.7, 101553.1, 101621.4, 101716.4,
  99238.27, 99092.09, 99960.76, 101211, 101333.2, 101375.7, 101429.8, 
    101476.6, 101517.6, 101541.6, 101544.3, 101524.8, 101534, 101604, 101715.1,
  99162.2, 98571.64, 98535.73, 100238.9, 101310.8, 101372.1, 101414, 
    101466.5, 101506.3, 101532.6, 101539.6, 101513.1, 101536.4, 101611.3, 
    101712.3,
  99405.19, 98723.1, 99146.84, 99638.83, 101200.1, 101352.1, 101403.9, 
    101456.5, 101501.5, 101531.6, 101541.5, 101530, 101541.6, 101618.9, 
    101713.6,
  98249.83, 98110.36, 99361.49, 99725.96, 100327.9, 101284.9, 101389.4, 
    101440.8, 101493.9, 101538.8, 101552.3, 101551.4, 101569.3, 101642.9, 
    101724.3,
  98289.62, 96890.41, 96736.71, 97864.78, 99526.36, 100278.5, 101367.4, 
    101450.8, 101484.5, 101546.5, 101570.7, 101588.5, 101606.9, 101666.6, 
    101746.6,
  101785.6, 101795.7, 101769.7, 101731.7, 101707, 101669.2, 101628.5, 
    101589.9, 101547.5, 101503.8, 101466.4, 101427.8, 101389.2, 101348.2, 
    101301.9,
  100304.9, 101679.9, 101713.2, 101690.3, 101681.1, 101666.7, 101647.6, 
    101621.3, 101588.5, 101557.1, 101527.1, 101500.1, 101477, 101447.5, 101404,
  100353.1, 101334.3, 101661.8, 101647.4, 101652.9, 101645.9, 101639.6, 
    101634.8, 101614.5, 101595.8, 101578.2, 101560.3, 101538.6, 101515.9, 
    101489.7,
  99964.41, 101221, 101602, 101611.8, 101615.7, 101623.7, 101630.3, 101634.4, 
    101628.5, 101621.2, 101618.5, 101612.2, 101604.2, 101591.2, 101573.7,
  99863.88, 100544.7, 101397.1, 101569.2, 101581, 101598.2, 101610.1, 
    101625.4, 101635.6, 101638.8, 101643.5, 101645.2, 101651.6, 101651.1, 
    101645.4,
  99528.8, 99372.83, 100240.4, 101467.8, 101539, 101560.1, 101587.2, 
    101610.9, 101637.6, 101651.3, 101667.1, 101685.5, 101696.5, 101700, 
    101704.3,
  99427.82, 98812.01, 98774.98, 100473.8, 101503, 101517.9, 101552.5, 
    101584.2, 101626.3, 101658.6, 101687.5, 101707.9, 101730.2, 101742.7, 
    101766.6,
  99662.36, 98957.85, 99368.42, 99852.97, 101395.5, 101495.8, 101528.1, 
    101567.4, 101620.9, 101670.3, 101706.8, 101735.4, 101765.6, 101785.9, 
    101812,
  98502.64, 98359.49, 99602.28, 99932.74, 100521.1, 101427.7, 101511, 
    101554.6, 101627.8, 101671.7, 101726, 101765.5, 101798.4, 101834.6, 
    101864.8,
  98544.56, 97142.5, 96992.23, 98119.38, 99766.29, 100486.7, 101497.3, 
    101565.1, 101624.7, 101679.9, 101736.1, 101788.7, 101824.6, 101864.8, 
    101901.7,
  101852.8, 101895.4, 101941.2, 102000.6, 102060.9, 102102.1, 102123.5, 
    102145.4, 102151.9, 102156.5, 102151.1, 102136.1, 102107.5, 102071.5, 
    102034,
  100389.4, 101846.8, 101889.4, 101925.5, 101981.6, 102040.1, 102079.6, 
    102117.2, 102138.9, 102146.4, 102162.2, 102167.8, 102152.8, 102130.6, 
    102101.8,
  100406.9, 101442.6, 101846, 101904, 101915.9, 101964.9, 102012.4, 102055.9, 
    102089.9, 102123, 102146.6, 102155.5, 102154, 102150.1, 102129.6,
  100004.5, 101287.2, 101716, 101785.6, 101870.6, 101920.6, 101969.7, 
    102002.3, 102034.1, 102064.4, 102093.1, 102117.5, 102136.7, 102139.1, 
    102132.5,
  99861.68, 100587.7, 101492.1, 101715.3, 101755, 101810, 101873, 101934.3, 
    101984.4, 102027.4, 102060.8, 102073.9, 102094.3, 102107.7, 102110.9,
  99523.51, 99383.31, 100274, 101567.6, 101683.7, 101754.3, 101815.4, 
    101865.7, 101905.1, 101945.8, 101998, 102037.3, 102062.9, 102081.5, 
    102082.6,
  99421.09, 98818.23, 98811.91, 100533.6, 101592, 101639.5, 101718.9, 
    101790.5, 101848.7, 101913.1, 101952.4, 101994.1, 102022.8, 102046.4, 
    102058.2,
  99650.72, 98952.27, 99385.91, 99888.51, 101462.1, 101599.1, 101659.9, 
    101738.3, 101800.5, 101852.2, 101911, 101944.4, 101983.3, 102012.5, 
    102024.2,
  98495.12, 98345.2, 99609.55, 99959.77, 100556, 101483.1, 101619.3, 101696, 
    101780.5, 101842.1, 101897.3, 101935.1, 101974.8, 101998.7, 102018.5,
  98549.57, 97122.11, 96977.2, 98122.38, 99760.98, 100487.4, 101567.2, 
    101672.6, 101751.8, 101824.4, 101891.9, 101942.2, 101984, 102018.4, 
    102045.4,
  101647.1, 101747.5, 101785.3, 101831.3, 101875.9, 101923.9, 101967.3, 
    101996.5, 102025.9, 102038, 102067, 102068.1, 102051.6, 102026.4, 101999,
  100197.6, 101634.1, 101704, 101768, 101821.9, 101869.8, 101908.4, 101942.7, 
    101972.2, 102004.5, 102038.2, 102064.8, 102084.9, 102093.3, 102077.6,
  100204.2, 101229.4, 101609.7, 101657.6, 101710.8, 101757.1, 101818.8, 
    101873.4, 101922.3, 101964.3, 102002.2, 102028.7, 102056.3, 102084.1, 
    102098.9,
  99835.1, 101096.8, 101528.7, 101578.4, 101643.1, 101692.9, 101737.8, 
    101766, 101819.6, 101864, 101926.5, 101986.1, 102030.5, 102059.1, 102078.5,
  99754.6, 100416.4, 101321.7, 101516.1, 101563.6, 101618.7, 101689.2, 
    101757.3, 101813.1, 101857.1, 101891.9, 101930.3, 101973, 102027.1, 
    102063.6,
  99467.46, 99291.48, 100148.5, 101410.9, 101510.9, 101567.2, 101634.4, 
    101700.5, 101762.8, 101819.9, 101881.3, 101928.5, 101957.4, 101982, 
    102014.3,
  99383.97, 98761.96, 98717.36, 100410, 101447.9, 101504.7, 101588.3, 
    101681.2, 101757.5, 101825.8, 101873.8, 101912.8, 101952, 101996.6, 
    102027.6,
  99636.6, 98921.55, 99329.77, 99808.88, 101337.9, 101463.5, 101540.2, 
    101644, 101730.1, 101807.5, 101874, 101920, 101960, 101986.7, 102012.2,
  98495.21, 98334.12, 99573.78, 99902.76, 100482.2, 101408.9, 101514.9, 
    101623, 101722.5, 101804, 101876.7, 101931.3, 101975.8, 102016.3, 102043.2,
  98571.84, 97120.39, 96965.94, 98092.29, 99757.84, 100472.2, 101497.9, 
    101618.5, 101712.2, 101796.2, 101870.8, 101930, 101978.9, 102025, 102061.1,
  101095.7, 101247.4, 101368.9, 101460.7, 101544.8, 101620.4, 101699.9, 
    101768.6, 101819.7, 101872.5, 101920.2, 101963.3, 101987.4, 101993, 
    101991.4,
  99689.04, 101122.6, 101265.7, 101364.8, 101451.7, 101539.1, 101611.4, 
    101685, 101750.2, 101808.8, 101868.2, 101926.2, 101971.6, 102008.6, 
    102025.2,
  99746.63, 100756.6, 101194.2, 101271.8, 101373.1, 101445.9, 101538.9, 
    101631.8, 101700, 101743.6, 101808.2, 101875.8, 101932.8, 101979.8, 
    102023.3,
  99475.31, 100724, 101170.9, 101240.3, 101316.3, 101414, 101482.6, 101572.8, 
    101659.2, 101711.8, 101769.9, 101823.3, 101889, 101947.9, 102000.3,
  99494.36, 100142.2, 101022.2, 101239.6, 101296.8, 101384.4, 101472.7, 
    101564, 101640.9, 101712.6, 101771.4, 101826.3, 101874.1, 101907.5, 
    101959.8,
  99274.02, 99099.81, 99947.37, 101204.5, 101311, 101367.4, 101455.3, 
    101534.2, 101624.4, 101690.9, 101765.5, 101824.5, 101884.8, 101919.7, 
    101958,
  99232.76, 98614.34, 98576.55, 100272.2, 101335.1, 101385, 101457.2, 
    101535.5, 101618.3, 101700.9, 101770.2, 101828.6, 101887.9, 101929.2, 
    101972.1,
  99511.27, 98798.55, 99226.24, 99715.9, 101276.7, 101403.3, 101466.4, 
    101537.9, 101623.8, 101698.9, 101771.5, 101832.6, 101891.5, 101941.7, 
    101986.2,
  98375.95, 98212.84, 99471.74, 99829.93, 100448.8, 101378, 101470.6, 
    101531.5, 101628.5, 101707.1, 101781.7, 101845.7, 101905.9, 101954.8, 
    101996,
  98456.34, 97027.77, 96887.04, 98009.3, 99715.49, 100461.3, 101488, 
    101542.7, 101629.7, 101713.2, 101783.8, 101847.9, 101906.5, 101959.5, 
    102006.3,
  101005.1, 100914.3, 100822.9, 100695.2, 100562.7, 100422, 100293.1, 
    100197.6, 100149.7, 100124.4, 100106.1, 100177.1, 100374.2, 100607.8, 
    100832.6,
  99614.95, 100864.1, 100801.7, 100653, 100524.8, 100409.7, 100306.5, 
    100241.8, 100204.7, 100189, 100188.9, 100245.4, 100407.3, 100612.7, 
    100823.6,
  99794.1, 100684.7, 100940.9, 100809.6, 100693.4, 100585.4, 100478.9, 
    100399, 100343.9, 100299.8, 100281.4, 100302.6, 100407.9, 100584.6, 
    100778.7,
  99547.86, 100681.1, 100986.6, 100903, 100810.6, 100713, 100635.8, 100568.7, 
    100529.1, 100505.6, 100501.3, 100516.7, 100589.6, 100717.4, 100869.8,
  99547.04, 100127.2, 100916, 101015.5, 100945.3, 100869.8, 100808.1, 
    100748.4, 100715, 100693.4, 100691.5, 100708.2, 100757.5, 100845.6, 
    100963.5,
  99283.68, 99047.03, 99843.25, 101010.9, 101037.1, 100976, 100931.2, 
    100891.8, 100876.5, 100871.2, 100880.6, 100903.8, 100951.2, 101021.7, 
    101102.5,
  99189.57, 98532.81, 98451.99, 100091.7, 101100.1, 101078.8, 101046.7, 
    101019.9, 101008.2, 101008.6, 101023.2, 101044.6, 101086.3, 101141.1, 
    101218.1,
  99497.82, 98736.48, 99096.03, 99549.48, 101075.5, 101147, 101129, 101118.8, 
    101114.7, 101123.2, 101138.6, 101162.6, 101200, 101249.3, 101310.7,
  98369.92, 98179.75, 99388.34, 99698.48, 100261.6, 101165.2, 101194.4, 
    101191.1, 101196.4, 101211.1, 101228.6, 101256.2, 101292.1, 101338.8, 
    101396.7,
  98466.55, 96989.88, 96809.87, 97904.8, 99534.41, 100263.9, 101251.4, 
    101277.4, 101263.1, 101297.4, 101314.9, 101347.3, 101379.6, 101425.1, 
    101480,
  101683.1, 101771.8, 101778.9, 101756.2, 101717.8, 101679.7, 101633.8, 
    101586.3, 101519.6, 101427.9, 101294.6, 101099.3, 100882.5, 100674.8, 
    100497,
  100306.3, 101727.1, 101778.1, 101763.2, 101734.2, 101699.7, 101652, 
    101605.3, 101535.6, 101429.5, 101294.8, 101112.8, 100865.2, 100621.9, 
    100425.7,
  100391.3, 101406.9, 101778.2, 101785.8, 101765.6, 101730.4, 101683.4, 
    101634.1, 101564.7, 101472.2, 101337.1, 101154.9, 100892.4, 100615.7, 
    100380,
  100051.8, 101330.9, 101740.7, 101783, 101772.8, 101747.9, 101709.2, 
    101663.9, 101602.7, 101514.1, 101395.5, 101229.9, 101000.5, 100725.7, 
    100469.5,
  99991.49, 100683.9, 101578.3, 101769.3, 101784.8, 101767.7, 101734.9, 
    101689.2, 101634.1, 101557.8, 101455.9, 101313.2, 101120.1, 100881.8, 
    100631.2,
  99671.03, 99509.54, 100419.2, 101686.8, 101773.7, 101772.4, 101754.4, 
    101717.6, 101668.3, 101601, 101511, 101392.3, 101237.8, 101045.2, 100827.9,
  99543.52, 98960.98, 98934.74, 100691.2, 101750.8, 101775.3, 101761.6, 
    101738.7, 101699.2, 101640.2, 101563.5, 101466.6, 101340, 101183.5, 
    101002.9,
  99742.65, 99083.76, 99538.31, 100048.6, 101643.6, 101759.3, 101767.8, 
    101749.4, 101716.1, 101671.9, 101612.1, 101529.4, 101428.2, 101302.9, 
    101154.5,
  98529.41, 98416.83, 99744.62, 100118.8, 100745.3, 101703.2, 101747.4, 
    101745.4, 101729, 101696.8, 101644.8, 101583.4, 101501.2, 101401.6, 101281,
  98566.01, 97124.18, 97012.63, 98216.9, 99935.86, 100725.2, 101749, 
    101743.6, 101716.6, 101703.5, 101661.2, 101614.9, 101546.9, 101471.3, 
    101376.7,
  101175.2, 101296, 101407, 101513, 101604.6, 101683.8, 101764.3, 101854.8, 
    101915.4, 101959.9, 102007.6, 102037.9, 102066.5, 102083.7, 102078.5,
  99791.94, 101265.8, 101392.3, 101483.3, 101588.6, 101667, 101746.5, 
    101835.1, 101906.1, 101952.2, 101994.4, 102028.8, 102043, 102056, 102052.5,
  99893.38, 100947.4, 101381.9, 101475, 101574.3, 101653.5, 101730.5, 
    101815.3, 101893, 101952.1, 101984.9, 102012.2, 102017.4, 102029.3, 
    102018.1,
  99606.27, 100899.6, 101362.4, 101467.2, 101561.9, 101646.5, 101719.6, 
    101795.6, 101873.9, 101936.4, 101974.6, 101995.7, 101998.6, 102005.3, 
    101994.4,
  99605.3, 100280.8, 101191.9, 101450.8, 101550.9, 101635.9, 101713.2, 
    101777.8, 101851.1, 101917.3, 101953.4, 101966.6, 101978.1, 101980.5, 
    101968.4,
  99318.69, 99154.88, 100055.1, 101357.5, 101521.4, 101617.4, 101693.3, 
    101765.4, 101832.8, 101895.8, 101933.8, 101945.1, 101956.5, 101962.3, 
    101946.4,
  99240.19, 98634.38, 98621.36, 100368.9, 101478.9, 101588, 101673.2, 
    101746.9, 101809.9, 101873.1, 101911.1, 101929.1, 101935, 101939.3, 101925,
  99472.91, 98778.62, 99231.88, 99750.8, 101361.4, 101550.6, 101643.9, 
    101722.7, 101791.2, 101840.9, 101887.9, 101912.1, 101916.8, 101918.5, 
    101903.7,
  98299.23, 98152.91, 99438.1, 99822.92, 100476.3, 101482.2, 101620, 
    101688.7, 101771, 101818.6, 101856.5, 101885.9, 101895.9, 101900.2, 
    101886.8,
  98347.31, 96926.85, 96787.71, 97936.86, 99665.66, 100460.1, 101608.3, 
    101681.7, 101734, 101803.5, 101826.8, 101858.1, 101873, 101876.6, 101864.5,
  100476.5, 100428.5, 100392.9, 100369.6, 100385.8, 100453.1, 100585.7, 
    100775, 100991.1, 101218.1, 101416.3, 101585.5, 101737.4, 101855.6, 
    101955.3,
  99129.43, 100419.3, 100456, 100446, 100465.6, 100518.3, 100613.2, 100757.6, 
    100949.3, 101165.4, 101375.9, 101543.6, 101699.5, 101840, 101933.1,
  99281.48, 100198.2, 100528, 100536.2, 100547.7, 100589.4, 100663.4, 100768, 
    100910.5, 101095.1, 101296.9, 101494.8, 101637.1, 101790.1, 101896.1,
  99029.38, 100199.1, 100566.5, 100580.5, 100604.5, 100655, 100728.4, 
    100821.8, 100940.2, 101081, 101251.9, 101438.4, 101588.5, 101728.5, 
    101860.7,
  99074.48, 99657.02, 100482.1, 100654.2, 100676, 100720.6, 100789.8, 
    100885.7, 100994.4, 101111, 101243.6, 101400, 101553.6, 101665.4, 101788.5,
  98824.59, 98605.99, 99421.62, 100632.4, 100728.8, 100774.9, 100853.3, 
    100943.1, 101051.3, 101158.7, 101274.5, 101398.1, 101529.8, 101649.3, 
    101741.4,
  98792.74, 98144.38, 98079.6, 99738.77, 100774.5, 100822, 100897, 100989.4, 
    101094.9, 101206.9, 101308.1, 101418.3, 101522.1, 101624.5, 101714.4,
  99081.79, 98344.59, 98728.7, 99199.22, 100722.7, 100853.6, 100932.5, 
    101031.1, 101131.1, 101240.1, 101339.5, 101440.6, 101530.7, 101623.5, 
    101692.6,
  97972.69, 97786.28, 98993.91, 99336.95, 99913.16, 100845.8, 100957.5, 
    101056.9, 101155.7, 101267.5, 101360.9, 101455.7, 101541.6, 101620.6, 
    101682.2,
  98075.14, 96619.55, 96453.29, 97542.97, 99194.54, 99939.22, 100980.1, 
    101101.7, 101171.3, 101286.9, 101373.1, 101460.4, 101541.9, 101621.2, 
    101675,
  100945.1, 100929.3, 100865.9, 100749.1, 100616.2, 100465.4, 100304.8, 
    100129.1, 99950.19, 99799.73, 99732.64, 99805.54, 99964.17, 100172, 
    100400.3,
  99550.58, 100888.9, 100887.1, 100793.1, 100679.5, 100549.8, 100410.7, 
    100263.6, 100114.5, 99986.91, 99920.59, 99946.53, 100040.7, 100184.1, 
    100355.8,
  99620.5, 100579.3, 100907.8, 100833.5, 100746.7, 100642.5, 100524.7, 
    100400.8, 100272.5, 100150.7, 100062.6, 100044.5, 100107.8, 100213.8, 
    100352,
  99296.6, 100503.8, 100873.6, 100841.8, 100780, 100697.8, 100601.3, 
    100497.5, 100390, 100284.2, 100202, 100160.8, 100195.7, 100267.4, 100367.2,
  99238.63, 99876.74, 100715.9, 100855.6, 100809.6, 100744.5, 100671.9, 
    100581.6, 100492.7, 100400.6, 100317.1, 100263.1, 100255.4, 100312.6, 
    100378.5,
  98900.24, 98707.85, 99555.34, 100770.8, 100813.9, 100761.5, 100707, 100641, 
    100568.6, 100492.4, 100419.9, 100362.7, 100340.2, 100367.4, 100410.2,
  98774.34, 98157.68, 98089.69, 99773.77, 100790.2, 100770.4, 100722.1, 
    100677.4, 100627.5, 100568, 100505.9, 100455.6, 100428, 100431.3, 100472.3,
  99021.45, 98292.27, 98679.35, 99169.15, 100691.1, 100763, 100735.9, 
    100708.9, 100674.2, 100632.5, 100589.5, 100546, 100521.8, 100519.8, 
    100538.7,
  97872.65, 97679.95, 98897.2, 99228.52, 99819.95, 100718.7, 100733, 
    100710.8, 100699.7, 100679.9, 100655, 100632.5, 100610.1, 100609.6, 
    100626.4,
  97947.09, 96481.71, 96319.21, 97410.48, 99046.72, 99776.12, 100750.3, 
    100737.1, 100712.6, 100719, 100703.7, 100701.7, 100692.5, 100699.8, 
    100709.4,
  100871.3, 100933, 100945.5, 100905.1, 100864.4, 100801.8, 100716.4, 
    100616.9, 100522.3, 100458.7, 100431, 100450.6, 100507.5, 100587.2, 
    100674.1,
  99486.52, 100888.3, 100931.2, 100896.2, 100865.7, 100814, 100734.5, 
    100640.1, 100547.4, 100465.3, 100409.2, 100400, 100421.3, 100478.1, 100555,
  99548.42, 100555.6, 100916.4, 100910.6, 100882.5, 100844.1, 100781.9, 
    100691.8, 100589.3, 100491.4, 100404.3, 100352.9, 100342.4, 100377.7, 
    100435.3,
  99210.64, 100478.4, 100865.5, 100894.2, 100886.3, 100855.5, 100809.5, 
    100743, 100653.5, 100552.3, 100459.1, 100383, 100337.7, 100336.4, 100373.4,
  99126.31, 99836.02, 100708.3, 100890.9, 100892.6, 100872.9, 100844.3, 
    100791, 100720.3, 100629.2, 100528.7, 100442.2, 100373.8, 100337.3, 
    100340.4,
  98793.7, 98667.98, 99551.23, 100815.8, 100885.4, 100877.9, 100861.4, 
    100830.1, 100774.4, 100701.8, 100615.2, 100528.5, 100452.7, 100399, 
    100369.7,
  98665.95, 98086.08, 98066.02, 99812.1, 100858.5, 100881.6, 100869.2, 
    100856.3, 100822.1, 100768.9, 100694.9, 100617.2, 100540.5, 100479.5, 
    100432,
  98856.56, 98189.44, 98645.75, 99146.31, 100736.7, 100858.9, 100867.2, 
    100865.4, 100847.5, 100814.6, 100763.6, 100699.1, 100634.5, 100573.6, 
    100521.2,
  97658.21, 97515.83, 98827.88, 99194.43, 99815.61, 100786.7, 100857.2, 
    100864.7, 100863.7, 100847.6, 100808.8, 100764, 100709.7, 100658.6, 
    100610.1,
  97722.73, 96287.2, 96142.46, 97323.84, 99007.84, 99789.4, 100840.3, 
    100858.4, 100856.7, 100863.5, 100835.3, 100809.6, 100765.6, 100726.8, 
    100682.1,
  100810.9, 100819.4, 100819.6, 100813.2, 100817.6, 100793.8, 100759.9, 
    100737.9, 100727.7, 100736.4, 100762.7, 100821.4, 100920.3, 101053.3, 
    101171.6,
  99394.36, 100761.7, 100803.8, 100800, 100796.3, 100803.1, 100781.2, 
    100758.6, 100742.7, 100740.7, 100757.1, 100804.8, 100875.3, 100978.5, 
    101093.8,
  99456.19, 100439.4, 100782.4, 100787.5, 100788.2, 100803.3, 100799.3, 
    100775.7, 100759.2, 100752, 100756.9, 100779.9, 100828.7, 100913.2, 
    101023.8,
  99107.08, 100343.7, 100725.5, 100750.9, 100756.2, 100766.5, 100784.3, 
    100778.3, 100769.4, 100757.2, 100759, 100776.7, 100814, 100869.6, 100955,
  99024.03, 99682.71, 100516.1, 100698.2, 100717.7, 100729.7, 100745, 
    100760.8, 100776.6, 100784.3, 100788, 100796.5, 100814.3, 100842.4, 
    100896.5,
  98717.74, 98519.17, 99384.57, 100604.7, 100674.3, 100692.7, 100727.6, 
    100751.9, 100766.4, 100775.3, 100786.1, 100797.3, 100811.5, 100844.7, 
    100878.1,
  98560.25, 97917.38, 97857.88, 99574.4, 100603.9, 100637.5, 100673.1, 
    100724.7, 100772, 100815.2, 100841.3, 100847.8, 100854.2, 100874, 100897.1,
  98799.84, 98063.11, 98426.59, 98899.2, 100435.5, 100515.8, 100542.1, 
    100596.8, 100672.1, 100746.9, 100801.7, 100847.7, 100875.2, 100900.8, 
    100920.9,
  97617.48, 97418.2, 98622.19, 98959.66, 99511.01, 100397.4, 100420.6, 
    100419.5, 100475.8, 100572.3, 100654.6, 100734.5, 100804.4, 100867.1, 
    100903.8,
  97706.06, 96260.55, 96062.88, 97132.32, 98748.89, 99464.36, 100436.6, 
    100449.8, 100432.2, 100494.8, 100545.1, 100628, 100706, 100799.9, 100874.8,
  101498.8, 101536.1, 101528.7, 101500.8, 101481.6, 101441.4, 101404.9, 
    101382, 101344.9, 101306.7, 101262.5, 101225.5, 101195, 101161.7, 101131.3,
  100070.5, 101465, 101505.7, 101469, 101455.6, 101429.4, 101401.4, 101378, 
    101343.8, 101304.8, 101264, 101225, 101192.3, 101163.7, 101140,
  100141, 101129.3, 101473.6, 101452, 101444.5, 101422.1, 101391.3, 101366.8, 
    101332.7, 101296.6, 101259.3, 101225.2, 101194.6, 101160.9, 101131.9,
  99789.46, 101036, 101412.7, 101427.7, 101413.2, 101394.6, 101372.3, 
    101349.5, 101319.5, 101286.5, 101250.4, 101216.7, 101182, 101154.9, 
    101127.3,
  99707.25, 100369.2, 101221, 101396.3, 101386.8, 101372.2, 101351.1, 
    101329.1, 101301.1, 101268, 101236.3, 101205.7, 101180.2, 101158.4, 
    101136.7,
  99386.8, 99205.13, 100068.5, 101296, 101361.6, 101344.7, 101327.7, 
    101308.3, 101282.8, 101250.7, 101217.1, 101186.2, 101158.1, 101134, 
    101111.5,
  99224.12, 98604.95, 98566.68, 100303.4, 101316.3, 101321.5, 101302.9, 
    101280.7, 101252.3, 101219.4, 101179.1, 101140.8, 101102.8, 101073.4, 
    101061.1,
  99425.5, 98727.74, 99147.05, 99649.37, 101207.3, 101289.6, 101271.4, 
    101245.7, 101208.5, 101164.7, 101118.9, 101074.9, 101037.3, 101007.3, 
    100983.8,
  98186.09, 98070.23, 99334.88, 99683.43, 100292.1, 101222.5, 101248.3, 
    101204.5, 101168.3, 101122.5, 101063.5, 101002.6, 100944.1, 100905.1, 
    100871.9,
  98146.32, 96741.27, 96635.67, 97814.16, 99485.74, 100244.5, 101213.2, 
    101189.4, 101113.6, 101054.1, 100972.7, 100894.9, 100813, 100763.1, 
    100721.8,
  101519, 101587.1, 101626.5, 101649.6, 101686.2, 101709.7, 101710.7, 
    101714.9, 101726.4, 101731.2, 101726.5, 101724.4, 101720.1, 101716.4, 
    101692.5,
  100129.9, 101544.4, 101618.5, 101655.4, 101685, 101704.8, 101714.9, 
    101726.4, 101743.2, 101740.2, 101741.9, 101735.4, 101734, 101696.2, 
    101660.5,
  100209.5, 101221.8, 101601.5, 101646.3, 101680.7, 101707.4, 101725.1, 
    101750.2, 101753.8, 101749, 101740.2, 101739.3, 101726.3, 101696.6, 
    101646.8,
  99871.48, 101149.1, 101557.6, 101625.4, 101663.8, 101687.6, 101716.7, 
    101735.5, 101734.4, 101734.5, 101724, 101723.4, 101704.5, 101674.3, 
    101614.9,
  99800.19, 100492.7, 101377.6, 101590.5, 101636.5, 101671, 101696.8, 
    101710.1, 101717.3, 101712.4, 101702.7, 101697.4, 101677.1, 101645.4, 
    101584.8,
  99474.88, 99312.58, 100222.1, 101492.1, 101598.8, 101638.8, 101665.4, 
    101685.5, 101686.7, 101682.2, 101675.9, 101660.5, 101640.8, 101612.1, 
    101556.5,
  99330.27, 98731.28, 98725.23, 100485, 101550.1, 101600.8, 101629.4, 
    101644.2, 101653.7, 101647.6, 101638.7, 101622.9, 101603.7, 101577.6, 
    101534.1,
  99509.38, 98843.84, 99299.12, 99823.12, 101433.1, 101551.7, 101589.4, 
    101608.3, 101615.5, 101617.2, 101605.5, 101594.2, 101571.7, 101545.9, 
    101507.2,
  98248.45, 98149.29, 99471.77, 99866.55, 100514.8, 101484.4, 101552, 
    101570.6, 101585.4, 101584.7, 101574.1, 101561.2, 101537.3, 101514.4, 
    101484,
  98229.65, 96829.37, 96731.27, 97948.38, 99678.57, 100478.4, 101532.4, 
    101548.1, 101550, 101557.6, 101542.5, 101530, 101504.5, 101484.2, 101453.4,
  101601.1, 101662.2, 101690.6, 101706.3, 101724.5, 101739.2, 101752.1, 
    101759.7, 101763.4, 101757.8, 101750.9, 101734.6, 101718.5, 101693.3, 
    101677.8,
  100183, 101604, 101684.2, 101723.8, 101757.9, 101783.3, 101799.2, 101813.4, 
    101829.2, 101827.4, 101830, 101818.7, 101807.1, 101787.3, 101765.8,
  100261.3, 101268.7, 101641.5, 101684.2, 101725.2, 101768.7, 101811.5, 
    101851.8, 101877.3, 101886, 101889.8, 101883.4, 101877, 101860.6, 101842.6,
  99916.95, 101179.9, 101607.6, 101675.2, 101718.2, 101768.5, 101810.3, 
    101846.9, 101872.7, 101898.3, 101916.7, 101917.8, 101920.7, 101907, 
    101888.4,
  99834.78, 100502.7, 101393.9, 101603.3, 101652.7, 101706.3, 101769.6, 
    101831.7, 101880.5, 101903.5, 101921.6, 101934.2, 101938.4, 101942.2, 
    101916.9,
  99517.83, 99329.35, 100226.7, 101489.8, 101617.8, 101672.2, 101718.3, 
    101768.6, 101828.2, 101875.6, 101918.2, 101936.4, 101949.8, 101949.1, 
    101922.2,
  99362.08, 98705.48, 98707.35, 100472.6, 101566.2, 101645.6, 101693.8, 
    101737.4, 101785.7, 101834.7, 101877.9, 101899.7, 101921.1, 101923, 
    101905.4,
  99522.41, 98794.33, 99200.07, 99715.77, 101332.7, 101511.4, 101599.6, 
    101675.6, 101728.2, 101779.6, 101824.9, 101861.6, 101879.1, 101883.4, 
    101872.2,
  98262.81, 98126.94, 99336.77, 99691.75, 100342.7, 101378.4, 101516.4, 
    101588.6, 101669.6, 101726.4, 101764.6, 101801.3, 101821.2, 101834.5, 
    101829.2,
  98254.45, 96824.65, 96639.62, 97756.74, 99438.53, 100230.9, 101438.3, 
    101521.8, 101591.5, 101674.1, 101709.3, 101749.9, 101766.8, 101782.7, 
    101791.6,
  101485.5, 101585.4, 101632.3, 101668.3, 101723.1, 101771.5, 101819.2, 
    101862.9, 101900.4, 101923.9, 101945.8, 101952.7, 101969.5, 101990.8, 
    102016.2,
  100081.7, 101498.2, 101573.6, 101617.3, 101685.4, 101748.1, 101807.9, 
    101864.8, 101908.4, 101943.5, 101969.2, 101984.5, 102002.6, 102012.5, 
    102017.3,
  100136.7, 101121.4, 101499, 101559.1, 101624.9, 101705.2, 101775.1, 
    101842.5, 101899.3, 101949.7, 101984.6, 102011.9, 102028, 102041.9, 102049,
  99773.53, 101004.3, 101425.1, 101489.2, 101554, 101632.2, 101716.9, 
    101794.3, 101857.8, 101919.2, 101966.5, 102007.7, 102040.1, 102062.8, 
    102074.2,
  99697.15, 100313.5, 101181.6, 101397.6, 101483.9, 101560.2, 101636.4, 
    101723.4, 101795.3, 101875, 101938.5, 101992, 102033.9, 102068.4, 102091.9,
  99361.09, 99112.79, 99975.74, 101223, 101372.9, 101467.8, 101558.8, 
    101644.8, 101723.5, 101802.9, 101882, 101947.3, 102003.4, 102046.7, 
    102081.2,
  99237.52, 98541.34, 98453.64, 100148.6, 101256.3, 101365.2, 101466.9, 
    101569, 101652.2, 101736.3, 101809.3, 101886.9, 101946.3, 102002.3, 
    102047.2,
  99473.98, 98693.17, 99029.33, 99471.91, 101051.6, 101263.6, 101377.7, 
    101481.5, 101578.8, 101665, 101739.1, 101821.6, 101885.5, 101942.9, 101995,
  98282.14, 98088.12, 99275.05, 99574.55, 100128.6, 101121.6, 101286.8, 
    101405.2, 101509.8, 101607.3, 101669, 101747.4, 101816.7, 101884.1, 
    101929.2,
  98317.53, 96854.49, 96655.52, 97751.51, 99383.91, 100135.6, 101245.6, 
    101365.6, 101442.8, 101568.9, 101629.1, 101693.4, 101739.5, 101800.6, 
    101853.6,
  101350.4, 101289.5, 101222.3, 101141.6, 101111.1, 101079.4, 101080.1, 
    101106.7, 101168.3, 101253.8, 101353.7, 101459.6, 101559.1, 101643.4, 
    101711.1,
  99918.16, 101216.9, 101205.4, 101142, 101096.8, 101077.1, 101083.6, 
    101113.5, 101165.2, 101248, 101345.5, 101450.6, 101548.9, 101637.5, 
    101718.5,
  100018.2, 100922.7, 101220.1, 101148.1, 101104.1, 101082.7, 101077.2, 
    101100, 101145.8, 101229, 101330, 101432.8, 101530.3, 101619.4, 101708.7,
  99703.23, 100867, 101200.2, 101148.3, 101104.3, 101080.4, 101073.8, 
    101099.7, 101152.7, 101240.7, 101336.6, 101438, 101534.9, 101618.2, 
    101699.9,
  99678.26, 100267.9, 101059.3, 101170.9, 101124.8, 101094.8, 101093.9, 
    101117.8, 101172.6, 101249.3, 101340.3, 101438.9, 101532.3, 101624.9, 
    101709.4,
  99404.73, 99155.81, 99964.16, 101136.5, 101164.7, 101133.3, 101130.7, 
    101150.3, 101188.4, 101244.8, 101325.2, 101418.4, 101509.3, 101598, 
    101681.9,
  99308.47, 98630.73, 98538.59, 100190.3, 101194.9, 101183.4, 101166.2, 
    101174.2, 101203.9, 101253.4, 101322.4, 101402.1, 101485.5, 101571.1, 
    101660.2,
  99546.24, 98789.24, 99148.21, 99606.74, 101135.6, 101212.3, 101203.4, 
    101208.6, 101225.5, 101266.1, 101320.2, 101390, 101462.4, 101535.2, 
    101612.1,
  98350.65, 98176.05, 99391.47, 99707.77, 100275.3, 101180.9, 101210.2, 
    101214, 101235.8, 101275.9, 101320.7, 101381.8, 101440.2, 101502.4, 
    101567.8,
  98370.97, 96923.39, 96760.77, 97874.95, 99511.62, 100250.3, 101227.1, 
    101249.5, 101242.9, 101285.2, 101321.6, 101373.9, 101414.9, 101463.3, 
    101514.6,
  101850.2, 101730, 101574.4, 101354.9, 101135.7, 100910.2, 100679.7, 
    100454.5, 100229.5, 100054.3, 99957.51, 99943.86, 99996.04, 100075.6, 
    100165.3,
  100408.3, 101687.5, 101607, 101425, 101227.9, 101024.8, 100820.8, 100623.2, 
    100440.3, 100296.4, 100208.1, 100174.4, 100190.1, 100237.6, 100308.6,
  100529.6, 101434.2, 101670, 101509.8, 101339.1, 101162.1, 100987.9, 
    100819.9, 100664, 100532.7, 100434.5, 100378, 100368.4, 100389, 100429.9,
  100204.4, 101362.6, 101660.9, 101547.8, 101403.1, 101250.4, 101094.9, 
    100949.1, 100815.7, 100701.5, 100612.7, 100556.2, 100535.2, 100536.9, 
    100557.7,
  100145.9, 100748.1, 101527.8, 101596.5, 101472.9, 101341.7, 101209.5, 
    101077.5, 100959.5, 100854.5, 100767.3, 100704.8, 100669, 100656.3, 
    100667.1,
  99809.48, 99559.05, 100364.2, 101527.4, 101497, 101385, 101271, 101159.7, 
    101052.2, 100960.5, 100880.6, 100822.7, 100791, 100771.9, 100769.8,
  99649.37, 98942.59, 98840.8, 100530.6, 101492.9, 101419.3, 101318, 
    101226.4, 101135.4, 101059.8, 100987.7, 100926.1, 100882.5, 100855.5, 
    100847.2,
  99849.46, 99048.73, 99407.62, 99873.58, 101393.4, 101411.2, 101329.9, 
    101254, 101176.9, 101108.2, 101047.2, 100993.6, 100955.2, 100931.8, 
    100914.1,
  98589.96, 98388.38, 99619.65, 99925.6, 100491.6, 101361.7, 101324.1, 
    101245.4, 101180.5, 101129.5, 101072.1, 101028.6, 100992.2, 100963.3, 
    100945.1,
  98547.88, 97050.5, 96868.13, 98004.77, 99653.44, 100381.8, 101318.7, 
    101252.2, 101169.4, 101137.9, 101080.9, 101048.5, 101012, 100989.9, 
    100967.2,
  102204.8, 102143, 102041.5, 101881.2, 101772.6, 101645.7, 101495.2, 
    101321.9, 101128.5, 100902, 100647.6, 100385.7, 100149.7, 99972.74, 
    99831.56,
  100752.5, 102100.3, 102046.7, 101883.6, 101761.3, 101635.9, 101481.8, 
    101314.9, 101129.2, 100914.2, 100670.7, 100402.9, 100166.7, 99978.92, 
    99833.29,
  100838.9, 101793.9, 102052.8, 101900.2, 101779.6, 101652.6, 101511.8, 
    101351.7, 101174.8, 100969.5, 100737.8, 100482, 100238.6, 100030.8, 
    99865.65,
  100536, 101740.4, 102047.8, 101923.8, 101789.1, 101669.2, 101533.1, 
    101385.8, 101222, 101034.3, 100824.2, 100588.9, 100348.1, 100134.7, 
    99956.77,
  100493.7, 101113.3, 101884.2, 101944, 101814.6, 101691.6, 101566.7, 
    101428.2, 101279.8, 101111.8, 100923.3, 100713.5, 100494.1, 100279.8, 
    100096.6,
  100199.1, 99940.38, 100758.6, 101900.7, 101840.7, 101720.1, 101600, 101471, 
    101333.7, 101181.4, 101013.1, 100829.2, 100632, 100438.8, 100260.3,
  100085.4, 99367.87, 99240.93, 100930.4, 101859.2, 101753.8, 101631.3, 
    101511.5, 101385.1, 101249.5, 101099.5, 100940.1, 100767.4, 100593.2, 
    100425.9,
  100322.6, 99520.88, 99867.6, 100313.6, 101815.5, 101786.2, 101667, 
    101551.8, 101428.3, 101305.2, 101171.9, 101030.9, 100882.2, 100728.6, 
    100580.3,
  99071.19, 98871.14, 100113.3, 100398.6, 100953.5, 101778, 101700.1, 
    101581.8, 101472, 101360.3, 101240.7, 101117.3, 100986.2, 100854.6, 
    100724.5,
  99063.65, 97540.96, 97372.9, 98525.99, 100155.2, 100877, 101740.2, 
    101644.9, 101501.4, 101412.6, 101295, 101190.2, 101073.4, 100960.6, 
    100848.8,
  102510, 102544.1, 102508.4, 102470.9, 102446.3, 102404.8, 102351.5, 
    102289.6, 102221.8, 102137.3, 102040.6, 101922.9, 101780.5, 101616.2, 
    101431.5,
  101057.9, 102483.8, 102499.3, 102452.5, 102432.3, 102395.3, 102344.3, 
    102285.3, 102221.2, 102141.6, 102047.6, 101935.5, 101797.2, 101634.4, 
    101451.7,
  101138.2, 102135.6, 102466.3, 102440.6, 102423.3, 102386.8, 102341.2, 
    102294.3, 102234, 102157.3, 102065.4, 101957.8, 101826.8, 101674.5, 101503,
  100790.2, 102060.7, 102420.5, 102417.5, 102401.6, 102373.3, 102332.4, 
    102288.6, 102237.2, 102164.4, 102080.1, 101978.7, 101856.3, 101713.3, 
    101551.2,
  100719.2, 101387.8, 102218.9, 102388, 102383.7, 102356.8, 102323.7, 
    102283.7, 102241.6, 102175.1, 102095.7, 101999.9, 101887.5, 101755.7, 
    101606.2,
  100385.7, 100189.4, 101064.7, 102295.3, 102359.2, 102338.5, 102313.9, 
    102282.5, 102241.9, 102181.1, 102109.5, 102021.8, 101918, 101798.4, 101660,
  100249.4, 99589.39, 99534.56, 101283.6, 102316, 102323.6, 102300, 102276.9, 
    102239.9, 102188, 102123.2, 102042.6, 101949.5, 101839.3, 101713.2,
  100440.4, 99717.45, 100141.7, 100637.6, 102223.9, 102297.5, 102286, 
    102266.7, 102231.7, 102189.8, 102132.3, 102059.4, 101973.6, 101876.2, 
    101761.9,
  99164.75, 99040.35, 100342.9, 100684.8, 101297.2, 102236.1, 102270.3, 
    102246.4, 102220.1, 102187.2, 102135.9, 102071.8, 101993.3, 101904.8, 
    101803.2,
  99130.55, 97673.1, 97564.01, 98781.64, 100503.4, 101258.4, 102246.4, 
    102244.8, 102204.3, 102182.7, 102132.4, 102078.9, 102005.5, 101928.5, 
    101838.3,
  102447.8, 102513.4, 102549.2, 102555.9, 102604.7, 102622.6, 102617.8, 
    102615.7, 102620.9, 102607.6, 102574.1, 102533, 102486.7, 102422.3, 
    102341.9,
  100988.1, 102436.1, 102509.3, 102523.1, 102562, 102581.9, 102605.3, 
    102625.8, 102625.4, 102622.1, 102601.7, 102564.9, 102519.6, 102459.1, 
    102389.5,
  101048.6, 102073.6, 102451.9, 102485.2, 102532.5, 102566.5, 102596.7, 
    102616.6, 102632.3, 102639.1, 102625.6, 102594.3, 102555, 102503.4, 
    102436.8,
  100674.9, 101977.8, 102391.9, 102440.1, 102492.9, 102540.4, 102574.6, 
    102611.1, 102628.3, 102629.1, 102632.1, 102604.2, 102566.9, 102520.8, 
    102468.1,
  100604.5, 101296.3, 102194.1, 102401.5, 102449.1, 102513.4, 102556.2, 
    102593.8, 102622, 102627.5, 102623.4, 102609.1, 102576.7, 102538.6, 
    102487.4,
  100263.8, 100089.6, 101004.7, 102302.9, 102407.9, 102469.3, 102527, 102566, 
    102600.9, 102613.6, 102616.6, 102605.2, 102580.5, 102546.5, 102505.1,
  100115.6, 99498.67, 99485.37, 101267.6, 102369.3, 102424, 102482.5, 
    102529.5, 102560.4, 102587.2, 102596.3, 102593.4, 102579.6, 102551.2, 
    102510.7,
  100310.7, 99617.81, 100073.4, 100597.9, 102243.8, 102379.6, 102439.9, 
    102492.7, 102529.7, 102556.2, 102569.1, 102572.2, 102563.2, 102543.5, 
    102507,
  99050.44, 98916.99, 100241.1, 100641.7, 101298.1, 102306.1, 102397.4, 
    102445.9, 102498.6, 102528.5, 102543.3, 102547.8, 102543.2, 102529, 
    102501.2,
  99062.22, 97607.82, 97492.07, 98691.7, 100469.3, 101265.4, 102367.1, 
    102412.2, 102457.1, 102493.6, 102512.1, 102520.3, 102516.1, 102508.3, 
    102487.3,
  101957.5, 101987.8, 102081.5, 102085.5, 102171.9, 102212.3, 102292.9, 
    102376.3, 102463.7, 102527.9, 102561.4, 102564.2, 102572.5, 102569.5, 
    102562.9,
  100517.1, 101929.9, 102015, 102041.8, 102123.6, 102205.8, 102284.4, 
    102371.7, 102443.4, 102506.4, 102553.5, 102578.8, 102583.5, 102584.6, 
    102585.9,
  100597.8, 101590.8, 101979.4, 102031.1, 102078.8, 102160.7, 102233.5, 
    102334.1, 102428.6, 102506.2, 102560.2, 102596.3, 102608.9, 102607.2, 
    102597.3,
  100246, 101509.9, 101926.5, 101985.1, 102054.2, 102143.9, 102229.4, 
    102313.1, 102399.4, 102474.5, 102538.3, 102584.3, 102611.7, 102620.5, 
    102615.6,
  100192.1, 100860.1, 101746.1, 101958.3, 102016.1, 102098.7, 102191.7, 
    102281.9, 102366.5, 102447.2, 102512.1, 102565, 102600.3, 102622.7, 
    102624.9,
  99856.45, 99673.93, 100577.5, 101870.3, 101983.8, 102064.5, 102155.4, 
    102252.2, 102328.9, 102411.3, 102479.9, 102537.8, 102579.6, 102605.9, 
    102616.3,
  99729.93, 99113.2, 99089.17, 100856.8, 101957.5, 102028.3, 102106.9, 
    102202.4, 102290.4, 102367.3, 102438.9, 102501.2, 102548, 102581.5, 
    102599.2,
  99962.05, 99233.59, 99693.09, 100221.5, 101850, 102000.9, 102071.9, 
    102161.1, 102250.3, 102322.7, 102394.3, 102453.7, 102504.3, 102539.9, 
    102571.7,
  98738.12, 98583.16, 99894.37, 100298.6, 100950.7, 101944, 102041.5, 102116, 
    102201.4, 102285, 102345.4, 102407.7, 102458.5, 102505.3, 102539.8,
  98812.39, 97345.66, 97184.8, 98381.79, 100131.3, 100923, 102011.9, 
    102090.2, 102151.9, 102248.9, 102296.2, 102365, 102409.3, 102457.3, 
    102495.4,
  101372.7, 101426.8, 101455, 101446.1, 101456.9, 101477.3, 101519.4, 
    101582.3, 101677.8, 101814.4, 101968.3, 102112, 102228.5, 102306.2, 
    102379.6,
  99990.09, 101390.5, 101454.9, 101442.9, 101452.9, 101464.7, 101510, 
    101573.9, 101663, 101788.5, 101939.1, 102095.1, 102214.8, 102310.5, 
    102382.9,
  100097.2, 101076.3, 101450.1, 101461.1, 101466.1, 101489.8, 101517, 
    101590.2, 101669.9, 101774.6, 101914, 102075.5, 102202.3, 102310.3, 
    102387.1,
  99779.64, 101032.8, 101438.5, 101460, 101473.3, 101497.9, 101528.2, 
    101602.7, 101683.1, 101791, 101912.5, 102054.5, 102176.7, 102287.4, 
    102375.9,
  99752.26, 100416.2, 101278.8, 101474.9, 101486.8, 101515.1, 101549.9, 
    101624.4, 101711.2, 101806.1, 101906.1, 102025.5, 102151.6, 102268.4, 
    102366.6,
  99462.81, 99282.99, 100138.6, 101410.7, 101504.5, 101524.4, 101572.2, 
    101645.5, 101724.1, 101807.6, 101910.9, 102022.8, 102139, 102248.8, 
    102348.4,
  99365.98, 98734.52, 98690.3, 100422.3, 101498.7, 101535.7, 101576, 
    101659.7, 101736.4, 101836.3, 101921.5, 102021.4, 102130, 102242.2, 102338,
  99602.8, 98883.72, 99311.59, 99809.64, 101397.2, 101535.6, 101582.8, 
    101676, 101754.2, 101846.5, 101938.5, 102034.9, 102130.9, 102230.2, 
    102324.5,
  98423.12, 98268.88, 99523.58, 99907.41, 100517.8, 101495.3, 101604.5, 
    101691.7, 101775.5, 101862.6, 101939.3, 102039, 102127.6, 102219.7, 102307,
  98484.22, 97054.5, 96898.65, 98038.69, 99735.44, 100527, 101601, 101720.3, 
    101781.7, 101889.1, 101954.1, 102032.6, 102112.3, 102196.7, 102278.2,
  101658.4, 101666.9, 101669.8, 101655.8, 101650.2, 101641.3, 101628.9, 
    101617.5, 101607.5, 101598.6, 101604.9, 101638.9, 101691.6, 101756.3, 
    101815.8,
  100221.7, 101596.1, 101663.2, 101662.1, 101663.2, 101664.3, 101664.5, 
    101665, 101661.8, 101663.8, 101670.4, 101705.5, 101761.2, 101826, 101894.9,
  100325.6, 101295.3, 101648.8, 101651.7, 101663.1, 101670.4, 101682.6, 
    101696.4, 101714.6, 101722.1, 101730.8, 101767.7, 101831, 101906.1, 
    101986.1,
  99982.9, 101188.7, 101603.7, 101625, 101639.1, 101668.1, 101693.5, 
    101719.3, 101757.7, 101788.9, 101820, 101864.4, 101931.9, 102006.1, 
    102081.6,
  99922.79, 100559.3, 101418.4, 101596.4, 101624.5, 101656.2, 101706.1, 
    101755.9, 101804.3, 101851.7, 101893, 101944.8, 102008.5, 102076.2, 
    102150.6,
  99603.03, 99411.38, 100261.1, 101504.4, 101617.8, 101648.7, 101707.7, 
    101775.7, 101832.6, 101893.5, 101954.2, 102014.7, 102077.3, 102146.8, 
    102219.2,
  99528.03, 98884.12, 98846.76, 100534.8, 101601.1, 101643.8, 101707.5, 
    101789.8, 101862.2, 101930.6, 101997.5, 102062.9, 102128.1, 102194.9, 
    102268.9,
  99777.09, 99046.23, 99467.31, 99950.15, 101520.9, 101642.9, 101720.2, 
    101804.5, 101879, 101958.6, 102027.7, 102097.8, 102163.3, 102236.3, 
    102310.7,
  98618.16, 98452.98, 99704.39, 100055.8, 100663, 101604.7, 101725, 101813.7, 
    101894.2, 101975.5, 102051, 102121.7, 102190.2, 102262.7, 102335.8,
  98684.96, 97245.65, 97091.88, 98221.13, 99910.75, 100655.1, 101726.2, 
    101838.7, 101910.3, 101991.6, 102066.3, 102134.8, 102203.7, 102272, 
    102344.2,
  102091.9, 102137.8, 102150.2, 102134.8, 102129.3, 102107.9, 102084.9, 
    102057.2, 102025.9, 101988.9, 101955.8, 101919, 101883.4, 101852.6, 
    101813.5,
  100637, 102067.3, 102111.7, 102103.9, 102097.9, 102083.5, 102065.4, 
    102040.1, 102013, 101982.9, 101954.8, 101926.2, 101900.1, 101872.6, 
    101849.4,
  100683.5, 101693.6, 102055, 102054.6, 102058, 102054.7, 102048.1, 102038.9, 
    102023.3, 101995.9, 101969.1, 101939.2, 101910.8, 101883.5, 101862.4,
  100329.5, 101581.3, 101994.5, 102001.1, 102001.2, 102004.4, 101999, 
    102000.1, 101991.1, 101978.5, 101965.3, 101951, 101937.6, 101923.1, 
    101906.8,
  100235.1, 100905.1, 101787.8, 101950, 101953.5, 101961.3, 101967.4, 
    101986.3, 101989.4, 101987.5, 101976.7, 101968.4, 101954.3, 101945.3, 
    101934.1,
  99892.06, 99733.84, 100601.1, 101835.6, 101890.3, 101895.1, 101917.2, 
    101939.1, 101964.7, 101978.6, 101979.2, 101974, 101969.2, 101966.9, 
    101973.6,
  99769.07, 99126.62, 99090.86, 100797.4, 101849.3, 101859.7, 101883, 
    101923.5, 101953.5, 101981.3, 101999.1, 102010.5, 102018.5, 102031.2, 
    102051.5,
  100032.7, 99287.59, 99695.7, 100168.4, 101754.3, 101842.4, 101864.1, 
    101914.7, 101958.3, 101995.2, 102025.1, 102046.1, 102067.9, 102091.8, 
    102121.5,
  98859.01, 98683.06, 99937.63, 100273.4, 100866, 101784, 101855.7, 101915.2, 
    101970.5, 102023.2, 102065.4, 102098, 102128.3, 102158.8, 102194.1,
  98930.62, 97470.84, 97312.3, 98425.78, 100104.8, 100839.8, 101849.4, 
    101928.6, 101984.3, 102038.2, 102086.8, 102130.5, 102164.2, 102205.1, 
    102240.4,
  101955.2, 102000, 102015.1, 102021.5, 102018.6, 102006.7, 101989.2, 
    101964.5, 101933.6, 101893.4, 101846, 101797.5, 101745, 101689.4, 101636.4,
  100498.2, 101918.2, 101987.8, 102004.7, 102017.2, 102026.3, 102019.5, 
    102004.4, 101982.8, 101954.2, 101920.4, 101879.7, 101834.5, 101784.6, 
    101738.4,
  100558.5, 101573.7, 101943.8, 101959.4, 101983.4, 102006.5, 102015.3, 
    102019.6, 102015.9, 102000.3, 101978.9, 101950.3, 101915.6, 101875.7, 
    101832,
  100178.5, 101449.6, 101895.4, 101926.4, 101954.9, 101976.1, 102001.9, 
    102012.5, 102016.8, 102012.6, 101999.5, 101982.4, 101958.8, 101932.4, 
    101901.6,
  100127.7, 100807.1, 101682, 101875.6, 101907.8, 101926, 101949.5, 101970.2, 
    101991.3, 101996.9, 102000.5, 101999.3, 101987.9, 101970.4, 101945.8,
  99777.79, 99618.43, 100515.5, 101770.7, 101857.6, 101878.9, 101905.8, 
    101924.5, 101942.2, 101957.9, 101966.7, 101970.3, 101971.8, 101969.7, 
    101958,
  99690.3, 99011.13, 99018.18, 100761, 101800.2, 101809.2, 101824.4, 
    101856.4, 101877.5, 101899.9, 101920.2, 101943.1, 101954.6, 101957.5, 
    101952.1,
  99970.77, 99215.75, 99580.57, 100067.9, 101698.4, 101781.6, 101784.7, 
    101802.1, 101822.9, 101849.5, 101867.5, 101884.6, 101902.3, 101909, 
    101924.7,
  98806.85, 98614.73, 99847.31, 100176.8, 100756.1, 101719.7, 101751.9, 
    101760.7, 101812.5, 101843.5, 101866, 101901.2, 101905.6, 101921.4, 
    101930.6,
  98893.12, 97401.4, 97228.85, 98342.07, 100007.9, 100759.7, 101761.1, 
    101757.9, 101802.7, 101856.6, 101899.8, 101924.5, 101943.1, 101957.7, 
    101972.1,
  101801.9, 101877.5, 101908.1, 101926.9, 101938.6, 101947.1, 101948.9, 
    101945.7, 101933.5, 101917.6, 101895.2, 101873, 101843.5, 101817, 101781.5,
  100363.9, 101805.5, 101879, 101906.9, 101928.5, 101951.8, 101961.4, 
    101969.4, 101970.7, 101966.2, 101956.3, 101940.8, 101918.7, 101891.3, 
    101864.7,
  100443.5, 101468.8, 101846.2, 101874.5, 101900.6, 101934.1, 101956.8, 
    101984.3, 102002.2, 102007.9, 102007.3, 102000.2, 101988.3, 101969.2, 
    101944.5,
  100078.7, 101371.4, 101791.4, 101837.3, 101867, 101903, 101931.9, 101961.3, 
    101985.7, 102004.4, 102019.8, 102026.2, 102028.4, 102022, 102011.1,
  100007.9, 100694.8, 101585.4, 101783.5, 101812.5, 101844.9, 101874.1, 
    101910.5, 101941, 101969.8, 101996.4, 102019.7, 102037.3, 102046.9, 
    102046.3,
  99667.91, 99511.98, 100399.8, 101662.2, 101758.1, 101779.5, 101810.2, 
    101841.9, 101876, 101910, 101943, 101975.9, 102008.4, 102033.7, 102051,
  99516.41, 98912.62, 98916.7, 100634.2, 101681.1, 101711.1, 101738.4, 
    101770, 101802.4, 101834.7, 101875.1, 101913.4, 101950.1, 101987.9, 
    102017.1,
  99746.79, 99019.29, 99464.73, 99974.05, 101559.4, 101641.7, 101669.2, 
    101702.9, 101746.5, 101791, 101819.3, 101852.7, 101887.4, 101926.5, 
    101973.7,
  98604.83, 98389.8, 99657.16, 99987.13, 100595.6, 101572, 101617, 101662.6, 
    101711.7, 101771.2, 101802, 101838.5, 101861.2, 101882.7, 101913.3,
  98667.55, 97180.37, 97018.51, 98113.52, 99804.11, 100563.2, 101594.5, 
    101634.9, 101700.9, 101761.8, 101802.3, 101838.2, 101864.9, 101895.7, 
    101912.6,
  101487.1, 101592.7, 101670.5, 101741.1, 101803.7, 101877.3, 101947.9, 
    102017.6, 102077.5, 102129.6, 102166.7, 102197.9, 102220.6, 102235.3, 
    102231.6,
  100087.4, 101528, 101634.1, 101697.8, 101765.3, 101838.7, 101909.8, 
    101985.1, 102051.7, 102115, 102167.1, 102205.7, 102234.2, 102254.8, 
    102261.7,
  100167.6, 101198.8, 101597.6, 101663.9, 101724.3, 101791.8, 101860.2, 
    101935.6, 102005.4, 102076.1, 102139.1, 102189, 102232.4, 102268.6, 
    102285.6,
  99827.43, 101116.4, 101545.3, 101618.9, 101677.8, 101742.5, 101805.8, 
    101877.2, 101947.4, 102017.5, 102090.6, 102150.6, 102200.4, 102241.3, 
    102272.8,
  99780.17, 100455.4, 101357.4, 101573.5, 101634.3, 101694.9, 101760.4, 
    101823.1, 101887.2, 101948.9, 102014.6, 102091.9, 102154.7, 102207.3, 
    102248.8,
  99474.36, 99305.24, 100201.1, 101471.1, 101592.2, 101646.1, 101715.9, 
    101780.2, 101842, 101900.7, 101951.2, 102011.2, 102085.6, 102145.3, 
    102194.8,
  99370.8, 98751.2, 98732.22, 100463, 101542.4, 101607.3, 101672.2, 101741.1, 
    101804.3, 101856.7, 101914.9, 101957.7, 102010, 102068.4, 102125.7,
  99597.21, 98884.59, 99318.79, 99819.8, 101423.6, 101562.5, 101635.8, 
    101705.2, 101775.8, 101829.2, 101877, 101923.2, 101961.5, 102007, 102061.1,
  98415.85, 98260.52, 99534.09, 99866.21, 100492.6, 101480.9, 101598.9, 
    101665.3, 101738.6, 101798.1, 101849, 101895.3, 101932.3, 101971, 102008,
  98459.23, 97014.77, 96864.91, 98015.23, 99704.26, 100461.4, 101558.8, 
    101633.2, 101699, 101766.4, 101814.2, 101857.7, 101896.6, 101937.4, 
    101971.9,
  101088, 101217, 101342, 101439.7, 101538.3, 101645.9, 101757, 101866.5, 
    101980.9, 102097.6, 102207.4, 102309.2, 102404.4, 102487, 102554.8,
  99734.55, 101176.4, 101330.7, 101425.2, 101524, 101631.4, 101740.9, 101849, 
    101958.1, 102063.1, 102164.7, 102263, 102354.7, 102441.8, 102514.5,
  99851.93, 100875.2, 101311.9, 101412.1, 101512.2, 101617.1, 101724.2, 
    101829.3, 101933.9, 102031.9, 102131.3, 102225.6, 102311.9, 102396.2, 
    102469.1,
  99560.08, 100822.1, 101281.2, 101387.3, 101488.8, 101593.7, 101703.6, 
    101808.7, 101907.2, 101994.9, 102082.7, 102169.8, 102252.1, 102331.7, 
    102405.2,
  99547.4, 100218.5, 101114.3, 101369.7, 101467.7, 101570.5, 101680.9, 
    101782.9, 101880.7, 101965.5, 102040, 102117.4, 102195.2, 102267.4, 
    102332.8,
  99281.84, 99116.75, 100001.5, 101287.4, 101446.4, 101542.1, 101650.9, 
    101754, 101849.7, 101931.3, 101999.4, 102062.3, 102126.1, 102195, 102255.8,
  99220.41, 98599.38, 98588.85, 100316.3, 101419.6, 101520.5, 101622.8, 
    101724.7, 101819.7, 101898.2, 101961.4, 102017.7, 102063.6, 102116.9, 
    102170.8,
  99471.28, 98760.16, 99206.35, 99715.57, 101316.3, 101492, 101596.8, 
    101695.9, 101785.7, 101864.5, 101920.1, 101972, 102011.2, 102052.2, 
    102090.1,
  98318.32, 98160.12, 99438.73, 99801.91, 100441.1, 101430.8, 101577, 
    101667.3, 101755.9, 101833.7, 101882.9, 101927.9, 101962.3, 102000.5, 
    102030.6,
  98376.93, 96950.11, 96804.3, 97956.41, 99666.65, 100442.4, 101551.7, 
    101652.1, 101719.1, 101801.8, 101843.9, 101883.2, 101910.9, 101941.4, 
    101969.9,
  101051, 101146.3, 101241.1, 101342.2, 101445.5, 101551.8, 101660.8, 
    101768.1, 101867, 101960.7, 102055.4, 102136.4, 102211.4, 102270.2, 
    102317.7,
  99701.31, 101109.3, 101245.8, 101346.2, 101447.8, 101551.6, 101655.1, 
    101755.7, 101851, 101940.6, 102029.6, 102103, 102165.5, 102220.9, 102260.8,
  99830.67, 100830.8, 101243.2, 101334.3, 101437.4, 101538.1, 101641.9, 
    101741.2, 101834.4, 101919.1, 102000, 102067.9, 102118, 102154.3, 102179.1,
  99534.62, 100782.3, 101227.3, 101325.8, 101428.6, 101528.3, 101625.8, 
    101719.8, 101807.4, 101887, 101962.2, 102027.6, 102073.6, 102096.8, 
    102100.7,
  99525.31, 100184, 101073.1, 101316.4, 101411.4, 101507.4, 101606.4, 
    101697.8, 101782.7, 101858.2, 101926.4, 101986.1, 102028.2, 102039.1, 
    102027.8,
  99254.2, 99084.95, 99967.41, 101241.5, 101394, 101485.5, 101582.8, 
    101670.8, 101752.9, 101825.3, 101891.1, 101945.8, 101991.7, 101999.7, 
    101972.9,
  99184.3, 98573.38, 98558.59, 100277.6, 101370, 101462.9, 101558.4, 
    101643.8, 101727.8, 101796.1, 101857.9, 101908.5, 101945.1, 101965.5, 
    101939.4,
  99428.62, 98733.72, 99178.45, 99679.87, 101269.3, 101433.4, 101536.7, 
    101621.9, 101700.7, 101768.4, 101826.4, 101879.8, 101917.4, 101940.5, 
    101928.8,
  98275.1, 98130.82, 99404.38, 99769.48, 100395.8, 101369.4, 101510.3, 
    101599.8, 101675.5, 101745.1, 101795.2, 101847.8, 101889.9, 101921.2, 
    101926.2,
  98333.4, 96917, 96778.88, 97931.25, 99634.16, 100385.7, 101480.1, 101591.3, 
    101648.2, 101723.3, 101765.2, 101807, 101849.4, 101887.6, 101910.7,
  100970.2, 100968.1, 100976.9, 100992.7, 101010.6, 101039.1, 101078.4, 
    101130.3, 101193, 101265, 101342.6, 101402.7, 101441.5, 101462.1, 101482.2,
  99587.86, 100947.6, 100992.2, 100995.5, 101021.8, 101054.3, 101105.6, 
    101167.4, 101235.3, 101306.1, 101378.5, 101435.8, 101474.4, 101484.1, 
    101485.5,
  99683.16, 100650.6, 100992.9, 101008.9, 101033.4, 101071.1, 101127.1, 
    101188.3, 101257.5, 101334.4, 101407.5, 101469.9, 101502.9, 101500.8, 
    101485.5,
  99355.02, 100596.6, 100990.9, 101007.7, 101037.2, 101088.8, 101147.5, 
    101215.4, 101289.4, 101365.9, 101430.8, 101501.2, 101535.7, 101532.2, 
    101507.2,
  99313.94, 99974.17, 100828.9, 101021.1, 101050.7, 101097.3, 101159, 
    101230.2, 101304.7, 101382, 101452.9, 101521.8, 101568.6, 101568.9, 
    101545.3,
  99041.1, 98863.98, 99717.1, 100956.2, 101059.9, 101107.1, 101172.5, 
    101246.8, 101322, 101398.3, 101469.8, 101536.4, 101593.9, 101611.7, 
    101597.1,
  99013.84, 98378.81, 98329.62, 100020.8, 101073, 101123.4, 101185.8, 101258, 
    101334.7, 101410.6, 101482.8, 101542.2, 101604.1, 101648.6, 101661.5,
  99276.59, 98556.46, 98974.41, 99458.62, 101006.8, 101131.8, 101197.1, 
    101274.8, 101346, 101418.7, 101489.8, 101549.7, 101613.5, 101656.4, 
    101696.7,
  98142.14, 97987.3, 99228.24, 99568.97, 100167.7, 101104.2, 101208.9, 
    101284.2, 101356.4, 101430.8, 101494.8, 101552.2, 101614.5, 101668.5, 
    101719.6,
  98205.45, 96778.62, 96624.41, 97747.22, 99430.25, 100162.1, 101212.3, 
    101297.4, 101355.8, 101437.8, 101498.2, 101554.6, 101605.8, 101653.8, 
    101709.8,
  101584.2, 101575.2, 101545, 101481, 101400.3, 101328.2, 101263.1, 101210.1, 
    101155.8, 101097.3, 101036.2, 100975.9, 100920.3, 100871.1, 100834.4,
  100136.2, 101513.5, 101525.7, 101448.6, 101382.1, 101325.8, 101266.3, 
    101208.6, 101153, 101098.8, 101049, 101002.6, 100962.1, 100927.2, 100893.4,
  100206.1, 101187.9, 101495.8, 101425.1, 101367.5, 101306.4, 101244.4, 
    101202.5, 101162.5, 101109.1, 101059.5, 101012.1, 100975.5, 100945.2, 
    100921.2,
  99845.29, 101072.1, 101427.5, 101378.7, 101320.5, 101271.1, 101225.8, 
    101180.4, 101132.5, 101081.1, 101044.6, 101009.4, 100978.1, 100954.4, 
    100933,
  99759.21, 100406.6, 101221.6, 101345.2, 101283.8, 101226, 101175.1, 
    101133.4, 101103.2, 101070.5, 101039.8, 101009.1, 100987.8, 100972.1, 
    100958.3,
  99396.12, 99183.43, 100030.5, 101215.7, 101227.2, 101170.8, 101133.4, 
    101107.9, 101090.7, 101070.9, 101058.6, 101042, 101035.1, 101028.3, 
    101026.8,
  99241.53, 98564.3, 98503.7, 100191.6, 101173.9, 101138.4, 101099, 101084.8, 
    101079.6, 101079, 101071.8, 101070.7, 101075.3, 101081.6, 101094.7,
  99409.61, 98636.34, 99010.31, 99507.77, 101060.1, 101096.5, 101063.7, 
    101065.4, 101067.6, 101085, 101098.5, 101108.8, 101122.4, 101131.7, 
    101154.6,
  98169.37, 97987.32, 99227.75, 99550.88, 100112.2, 101007.5, 101027.8, 
    101033.1, 101057.5, 101089, 101105.2, 101131.9, 101149.3, 101175.7, 
    101214.8,
  98170.79, 96698.02, 96533.66, 97667.65, 99302.55, 100026.9, 100960.4, 
    100988.8, 101020.6, 101090.7, 101125.4, 101161.8, 101189.4, 101220, 
    101253.7,
  101778.1, 101797.8, 101778.3, 101730, 101657.8, 101572.6, 101486.1, 
    101396.8, 101305.4, 101213.1, 101125.5, 101043.1, 100965.9, 100896.6, 
    100837.7,
  100362.9, 101758.4, 101777.3, 101731, 101676.2, 101610.3, 101535.9, 
    101460.8, 101383.8, 101303.9, 101225.9, 101151.1, 101080.9, 101016.6, 
    100958.9,
  100458.4, 101441.7, 101770.5, 101730.6, 101680, 101624.9, 101564, 101502.2, 
    101440.7, 101375.5, 101309.4, 101244.2, 101179.2, 101116, 101057.8,
  100122, 101378.5, 101737.5, 101719.1, 101673, 101627.2, 101575.9, 101525.8, 
    101475, 101423.1, 101365.9, 101308.1, 101249.2, 101195.2, 101140.8,
  100042.6, 100714, 101543.2, 101694.6, 101656.3, 101617, 101572.5, 101531.4, 
    101488.8, 101445.7, 101396.9, 101347.3, 101295.8, 101247.2, 101200.2,
  99709.84, 99510.34, 100383.9, 101596.9, 101632.9, 101591.1, 101557.5, 
    101521.7, 101484.7, 101446.8, 101405.9, 101360.9, 101318.7, 101276.1, 
    101232.2,
  99560.12, 98900.19, 98844.64, 100576.3, 101580.2, 101556.7, 101517.8, 
    101482.9, 101452.9, 101423.8, 101390.4, 101349.7, 101311, 101272.5, 
    101235.1,
  99750.94, 99023.47, 99420.84, 99913.7, 101464, 101511.2, 101469.7, 
    101436.2, 101401, 101371, 101339.7, 101308.6, 101286.8, 101257, 101221,
  98509.94, 98363.19, 99626.35, 99945.66, 100523.3, 101422.4, 101417.5, 
    101364.9, 101330.3, 101307.8, 101285.3, 101261.2, 101231.1, 101192.2, 
    101172.2,
  98481.94, 97022.27, 96882.77, 98054.7, 99703.4, 100438.7, 101357.6, 
    101312.1, 101235.9, 101230.8, 101197, 101188.6, 101178.9, 101181.2, 
    101162.5,
  102123.1, 102153.8, 102100, 101991.8, 101880.6, 101783.5, 101682.8, 
    101572.5, 101463.4, 101336.8, 101209.1, 101072.1, 100935.1, 100818.6, 
    100730.8,
  100680, 102076.2, 102092.9, 102010.4, 101904.9, 101803.3, 101698.8, 
    101593.1, 101486, 101370.2, 101252.5, 101135.8, 101020.1, 100919.4, 
    100838.8,
  100747.7, 101752.1, 102089.4, 102023.4, 101924, 101826.5, 101729, 101630.5, 
    101534.2, 101431.1, 101324.1, 101217.4, 101111, 101012.8, 100930.5,
  100422.5, 101669.4, 102051.6, 102020.7, 101936, 101848.1, 101753.6, 
    101658.6, 101566.3, 101472.7, 101375, 101279.9, 101185.8, 101098.5, 
    101024.2,
  100358.4, 101014, 101852.3, 102009.5, 101939.1, 101859.4, 101776, 101688, 
    101602.1, 101518, 101428.8, 101341.1, 101254.8, 101172.1, 101096.3,
  100047.8, 99829.91, 100690.9, 101912.7, 101935.1, 101869.8, 101794.7, 
    101713.1, 101630.5, 101548, 101466.8, 101384.4, 101304.9, 101231.1, 
    101163.4,
  99905.55, 99239.37, 99161.7, 100903.3, 101906, 101865.4, 101799.9, 
    101729.8, 101653.9, 101578.1, 101499.9, 101424.4, 101349.8, 101277.6, 
    101204.5,
  100110, 99374.97, 99767.98, 100257, 101819.4, 101864.2, 101802.4, 101742.1, 
    101667.7, 101597.6, 101523.9, 101447, 101373, 101304.6, 101242.6,
  98853.67, 98692.91, 99973.92, 100307.3, 100901.6, 101799.7, 101795.3, 
    101733.2, 101671.6, 101606.4, 101533.7, 101461.7, 101388.7, 101318.4, 
    101240.4,
  98825.69, 97362.5, 97231.09, 98412.02, 100083.8, 100840.1, 101782.4, 
    101749.9, 101663.2, 101613.1, 101531.4, 101463.6, 101381.2, 101302.8, 
    101241.1,
  102315.1, 102302.3, 102267.1, 102214.6, 102167.8, 102100.7, 102022.7, 
    101928.2, 101818.6, 101688, 101534, 101350.9, 101165.1, 100984.1, 100834.9,
  100869.2, 102266.3, 102261.7, 102191.2, 102144.3, 102085.9, 102004.5, 
    101914.1, 101800.7, 101666.8, 101516.4, 101338, 101148.2, 100972, 100824.4,
  100943, 101934.3, 102250.1, 102177.3, 102122.9, 102065.1, 101991.5, 
    101909.3, 101805.6, 101684.4, 101543.4, 101377, 101191.3, 101014, 100857,
  100616.1, 101878.4, 102231.4, 102176.6, 102106.8, 102052.6, 101982.4, 
    101906.4, 101811.7, 101696, 101562.8, 101409.4, 101236.5, 101068, 100910.4,
  100553.7, 101219.5, 102060.3, 102172.5, 102105.8, 102043.7, 101978.2, 
    101906.2, 101822.7, 101722, 101600.8, 101466.6, 101308.4, 101148.4, 
    100997.8,
  100246.5, 100035.7, 100914.4, 102110, 102108.2, 102046.8, 101982.8, 
    101912.8, 101833.7, 101742.6, 101631.5, 101509, 101371.8, 101227.7, 101085,
  100119.2, 99454.41, 99378.12, 101124, 102100.1, 102048.4, 101983.6, 
    101920.2, 101846, 101763.8, 101668.1, 101557.4, 101437.5, 101311.5, 
    101181.9,
  100341, 99600.07, 99990.66, 100486.5, 102045.5, 102064, 101996.3, 101932.5, 
    101859.4, 101783.4, 101697.1, 101597, 101491, 101379.1, 101264.7,
  99087.24, 98936.91, 100225.3, 100553.7, 101147.8, 102028.1, 102005.6, 
    101937.5, 101872, 101804.8, 101723.1, 101638.5, 101541.8, 101444.1, 
    101342.7,
  99066.3, 97591.97, 97465.05, 98651.73, 100335.6, 101102.3, 102015.4, 
    101976.1, 101880.8, 101829.2, 101746.7, 101670.5, 101583.5, 101497, 
    101408.3,
  102194.9, 102251.4, 102270.5, 102264.6, 102231.9, 102207.2, 102172.6, 
    102133.2, 102068.6, 101967.7, 101840.5, 101699.8, 101551.8, 101436.4, 
    101357.6,
  100742.8, 102204, 102259.2, 102243.5, 102228.2, 102208.2, 102162.6, 
    102123.4, 102063.3, 101973.2, 101850.7, 101713, 101563.7, 101438, 101335.3,
  100830.4, 101873.2, 102243.8, 102233.7, 102211.4, 102195.2, 102160.4, 
    102124, 102073, 101996.9, 101889.2, 101751.8, 101591.9, 101438.3, 101305.7,
  100496.3, 101798.4, 102201.8, 102225.4, 102207.9, 102186.7, 102155.2, 
    102121.8, 102078.1, 102011.3, 101917.3, 101797.5, 101644.9, 101486.6, 
    101338.3,
  100451.4, 101131.3, 102021.2, 102191.3, 102192.8, 102178.2, 102150.1, 
    102115.9, 102080.6, 102027.8, 101944.2, 101842.5, 101704.6, 101546.3, 
    101384.3,
  100141.8, 99945.81, 100845, 102120.3, 102189.4, 102175.9, 102153.9, 
    102124.4, 102083.7, 102036, 101966.9, 101877.3, 101759.2, 101617.7, 
    101461.1,
  100010.4, 99381.44, 99323.34, 101094, 102144.3, 102163, 102143.4, 102120.9, 
    102085.8, 102047, 101983.2, 101910.2, 101810.1, 101682.6, 101538.2,
  100220.5, 99515.85, 99950.12, 100456.8, 102059.1, 102147.9, 102139.9, 
    102125.7, 102091.3, 102052.3, 102000.1, 101932, 101851.6, 101739.1, 
    101613.4,
  98967.32, 98830.59, 100153.1, 100523.6, 101142.6, 102084, 102129.3, 
    102121.1, 102095.9, 102062.9, 102014.2, 101955.9, 101884.1, 101793.9, 
    101677.3,
  98964.74, 97503.95, 97385.71, 98598.14, 100338.3, 101131.8, 102119.4, 
    102129.2, 102092.1, 102073.3, 102024, 101973.8, 101906.1, 101832.7, 101740,
  101933.8, 102042, 102099.8, 102147.2, 102184.7, 102232.9, 102262.1, 
    102284.1, 102246.3, 102208.6, 102204.2, 102255.8, 102306.8, 102340.6, 
    102349.5,
  100507.2, 101982.3, 102083.9, 102133.3, 102169.7, 102222.5, 102252.7, 
    102266.6, 102243.9, 102211.5, 102205.5, 102218.9, 102253.7, 102282.4, 
    102313.5,
  100601.9, 101657.4, 102059.9, 102113.9, 102155.5, 102210.8, 102250.5, 
    102275.8, 102260.1, 102214.4, 102182.6, 102177.8, 102211.9, 102246.3, 
    102251.1,
  100267.3, 101582.9, 102023.9, 102099.4, 102147.5, 102192.8, 102233.2, 
    102275.4, 102269.7, 102236.9, 102187.1, 102159.6, 102154.6, 102190.7, 
    102207.3,
  100230.6, 100928.2, 101843, 102072.9, 102129.7, 102176.7, 102212.8, 
    102251.8, 102276.1, 102253.9, 102199.9, 102155.7, 102122.8, 102136.2, 
    102153.6,
  99925.59, 99762.03, 100689.3, 101990, 102114.7, 102159.1, 102197.2, 
    102243.6, 102276.3, 102261.5, 102224, 102164.6, 102120, 102101.9, 102114.8,
  99822.5, 99201.03, 99194.35, 100985.3, 102082.6, 102140.5, 102181.3, 
    102215.3, 102254.4, 102266.7, 102236.1, 102182.9, 102129.2, 102083.9, 
    102079.2,
  100046, 99342.13, 99813.12, 100339.9, 101985.9, 102116.5, 102164.1, 
    102200.3, 102227.6, 102251.4, 102246, 102204, 102147.9, 102091.7, 102053.8,
  98832.13, 98691.58, 100015.4, 100393.3, 101059.7, 102057.5, 102153.1, 
    102184, 102212.8, 102236.8, 102244.5, 102218.1, 102170.2, 102111.2, 
    102055.7,
  98862.75, 97409.41, 97287.34, 98489.23, 100236.2, 101035.4, 102122, 
    102177.5, 102199.6, 102221.9, 102229.1, 102226.3, 102185.6, 102134.7, 
    102073.6,
  101713.1, 101767.3, 101831.3, 101897.8, 101955.9, 102030.8, 102109.9, 
    102195.9, 102269, 102319.2, 102364.7, 102448.4, 102547.4, 102610.7, 102676,
  100335.3, 101757.5, 101863.3, 101919.6, 101974.4, 102044, 102131.4, 
    102218.8, 102292.6, 102335.1, 102388.6, 102440, 102538.1, 102588.5, 
    102657.5,
  100468.7, 101486.2, 101882.9, 101939.7, 102001.6, 102065.3, 102144.7, 
    102229.8, 102307.6, 102355.6, 102392.6, 102430, 102531.9, 102580, 102633.8,
  100177.1, 101444.3, 101877.1, 101942.4, 102012.7, 102074.5, 102153.8, 
    102239.3, 102315.1, 102368.3, 102391.2, 102430.9, 102502.9, 102580.8, 
    102609.1,
  100177.2, 100840.9, 101733.4, 101955.3, 102020, 102084.9, 102156.4, 
    102239.9, 102317, 102375.3, 102397.8, 102422.9, 102465.9, 102563.3, 
    102591.2,
  99898.67, 99712.53, 100597, 101896.3, 102025.1, 102086.4, 102157.9, 
    102235.1, 102316.7, 102376.7, 102405.3, 102420.7, 102459, 102532.7, 
    102582.8,
  99829.7, 99184.95, 99163.05, 100910.1, 102029.8, 102088.6, 102154.2, 
    102220.6, 102306.8, 102370.9, 102408.1, 102412.8, 102444.9, 102486.7, 
    102567.9,
  100075.4, 99346.95, 99792.73, 100304.7, 101938.2, 102082.4, 102153, 
    102217.8, 102291, 102368.4, 102404.7, 102415.4, 102431.9, 102461, 102532.3,
  98889.7, 98725.8, 100026.3, 100403.6, 101052.1, 102043.9, 102148.6, 102203, 
    102277.7, 102361.2, 102405, 102426.1, 102424.9, 102446.7, 102479.7,
  98941.2, 97478.39, 97333.26, 98506.07, 100266.1, 101023.1, 102136, 
    102202.3, 102251.1, 102344.4, 102398.4, 102423.7, 102419.2, 102435.5, 
    102456.8,
  101525.7, 101455, 101400.3, 101334.5, 101280.9, 101243.4, 101228.5, 
    101228.7, 101262, 101312.1, 101413.5, 101522.2, 101661.5, 101818.4, 101985,
  100174.5, 101464.5, 101462.5, 101406.8, 101363.5, 101325.7, 101310.6, 
    101312.7, 101348.6, 101403.5, 101478, 101566, 101687.3, 101840.7, 101998,
  100318.9, 101230.3, 101527.4, 101477.4, 101434.6, 101404.6, 101392.2, 
    101395.5, 101427.8, 101480.1, 101547.4, 101634.3, 101742.5, 101882.6, 
    102017.3,
  100062.1, 101217.7, 101564.4, 101537, 101504.6, 101482.3, 101473.6, 101483, 
    101511.9, 101569.5, 101623.8, 101705.3, 101793.4, 101916.9, 102045.6,
  100076.8, 100643.8, 101452.6, 101590.2, 101564.6, 101543.8, 101547.2, 
    101554.2, 101584.3, 101644.9, 101702.9, 101774.3, 101857.3, 101965.5, 
    102082.5,
  99821.42, 99558.23, 100368.3, 101587.5, 101630.7, 101608.7, 101609.8, 
    101627, 101657.2, 101718.9, 101774.4, 101839.9, 101919.4, 102012.1, 
    102119.3,
  99763.82, 99055.29, 98951.55, 100635.6, 101666.8, 101666.1, 101661.5, 
    101681.9, 101716.7, 101781.3, 101839.6, 101907.6, 101977.9, 102054.4, 
    102157.7,
  100046.8, 99247.94, 99615.14, 100075.9, 101621.8, 101710.5, 101714.8, 
    101747.2, 101782.6, 101844.6, 101900.2, 101961.5, 102025.1, 102099.9, 
    102192.2,
  98865.11, 98652.41, 99883.27, 100211.3, 100780.5, 101710.8, 101757.8, 
    101793.2, 101839.4, 101901, 101958.9, 102016.3, 102073.6, 102140.5, 102220,
  98940.77, 97448.15, 97260.09, 98370.85, 100045, 100781.5, 101814, 101869.9, 
    101882.4, 101956.4, 102008.9, 102061.9, 102111.6, 102172.5, 102239.4,
  101323.1, 101256.3, 101193.2, 101082.7, 100943.1, 100796.1, 100661.4, 
    100551.6, 100456.5, 100383.9, 100349.6, 100351.8, 100382.6, 100430.8, 
    100482.4,
  99984.71, 101290.5, 101266.8, 101164.2, 101059.5, 100946, 100825.7, 
    100713.8, 100618.9, 100540.6, 100494.3, 100476.1, 100486, 100507.3, 
    100549.2,
  100134.1, 101075.3, 101360, 101268.5, 101163.5, 101061.7, 100960.6, 
    100863.4, 100775.5, 100708, 100654.1, 100614.8, 100602.1, 100601.2, 
    100625.9,
  99894.61, 101082.7, 101417, 101358.9, 101270.3, 101171, 101083.5, 100997.3, 
    100916.2, 100844.9, 100785.7, 100740.3, 100716.9, 100703.2, 100713.6,
  99916.95, 100518.7, 101327.9, 101432.8, 101362.4, 101281.7, 101195.8, 
    101113.8, 101036.2, 100968.5, 100910.6, 100870.1, 100830.6, 100804, 
    100802.9,
  99679.63, 99423.52, 100241.3, 101439.6, 101439.1, 101363.6, 101292.1, 
    101219, 101147.1, 101081.9, 101028.3, 100983.7, 100947.5, 100923.8, 
    100924.2,
  99611.18, 98912.45, 98801.78, 100489.9, 101495.7, 101444.8, 101372.8, 
    101307.1, 101238.7, 101179.8, 101129.6, 101085.7, 101050.2, 101030.1, 
    101023,
  99896.81, 99112.89, 99465.55, 99919.41, 101460.1, 101505.9, 101440.9, 
    101391.6, 101331.3, 101276.5, 101225.1, 101186.4, 101158.9, 101139.6, 
    101136.5,
  98683.25, 98485.88, 99732.92, 100065.5, 100621.5, 101509.4, 101492.3, 
    101436.6, 101390.4, 101347.4, 101309.2, 101279.9, 101254.8, 101247.5, 
    101248.9,
  98728.83, 97226.79, 97042.1, 98172.03, 99833.33, 100583.3, 101561, 
    101523.8, 101448.3, 101428, 101380.1, 101364.3, 101349.1, 101352, 101365.4,
  100752.8, 100805.4, 100859.1, 100914.5, 100956.9, 100928.1, 100877.1, 
    100815, 100750.9, 100672.2, 100598.4, 100532.8, 100462.1, 100394.5, 
    100330.4,
  99296.35, 100724.8, 100789.1, 100798.8, 100830, 100872.3, 100896.2, 
    100875.6, 100827.5, 100758.4, 100685.1, 100610.7, 100527.2, 100452.4, 
    100388,
  99388.59, 100379.4, 100697.8, 100692.7, 100764.8, 100825.7, 100881.3, 
    100904.5, 100893.9, 100864.6, 100806.8, 100736.6, 100655.6, 100569.7, 
    100493.9,
  99070.61, 100261.3, 100602.2, 100542, 100608.7, 100721.7, 100816.4, 
    100878.7, 100912.8, 100925.8, 100906.4, 100863.7, 100796.2, 100719, 
    100643.2,
  99060.34, 99653.69, 100431, 100501.8, 100533.1, 100645.9, 100763.5, 
    100845.8, 100908.3, 100955, 100971.3, 100964.4, 100930.2, 100874.9, 100807,
  98788.7, 98526.05, 99313.8, 100506.8, 100592.1, 100654.9, 100733.2, 
    100816.6, 100898.7, 100970.2, 101007.5, 101022.4, 101016.6, 100989.3, 
    100948.3,
  98720.01, 98011.15, 97907.02, 99587.09, 100630.1, 100673.5, 100733.4, 
    100814.4, 100898.2, 100981.8, 101040.6, 101074.4, 101082.9, 101076.4, 
    101056.9,
  99006.1, 98211.91, 98581.91, 99040.92, 100585.9, 100697.4, 100747.1, 
    100824.8, 100907.3, 100992.8, 101057, 101106.7, 101130.7, 101137.6, 101134,
  97847.44, 97614.5, 98833.2, 99173.45, 99763.1, 100684.8, 100768.8, 
    100845.3, 100934.9, 101024.5, 101092.6, 101146.8, 101177.6, 101197.4, 
    101201.7,
  97943.91, 96435.85, 96228.7, 97326.3, 98996.76, 99735.11, 100807.1, 100892, 
    100954.5, 101057.4, 101124.6, 101185.2, 101219.8, 101245.9, 101258,
  100113.7, 100060.7, 100053.3, 100085.7, 100153.9, 100236.4, 100377.6, 
    100557.3, 100720.7, 100867.6, 100973, 101070.1, 101153.7, 101223.4, 
    101271.9,
  98473.77, 99769.23, 99791.98, 99864.82, 99947.13, 100047.8, 100185.1, 
    100345.1, 100496.7, 100639.5, 100787.7, 100921.3, 101030.4, 101124.8, 
    101194.9,
  98376.46, 99331.47, 99611.84, 99721.31, 99790.67, 99915.77, 99981.77, 
    100123.7, 100281.7, 100435.4, 100594.3, 100756.4, 100892.8, 101011.4, 
    101100.4,
  98091, 99336.88, 99602.75, 99658.51, 99744.88, 99870.75, 99909.6, 100036.1, 
    100122.9, 100266.9, 100417.5, 100602.8, 100772.5, 100911.9, 101019,
  98143.6, 98815.19, 99574.2, 99771.6, 99790.73, 99890.3, 99914.69, 99980.3, 
    100058.2, 100131.8, 100256.6, 100443.6, 100623.5, 100813.2, 100958.5,
  98054.24, 97781.38, 98590.58, 99835.23, 99916.02, 99957.88, 99981.59, 
    100016.8, 100019.9, 100106.1, 100172, 100319.8, 100489.2, 100673.3, 
    100860.8,
  98205.02, 97390.43, 97246.54, 98966.12, 100027.5, 100052.2, 100049.6, 
    100075.3, 100075, 100117.2, 100172.1, 100265.9, 100409.9, 100569.5, 
    100761.6,
  98711.05, 97784.21, 98055.39, 98499.7, 100081, 100174, 100155.8, 100147.1, 
    100149.7, 100152.9, 100207.4, 100271, 100375.3, 100518.3, 100689,
  97727.66, 97344.8, 98489.63, 98768.38, 99340.39, 100263.4, 100271.3, 
    100233, 100225.6, 100222, 100253.6, 100299, 100382, 100493.2, 100648.9,
  97990.15, 96296.13, 95975.84, 97008.36, 98671.59, 99415.79, 100410.8, 
    100367.9, 100309.7, 100306.3, 100311.3, 100342.7, 100412.8, 100493.7, 
    100624.5,
  100748.9, 100630.9, 100502.5, 100369.9, 100287.4, 100228, 100183.6, 
    100186.7, 100174, 100162.8, 100137.7, 100100.2, 100050.7, 100052.8, 
    100079.7,
  99320.95, 100583.3, 100524.7, 100403.4, 100325.8, 100260.8, 100164.9, 
    100155.3, 100134.9, 100120, 100084.7, 100031.8, 100002.2, 100009, 100046.8,
  99376.8, 100292.2, 100516.8, 100361.1, 100281, 100239.7, 100213.1, 
    100205.6, 100184.1, 100162.7, 100135.8, 100093.5, 100062.6, 100055.2, 
    100075.4,
  99106.48, 100244.7, 100491.5, 100394, 100313, 100265.2, 100220.1, 100206.5, 
    100199, 100179.7, 100159.4, 100132.6, 100105.5, 100091.9, 100118.8,
  99113.3, 99641.66, 100357.7, 100424.2, 100320.3, 100270.4, 100254.8, 
    100264.3, 100258.4, 100250.8, 100245.9, 100210.4, 100205.3, 100182.1, 
    100199.3,
  98890.34, 98542.32, 99286.12, 100379.3, 100328.9, 100267.3, 100252.4, 
    100261.1, 100264.8, 100271, 100276.7, 100264.9, 100275.8, 100263.5, 
    100272.6,
  98865.53, 98049.01, 97849.72, 99463.78, 100360.9, 100299, 100266.7, 100266, 
    100280.2, 100298.1, 100320.2, 100319.4, 100330.2, 100341.5, 100338.7,
  99225.45, 98325.94, 98535.51, 98915.84, 100350.8, 100333.1, 100281.2, 
    100270.4, 100279.9, 100297.5, 100330.5, 100350.2, 100371.1, 100397.6, 
    100408,
  98117.52, 97803.01, 98927.96, 99125.89, 99600.38, 100407, 100349.9, 
    100292.2, 100297.9, 100311.9, 100348.6, 100371.8, 100404.3, 100436.6, 
    100456.1,
  98248.57, 96633.95, 96334.34, 97360.83, 98907.91, 99599.52, 100471, 
    100419.8, 100329.5, 100351.7, 100372.4, 100401.3, 100431.4, 100475.6, 
    100493.9,
  101565.6, 101543.2, 101526.6, 101480.6, 101417.6, 101361.2, 101304.6, 
    101249, 101203, 101154.1, 101106.1, 101055.5, 101009.1, 100960.8, 100916.4,
  100227.9, 101564.6, 101592.4, 101538.6, 101477.2, 101415, 101355.9, 
    101300.4, 101248.6, 101198.2, 101149.1, 101102.6, 101058.2, 101011, 
    100964.7,
  100367.4, 101330.2, 101652, 101594.8, 101527.4, 101459.2, 101398.8, 
    101340.9, 101289.4, 101242.6, 101194, 101150.6, 101102.2, 101056.7, 
    101006.2,
  100127.2, 101336.8, 101691.9, 101655.4, 101577.8, 101502.4, 101435.9, 
    101371.8, 101318.9, 101274.3, 101227.9, 101185, 101144.4, 101101.2, 
    101057.6,
  100152.5, 100766.2, 101573.5, 101698.7, 101628.4, 101541.5, 101463.6, 
    101398.2, 101342.6, 101298, 101253.4, 101210.7, 101168.9, 101129.2, 
    101089.9,
  99911.36, 99661.69, 100484.8, 101669.7, 101673.9, 101577.9, 101489.6, 
    101427.3, 101369.2, 101320.9, 101271.9, 101225.7, 101185.8, 101150, 
    101117.3,
  99860.15, 99149.25, 99033.7, 100717.1, 101707.4, 101626.3, 101521.3, 
    101446.1, 101389.2, 101335.3, 101281.9, 101234.7, 101194, 101160.3, 
    101131.3,
  100149.6, 99356.91, 99699.11, 100150.2, 101685.5, 101672.8, 101556.7, 
    101479.9, 101408.6, 101348.2, 101294.5, 101241.5, 101201.1, 101163.4, 
    101139.2,
  98962.1, 98758.56, 99994.33, 100288, 100854.8, 101716.2, 101616.8, 101497, 
    101427.5, 101362.5, 101299.4, 101249.9, 101196.1, 101164.1, 101141.5,
  99021.88, 97488.12, 97316.48, 98439.9, 100075.9, 100802.2, 101710.1, 
    101595.3, 101444.7, 101387.8, 101309.6, 101254.2, 101199, 101163.7, 
    101144.9,
  101865.3, 101867, 101858.8, 101836.5, 101805.5, 101772, 101741.6, 101707.5, 
    101676.7, 101645.9, 101615.9, 101588.8, 101565.9, 101540.5, 101516.6,
  100506.7, 101866.2, 101929.7, 101911, 101884.6, 101847.2, 101818.6, 
    101789.9, 101766.1, 101743, 101721.4, 101698.7, 101674.5, 101652.9, 
    101631.4,
  100651.6, 101633.7, 101994.6, 101980.2, 101958.6, 101932.8, 101905.7, 
    101881.4, 101859.1, 101839.9, 101821.9, 101802.8, 101782.1, 101759.3, 
    101737.6,
  100390.2, 101621.6, 102027.8, 102035.4, 102018.9, 102000.6, 101975.9, 
    101956.5, 101938.5, 101924.4, 101911.3, 101895.9, 101879.7, 101860, 
    101838.4,
  100401.6, 101043.4, 101910.5, 102089.8, 102077.6, 102059.9, 102045.2, 
    102030.6, 102016, 102003.4, 101991.6, 101980.5, 101968.5, 101951.7, 
    101933.2,
  100134.8, 99918.76, 100777, 102036.5, 102119.6, 102108.2, 102099.7, 
    102090.8, 102079.6, 102071.9, 102059.2, 102051.3, 102040.1, 102029.2, 
    102012.5,
  100072.5, 99396.06, 99342.45, 101064.1, 102148.4, 102158.5, 102151.6, 
    102146.7, 102139.5, 102132.5, 102121.8, 102114.5, 102102.6, 102091.6, 
    102076.4,
  100310.9, 99557.85, 99987.48, 100482.3, 102082.5, 102180.7, 102188.4, 
    102188.4, 102186.2, 102179, 102173, 102163, 102157.4, 102141.2, 102129.4,
  99109.68, 98932.84, 100218.2, 100570.6, 101204.8, 102172.7, 102227.5, 
    102223.3, 102226.4, 102219, 102212.1, 102202, 102197.5, 102185.1, 102171.4,
  99151.21, 97669.95, 97510.26, 98674.4, 100407, 101152.2, 102240, 102255.8, 
    102243.9, 102249.2, 102237.7, 102235.3, 102234.3, 102215.5, 102193.2,
  102164.9, 102160.6, 102143.2, 102107.5, 102055.3, 102014.6, 101969.3, 
    101918.3, 101869.2, 101816.5, 101762.5, 101714.5, 101667.3, 101626.4, 
    101588.2,
  100749.4, 102117.1, 102158.8, 102129.2, 102087.2, 102044.3, 102009.4, 
    101970, 101928.4, 101882.4, 101836.8, 101792.8, 101751.2, 101709.2, 
    101673.6,
  100854, 101833.2, 102183.6, 102159.6, 102126, 102084.8, 102054, 102021.5, 
    101988.7, 101954.7, 101918.6, 101880.7, 101842.4, 101806.8, 101769.1,
  100555.3, 101783.4, 102176.5, 102175.3, 102151.9, 102118.9, 102090.5, 
    102064.6, 102039.8, 102014.9, 101986, 101957.1, 101926.1, 101895.8, 
    101864.5,
  100530.3, 101161.7, 102025.4, 102191.2, 102177.2, 102145.3, 102125.3, 
    102106.7, 102090.9, 102073, 102053.7, 102029.6, 102006.6, 101981.2, 
    101957.5,
  100240.7, 100021.5, 100871.4, 102122, 102187.6, 102161, 102147, 102136, 
    102127.9, 102117.7, 102109.4, 102094.3, 102078.5, 102062.2, 102046.9,
  100142.9, 99470.06, 99403.64, 101117.8, 102185.4, 102175.8, 102164.4, 
    102163.1, 102162.2, 102161.4, 102157.5, 102151.1, 102147.3, 102142.6, 
    102129.9,
  100384.9, 99613.27, 100014.6, 100498.1, 102079, 102163.3, 102166.2, 
    102171.3, 102180.1, 102190.1, 102197.9, 102203.7, 102207.2, 102203.2, 
    102196.3,
  99171.26, 98978.76, 100243, 100575.9, 101178.7, 102121.4, 102163.7, 102171, 
    102199.7, 102215.8, 102227.1, 102241.7, 102250.1, 102259.2, 102261.4,
  99220.04, 97726.09, 97551.36, 98689.17, 100396.6, 101130.7, 102161.6, 
    102183.2, 102197, 102231.7, 102249.5, 102268.6, 102289.7, 102308.1, 
    102308.6,
  102472.2, 102495.7, 102504.3, 102483.5, 102440.1, 102412.2, 102382.8, 
    102337.4, 102290.4, 102230.1, 102164.4, 102091.2, 102014.1, 101928.7, 
    101839.1,
  101040.4, 102462.6, 102517.3, 102497.2, 102451.6, 102432.4, 102409.4, 
    102379.8, 102342.9, 102295.1, 102238, 102175, 102109.1, 102032.4, 101950.6,
  101129.4, 102145.4, 102506.8, 102497.5, 102465.6, 102443.3, 102430.6, 
    102410.9, 102383.3, 102347.7, 102300.2, 102246.2, 102185.2, 102118.6, 
    102046.7,
  100796.7, 102076.9, 102481.4, 102500.4, 102475.6, 102441.6, 102431, 
    102417.9, 102402, 102377.5, 102341, 102297.3, 102247.4, 102187.6, 102124.6,
  100741.8, 101426.1, 102304.9, 102491.2, 102466.1, 102426.3, 102419.2, 
    102420, 102402.9, 102389.2, 102363.9, 102326.9, 102284.6, 102235.3, 
    102180.8,
  100428.7, 100238.3, 101123, 102410.4, 102453.7, 102422.8, 102408.4, 
    102399.2, 102393.5, 102383.5, 102366.2, 102342.5, 102310.4, 102270, 
    102224.2,
  100316.4, 99666.29, 99606.33, 101376.2, 102435.7, 102418.1, 102396.7, 
    102387.4, 102378.4, 102376.3, 102363.6, 102343.1, 102318.3, 102290.7, 
    102253.2,
  100547.1, 99809.22, 100226.4, 100739.8, 102347.4, 102404.5, 102389.1, 
    102375.6, 102367.9, 102364.5, 102353.6, 102340.8, 102324, 102298.3, 
    102268.9,
  99313.55, 99147.48, 100453, 100785.6, 101409.8, 102353.3, 102376.1, 
    102357.2, 102351.9, 102348, 102337.9, 102327.2, 102318, 102302.4, 102282.1,
  99325.14, 97837.75, 97694.23, 98891.05, 100607, 101367.6, 102359.7, 
    102354.9, 102331.4, 102333.5, 102327.5, 102323.7, 102309.8, 102299.8, 
    102288.5,
  102436.7, 102530.1, 102574.9, 102595, 102601.4, 102595, 102590.1, 102577.6, 
    102555.6, 102522.4, 102475.3, 102422.8, 102363.2, 102297.9, 102234.2,
  101039.5, 102494, 102579.3, 102607, 102630.5, 102621.4, 102625.8, 102622.7, 
    102611.6, 102589.5, 102553, 102507.5, 102454.4, 102394.1, 102329.5,
  101145.1, 102186.3, 102585.1, 102615.6, 102655.3, 102644.6, 102657.9, 
    102662.2, 102659.3, 102645, 102620.2, 102585.9, 102540.9, 102488.2, 
    102427.2,
  100818.9, 102117.7, 102554.7, 102609.3, 102650.8, 102650.5, 102678.1, 
    102694.6, 102698.6, 102694.2, 102677.2, 102649.4, 102614.4, 102570.1, 
    102516.3,
  100779.3, 101469.8, 102376.9, 102592.7, 102630.5, 102650.6, 102681.9, 
    102718.6, 102734.1, 102737.1, 102725.5, 102704, 102674.3, 102639.7, 
    102595.1,
  100464.9, 100290.9, 101196.7, 102494.2, 102596.2, 102627.3, 102658.3, 
    102712.9, 102731.7, 102756.4, 102759.3, 102744.4, 102721.4, 102692.2, 
    102658.4,
  100353.2, 99725.7, 99705.45, 101475.9, 102561.7, 102599.9, 102627.3, 
    102687, 102723.4, 102746.2, 102755.1, 102754.1, 102744.9, 102729.1, 
    102702.3,
  100556.5, 99850.83, 100309.1, 100834.3, 102454.6, 102565.1, 102597.6, 
    102642.9, 102700.3, 102732, 102751.3, 102754.4, 102753.6, 102745.6, 
    102729.2,
  99330.56, 99189.34, 100507.8, 100875, 101536.4, 102516.6, 102579.8, 
    102608.8, 102647.5, 102684.8, 102718.8, 102748.3, 102745.5, 102748, 
    102740.1,
  99327.8, 97877.21, 97750.21, 98964.04, 100701.1, 101489.4, 102549.2, 
    102588.6, 102613.8, 102647.2, 102668.8, 102697.6, 102721.8, 102739.4, 
    102734.7,
  102102.7, 102203.9, 102271.6, 102314.7, 102363.9, 102384.3, 102427.7, 
    102468.5, 102511, 102541.4, 102564, 102574.7, 102578.7, 102577.5, 102571.3,
  100743.1, 102179.9, 102293.6, 102350.5, 102413.3, 102441.9, 102494, 
    102545.3, 102596.1, 102632.8, 102659.9, 102676.2, 102687.1, 102690.5, 
    102685.5,
  100876.1, 101908.6, 102322.8, 102382, 102447, 102487.6, 102547.5, 102605.5, 
    102664.4, 102706.4, 102738.3, 102760.8, 102777.5, 102785.9, 102786.8,
  100588.9, 101874.9, 102328, 102402.6, 102471.2, 102525.1, 102587.6, 
    102655.5, 102715.5, 102763.2, 102806, 102835.9, 102855.4, 102865.7, 
    102870.9,
  100582.7, 101265.5, 102180.6, 102421.6, 102485.5, 102545.8, 102612.4, 
    102685.8, 102750.6, 102805.2, 102858.2, 102895.1, 102919.9, 102930.8, 
    102941.3,
  100300.5, 100132.9, 101040.6, 102348.4, 102493.3, 102553.8, 102619.3, 
    102697.4, 102765.7, 102829.7, 102890.5, 102931.6, 102962.5, 102983.9, 
    102997.8,
  100239.1, 99602.89, 99603.34, 101359.6, 102482.8, 102556.9, 102625.2, 
    102696.5, 102773.8, 102840.2, 102899.1, 102949.1, 102983.4, 103011.7, 
    103031.4,
  100464.1, 99754.51, 100234.7, 100763.2, 102389.3, 102542.7, 102616.4, 
    102687.8, 102765.2, 102834.7, 102902.7, 102957.7, 102995.9, 103026.9, 
    103049.2,
  99272.58, 99129.86, 100437.1, 100821.9, 101498.1, 102507.8, 102617.5, 
    102675, 102751.1, 102822.2, 102886.3, 102954.8, 102995.3, 103031.9, 103057,
  99299.57, 97854, 97726.81, 98930.47, 100669.3, 101441.9, 102594.3, 
    102668.9, 102721.1, 102804.4, 102855.8, 102926.7, 102983.9, 103021.1, 
    103050.7,
  102143.5, 102192.1, 102221.7, 102241.5, 102258.5, 102261.6, 102266.9, 
    102265.9, 102270.1, 102273.2, 102272.4, 102269.2, 102263.3, 102251.6, 
    102238.3,
  100759.7, 102166.9, 102254.4, 102283.4, 102312.3, 102325.2, 102340.2, 
    102354.2, 102369, 102385.2, 102395.4, 102403.4, 102408.2, 102408.1, 
    102404.5,
  100887.6, 101897.6, 102291.5, 102322.3, 102354.8, 102379.4, 102400.4, 
    102423, 102448.4, 102476.4, 102498.9, 102518, 102531.8, 102539.9, 102542.4,
  100592.2, 101851.8, 102286.6, 102338.7, 102378.4, 102416.7, 102449.5, 
    102482.3, 102517.9, 102553.5, 102584.4, 102614.2, 102637, 102654.5, 
    102664.8,
  100583.7, 101242.5, 102142.8, 102361.1, 102400.6, 102442.2, 102486.9, 
    102530.7, 102574.7, 102620.2, 102660.9, 102696.1, 102726.5, 102751.4, 
    102768,
  100302.4, 100115.8, 101006.6, 102292.7, 102415, 102460.9, 102514.7, 
    102569.1, 102618.8, 102675.9, 102718.5, 102760.9, 102798.7, 102827.2, 
    102848.6,
  100230.1, 99582.91, 99564.7, 101304.1, 102412.1, 102474.7, 102535, 
    102596.7, 102652.8, 102716.5, 102760.9, 102811.6, 102852.1, 102884.5, 
    102911.6,
  100459.7, 99737.57, 100190.3, 100707.8, 102329, 102471.7, 102543.3, 
    102607.6, 102673.4, 102739.8, 102786.3, 102845.5, 102885.1, 102923.4, 
    102951.7,
  99269.02, 99116.99, 100411.7, 100767.8, 101440.3, 102433.1, 102554.5, 
    102605, 102679.2, 102747.8, 102799.7, 102857.5, 102903.2, 102942.5, 
    102973.7,
  99298.84, 97844.42, 97709.99, 98891.93, 100644.1, 101397.1, 102545, 
    102598.1, 102657.5, 102739.7, 102796.8, 102849.8, 102902.6, 102949, 
    102981.5,
  101917.1, 102014.5, 102075.4, 102121.8, 102169.7, 102201.5, 102234.8, 
    102265.3, 102298.7, 102326.9, 102352.1, 102376.9, 102394.8, 102404.9, 
    102409.2,
  100565.7, 101998.9, 102111.8, 102162.9, 102213.3, 102244.2, 102280, 
    102321.4, 102363.6, 102408, 102445.2, 102476, 102496.1, 102510.3, 102518.9,
  100697.3, 101718.8, 102135.1, 102185.3, 102243.9, 102285.9, 102332.9, 
    102384, 102438.3, 102490, 102529.6, 102559.7, 102586.9, 102607.1, 102620.5,
  100408.3, 101679.4, 102134, 102197.8, 102256.7, 102307.4, 102365.6, 
    102428.3, 102494, 102549.2, 102596.7, 102636.2, 102671.2, 102694.9, 
    102713.4,
  100400.1, 101070.8, 101976.1, 102205.9, 102262.6, 102322.7, 102391, 102462, 
    102535, 102598.5, 102655.2, 102700.8, 102737.5, 102766.7, 102792.5,
  100121.1, 99949.48, 100842.2, 102126.8, 102258.1, 102319.8, 102401, 
    102480.7, 102562.7, 102635.2, 102691.8, 102743.9, 102787.9, 102827, 
    102860.1,
  100054.3, 99424.84, 99411.39, 101141.9, 102241.6, 102317.2, 102408.2, 
    102488.5, 102579.4, 102653.6, 102713.3, 102774.1, 102823.2, 102866.3, 
    102903.8,
  100282.2, 99573.27, 100033.5, 100543.4, 102147.6, 102297.5, 102405.7, 
    102489.3, 102586.6, 102664.9, 102726.5, 102786.9, 102840.3, 102888.4, 
    102933.2,
  99109.03, 98958.66, 100246.4, 100601.3, 101256.4, 102246.6, 102407.1, 
    102492.5, 102579.9, 102666.5, 102726.6, 102790.2, 102845.5, 102897.6, 
    102945.2,
  99141.74, 97701.03, 97567.41, 98740.08, 100471.2, 101212.3, 102378.8, 
    102492.2, 102561.6, 102660.1, 102717.9, 102780.7, 102837.9, 102896.5, 
    102949.6,
  101947.1, 102012, 102060.8, 102094.1, 102123.8, 102147.3, 102166.3, 
    102185.1, 102204.8, 102216.8, 102225.2, 102226, 102223.1, 102212.3, 102196,
  100577.5, 101985.2, 102086.1, 102126.3, 102169.4, 102198.6, 102226, 
    102255.9, 102285.2, 102312.1, 102331.9, 102343.9, 102350, 102349.1, 102343,
  100703.8, 101706.2, 102100.8, 102146.6, 102188.5, 102231.6, 102276.6, 
    102319.6, 102360.2, 102400.2, 102430.6, 102450.7, 102464.2, 102472.6, 
    102475.1,
  100412.7, 101662.1, 102094.2, 102149.7, 102201.2, 102255.4, 102310.8, 
    102364, 102414.7, 102463.1, 102500.9, 102532.4, 102556.6, 102576.1, 
    102588.7,
  100401.4, 101054.2, 101935.2, 102155.9, 102205.7, 102268.2, 102330.2, 
    102397.2, 102456, 102514.5, 102560.2, 102601.7, 102633.8, 102662.2, 
    102684.4,
  100121.6, 99937.87, 100810.3, 102085.9, 102207.2, 102272.1, 102344.9, 
    102418.7, 102485.8, 102551.1, 102604.9, 102651.5, 102694.7, 102732.3, 
    102763.4,
  100055.1, 99413.33, 99381.64, 101106.1, 102202.3, 102272.6, 102355, 
    102433.3, 102505.6, 102576.9, 102635.7, 102690.3, 102739.8, 102783.7, 
    102823,
  100292.6, 99570.73, 100010.2, 100514.8, 102124.4, 102268.7, 102358.6, 
    102440.8, 102514.2, 102592.3, 102650.9, 102713.8, 102769.5, 102819.9, 
    102868.7,
  99117.7, 98960.31, 100242, 100593.2, 101246.6, 102228.9, 102361.8, 
    102444.8, 102515.9, 102596.3, 102654.6, 102724.7, 102783.4, 102840.8, 
    102893.7,
  99166.12, 97716.99, 97573.07, 98739.06, 100480.1, 101217.3, 102342.3, 
    102445.7, 102504.7, 102591.3, 102650.8, 102721.6, 102781.8, 102844.9, 
    102901.9,
  102117.1, 102129.9, 102134.1, 102133.5, 102124.9, 102118.8, 102112.5, 
    102108.1, 102112.6, 102109.9, 102111.9, 102107.1, 102105.4, 102096.8, 
    102085.9,
  100716.7, 102096.1, 102155.7, 102163.5, 102164.1, 102168.9, 102170.1, 
    102174.7, 102185, 102192.7, 102203.9, 102210.3, 102212.8, 102211.9, 
    102209.8,
  100840.9, 101816.6, 102174.4, 102183.9, 102195.2, 102205.5, 102218.1, 
    102236.9, 102253.7, 102274.6, 102295.3, 102311, 102324.3, 102333.9, 
    102333.9,
  100556.7, 101783.4, 102181.5, 102206.5, 102225.2, 102239.8, 102259.2, 
    102283.4, 102307.2, 102333.9, 102361, 102384.9, 102404.6, 102422.3, 
    102435.2,
  100554.2, 101187.2, 102047.1, 102232.7, 102249, 102269.8, 102292.2, 
    102327.3, 102358.2, 102391.7, 102422.5, 102453, 102477.6, 102504.8, 
    102526.2,
  100285.1, 100079.5, 100930.6, 102179.2, 102269.1, 102285, 102318, 102358.6, 
    102397.6, 102436.9, 102473.9, 102510.4, 102544.6, 102578.6, 102605.4,
  100209.9, 99549.3, 99494.05, 101205.4, 102274.1, 102299.2, 102329.2, 
    102383.4, 102425.1, 102472.7, 102515.2, 102559.5, 102602.3, 102639.3, 
    102674,
  100465, 99711.33, 100127.3, 100610.4, 102196.3, 102295.9, 102333, 102397.4, 
    102443.3, 102495.1, 102544.8, 102596.7, 102644.4, 102687.2, 102726.7,
  99271.34, 99098.12, 100370.2, 100701.9, 101309.9, 102259.7, 102331, 
    102406.3, 102451.4, 102511.2, 102564.2, 102623.3, 102669.8, 102717.4, 
    102763.4,
  99323.77, 97848.24, 97690.14, 98838, 100551.4, 101289.2, 102322, 102412.5, 
    102450.1, 102516.3, 102570.7, 102635.4, 102681.8, 102735.8, 102783.1,
  102217.8, 102286.4, 102307.5, 102337.3, 102363.1, 102374.9, 102364.5, 
    102341.8, 102314.5, 102269.6, 102217.2, 102157.7, 102082.5, 101994.3, 
    101893,
  100775, 102219.3, 102287, 102291.2, 102302.8, 102322.4, 102327.9, 102320.9, 
    102306.7, 102273.6, 102225.5, 102173.2, 102111.7, 102041.8, 101959.1,
  100858, 101884.7, 102258.4, 102271.3, 102273.8, 102277.7, 102289.1, 
    102292.8, 102287.9, 102265.3, 102234.4, 102195.9, 102145.9, 102086.8, 
    102017.2,
  100524.4, 101781.4, 102214.7, 102247.1, 102258, 102253.3, 102261.4, 
    102267.2, 102263.3, 102253.2, 102232.4, 102203.8, 102167.5, 102123.2, 
    102067.3,
  100499.2, 101143.1, 102021.6, 102224.5, 102242.4, 102246.3, 102248.7, 
    102240.9, 102240.2, 102239.5, 102233, 102211, 102189.1, 102151.3, 102110,
  100208.5, 100008.2, 100874.7, 102141.5, 102230.1, 102238.5, 102240.8, 
    102248.7, 102243.5, 102241.8, 102231.8, 102216.4, 102199.4, 102180.6, 
    102150.3,
  100122.3, 99466.45, 99409.19, 101138.7, 102206.5, 102225.7, 102233.3, 
    102235.1, 102245.5, 102238.7, 102241.6, 102231.4, 102222.8, 102208, 
    102190.4,
  100374.6, 99623.02, 100037.2, 100518, 102117.1, 102211, 102220.1, 102241.2, 
    102256.6, 102264.5, 102259, 102255.2, 102250.8, 102245.3, 102233,
  99183.8, 99001.98, 100278.9, 100605.6, 101206.7, 102163.3, 102204.3, 
    102225.2, 102246.8, 102267.2, 102278.2, 102290.7, 102286.8, 102289.4, 
    102282.1,
  99239.23, 97750.84, 97587.84, 98739.01, 100436.6, 101200.3, 102191.7, 
    102218.9, 102245.8, 102273.7, 102292.2, 102307.6, 102318.6, 102328.2, 
    102330.6,
  101798.7, 101892, 101962, 102015.3, 102071.1, 102139.1, 102220, 102282.8, 
    102339.9, 102384.5, 102407.7, 102420.3, 102405.1, 102366, 102336.9,
  100416.7, 101858.5, 101968.5, 102017.9, 102068.8, 102119.3, 102197.4, 
    102263.8, 102318.8, 102366.5, 102398.6, 102411.4, 102401.9, 102369.1, 
    102339.4,
  100532.3, 101558.8, 101972.3, 102018.9, 102064.4, 102098.4, 102180.4, 
    102247.1, 102302.8, 102350.1, 102384.8, 102405.9, 102411.2, 102387.4, 
    102350.4,
  100231.4, 101507.2, 101956, 102019.8, 102060.1, 102087.9, 102144, 102223.4, 
    102280.1, 102322.5, 102358.1, 102381.7, 102392.6, 102383.7, 102352,
  100219, 100876.5, 101781.8, 102015.3, 102060.2, 102090.6, 102116.5, 
    102178.7, 102254.2, 102294.9, 102336.5, 102358.5, 102376.6, 102372, 
    102352.5,
  99938.63, 99751.45, 100637.2, 101933.1, 102048.4, 102082.3, 102116, 
    102152.2, 102203.9, 102267.8, 102303, 102325.8, 102345.4, 102352, 102348.1,
  99863.59, 99219.47, 99192.94, 100929.4, 102024, 102065.8, 102098.3, 
    102130.3, 102165.7, 102204.9, 102252.2, 102289.2, 102312.6, 102318.5, 
    102319.5,
  100106.1, 99372.06, 99812.78, 100317.3, 101923.2, 102045.8, 102082.4, 
    102116.7, 102153.8, 102181.8, 102205.7, 102233.9, 102267.8, 102279.1, 
    102294.7,
  98922.11, 98751.22, 100036.9, 100384.2, 101009.4, 101981.6, 102054.7, 
    102089.3, 102133.2, 102160.8, 102178.7, 102191.5, 102214.5, 102238.4, 
    102247.8,
  98973.6, 97502.82, 97345.07, 98504.12, 100221.5, 100987.6, 102040.3, 
    102071.4, 102119.4, 102161.7, 102179.1, 102179.9, 102190.4, 102198.7, 
    102212.6,
  101730.2, 101753.6, 101769.2, 101784.4, 101793.1, 101794.3, 101805.8, 
    101820.4, 101847.2, 101880, 101920.6, 101959.7, 102005.8, 102049.4, 
    102086.8,
  100356.6, 101724.2, 101805.4, 101831.4, 101851.6, 101861.9, 101878.2, 
    101903.5, 101934.8, 101971.8, 102016.8, 102064, 102115.1, 102159.4, 
    102196.5,
  100493, 101461.6, 101839.3, 101861.4, 101888.7, 101905, 101932.8, 101961.3, 
    101996.5, 102040, 102090.3, 102141.5, 102192.9, 102242, 102278.6,
  100217.8, 101440.4, 101855.2, 101890, 101924.9, 101949.4, 101980.8, 
    102011.8, 102051.8, 102097, 102146.3, 102198.1, 102255.2, 102304.8, 
    102347.5,
  100219.3, 100857.2, 101721.3, 101919.7, 101952.5, 101984.6, 102015, 
    102049.6, 102092.7, 102136.9, 102186.4, 102241, 102300.9, 102352.6, 
    102401.8,
  99950.33, 99749.55, 100607.4, 101869, 101970.5, 102000.4, 102038.6, 102078, 
    102119.7, 102167.9, 102218.4, 102270.4, 102334.7, 102386.5, 102435,
  99887.48, 99231.67, 99187.79, 100892.7, 101971.3, 102009.8, 102049.4, 
    102097.2, 102143.2, 102187.7, 102236.2, 102286.9, 102350.3, 102406.8, 
    102453.9,
  100139.3, 99392.91, 99817.23, 100305, 101887.7, 102005.7, 102052.9, 
    102105.3, 102158.8, 102203.7, 102250.4, 102296.4, 102360.4, 102411.6, 
    102464.4,
  98960.27, 98785.77, 100057.1, 100390.7, 100995.9, 101955.7, 102050.9, 
    102108.7, 102167.7, 102215.4, 102263.4, 102293.9, 102352, 102413.6, 
    102458.9,
  99018.96, 97552.92, 97395.91, 98536.1, 100246.1, 100974.1, 102037.2, 
    102111.9, 102168.1, 102227.2, 102273, 102303.7, 102336.2, 102394.9, 
    102446.8,
  102406.6, 102447.6, 102423.8, 102388.2, 102325, 102270.2, 102204, 102130.9, 
    102052.1, 101980.2, 101903.1, 101816.4, 101730.3, 101651.9, 101573.5,
  100921.8, 102364.6, 102396.2, 102363.5, 102313.6, 102263.2, 102213.9, 
    102153.4, 102090.9, 102023.4, 101949.6, 101876.3, 101800.8, 101727.3, 
    101659.2,
  100978.4, 102001.1, 102354.5, 102329.1, 102293.9, 102255.1, 102215.3, 
    102169.4, 102116.7, 102060.5, 102002.4, 101940.6, 101875.2, 101812.3, 
    101749.4,
  100607.1, 101886.9, 102289.1, 102285.6, 102258.7, 102229.3, 102198, 102163, 
    102124.2, 102082.1, 102035.9, 101988.8, 101935.2, 101883.8, 101836.7,
  100548, 101223.9, 102090, 102241.8, 102233.3, 102210, 102191.5, 102165.6, 
    102132.7, 102101.9, 102064.5, 102022.1, 101988.4, 101947.2, 101906,
  100250.9, 100037.5, 100929.2, 102162.1, 102205.6, 102189.7, 102177.5, 
    102156.7, 102139.3, 102116.8, 102093.2, 102060.9, 102030.2, 102000.3, 
    101974.3,
  100157.9, 99495.45, 99430.35, 101148.2, 102190.9, 102178.3, 102166.6, 
    102160.4, 102148.6, 102136.2, 102117.1, 102095.8, 102074.1, 102051.7, 
    102033.1,
  100409, 99655.8, 100051.5, 100525.1, 102105.5, 102176.5, 102165.3, 
    102165.6, 102159.9, 102155.5, 102150.5, 102136.2, 102119.7, 102105.3, 
    102093.6,
  99214.04, 99036.05, 100295.2, 100625.8, 101204.7, 102137, 102165, 102164.7, 
    102177.6, 102181.5, 102180.1, 102175.3, 102166.2, 102157.3, 102150.1,
  99269.88, 97785.73, 97626.26, 98762.41, 100442.2, 101183.5, 102171.3, 
    102180.3, 102187.4, 102208.8, 102219, 102226.6, 102224.8, 102218.5, 
    102211.1,
  102354.7, 102411.5, 102388.9, 102338.5, 102262.6, 102187.4, 102110.1, 
    102017, 101924.3, 101828.4, 101731.7, 101638.6, 101542.3, 101456.9, 
    101375.4,
  100891, 102337.3, 102377.8, 102342.1, 102284.3, 102215.3, 102139.4, 102058, 
    101970, 101882.3, 101784.3, 101693.7, 101603, 101514.8, 101429.9,
  100958.5, 101994.3, 102353.7, 102333.3, 102290.9, 102230.9, 102173.2, 
    102099.8, 102024.1, 101937.4, 101846.7, 101753.6, 101665, 101575.6, 
    101488.5,
  100575.9, 101888.3, 102299.6, 102310, 102276.7, 102240.6, 102190.8, 
    102134.1, 102069, 101995.8, 101916.4, 101827.1, 101738.5, 101649.5, 
    101560.6,
  100527.6, 101200.4, 102093.8, 102269.3, 102258.3, 102225.9, 102193.7, 
    102144.9, 102090.1, 102035.1, 101968.1, 101891.5, 101806.5, 101722.9, 
    101636,
  100201.8, 100026.9, 100908.1, 102177.6, 102232.1, 102212.2, 102189.9, 
    102155.7, 102110.9, 102061.2, 102004, 101937.8, 101869.5, 101790.9, 
    101712.1,
  100115.7, 99439.85, 99394.66, 101148, 102191.1, 102181.9, 102159.6, 
    102139.6, 102113.8, 102075.2, 102031, 101974.3, 101909.7, 101841.7, 
    101772.1,
  100388, 99609.33, 99997.99, 100498, 102091.8, 102165.8, 102142, 102128.7, 
    102102.9, 102074.7, 102036.7, 101995.3, 101941.3, 101882.7, 101817.7,
  99196.7, 99001.86, 100249.5, 100571.9, 101167.4, 102094.6, 102114, 
    102093.1, 102089.4, 102066, 102029.2, 101997.4, 101951.3, 101903.1, 
    101851.1,
  99242.07, 97745.9, 97577.77, 98711.75, 100373.6, 101147.5, 102121.7, 
    102106.5, 102064.5, 102060.4, 102019.9, 101994.1, 101955.2, 101910.8, 
    101860.3,
  102053, 102071.3, 102049.5, 102007.6, 101957.4, 101905.1, 101852.4, 
    101790.3, 101733.1, 101674.5, 101613.7, 101558.3, 101506.5, 101452.8, 
    101406.6,
  100624.9, 102023.3, 102052.3, 102039.1, 101988.9, 101933.7, 101892, 
    101842.2, 101794.8, 101746.9, 101696.1, 101647.1, 101598.2, 101551, 
    101501.1,
  100687.3, 101701.7, 102045.1, 102027.2, 101990.2, 101947.8, 101904.3, 
    101866.3, 101836, 101791.3, 101753, 101713.9, 101677.6, 101627.3, 101581.4,
  100367.8, 101614.7, 102012.4, 102012.4, 101993.2, 101971, 101937.9, 
    101898.2, 101864.3, 101838.1, 101805.9, 101773.2, 101738.7, 101696.2, 
    101649.8,
  100332.4, 100971, 101832.4, 101993.9, 101977.5, 101966.7, 101942.9, 
    101911.8, 101882.6, 101857.5, 101828.9, 101806.2, 101780.2, 101742.1, 
    101698.7,
  100022.9, 99817.59, 100671.8, 101928, 101974.9, 101955.9, 101940.4, 
    101923.3, 101900.9, 101881.5, 101856.6, 101832.5, 101809.9, 101784.3, 
    101741.6,
  99934.81, 99271.48, 99192.58, 100914.2, 101952.7, 101958.9, 101940, 
    101925.6, 101908, 101892.4, 101874.4, 101854.4, 101829.6, 101808.1, 
    101775.3,
  100226.9, 99438.91, 99833.09, 100304.5, 101878.4, 101950, 101942.5, 101928, 
    101927.1, 101909.9, 101893.1, 101870.7, 101843.9, 101819, 101793.7,
  99044.8, 98839.99, 100086, 100407.6, 100980.1, 101910.3, 101930.8, 101932, 
    101925.1, 101919.1, 101905.1, 101886.2, 101861.6, 101836, 101810.9,
  99100.62, 97593.44, 97420.7, 98543.6, 100209.4, 100972.5, 101941.3, 
    101952.7, 101915.8, 101925.6, 101917.9, 101903.2, 101880.9, 101859.3, 
    101828.6,
  102127, 102163, 102157.4, 102121.2, 102060.9, 102000.5, 101938.8, 101863.7, 
    101776.8, 101681.4, 101572.8, 101456.6, 101333.1, 101202.1, 101061.2,
  100749.3, 102158.5, 102191, 102171, 102122, 102064.3, 102005.9, 101939.9, 
    101860.1, 101771.8, 101669.9, 101557.5, 101445, 101319.1, 101185.4,
  100873.5, 101884.5, 102223.7, 102206.6, 102163.6, 102109.9, 102056.3, 
    101996.8, 101932.1, 101852.3, 101762.6, 101656.9, 101541.9, 101421.6, 
    101291.7,
  100580, 101847.2, 102235.3, 102239.5, 102199.2, 102148.5, 102103.9, 
    102049.6, 101987.3, 101918.7, 101836.9, 101739.7, 101637.2, 101520.8, 
    101398.2,
  100546.2, 101213.9, 102083.3, 102252.1, 102227.1, 102174.8, 102133, 
    102085.8, 102028.1, 101966.1, 101897.7, 101812.4, 101715, 101610.2, 
    101494.9,
  100256.1, 100048.8, 100935, 102195.6, 102243.8, 102196.6, 102159.6, 
    102116.6, 102064.9, 102006.8, 101944, 101868.2, 101783.4, 101687.6, 
    101587.4,
  100151.6, 99495.32, 99437.48, 101192.8, 102231, 102207.1, 102171, 102130.6, 
    102081, 102031.5, 101977, 101912.4, 101839.8, 101753.1, 101661.4,
  100367, 99643.5, 100041.9, 100560.5, 102155.1, 102214.8, 102181.1, 
    102144.8, 102096.5, 102042.8, 101990.5, 101936.4, 101875.3, 101807.3, 
    101724.2,
  99158.15, 98993.6, 100275.1, 100623.9, 101237.5, 102169.1, 102185, 
    102142.3, 102100.4, 102052.6, 101997.2, 101946.7, 101894.3, 101834.2, 
    101767.3,
  99186.51, 97693.64, 97553.85, 98721.9, 100422, 101194.9, 102171.1, 
    102164.7, 102100.6, 102060.5, 101998.3, 101941.4, 101886.6, 101839.8, 
    101787.9,
  101716.8, 101722.9, 101705.6, 101681.1, 101640.7, 101584.8, 101525, 
    101460.6, 101399.3, 101338.5, 101269.4, 101199.5, 101119.2, 101040.5, 
    100966.4,
  100379, 101732.3, 101772.7, 101755.7, 101732, 101684.3, 101633.1, 101576.2, 
    101516.3, 101456.7, 101388.1, 101317.6, 101250.4, 101186.5, 101121.1,
  100538.5, 101506.2, 101849.7, 101837.3, 101820.4, 101783, 101739.8, 
    101682.9, 101628, 101566.8, 101508.8, 101447.9, 101384.9, 101320.3, 
    101255.6,
  100288.9, 101507, 101902, 101909.1, 101902.6, 101876.1, 101843.5, 101800.6, 
    101753.6, 101700.1, 101649.3, 101594.5, 101536.2, 101475.2, 101410.4,
  100303.9, 100936.4, 101794.6, 101969.1, 101973.9, 101960.2, 101938.3, 
    101907.1, 101870.9, 101827.8, 101782.4, 101733.7, 101683.1, 101628, 
    101569.1,
  100049.7, 99835.72, 100690.5, 101946.7, 102026.6, 102025.3, 102015.8, 
    101999, 101975.7, 101947.4, 101913.1, 101873.9, 101829.4, 101780.9, 
    101729.1,
  99976.09, 99324.65, 99261.05, 100985.8, 102054.1, 102072.7, 102065.4, 
    102061.6, 102052.9, 102039.2, 102016.5, 101988.9, 101955.6, 101917.2, 
    101872,
  100239.2, 99500.89, 99914.73, 100410, 102000.3, 102102.5, 102107.7, 
    102115.1, 102117.1, 102114.3, 102105.4, 102088.4, 102066.9, 102036, 
    102001.9,
  99045.22, 98883.27, 100162.9, 100504.6, 101106.5, 102068.4, 102124.4, 
    102138.2, 102155.2, 102170.1, 102169.5, 102166.8, 102152.2, 102133.8, 
    102106.4,
  99101.91, 97640.21, 97483.77, 98637.88, 100336.2, 101092.4, 102138.5, 
    102177, 102182.9, 102217.8, 102220.2, 102229, 102223.8, 102214.2, 102192,
  102217, 102274.4, 102262.5, 102236.6, 102197.4, 102158.4, 102116.6, 
    102048.9, 101983.1, 101904.1, 101825, 101739, 101661.1, 101577.6, 101485.3,
  100757.3, 102186, 102230.2, 102202.8, 102169.5, 102138.9, 102109, 102052.5, 
    101993.9, 101928.6, 101852.6, 101782.6, 101704.5, 101627.5, 101539.2,
  100815.1, 101824.6, 102186, 102161.6, 102136.5, 102114.5, 102084.6, 
    102045.4, 101996.5, 101949.7, 101882.1, 101812, 101743.6, 101671.1, 
    101590.5,
  100473.1, 101730.2, 102132.9, 102126.6, 102101.8, 102086.6, 102066.5, 
    102032.8, 101992.1, 101950.5, 101897.8, 101840.7, 101775.9, 101711.1, 
    101642.1,
  100415.8, 101078, 101942.1, 102102.8, 102088, 102067.8, 102050.8, 102020.2, 
    101985.8, 101946.5, 101902.4, 101852.8, 101798, 101732.1, 101665,
  100111.1, 99912.7, 100788.2, 102028.2, 102076.4, 102057.4, 102044.7, 
    102022.4, 101992.5, 101958.4, 101921.2, 101873.2, 101821.8, 101764.9, 
    101705.4,
  100020.2, 99356.64, 99302.92, 101024.6, 102059.7, 102051.7, 102037.6, 
    102023.9, 102001.1, 101973.5, 101940.8, 101896.2, 101853.1, 101797.6, 
    101741.2,
  100266, 99510.25, 99917.36, 100401.2, 101991.6, 102060.7, 102042.8, 
    102032.4, 102015.8, 101994.2, 101965.6, 101928.5, 101886.7, 101840.9, 
    101788.6,
  99060.41, 98893.62, 100166.6, 100490.5, 101083.7, 102023, 102051.1, 
    102038.5, 102028.4, 102016.1, 101990.2, 101964.3, 101929.5, 101889.3, 
    101844.9,
  99108.91, 97640.45, 97478.5, 98637.46, 100329.3, 101070.5, 102062.6, 
    102066.2, 102043.4, 102044.1, 102020.8, 102000.9, 101971.4, 101940.5, 
    101904.2,
  101916.8, 101994.4, 102032.6, 102054.4, 102055.8, 102047, 102043.8, 
    102026.8, 101998.1, 101959.3, 101906.6, 101848.8, 101785.4, 101717.8, 
    101643.7,
  100501.1, 101941.2, 102022.9, 102046.9, 102061.9, 102074.2, 102085, 
    102074.8, 102060.9, 102032, 101992.4, 101944.7, 101890.1, 101831.6, 
    101763.8,
  100583.5, 101621.8, 102009.9, 102038.3, 102058.7, 102084.6, 102096.1, 
    102103.6, 102101.9, 102085.3, 102061.8, 102024.4, 101980, 101929.1, 
    101871.6,
  100241.5, 101544, 101974.2, 102021, 102051.3, 102085, 102106, 102111.3, 
    102111.3, 102116.4, 102109.8, 102081.9, 102047, 102008.4, 101960,
  100187.2, 100879, 101789.1, 102005.4, 102034.3, 102062.1, 102084.8, 
    102109.3, 102120.7, 102132, 102133.7, 102123.8, 102103.8, 102071.2, 
    102031.3,
  99872.9, 99710.23, 100615.7, 101910, 102017.1, 102047.1, 102067.5, 
    102095.6, 102115.6, 102136.6, 102137.8, 102138.5, 102132.4, 102118.7, 
    102097.3,
  99782.24, 99138.68, 99128.16, 100879.5, 101968.2, 102007.3, 102042.7, 
    102092.6, 102106, 102110.8, 102129, 102134.6, 102151.6, 102147.5, 102139.8,
  100013.9, 99291.52, 99739.49, 100246.8, 101867.1, 101978.5, 101997.8, 
    102048.1, 102075.2, 102115.8, 102122.1, 102118, 102136.3, 102146.6, 
    102154.8,
  98811.1, 98654.23, 99952.87, 100307.4, 100941, 101907.5, 101974.2, 
    101998.2, 102039.5, 102062.2, 102082.8, 102110.3, 102118.2, 102135.7, 
    102139.9,
  98857.86, 97398.3, 97241.72, 98423.39, 100162, 100909.6, 101966.9, 
    101972.1, 101989, 102028.7, 102045.3, 102078.3, 102101.8, 102115.7, 
    102127.2,
  101616.1, 101688.8, 101726.5, 101753.8, 101771.9, 101768, 101764.3, 
    101739.9, 101711, 101680.9, 101643.4, 101598.5, 101558.1, 101505.7, 
    101445.4,
  100187.4, 101627.4, 101698.9, 101734, 101776.9, 101783.7, 101789.2, 
    101779.3, 101762.3, 101740.1, 101709, 101673.5, 101636.7, 101592.9, 
    101541.4,
  100270.8, 101287.8, 101675, 101714.7, 101756.1, 101773.1, 101799.2, 
    101810.6, 101804.4, 101791.4, 101768.5, 101742.5, 101711.2, 101680, 
    101634.2,
  99940.81, 101198, 101629, 101682, 101730, 101743.4, 101780.5, 101814.4, 
    101826.7, 101826.9, 101820.6, 101804.6, 101786.5, 101760.2, 101726.8,
  99908.41, 100566.1, 101451.2, 101652.1, 101696.5, 101732.6, 101759.4, 
    101799.2, 101829.9, 101848.2, 101859.8, 101855.6, 101849.1, 101831.8, 
    101811.5,
  99630.29, 99423.8, 100292.6, 101572.4, 101671.9, 101703.5, 101745, 
    101779.3, 101814.8, 101857.8, 101875.4, 101878.9, 101880.5, 101878, 
    101874.7,
  99544.24, 98886.66, 98844.8, 100571.8, 101641.9, 101679.4, 101713.4, 
    101757, 101796.1, 101828.7, 101863.1, 101880.6, 101896.9, 101911, 101912,
  99795.41, 99048.7, 99465.74, 99961.26, 101551.1, 101648.1, 101690.7, 
    101733.7, 101781.1, 101814.6, 101846.3, 101866.8, 101884.4, 101905.7, 
    101926.4,
  98596.12, 98427.95, 99705.69, 100050.6, 100661.9, 101606.9, 101668.9, 
    101703.6, 101753.5, 101800.6, 101832.3, 101858.9, 101881.5, 101904.9, 
    101939.7,
  98658.69, 97184.15, 97038.59, 98185.88, 99886.29, 100633.2, 101655.9, 
    101700, 101736.8, 101798.8, 101828.6, 101864.5, 101883.4, 101909.6, 101935,
  101876.8, 101984.4, 102042.8, 102091, 102130.3, 102161.1, 102202.6, 
    102235.7, 102286.3, 102327.5, 102368.2, 102401, 102425, 102432.2, 102426,
  100481.7, 101930.7, 102021.7, 102065, 102105.9, 102142.2, 102186.8, 
    102222.2, 102251.1, 102306.9, 102350.5, 102387, 102418.5, 102426.2, 
    102424.5,
  100558.3, 101593.5, 101995.5, 102035.4, 102075.8, 102113.8, 102176.5, 
    102211.5, 102232.6, 102278.1, 102327.7, 102362.7, 102395.8, 102414.6, 
    102424.3,
  100225.1, 101514.9, 101950.3, 102008.9, 102039.3, 102081.5, 102134.3, 
    102183.3, 102227.5, 102246.6, 102281.3, 102322.1, 102354.2, 102380.3, 
    102397.6,
  100163.9, 100851, 101755.8, 101970.2, 102011.1, 102047.8, 102098.8, 
    102150.6, 102192.5, 102228.1, 102251.1, 102276.8, 102308.8, 102332.2, 
    102354.9,
  99852.22, 99673.82, 100578, 101858.8, 101959.6, 102002.2, 102048.2, 
    102109.8, 102166.2, 102211.1, 102236, 102255.9, 102269, 102288.9, 102312.7,
  99738.72, 99108.52, 99080.72, 100838.6, 101915.2, 101960.3, 102004.8, 
    102064.4, 102115.9, 102174.6, 102212.7, 102234.2, 102248, 102258, 102272.4,
  99947.94, 99234.77, 99672.89, 100182.8, 101787.9, 101898.4, 101946.1, 
    102004.2, 102064.5, 102113.7, 102165.7, 102202.2, 102220.8, 102234.8, 
    102240.2,
  98725.68, 98586.9, 99888.41, 100224, 100856.6, 101826.2, 101896.3, 
    101943.6, 102011.3, 102067, 102111.4, 102155.1, 102179.5, 102202.7, 102214,
  98741.73, 97284.52, 97158.44, 98348.05, 100060.8, 100814.6, 101848.2, 
    101891.2, 101947.6, 102019.6, 102067.7, 102108.3, 102130.7, 102154.7, 
    102159.1,
  102020.2, 102121.4, 102190.3, 102242.4, 102303.3, 102347.8, 102407.1, 
    102452.2, 102494.6, 102534.6, 102564.2, 102590.4, 102612.9, 102631.1, 
    102640.7,
  100621.4, 102073.7, 102185.9, 102243.1, 102309.6, 102362.6, 102428.9, 
    102478.2, 102525.7, 102570.2, 102609.7, 102640.8, 102672.1, 102699.6, 
    102716.5,
  100718.5, 101754.3, 102169.2, 102232.5, 102297.9, 102359.7, 102433.5, 
    102492.3, 102543.4, 102593.4, 102639.7, 102677.2, 102716.1, 102749.3, 
    102773.3,
  100391.1, 101679.4, 102133.1, 102212, 102284.9, 102351.4, 102425.5, 102492, 
    102545.8, 102602.9, 102645.9, 102690.6, 102734.6, 102773.4, 102812.2,
  100344.8, 101028.5, 101946.4, 102181.5, 102256.6, 102328.1, 102405.9, 
    102477.8, 102537.9, 102597.9, 102646.3, 102692.2, 102737.6, 102787.4, 
    102832.7,
  100026.5, 99861.86, 100775, 102080, 102226.8, 102297.2, 102377.8, 102455.7, 
    102517.1, 102580.4, 102630.7, 102681.3, 102728.7, 102781.7, 102830.4,
  99928.38, 99303.13, 99303.9, 101061.4, 102179.8, 102266, 102343.3, 
    102427.2, 102491.2, 102552.8, 102608.5, 102661.5, 102707.8, 102761.2, 
    102812.9,
  100130.2, 99432.97, 99903.31, 100431.4, 102053.6, 102217, 102297.1, 
    102388.3, 102461, 102517.6, 102571.6, 102623.5, 102672.8, 102719, 102767.9,
  98922.5, 98786.84, 100089.2, 100458.2, 101130.4, 102148.8, 102260.5, 
    102330.2, 102424.4, 102483.5, 102535, 102581.7, 102629.7, 102679.7, 
    102720.3,
  98930.55, 97495.08, 97361.45, 98564.32, 100288.1, 101079.6, 102207.4, 
    102282.2, 102360.1, 102442.9, 102497.2, 102543.7, 102581.2, 102623.9, 
    102660.5,
  101816.1, 101943.7, 102030.2, 102106.2, 102179.7, 102250.5, 102331.6, 
    102396, 102450.9, 102504.9, 102535.8, 102564, 102583.1, 102592.8, 102586.8,
  100437.9, 101888.3, 102024.8, 102108.4, 102189, 102266.1, 102349.8, 
    102416.2, 102475.3, 102532.5, 102574.2, 102613.9, 102640.3, 102657, 
    102661.7,
  100546.9, 101581.5, 102015.6, 102099.7, 102184, 102266.5, 102357.2, 
    102434.7, 102498.3, 102565, 102611.9, 102651.7, 102683.6, 102713, 102724.1,
  100230.1, 101524.3, 101988.2, 102084.9, 102174.2, 102262.8, 102355, 
    102441.7, 102511.3, 102578.8, 102626.7, 102674, 102716.8, 102750.3, 
    102774.1,
  100204.4, 100896, 101818.6, 102071.7, 102154.2, 102248.2, 102344, 102441, 
    102518, 102586.7, 102639.3, 102689, 102731.6, 102777.2, 102812.7,
  99907.41, 99758.41, 100665.1, 101984.6, 102136.1, 102224.1, 102320.1, 
    102423.5, 102510.8, 102580.1, 102637.7, 102691, 102738.4, 102790.2, 
    102830.7,
  99834.91, 99219.26, 99229.41, 100984.2, 102105.4, 102201.8, 102295.5, 
    102398.3, 102498.9, 102568.7, 102632, 102687, 102731.3, 102772.3, 102819.4,
  100054.7, 99366.43, 99847.69, 100382.2, 101996.5, 102164.9, 102263.8, 
    102359.1, 102471.5, 102548.1, 102614.4, 102676.5, 102724.1, 102763.3, 
    102802.1,
  98878.36, 98743.2, 100045, 100429.3, 101099.7, 102105.1, 102246, 102320.8, 
    102432.4, 102523.2, 102590, 102655.3, 102711.1, 102753.9, 102789.7,
  98921.2, 97492.22, 97364.61, 98551.25, 100291.9, 101055.1, 102213, 
    102295.7, 102379.1, 102487.2, 102556.2, 102622.1, 102686.1, 102740.6, 
    102779.8,
  101812.2, 101876.7, 101917.1, 101947.1, 101973.5, 101990.6, 101997.3, 
    102003.2, 101997.7, 101992.4, 101975.7, 101948.4, 101913.5, 101862.1, 
    101800.8,
  100411.2, 101825, 101916.6, 101947.7, 101983.4, 102006, 102026.3, 102036.5, 
    102043, 102044, 102034.7, 102018.7, 101993.3, 101956.5, 101908.5,
  100523.3, 101531.8, 101923.8, 101955.7, 101993.8, 102020, 102045.9, 102068, 
    102083, 102091.5, 102091.7, 102084.9, 102064.5, 102039, 101999.9,
  100215.9, 101475.6, 101904.3, 101954.1, 101989.5, 102025.8, 102061.3, 
    102093.3, 102118.2, 102135.5, 102146.3, 102148.7, 102137.2, 102121.5, 
    102087.4,
  100204.1, 100866.2, 101752.4, 101960.6, 101990.8, 102029.3, 102067.2, 
    102111.4, 102143.6, 102170.8, 102190.4, 102203.6, 102202.9, 102192.2, 
    102170.9,
  99924.17, 99748.64, 100622.5, 101893.7, 101992.5, 102029.2, 102072.2, 
    102120.6, 102159.2, 102198.2, 102227.1, 102248.7, 102256.2, 102257.4, 
    102251.2,
  99858.66, 99226.09, 99201.38, 100914, 101992.2, 102039.8, 102080.7, 
    102133.4, 102176.6, 102220.7, 102253, 102281.7, 102298.5, 102312.2, 
    102318.8,
  100097.6, 99384.3, 99826.91, 100322.2, 101914.2, 102044, 102088.5, 
    102147.6, 102191.2, 102237.3, 102273.5, 102306.8, 102332.8, 102354.6, 
    102366.5,
  98923.23, 98774.75, 100061.2, 100413.8, 101039.6, 102018, 102105.8, 
    102163.4, 102204.1, 102252.5, 102289.8, 102328.3, 102355.7, 102385.9, 
    102400.7,
  98972.16, 97537.35, 97393.82, 98557.35, 100279.5, 101027.3, 102098.6, 
    102174.2, 102202.3, 102264.2, 102302, 102344.6, 102372.4, 102404, 102427.6,
  102009, 102170.4, 102269.6, 102349.2, 102423.3, 102495.7, 102556, 102603, 
    102628.5, 102637.3, 102627.5, 102605.2, 102555.4, 102489, 102394,
  100552.9, 102041.6, 102172.5, 102254.9, 102331, 102406.7, 102463.7, 102510, 
    102537.9, 102551.7, 102549.7, 102533.8, 102497.3, 102439.8, 102355.1,
  100598.2, 101666.8, 102100.7, 102172.2, 102244, 102312.9, 102371.9, 
    102416.1, 102446.6, 102465.1, 102464.8, 102454, 102431, 102383, 102312.7,
  100236.8, 101550.7, 102011.7, 102097.6, 102163, 102233.1, 102286.3, 
    102331.7, 102361.4, 102378.7, 102380.3, 102371.4, 102351, 102317.5, 
    102257.3,
  100183.6, 100880.1, 101795.3, 102028.9, 102092.8, 102149.9, 102203.8, 
    102249.5, 102282.9, 102298.6, 102303.9, 102291.7, 102269.6, 102236.5, 
    102186.2,
  99877.96, 99715.7, 100627.6, 101915.9, 102030.9, 102082.9, 102129.2, 
    102178.3, 102205.1, 102227.5, 102229.7, 102221.6, 102195.9, 102164.6, 
    102120,
  99781.61, 99161.82, 99144.84, 100898.6, 101978.7, 102028.7, 102065.4, 
    102108.1, 102136.9, 102157.3, 102165.6, 102160.1, 102134.7, 102105.8, 
    102062,
  100011.5, 99303.65, 99752.12, 100259.5, 101864.4, 101976.9, 102011.1, 
    102050.1, 102072.9, 102099.8, 102106.2, 102102.3, 102081.5, 102054.8, 
    102011.6,
  98817.69, 98674.33, 99968.34, 100323.3, 100950.1, 101910.7, 101963.2, 
    102000.6, 102026.3, 102044.7, 102053.7, 102053.6, 102036.8, 102010.6, 
    101974.4,
  98857, 97418.6, 97275.76, 98447.55, 100156.2, 100929.1, 101938.6, 101954.1, 
    101975, 102010.1, 102018.5, 102019.7, 102004.5, 101980.8, 101944.8,
  101800.6, 101994.8, 102138.5, 102257.4, 102371.4, 102483.5, 102578.8, 
    102666.5, 102730.9, 102777.2, 102805.2, 102811.5, 102804.1, 102775.7, 
    102726.7,
  100386, 101898.5, 102076.9, 102199.6, 102322.3, 102446.2, 102540.2, 
    102631.1, 102700.9, 102750.5, 102786.8, 102803.4, 102800.6, 102781.1, 
    102739.1,
  100477.1, 101568.6, 102040.6, 102165.8, 102285.2, 102404.9, 102510.9, 
    102595.8, 102670.5, 102731.1, 102768.1, 102792.3, 102792.9, 102779.4, 
    102744.3,
  100148.6, 101479.5, 101974.8, 102108.1, 102231.7, 102361, 102466.5, 
    102556.5, 102633.1, 102694.6, 102736.1, 102767.7, 102777.5, 102765.7, 
    102737,
  100110.4, 100827.7, 101790.6, 102069.2, 102188.7, 102309.7, 102420.3, 
    102512.6, 102585, 102653.2, 102695.8, 102730, 102744.6, 102740.2, 102718.5,
  99801.27, 99657.75, 100604, 101953.6, 102128.8, 102253.2, 102369.5, 
    102464.1, 102536.4, 102606.2, 102647.3, 102680.2, 102697.3, 102702.1, 
    102694.6,
  99715.33, 99111.22, 99126.77, 100927, 102067.9, 102192.1, 102307.2, 
    102407.5, 102485.8, 102553.1, 102604.3, 102639.6, 102659, 102665.9, 
    102659.1,
  99944.05, 99246.5, 99723.6, 100280.1, 101939.8, 102122.2, 102238.6, 
    102344.7, 102430.2, 102493.5, 102547.3, 102586.5, 102612.1, 102620.5, 
    102618.3,
  98752.46, 98618.35, 99930.98, 100313.1, 101003.1, 102032.6, 102172.8, 
    102275, 102365.4, 102440.3, 102490.4, 102530.9, 102557.8, 102576.1, 
    102578.9,
  98798.12, 97358.04, 97224.56, 98416.01, 100182.9, 100985, 102116.1, 
    102202.6, 102296.9, 102373.4, 102432.8, 102471.9, 102500.3, 102518.1, 
    102528.7,
  101148.7, 101159.5, 101159.7, 101190.7, 101248.5, 101324.3, 101422.1, 
    101524, 101627.5, 101739.1, 101841.3, 101936.5, 102019.9, 102084.1, 
    102128.1,
  99790.12, 101159.6, 101240.8, 101273.3, 101329.4, 101395, 101490.7, 101598, 
    101696.5, 101803.5, 101901.9, 101999.7, 102081.9, 102149.1, 102191.2,
  99919.16, 100900.4, 101272.9, 101303.1, 101368.2, 101442.8, 101547.1, 
    101651.9, 101745.5, 101855.6, 101953.7, 102053.1, 102139.1, 102203.2, 
    102253.6,
  99657.43, 100899.8, 101327.8, 101371.3, 101429.6, 101505.7, 101602.1, 
    101704.2, 101794.4, 101900.2, 101996.9, 102092.4, 102185.7, 102250.5, 
    102303.2,
  99680.09, 100327.9, 101210, 101420.2, 101472.9, 101545.1, 101637.3, 
    101743.2, 101835.6, 101937.9, 102033.5, 102124.9, 102220.1, 102286.8, 
    102341.9,
  99447.74, 99244.15, 100116.7, 101399.5, 101522.5, 101588.4, 101677.7, 
    101780.1, 101873.8, 101968.9, 102060.4, 102153.6, 102241.3, 102315.3, 
    102374.2,
  99418.58, 98765.18, 98729.97, 100448.5, 101546.2, 101622.6, 101703.9, 
    101810.6, 101907.2, 101998.2, 102086.8, 102176.8, 102261.3, 102330.8, 
    102392.5,
  99706.78, 98966.09, 99391.2, 99899.79, 101495.7, 101652.8, 101730.9, 
    101838.8, 101933.6, 102023.2, 102106.6, 102189.7, 102276.7, 102344.8, 
    102405.7,
  98570.3, 98392.06, 99660.09, 100019.4, 100648.6, 101638.5, 101763.6, 
    101855.6, 101951.9, 102048.4, 102128.4, 102196.9, 102282.5, 102348.9, 
    102404.3,
  98659.99, 97197.95, 97034.06, 98180.57, 99896.32, 100665, 101768.9, 
    101885.1, 101959.6, 102067.6, 102143.4, 102207.3, 102279.5, 102348.7, 
    102405.7,
  101745.5, 101742.2, 101714.4, 101681.7, 101629.9, 101556.7, 101476.6, 
    101391, 101299.9, 101215.3, 101138.7, 101074.8, 101030.1, 100997.1, 
    100967.7,
  100372.7, 101750.6, 101768.7, 101729.7, 101681.6, 101616.9, 101539.3, 
    101454.5, 101378.4, 101304.1, 101241.8, 101187.9, 101144.1, 101112.8, 
    101091,
  100505.1, 101497.2, 101822.4, 101782.9, 101727.9, 101671.9, 101600.1, 
    101526.5, 101460.2, 101391, 101336.1, 101282.9, 101249.5, 101225.1, 
    101209.2,
  100214.3, 101469.5, 101842.3, 101817.9, 101769.4, 101710.3, 101649.7, 
    101586.1, 101521.6, 101467.4, 101418.6, 101379.2, 101345, 101322.4, 
    101313.3,
  100194.9, 100847.8, 101704.3, 101837.8, 101799.1, 101744, 101685.4, 
    101631.1, 101575.2, 101522.7, 101480.8, 101447.3, 101422.5, 101407.2, 
    101403.6,
  99897.77, 99687.48, 100562.7, 101794, 101819.3, 101766.9, 101719.9, 
    101672.1, 101617, 101571, 101537.8, 101510.8, 101490.9, 101483.9, 101488.7,
  99775.34, 99122.88, 99056.77, 100796.9, 101820.7, 101790.8, 101737.2, 
    101697.5, 101653.4, 101616, 101587.1, 101566.9, 101554.9, 101557.8, 
    101568.1,
  100016.8, 99270.19, 99668.45, 100160.3, 101742.1, 101806.2, 101765.3, 
    101734, 101694.9, 101660.2, 101636.9, 101621.3, 101613, 101619.9, 101638.4,
  98769.6, 98604.66, 99897.87, 100253.2, 100841.3, 101770.8, 101773.1, 
    101749.9, 101728.6, 101710.8, 101690.1, 101680.2, 101677.4, 101685.5, 
    101710.7,
  98804.97, 97334.21, 97180.69, 98343.17, 100044.9, 100816, 101797.9, 
    101791.1, 101751.8, 101754.3, 101739.9, 101742.5, 101745.2, 101757.6, 
    101781.9,
  101102.1, 101160.4, 101193.7, 101226.3, 101257.5, 101298.1, 101344.8, 
    101392.4, 101435.1, 101466.8, 101485.3, 101495.3, 101498.4, 101492.6, 
    101474.3,
  99742.37, 101159.8, 101257.1, 101291.1, 101332, 101375.1, 101426.8, 
    101478.1, 101520.6, 101552.5, 101577.4, 101594.2, 101598, 101596, 101583.7,
  99894.62, 100914.3, 101309.9, 101341.1, 101393.7, 101442.7, 101499.4, 
    101557.2, 101598.6, 101635.8, 101665.3, 101683.7, 101694.3, 101692.9, 
    101679.7,
  99631.84, 100905.2, 101350.7, 101403.3, 101457.3, 101509.4, 101566, 
    101624.1, 101669.6, 101712.7, 101742.9, 101764.3, 101774.5, 101774.9, 
    101765.5,
  99666.33, 100335.4, 101238.6, 101458.8, 101504.7, 101562.9, 101621.3, 
    101682.6, 101731.8, 101771.6, 101809, 101827.8, 101839.5, 101841.8, 
    101837.4,
  99415.5, 99243.88, 100129.3, 101432.1, 101548.9, 101596.9, 101661.6, 
    101723.3, 101771.2, 101818.1, 101853.6, 101874.9, 101888, 101893.4, 
    101888.1,
  99379.35, 98754.75, 98735.45, 100468, 101573.6, 101625.6, 101686.2, 
    101746.9, 101802.2, 101847.1, 101881.2, 101906.2, 101922.6, 101933.6, 
    101933.5,
  99653.89, 98935.53, 99387.2, 99898.31, 101509.2, 101645.4, 101707.4, 
    101762.3, 101818.6, 101865.8, 101903.1, 101928.9, 101946.4, 101959.8, 
    101957.2,
  98504.97, 98350.16, 99632.59, 100012.3, 100638.3, 101616.8, 101722.3, 
    101767.7, 101828.8, 101876.4, 101914.4, 101943.9, 101962.7, 101977.4, 
    101981.6,
  98587.09, 97140.83, 96989.61, 98143.82, 99862.7, 100633.7, 101725.9, 
    101783.8, 101820.2, 101885.3, 101920.1, 101950.8, 101963.9, 101982.1, 
    101992,
  101116.2, 101093, 101057.3, 101023.7, 100974.2, 100898.8, 100821.2, 
    100747.5, 100685.5, 100632.3, 100596, 100572.9, 100554, 100540.3, 100532.1,
  99682.87, 101075.1, 101085.8, 101039.3, 100982.4, 100913, 100858.8, 
    100812.1, 100772.6, 100732.2, 100702.6, 100675.9, 100661.1, 100654.1, 
    100654.8,
  99730.4, 100748.6, 101074.1, 101044.5, 101007.1, 100969.2, 100923.8, 
    100890.2, 100860, 100837.8, 100814.4, 100796.4, 100782.1, 100778.3, 
    100784.7,
  99346.04, 100601.8, 100995.1, 100996.7, 100972.1, 100958.9, 100945.1, 
    100930, 100918.4, 100913.1, 100906.1, 100899.5, 100895, 100900.5, 100910.7,
  99271.91, 99945.22, 100810.3, 100975.3, 100965.4, 100968.6, 100971.3, 
    100976.8, 100981.2, 100984.3, 100992.5, 100999.4, 101003.8, 101016.7, 
    101034.3,
  98999.19, 98778.59, 99636.75, 100900, 100976.7, 100981.6, 100999.4, 
    101018.3, 101032.7, 101048.1, 101067.3, 101085.3, 101106.6, 101130.3, 
    101151.3,
  98965.54, 98308.77, 98255.08, 99952.48, 101026.8, 101036.6, 101043.9, 
    101068.2, 101087.1, 101111.6, 101134.9, 101157.5, 101186.1, 101216.9, 
    101247.2,
  99271.27, 98519.24, 98928.96, 99411.75, 100989, 101102.6, 101111.2, 
    101129.8, 101149.8, 101173.4, 101196.3, 101224.7, 101257.7, 101295.7, 
    101331.5,
  98174.42, 97986.73, 99236.17, 99590.14, 100177.4, 101120.1, 101183.2, 
    101204.3, 101235.2, 101261.4, 101284.3, 101315.6, 101346.1, 101385.6, 
    101422.9,
  98294.73, 96834.4, 96660.64, 97777.74, 99463.51, 100206.5, 101243, 
    101281.1, 101288.5, 101336.4, 101357.5, 101394.2, 101425.4, 101458.5, 
    101498.1,
  101188, 101131.3, 101077.2, 101011.6, 100951.5, 100892.3, 100838.5, 100797, 
    100760.4, 100742.6, 100725.7, 100711.7, 100711.2, 100713.6, 100726.7,
  99764.34, 101103.3, 101102, 101052.3, 101006.8, 100946.3, 100893.9, 
    100847.6, 100804.8, 100772.6, 100742.4, 100723.9, 100720, 100720.4, 
    100725.2,
  99877.09, 100840.7, 101131.6, 101061.2, 100979.5, 100915.9, 100868.4, 
    100827.2, 100788.8, 100755.7, 100722.4, 100689.6, 100665.2, 100644.8, 
    100625.6,
  99553.15, 100756.3, 101103.6, 101035.8, 100954.2, 100885.4, 100832.2, 
    100779.2, 100742.2, 100709.8, 100663.2, 100626, 100590, 100548.8, 100515.3,
  99519.89, 100139.8, 100941, 101010.8, 100927.1, 100848.3, 100797.4, 
    100738.5, 100684.1, 100646.4, 100608.3, 100564.1, 100532.1, 100515.1, 
    100516.5,
  99198.53, 98954.7, 99771.26, 100927.1, 100896.9, 100801.3, 100747.5, 
    100701.8, 100650.1, 100626.5, 100606.9, 100593.3, 100590.3, 100593.1, 
    100603.9,
  99079.94, 98373.48, 98268.44, 99952.64, 100926, 100863.8, 100795.9, 
    100756.7, 100710.4, 100687.8, 100673.6, 100663.1, 100659.9, 100675, 
    100696.4,
  99283.91, 98506.52, 98888.06, 99346.55, 100838.3, 100872.6, 100826.2, 
    100810.5, 100781, 100762.3, 100748, 100748.4, 100758.6, 100778.5, 100803.2,
  98021.12, 97823.6, 99081.85, 99434.11, 99997.97, 100884.1, 100869.1, 
    100841, 100833.3, 100837.7, 100829.5, 100835.9, 100852.6, 100881.3, 
    100921.7,
  98080.45, 96593.8, 96383.75, 97492.65, 99164.12, 99914.26, 100931, 
    100923.8, 100888.6, 100916.1, 100918.3, 100942.9, 100963.6, 101002.9, 
    101048.9,
  101957.8, 101784.8, 101655.1, 101515.3, 101369.5, 101206.2, 101049.9, 
    100910.2, 100794.2, 100694.3, 100606.7, 100525.6, 100458.2, 100393.3, 
    100336.1,
  100577.8, 101852, 101750.6, 101603.6, 101459.9, 101292.4, 101146.4, 
    101013.5, 100892.9, 100788.5, 100695.9, 100614, 100534.9, 100472, 100415.1,
  100750.3, 101676.2, 101873.8, 101714.1, 101544.8, 101392.6, 101261, 
    101135.3, 101017.1, 100909.1, 100814.2, 100730.2, 100651.9, 100581.2, 
    100520.1,
  100517.9, 101683.4, 101957.1, 101819.5, 101648.1, 101481.6, 101344.6, 
    101222.8, 101107.5, 101005.8, 100913.9, 100832.2, 100752.9, 100686.5, 
    100624.4,
  100554.8, 101098.8, 101869.9, 101890.3, 101735.8, 101574.5, 101433, 
    101311.4, 101198.4, 101095.7, 101001.1, 100918.5, 100842.2, 100777, 
    100719.7,
  100305.6, 99960.88, 100740, 101878.2, 101799.7, 101640.8, 101504.6, 
    101379.8, 101264, 101161.6, 101071.4, 100989.7, 100918.5, 100852.2, 
    100791.7,
  100234.5, 99427.47, 99243.77, 100912.8, 101846.2, 101706.2, 101557.6, 
    101441.2, 101323.6, 101221.2, 101127.9, 101041.3, 100966.9, 100899.5, 
    100840.8,
  100520, 99632.98, 99904.58, 100304, 101807.2, 101773.6, 101623.8, 101499.5, 
    101380.3, 101279.4, 101190.9, 101106.5, 101029.1, 100962.9, 100905.9,
  99281.45, 98979.27, 100190.4, 100442.1, 100936, 101757.7, 101649.3, 
    101526.8, 101425.2, 101333.5, 101238.7, 101165, 101094.9, 101038.2, 
    100986.3,
  99290.1, 97679.45, 97427.3, 98513.41, 100143.9, 100841, 101710, 101587.8, 
    101441.1, 101378.9, 101276.7, 101206.5, 101137.7, 101078.3, 101022.5,
  102383, 102255.4, 102135.6, 101963.7, 101772.1, 101554.7, 101337.4, 
    101140.7, 100958.1, 100797.2, 100644.2, 100496, 100357.1, 100220.6, 100081,
  101028.6, 102315.5, 102240, 102090.9, 101914.1, 101691.3, 101470.7, 
    101268.5, 101082.9, 100909.3, 100749.9, 100597.5, 100459.8, 100325.3, 
    100190.6,
  101202.2, 102125.5, 102331.4, 102188.5, 102014, 101823.8, 101615.3, 
    101397.2, 101200.7, 101025, 100862.7, 100708.7, 100565.7, 100429.2, 
    100295.2,
  100999.8, 102180.1, 102434.8, 102303.8, 102122.2, 101934.4, 101746, 
    101543.8, 101336.5, 101151.2, 100986.7, 100833.3, 100687.2, 100548.2, 
    100414.7,
  101043.6, 101621.9, 102377.2, 102403.6, 102232.1, 102040, 101861.9, 
    101675.5, 101478.3, 101277.3, 101111.4, 100958.7, 100813, 100672.5, 100533,
  100838.4, 100500.4, 101297.5, 102445, 102339.8, 102151.9, 101968.9, 
    101798.2, 101616.3, 101423.5, 101242.9, 101082.7, 100935.5, 100796.8, 
    100659.7,
  100798.9, 100007, 99819.62, 101515, 102443.2, 102270.9, 102078.6, 101909.6, 
    101737.9, 101560.3, 101383.4, 101218.3, 101064.2, 100925.8, 100785.1,
  101147.1, 100265.5, 100536.6, 100957.2, 102474.8, 102391.6, 102194.6, 
    102031.2, 101857.3, 101692.7, 101519.6, 101351.6, 101195.3, 101047.3, 
    100912.4,
  99937.89, 99663.62, 100884.2, 101149.1, 101655.2, 102487.6, 102312.6, 
    102131.9, 101967.6, 101812.9, 101647.6, 101487.6, 101325.6, 101177.8, 
    101037.3,
  100006.5, 98372.25, 98127.38, 99253.83, 100864.4, 101588.2, 102446.5, 
    102290.5, 102057.6, 101932.1, 101756.1, 101612, 101447.7, 101302, 101164.3,
  101809.6, 101694.2, 101585.2, 101448.1, 101259.3, 101055.1, 100851.7, 
    100667.4, 100476.3, 100313.4, 100159.1, 100005.6, 99896.99, 99816.83, 
    99743.02,
  100455.3, 101757.4, 101696.1, 101561.6, 101401.6, 101200.9, 100995.5, 
    100810.6, 100624.7, 100452.6, 100292.2, 100145.1, 100019, 99910.16, 
    99813.91,
  100612.6, 101557.5, 101800.8, 101670.1, 101513.8, 101337.8, 101151.1, 
    100957.5, 100774.9, 100598.1, 100437.5, 100281.3, 100134.2, 100013.7, 
    99911.83,
  100395.8, 101588.2, 101890.5, 101798.1, 101644.2, 101462.5, 101291.1, 
    101113, 100933, 100757.1, 100591.5, 100437.7, 100289.4, 100156.4, 100037.2,
  100449.2, 101027.3, 101810.5, 101878.5, 101754.1, 101586.7, 101414.9, 
    101249, 101078.7, 100908.7, 100748.3, 100587.5, 100438.6, 100299.2, 
    100174.3,
  100234.4, 99927.62, 100724, 101909.4, 101855.3, 101707.1, 101544.1, 
    101382.9, 101221.4, 101060.3, 100902, 100749.7, 100597.8, 100458.6, 
    100324.5,
  100206.5, 99436.52, 99264.49, 100968, 101938.7, 101819, 101658, 101508.9, 
    101353.1, 101203.7, 101050.6, 100903.2, 100759.4, 100618.8, 100488.4,
  100548.1, 99699.35, 99989.47, 100424, 101963.3, 101934.7, 101780.8, 
    101636.3, 101487.6, 101339.3, 101196.3, 101051.6, 100916.5, 100779.7, 
    100651.9,
  99360.93, 99103.15, 100329.9, 100630.1, 101153.9, 102006.1, 101896.8, 
    101744.3, 101602.4, 101470.2, 101328.3, 101195.3, 101060.1, 100936.2, 
    100811.3,
  99447.52, 97831.85, 97607.68, 98737.16, 100376.9, 101117.1, 102020.2, 
    101914.6, 101719.9, 101599.4, 101450.7, 101329.8, 101197.1, 101077.9, 
    100961.5,
  101800.8, 101763.8, 101763.4, 101661.7, 101523.5, 101374.9, 101258.7, 
    101132.3, 100983.9, 100847.2, 100712.9, 100593.5, 100506.9, 100402.7, 
    100291.6,
  100426.3, 101765.3, 101774.1, 101708.9, 101600.4, 101438.9, 101306.2, 
    101190.7, 101052.9, 100913.5, 100773.5, 100643, 100533.6, 100432.4, 
    100325.2,
  100574.5, 101532.6, 101815.2, 101749.9, 101647.8, 101514.3, 101365.3, 
    101245.9, 101117.3, 100980.9, 100841.2, 100705.3, 100575.4, 100466.1, 
    100361.8,
  100288.2, 101528.3, 101860.1, 101805.5, 101696.6, 101576.6, 101443.7, 
    101317.6, 101192.1, 101059, 100924.4, 100785, 100651, 100524.2, 100406.9,
  100303.9, 100926, 101741.6, 101853.5, 101757.2, 101631.9, 101506.4, 
    101382.5, 101258.8, 101129.2, 101001.4, 100867.8, 100730.4, 100595.1, 
    100467.4,
  100062.5, 99784.17, 100625.6, 101838.4, 101815.5, 101694.5, 101572, 
    101453.4, 101334.9, 101212.4, 101084, 100953.1, 100818.6, 100681.2, 100547,
  100005.7, 99264.16, 99130.27, 100863.4, 101863.2, 101757.2, 101635.2, 
    101520, 101401, 101286.1, 101165.6, 101039.6, 100911.8, 100778.8, 100644.9,
  100308.9, 99494.9, 99831.84, 100279.7, 101848.9, 101830.9, 101706.7, 
    101597.4, 101477.9, 101364.8, 101247.1, 101127.4, 101002.9, 100878.1, 
    100746.5,
  99088.23, 98863.84, 100134, 100455.1, 101013.4, 101889.1, 101786.5, 
    101658.9, 101551.1, 101441.9, 101326.7, 101215.3, 101095.2, 100974.8, 
    100855.5,
  99145.89, 97576.23, 97384.09, 98548.28, 100204.6, 100976.8, 101894.2, 
    101789.8, 101619.1, 101530.5, 101405.6, 101303.1, 101185.5, 101070.4, 
    100953.8,
  102015, 102038.4, 102049.6, 102031.8, 101992.2, 101922.7, 101859.4, 
    101812.6, 101749.8, 101697.3, 101642.1, 101578.4, 101545.8, 101528.1, 
    101456,
  100603.1, 102040.1, 102068.2, 102060.5, 102023.4, 101963.5, 101891.8, 
    101847.6, 101793.1, 101728.1, 101677.1, 101627.1, 101576.6, 101538.4, 
    101495.4,
  100704.4, 101732.6, 102082.9, 102088.8, 102035.6, 101987.9, 101923.9, 
    101873.9, 101830.6, 101775, 101713.9, 101658.3, 101607.1, 101563.9, 
    101524.8,
  100390.4, 101685.3, 102086.2, 102105, 102059.7, 102003.8, 101956.8, 
    101904.1, 101852.7, 101807.9, 101756.8, 101703, 101650.3, 101602.6, 
    101552.9,
  100374, 101041.4, 101936.5, 102104.7, 102090.2, 102017.9, 101970.6, 
    101928.5, 101877.6, 101832.4, 101787.6, 101741.1, 101689.1, 101639.1, 
    101591.5,
  100091.6, 99866.11, 100757.2, 102031.8, 102096.9, 102041.2, 101984.7, 
    101942.6, 101903.3, 101860.5, 101814.8, 101770.3, 101725, 101675.7, 
    101627.5,
  100003, 99317.22, 99242.48, 101021.2, 102085.5, 102037.6, 102001.9, 
    101959.6, 101906.3, 101875.6, 101840.4, 101797.1, 101756.9, 101713.6, 
    101667.6,
  100262.9, 99495.86, 99908.22, 100397.3, 102016.6, 102059.2, 102002.1, 
    101982.4, 101932.5, 101882.3, 101851.9, 101818.5, 101781.1, 101741.8, 
    101703.3,
  98996.19, 98823.83, 100157.7, 100522.7, 101124.6, 102072.7, 102033.1, 
    101980.6, 101953.9, 101907.4, 101866.3, 101837.5, 101803.5, 101771.1, 
    101732.5,
  99022.74, 97503.23, 97344.27, 98559.11, 100301.9, 101092.1, 102108, 102039, 
    101959.7, 101933.4, 101883.7, 101858.1, 101821.8, 101790.3, 101756.9,
  102381.2, 102363.8, 102335.7, 102273.7, 102194.2, 102102.7, 102015.5, 
    101937.4, 101852.6, 101776.1, 101699.3, 101621.5, 101554.8, 101496.4, 
    101442.4,
  100922.5, 102326.2, 102353.1, 102306, 102240.2, 102154.3, 102064.9, 
    101990.7, 101914.4, 101842.9, 101773.5, 101701.9, 101638.4, 101578.3, 
    101523.2,
  101006.7, 102010.7, 102357.1, 102338.7, 102267.4, 102193.3, 102111, 
    102040.7, 101976.7, 101904.9, 101837.9, 101769.6, 101702.9, 101645.1, 
    101597.2,
  100664.6, 101940.5, 102341.8, 102342.5, 102298.7, 102217.4, 102150.1, 
    102087.9, 102025.5, 101965.7, 101905.8, 101844.1, 101783.8, 101728.1, 
    101675.6,
  100601.6, 101264.3, 102149.9, 102329.5, 102308.9, 102232.5, 102175, 102126, 
    102071.2, 102016.1, 101964.5, 101908.8, 101850.5, 101793.7, 101745.4,
  100275.9, 100050.1, 100939.5, 102216.5, 102281.3, 102230.1, 102185.3, 
    102156.8, 102113.8, 102062.6, 102013.9, 101962.9, 101914.1, 101860.7, 
    101808.5,
  100126.8, 99445.91, 99385.83, 101169.3, 102221.1, 102207, 102175.9, 
    102160.2, 102134.5, 102101.6, 102058.2, 102014.6, 101966.3, 101923, 
    101874.6,
  100331.8, 99573.14, 99992.04, 100483.7, 102107.5, 102169.4, 102163.4, 
    102161.4, 102146.1, 102118.8, 102088.4, 102049.1, 102011.1, 101970.8, 
    101929,
  99033.3, 98871.66, 100203, 100559, 101160, 102117.5, 102141.5, 102138.8, 
    102147.8, 102130.8, 102101.3, 102077.7, 102041.6, 102008.8, 101972.9,
  99050.2, 97539.84, 97377.19, 98587.18, 100293.7, 101090.6, 102146.2, 
    102136.9, 102124, 102137.7, 102105.9, 102091.4, 102060.2, 102035.6, 102004,
  102414.8, 102386.1, 102311.7, 102210, 102083.5, 101956.8, 101827.2, 
    101699.2, 101553.9, 101414.5, 101280.8, 101146.1, 101019.7, 100892.7, 
    100763.6,
  100999.9, 102379.6, 102357.2, 102276.2, 102164.4, 102036.1, 101910.2, 
    101790.6, 101663.6, 101531.7, 101400.6, 101265.4, 101138.5, 101014.9, 
    100891.4,
  101113.6, 102085.4, 102387.7, 102317.8, 102211.6, 102094.4, 101972.1, 
    101860, 101743.6, 101621.6, 101496.7, 101371.5, 101247.3, 101125.5, 
    101005.3,
  100808.4, 102044, 102402.5, 102357.7, 102255.2, 102136.6, 102026.9, 
    101919.1, 101807.5, 101697.4, 101582.2, 101466.2, 101347.3, 101229.3, 
    101111.1,
  100776.6, 101399.6, 102229.2, 102370.1, 102299.6, 102171.4, 102063, 
    101964.4, 101863.4, 101756.8, 101652.6, 101544.9, 101435.1, 101322.8, 
    101208,
  100465.9, 100222.8, 101071, 102301.5, 102325.4, 102218.7, 102094.4, 
    102005.1, 101909.6, 101810.6, 101710.5, 101609.3, 101506.2, 101401.5, 
    101292.4,
  100342.5, 99635.58, 99525, 101289, 102314, 102245.7, 102123.4, 102035.8, 
    101946.8, 101857.1, 101762.9, 101665.6, 101570.8, 101470.5, 101369,
  100564.2, 99784.77, 100166.6, 100649, 102240, 102255.5, 102147.2, 102063.4, 
    101979.4, 101896.2, 101807.7, 101717.5, 101624.5, 101531.3, 101434.9,
  99271.81, 99096.49, 100395.9, 100726.5, 101315.2, 102205.8, 102147, 
    102071.3, 102000.5, 101927.9, 101846, 101764.6, 101677.1, 101589.6, 
    101498.7,
  99235.97, 97729.62, 97570.84, 98777.46, 100478.8, 101245.3, 102153.9, 
    102088.6, 102006.1, 101957.6, 101876.2, 101806.5, 101723.5, 101640.9, 
    101555.1,
  101866.8, 101830.8, 101763.7, 101671.3, 101568.3, 101438, 101314.3, 
    101192.7, 101063.7, 100934.3, 100812.3, 100687.5, 100575.8, 100468.7, 
    100358.7,
  100516.1, 101874.3, 101848.7, 101775, 101687.3, 101575.1, 101449.6, 
    101324.6, 101200.7, 101074.5, 100951.7, 100826.2, 100704.6, 100594.2, 
    100483.2,
  100678.1, 101662.6, 101949.1, 101883.9, 101794.8, 101688.4, 101577.8, 
    101457.8, 101336.2, 101212.6, 101091.3, 100971.2, 100849.3, 100732.7, 
    100622.3,
  100441.9, 101664.2, 102019.1, 101972.3, 101892, 101788.1, 101685.1, 
    101582.2, 101467.8, 101349.1, 101229.2, 101112.1, 100997, 100883.2, 
    100772.2,
  100474.2, 101072.7, 101913.9, 102028.2, 101977.4, 101893.8, 101786.7, 
    101682.9, 101581.4, 101472.4, 101359.1, 101246.6, 101134.5, 101024.4, 
    100915.7,
  100182.9, 99926.97, 100770.3, 102013.2, 102042.6, 101972.5, 101885.3, 
    101783.2, 101688.8, 101584.7, 101481.5, 101372.5, 101263.1, 101158.1, 
    101052.2,
  100113.6, 99389.53, 99257.48, 100998, 102057.7, 102024.4, 101952.5, 
    101866.7, 101779.6, 101683.5, 101586.8, 101485.9, 101387.7, 101284.5, 
    101184.3,
  100389.7, 99578.86, 99934.98, 100404.3, 102004.5, 102052.6, 101994.2, 
    101930.6, 101857, 101768.1, 101677.4, 101585.2, 101494.8, 101401, 101307.1,
  99121.84, 98910.06, 100197.2, 100521.4, 101114.9, 102054.9, 102019.1, 
    101959.7, 101908.2, 101840.9, 101753.9, 101673.8, 101587.9, 101505.8, 
    101418.2,
  99150.22, 97566.31, 97389.3, 98568.49, 100302.6, 101076.6, 102067.9, 
    102004.7, 101931.6, 101892, 101817.1, 101750, 101669.4, 101594.1, 101515.8,
  101752.2, 101709.1, 101680.2, 101619.8, 101554.8, 101459.9, 101390.3, 
    101328.8, 101269.2, 101212.1, 101160.2, 101118.8, 101077.5, 101034.8, 
    100984.4,
  100373, 101728.2, 101747.5, 101700.5, 101637.8, 101539.9, 101439, 101369.3, 
    101311.6, 101260.2, 101205.8, 101155.6, 101116, 101077.6, 101034.9,
  100525.6, 101507, 101828.2, 101782.6, 101716.1, 101625.4, 101533.4, 
    101436.8, 101365.6, 101301.8, 101249.6, 101196.7, 101152.3, 101119.8, 
    101080.3,
  100286, 101510.1, 101883, 101848.8, 101792.7, 101707.4, 101619.4, 101532.4, 
    101442.5, 101368.6, 101302.7, 101249.2, 101199.2, 101159.3, 101121.5,
  100328.3, 100939.5, 101794.9, 101915.8, 101874.9, 101800.4, 101703.1, 
    101617, 101531.7, 101446.2, 101374.8, 101304.7, 101246.2, 101197.7, 
    101158.9,
  100074.3, 99820.95, 100668.7, 101913, 101945.4, 101890, 101802.5, 101712, 
    101625.8, 101541.6, 101459.3, 101386.1, 101312.9, 101249.6, 101201.2,
  100018.9, 99304.31, 99192.48, 100929, 101986.4, 101950.6, 101881.4, 
    101802.8, 101717.5, 101633.4, 101552.8, 101475.6, 101400.8, 101329.1, 
    101264.2,
  100312.4, 99510.44, 99879.8, 100355, 101948.1, 101989.5, 101936.5, 
    101878.7, 101807.1, 101726.4, 101646.1, 101569.1, 101496.7, 101423.5, 
    101354.7,
  99084.72, 98885.86, 100168.4, 100504.1, 101087.7, 102009.5, 101982.4, 
    101919.5, 101866.4, 101808.3, 101734.5, 101665.4, 101589.1, 101521.6, 
    101453.1,
  99147.15, 97585.91, 97397.14, 98566.6, 100276.4, 101051.3, 102050.6, 
    102001.9, 101908.3, 101872.4, 101807.9, 101744.5, 101679.5, 101614.2, 
    101550.6,
  102210.5, 102195.5, 102178.2, 102122.8, 102040.3, 101946.2, 101855, 
    101764.8, 101671.6, 101585.2, 101509.8, 101429.2, 101356, 101282.9, 
    101210.3,
  100795.8, 102183.8, 102208.7, 102166.4, 102115.3, 102022.5, 101927.3, 
    101832.2, 101746.9, 101663.4, 101581, 101503.4, 101426.1, 101361, 101296.4,
  100919.1, 101922.7, 102257.5, 102228.1, 102165.2, 102091.3, 102005.3, 
    101919.4, 101832.1, 101747.2, 101659.8, 101578, 101504.5, 101434.3, 
    101374.9,
  100635.6, 101896.6, 102277.2, 102269.2, 102222, 102145.1, 102072.2, 
    101993.7, 101914.2, 101828.8, 101751.1, 101667.5, 101589.3, 101518.9, 
    101453.1,
  100637.7, 101284, 102152.4, 102294.5, 102271.5, 102207.3, 102131.8, 
    102053.9, 101981.3, 101902.8, 101823.7, 101748.1, 101667.4, 101593.7, 
    101527.4,
  100369.5, 100133.1, 101012.4, 102267.6, 102313.4, 102272.4, 102196.7, 
    102128.7, 102051.8, 101979.6, 101904.6, 101824.8, 101752.2, 101674.4, 
    101602.3,
  100283.6, 99589.35, 99503.66, 101269.3, 102334.2, 102309.1, 102249.3, 
    102186.5, 102118.9, 102044.9, 101973.4, 101902.1, 101826.4, 101754.9, 
    101683.7,
  100557.3, 99779.36, 100173.2, 100657, 102277, 102341.8, 102284.5, 102245.4, 
    102186.5, 102117.9, 102046.2, 101973.7, 101905, 101834.3, 101766.3,
  99300.81, 99117.45, 100429.4, 100784.7, 101384.4, 102332.4, 102320.4, 
    102264.7, 102229.7, 102175.1, 102108.3, 102044.1, 101975, 101909.9, 
    101845.3,
  99337.59, 97818.7, 97642.96, 98831.09, 100555.1, 101356.2, 102373.5, 
    102338.8, 102262.2, 102233.1, 102166.7, 102113.2, 102045, 101983.5, 
    101919.7,
  102455.2, 102563.2, 102627.2, 102662.2, 102662.5, 102641.3, 102639.6, 
    102632.2, 102611.5, 102580.7, 102538.4, 102477.8, 102409.2, 102338.1, 
    102258.2,
  101036.8, 102530.8, 102633, 102677.9, 102685.9, 102676.2, 102673.3, 
    102670.7, 102658.3, 102640.4, 102600.7, 102548.7, 102481.4, 102411.1, 
    102332.9,
  101154.7, 102224.7, 102639.8, 102695.9, 102700.9, 102699.4, 102704.1, 
    102706.1, 102698, 102683.4, 102652.5, 102605.2, 102544.3, 102473.1, 
    102399.2,
  100833.6, 102169.9, 102623, 102696.2, 102735.4, 102711.6, 102722.7, 
    102734.5, 102726.8, 102714.1, 102690.8, 102652.3, 102600.8, 102535.5, 
    102463,
  100806, 101513.6, 102451.7, 102688.7, 102739.3, 102738.5, 102724.4, 
    102750.6, 102751.4, 102741.3, 102719.2, 102688.7, 102642.5, 102586.4, 
    102518.5,
  100496.8, 100320.9, 101257.2, 102595.4, 102730.8, 102752.4, 102737, 
    102753.5, 102763.3, 102759.5, 102741.1, 102715.7, 102679, 102625.8, 
    102566.6,
  100391.2, 99759.95, 99749.13, 101557.3, 102687, 102737.4, 102750.5, 
    102763.2, 102774.9, 102767.6, 102754.4, 102730.6, 102699.4, 102658.6, 
    102602.3,
  100614.1, 99901.66, 100379.6, 100912.7, 102585.1, 102712.6, 102746.5, 
    102762, 102771.3, 102767.7, 102761.3, 102743.5, 102717.7, 102680.9, 
    102631.1,
  99365.81, 99224.2, 100574.7, 100965.2, 101647.1, 102670.1, 102735.5, 
    102754, 102769.9, 102761.7, 102756.4, 102744.6, 102719.5, 102689.9, 
    102651.1,
  99387.19, 97909.98, 97773.15, 99000.35, 100780.3, 101611.8, 102726.3, 
    102748.6, 102750.5, 102760.1, 102746.2, 102743, 102721.5, 102696.7, 
    102659.9,
  101888, 101983.8, 102037.9, 102083.6, 102114.9, 102125.1, 102150.4, 
    102178.7, 102202.3, 102213.5, 102217.8, 102213.3, 102204.6, 102192.5, 
    102178.1,
  100511.9, 101965.5, 102077.2, 102130.7, 102171.2, 102200.7, 102237.6, 
    102274.3, 102306, 102327.2, 102339.7, 102345.8, 102345.8, 102338.5, 
    102328.4,
  100655.3, 101703.4, 102118.3, 102173.6, 102227.3, 102268, 102311.9, 
    102355.9, 102396.6, 102427, 102449.1, 102464, 102472.9, 102470.1, 102461.8,
  100374.9, 101672.4, 102137.8, 102207.9, 102276.4, 102327.2, 102376, 
    102425.9, 102478.2, 102516.9, 102546.2, 102565.1, 102578.5, 102584.8, 
    102583.7,
  100381.4, 101072.3, 101999.5, 102249.7, 102312.4, 102371.2, 102427.5, 
    102484.6, 102545.8, 102588.2, 102623, 102648.2, 102667.1, 102679.6, 
    102683.9,
  100106, 99947.2, 100860.2, 102193.6, 102341.5, 102398.6, 102466.8, 
    102530.4, 102596, 102645.1, 102687.4, 102719.2, 102748.3, 102764.2, 
    102774.1,
  100056.7, 99433.2, 99439, 101215.4, 102350.8, 102422.7, 102493, 102565.8, 
    102637.1, 102696, 102738.8, 102777, 102811, 102832.9, 102847.6,
  100305.4, 99604.79, 100091.7, 100630.4, 102271.2, 102427.6, 102507.2, 
    102586.2, 102665.5, 102729.7, 102778.6, 102823.7, 102858.6, 102889.9, 
    102907.3,
  99127.98, 98982.3, 100306.2, 100714, 101392.8, 102406.5, 102528.1, 
    102594.6, 102679.6, 102760.6, 102808.9, 102855.4, 102894.1, 102925.4, 
    102949.9,
  99182.17, 97728, 97598.06, 98791.74, 100573.6, 101345.1, 102524.9, 
    102610.9, 102676.5, 102778.6, 102828, 102876.4, 102918.1, 102954, 102979.6,
  100833.1, 100866.4, 100903.5, 100908.5, 100935.8, 100958, 100979, 101013.4, 
    101048.6, 101076.9, 101096, 101105.5, 101110.4, 101109.1, 101100,
  99511.9, 100898.5, 100997.5, 101012.3, 101038.1, 101068.3, 101101.7, 
    101139.2, 101175.2, 101207.5, 101234, 101254.4, 101267.2, 101278.3, 101281,
  99703.76, 100709.8, 101107.5, 101123.1, 101150.4, 101181.5, 101216.6, 
    101257.5, 101298.5, 101338.3, 101371.8, 101402.4, 101425.2, 101445.9, 
    101457.9,
  99486.51, 100745.4, 101189.2, 101223.4, 101256.6, 101285.9, 101330.1, 
    101372.8, 101418.5, 101463.1, 101503.8, 101540.6, 101569.4, 101596.2, 
    101620.3,
  99544.97, 100223, 101128.5, 101345.5, 101374.3, 101402.2, 101445.4, 
    101489.2, 101536.6, 101585.1, 101631, 101667.8, 101701.9, 101736.1, 
    101766.7,
  99326.86, 99169.48, 100063.2, 101359.4, 101477.5, 101506.4, 101544.6, 
    101599.4, 101652.6, 101706.4, 101754, 101795.1, 101834.4, 101872, 101906.2,
  99319.53, 98712.55, 98715.84, 100444.7, 101543, 101597.9, 101634.5, 
    101703.5, 101760.2, 101817.3, 101869.8, 101914.3, 101957, 101995.8, 
    102035.7,
  99628.76, 98924.55, 99393.33, 99919.68, 101526.4, 101681.1, 101714.7, 
    101791.1, 101849.7, 101910.9, 101970.2, 102021.4, 102068, 102110.2, 102154,
  98515.85, 98351.07, 99637.64, 100041.1, 100704, 101722.7, 101795.7, 
    101863.7, 101919.8, 101988.1, 102055.2, 102113.9, 102163.1, 102209.5, 
    102258.1,
  98628.6, 97175.6, 97004.71, 98159.95, 99905.02, 100710, 101842.9, 101936.6, 
    101961, 102044.4, 102117.5, 102186.6, 102239.6, 102294.1, 102345.6,
  101502, 101461.8, 101399.1, 101314.2, 101221.9, 101113.3, 100989.5, 
    100869.2, 100754.3, 100644.8, 100548.3, 100456.4, 100371.1, 100288.9, 
    100212.9,
  100167, 101499.4, 101495.6, 101423.7, 101347.4, 101251.2, 101141.5, 101036, 
    100940.2, 100845.1, 100757.9, 100673.1, 100593.8, 100519.7, 100450.3,
  100312.7, 101266.8, 101580.5, 101515.5, 101447.6, 101365.1, 101279.6, 
    101187.5, 101104.3, 101023.6, 100946.8, 100874.3, 100800.6, 100732.2, 
    100669,
  100058.6, 101256.5, 101625.2, 101584.1, 101535.1, 101470.2, 101396.2, 
    101321.7, 101251.6, 101179.7, 101113.2, 101049.4, 100985.2, 100924.6, 
    100869.4,
  100064.5, 100666.8, 101515.5, 101642.3, 101602.7, 101553.1, 101494.4, 
    101430.8, 101370.5, 101312.4, 101254.7, 101202.1, 101149.4, 101099.1, 
    101053.7,
  99775.09, 99543.02, 100383.4, 101619, 101659.5, 101618.6, 101574.9, 101525, 
    101477.6, 101431.1, 101383.6, 101339.5, 101298.3, 101258.3, 101221.1,
  99683, 99010.09, 98925.28, 100635, 101682, 101670.5, 101630.6, 101593.6, 
    101554.3, 101518.9, 101487.3, 101453.3, 101424.7, 101397.7, 101373,
  99933.91, 99174.61, 99564.84, 100034.8, 101616.8, 101701.9, 101677.9, 
    101656.5, 101629.5, 101601.9, 101576.9, 101558.5, 101540.9, 101524.6, 
    101510.9,
  98740.29, 98544.37, 99826.21, 100174.5, 100759.4, 101689.3, 101698.5, 
    101680.2, 101676.5, 101671.9, 101658.1, 101649.3, 101639.3, 101634.8, 
    101635,
  98837.78, 97344.41, 97157.56, 98286.98, 99992.7, 100769.2, 101777.5, 
    101757, 101717.1, 101733.8, 101725.7, 101732.1, 101728.4, 101731.2, 
    101741.6,
  101731.4, 101800.8, 101829.8, 101841.5, 101842.2, 101820.6, 101784.6, 
    101750.7, 101710.4, 101659.5, 101605, 101542.9, 101477.6, 101405.1, 
    101329.5,
  100339.2, 101794.6, 101871.2, 101892.1, 101899.8, 101885, 101861.3, 
    101837.6, 101810.9, 101772.9, 101729.5, 101671.7, 101609.9, 101545.9, 
    101477.1,
  100455, 101502.4, 101893.7, 101922.5, 101934.3, 101925, 101919.3, 101907.5, 
    101891.3, 101865.7, 101832.2, 101788.9, 101735.6, 101670.9, 101604.6,
  100144.9, 101449.6, 101889.5, 101937.9, 101962.7, 101965.3, 101955.2, 
    101956.3, 101953.6, 101942.4, 101920.6, 101887.6, 101844, 101792.3, 
    101735.3,
  100120.9, 100807.6, 101718.4, 101944.3, 101974, 101984.9, 101988.1, 
    101984.1, 101987.4, 101986.8, 101979.7, 101961.8, 101932.4, 101893.6, 
    101843.2,
  99816.48, 99654.16, 100545.9, 101850.3, 101959.1, 101982.6, 101999, 
    102016.8, 102027.7, 102032.5, 102026.9, 102013.7, 101994.1, 101966.8, 
    101933.3,
  99721.88, 99100.1, 99078.38, 100848.8, 101931, 101961.3, 101970.4, 
    101995.1, 102016.1, 102042.3, 102056.8, 102056.9, 102041.2, 102020.1, 
    101993.1,
  99985.19, 99240.29, 99697.38, 100219.4, 101844.2, 101962.8, 101986.2, 
    102016.2, 102032.9, 102040.9, 102043.4, 102064, 102069.5, 102061.1, 
    102044.3,
  98809.77, 98630.97, 99901.48, 100260, 100887.6, 101874, 101920.7, 101970.9, 
    102014.8, 102058.8, 102048.5, 102054.5, 102064.6, 102066.3, 102062.4,
  98884.46, 97410.9, 97244.37, 98393.27, 100106.4, 100868.6, 101934.6, 
    101955.1, 101972, 102036.9, 102064, 102078.2, 102079.8, 102085.1, 102080.9,
  101337.8, 101377.5, 101414.7, 101425.1, 101435.9, 101428.9, 101410.8, 
    101399.7, 101385.1, 101362.9, 101343.4, 101312.5, 101280.4, 101239, 
    101191.5,
  99943.66, 101353.7, 101452.2, 101475.8, 101494.1, 101488.1, 101475.1, 
    101474.9, 101472.1, 101466.1, 101454, 101434.7, 101408.2, 101376.9, 
    101338.4,
  100088.7, 101096, 101491.6, 101514.8, 101541.7, 101541.3, 101541, 101546, 
    101549.3, 101550.6, 101550.5, 101544.7, 101533.2, 101513.4, 101486,
  99820.12, 101080.4, 101514.8, 101551.6, 101584.6, 101595.8, 101601.7, 
    101611.8, 101621.3, 101632, 101642.1, 101645.6, 101642.9, 101632.6, 
    101617.7,
  99837.65, 100500.9, 101385.6, 101587.5, 101612.1, 101632.5, 101653.5, 
    101664.4, 101680.9, 101698.3, 101714.4, 101725.3, 101731.6, 101733.1, 
    101727.4,
  99582.54, 99397.13, 100265.8, 101546.9, 101641.8, 101661.2, 101680.6, 
    101698.5, 101718, 101744.8, 101767.1, 101790.5, 101808.4, 101818.8, 
    101821.4,
  99535.09, 98896.96, 98850.57, 100579.2, 101655.1, 101685.5, 101699.3, 
    101721.6, 101742.4, 101779.6, 101809.5, 101839.8, 101863.3, 101882.2, 
    101896.1,
  99815.76, 99080.27, 99505.16, 100003.8, 101595.5, 101708.5, 101719.9, 
    101743.6, 101770.7, 101801.3, 101838.7, 101875.7, 101904.7, 101928.1, 
    101948,
  98648.58, 98482.55, 99777.43, 100121.3, 100726.3, 101701.8, 101750.2, 
    101761.2, 101793.8, 101823.5, 101859.2, 101899, 101928.9, 101955.3, 
    101979.7,
  98727.11, 97264.12, 97111.95, 98263.18, 99984.73, 100723.2, 101763.2, 
    101789.2, 101804.1, 101839.2, 101867, 101906.5, 101940.3, 101974, 102000.9,
  100240.6, 100232.8, 100210.6, 100212.4, 100213.8, 100227.5, 100243.8, 
    100268.1, 100303.4, 100345.1, 100390.5, 100459.6, 100522.4, 100595.5, 
    100647.6,
  98775.59, 100146.2, 100163.4, 100183.1, 100222.3, 100252.5, 100281.9, 
    100325, 100371.1, 100424.9, 100471.4, 100512.7, 100551.8, 100607.8, 
    100657.7,
  98884.16, 99847.03, 100202.3, 100241.1, 100287.9, 100333.7, 100381.1, 
    100430.1, 100469.7, 100508, 100540.2, 100574.2, 100598.6, 100626.6, 
    100649.8,
  98656.7, 99846.62, 100271.3, 100316.1, 100367.4, 100428.7, 100483.6, 
    100529.5, 100575.5, 100620.7, 100661.3, 100700.4, 100732.7, 100760.1, 
    100781.2,
  98718.2, 99329.64, 100210.7, 100427.7, 100481.3, 100534.2, 100583.5, 
    100628.3, 100676.6, 100722.8, 100763.5, 100800.1, 100828.6, 100851.7, 
    100878,
  98527.48, 98325.95, 99185.14, 100462.2, 100581.4, 100620.4, 100665.4, 
    100714.2, 100760.8, 100809.1, 100851.4, 100887, 100923.7, 100959.5, 
    100993.2,
  98547.02, 97903.12, 97854.91, 99568.49, 100654.7, 100704, 100741.2, 
    100788.5, 100837.1, 100885.8, 100925.3, 100966.1, 101004.2, 101041.6, 
    101081.1,
  98885.86, 98147.46, 98572.3, 99062.95, 100640, 100769.8, 100805.9, 
    100852.6, 100903.5, 100949, 100995.3, 101038.6, 101081, 101123.2, 101166.2,
  97786.11, 97598.98, 98874.28, 99240.22, 99837.89, 100796.5, 100858.1, 
    100898.9, 100958.6, 101015, 101060.9, 101108.7, 101151.2, 101196.9, 
    101241.4,
  97915.29, 96456.5, 96268.93, 97411.95, 99117.42, 99865.71, 100923.9, 
    100965.3, 100995.2, 101075.4, 101120.1, 101177.7, 101221.5, 101268.7, 
    101318.6,
  100628.1, 100485.3, 100325.4, 100107.6, 99897.49, 99620.02, 99347.8, 
    99100.14, 98866.97, 98674.27, 98558.84, 98501.82, 98490.2, 98533.6, 
    98639.93,
  99306.17, 100547.2, 100430, 100216.6, 99997.88, 99759.85, 99526.88, 
    99323.46, 99156.34, 99022.34, 98912.28, 98831.58, 98804.28, 98834.84, 
    98911.55,
  99511.2, 100385.9, 100567.4, 100380, 100184.2, 99965.53, 99755.75, 
    99572.22, 99412.25, 99286.12, 99189.08, 99130.21, 99106.62, 99114.39, 
    99154.87,
  99328.7, 100449.9, 100682.6, 100525.6, 100345.5, 100155.7, 99972.94, 
    99813.09, 99673.01, 99559.17, 99470.37, 99403.87, 99372.36, 99372.96, 
    99407.86,
  99425.83, 99949.18, 100663.4, 100681.9, 100522.1, 100359.9, 100195.5, 
    100045.2, 99911.84, 99801.32, 99713.04, 99648.91, 99615.61, 99611.01, 
    99630.59,
  99237.09, 98907.49, 99632.77, 100752, 100677.8, 100535.2, 100391.5, 
    100258.9, 100134.6, 100033, 99944.99, 99880.33, 99840.2, 99828.43, 
    99838.91,
  99213.02, 98437, 98250.7, 99868.48, 100803, 100696.7, 100558, 100442.5, 
    100329, 100238.1, 100154.1, 100094.4, 100051.2, 100035.6, 100033.9,
  99532.91, 98677.01, 98946.85, 99342.8, 100820.4, 100816.4, 100692.7, 
    100598.8, 100499.1, 100418.3, 100345.2, 100288.8, 100247.6, 100225.7, 
    100221.7,
  98341.62, 98080.69, 99272.27, 99545.31, 100032.9, 100872.9, 100800.6, 
    100705.4, 100635.5, 100575.8, 100514.6, 100466.7, 100426.2, 100402.1, 
    100396.4,
  98390.32, 96836.79, 96588.91, 97680.15, 99286.79, 99986.79, 100911.6, 
    100854.6, 100743.9, 100719.1, 100654.2, 100617.4, 100581.2, 100556.9, 
    100551.6,
  101381.8, 101246.6, 101116.9, 100919.3, 100761.7, 100567.8, 100385.5, 
    100233.7, 100078.6, 99936.82, 99797.34, 99633.22, 99446.77, 99234.24, 
    99006.51,
  100065.5, 101337.5, 101235.6, 101061.4, 100887.2, 100705.1, 100522.7, 
    100349.6, 100190.3, 100055.3, 99921.28, 99777.05, 99620.49, 99463.27, 
    99316.87,
  100248, 101160.1, 101362.4, 101222.1, 101047, 100853.5, 100665.2, 100505.9, 
    100358.6, 100218, 100087.2, 99962.1, 99835.48, 99708.67, 99583.89,
  100048.2, 101212.8, 101462.3, 101348.8, 101187.8, 101007.1, 100831.9, 
    100674.9, 100522.5, 100386.7, 100266.5, 100152.4, 100044.9, 99935.7, 
    99842.56,
  100127.3, 100675.9, 101419.9, 101463.5, 101321.9, 101167.5, 101001.5, 
    100846.6, 100706.4, 100578.2, 100458.1, 100353.3, 100249.8, 100162.5, 
    100080.3,
  99944.98, 99602.08, 100355.4, 101512.9, 101446.8, 101302.3, 101158.5, 
    101016.2, 100884.5, 100760.3, 100647.7, 100543.8, 100453.3, 100376.8, 
    100307.5,
  99937.44, 99130.98, 98929.94, 100606.1, 101557.2, 101444.4, 101300.2, 
    101173.3, 101051.6, 100938.8, 100835.1, 100738.1, 100659.6, 100584.9, 
    100526.5,
  100286.5, 99395.88, 99658.21, 100073.8, 101583, 101569.9, 101432.9, 
    101322.8, 101204.5, 101101.7, 101000.7, 100916.3, 100841.5, 100778.8, 
    100724.4,
  99121.97, 98839.98, 100005.7, 100283.4, 100791, 101643.5, 101545, 101432.5, 
    101332, 101244.8, 101153, 101077.8, 101006.6, 100952.2, 100901.4,
  99219.62, 97592.54, 97331.79, 98433.78, 100047.5, 100764.5, 101674.4, 
    101581.7, 101428.6, 101368.2, 101273.1, 101213, 101145.8, 101092.4, 
    101043.9,
  102199, 102093.9, 101972.5, 101796.8, 101640.9, 101520.2, 101394.3, 
    101253.5, 101111.1, 100982.3, 100841.5, 100683.1, 100500.4, 100300.4, 
    100085.5,
  100774.2, 102113, 102044.9, 101877.5, 101684, 101527.5, 101388.2, 101262.1, 
    101123.1, 100987.6, 100852.2, 100702, 100532.6, 100349.8, 100152.4,
  100904.2, 101853, 102086.6, 101949.7, 101763, 101564.8, 101409.4, 101277.4, 
    101142.1, 101007.6, 100874.1, 100733.2, 100576, 100408.9, 100229.8,
  100649.7, 101855.2, 102125, 102028.1, 101844.6, 101621.7, 101436.6, 
    101298.6, 101161.9, 101026.6, 100899.8, 100769.5, 100623.4, 100473.4, 
    100311,
  100671.8, 101261.2, 102024, 102087.4, 101937.9, 101715.4, 101504.8, 
    101340.6, 101196.6, 101058.7, 100925.2, 100804.6, 100671.3, 100532.5, 
    100388.6,
  100436.3, 100128.8, 100924.2, 102078.9, 102004.5, 101813.6, 101593.4, 
    101410.9, 101251.1, 101100, 100964.8, 100836.9, 100712, 100586.6, 100453.8,
  100380.9, 99606.4, 99433.14, 101148.4, 102071.6, 101914.8, 101701, 
    101499.1, 101319.3, 101158.4, 101013.6, 100880.1, 100755.5, 100642.3, 
    100522.4,
  100694.3, 99847.03, 100134.6, 100564.7, 102083.4, 102014, 101811.8, 
    101619.2, 101428.3, 101251.2, 101086.9, 100946.6, 100820.2, 100704.8, 
    100597.8,
  99483.73, 99238.59, 100462.4, 100747.7, 101262.9, 102094.2, 101925.9, 
    101725.9, 101532, 101361.6, 101181.9, 101035.6, 100905.7, 100791.2, 
    100689.3,
  99553.94, 97945.26, 97727.31, 98861.34, 100479, 101200.8, 102047.4, 
    101891.1, 101636.9, 101483.3, 101297.1, 101151.2, 101009, 100895.4, 
    100794.1,
  102345.2, 102391.3, 102406.9, 102382.7, 102353.9, 102324.8, 102303.4, 
    102274.3, 102241.4, 102221.6, 102181.7, 102132, 102046.7, 101944, 101838.6,
  100908.5, 102381.4, 102432.6, 102422.1, 102381.2, 102332.7, 102307.8, 
    102285, 102248.8, 102226.4, 102182.8, 102126.9, 102051.8, 101950.9, 
    101840.9,
  101038, 102094.1, 102448.8, 102453.3, 102408.7, 102340.5, 102324.4, 102297, 
    102259.5, 102227.1, 102188.5, 102133.4, 102054.8, 101958.5, 101851.5,
  100735.3, 102052.6, 102455.9, 102478, 102441.2, 102351.6, 102325.9, 
    102301.8, 102265.9, 102230.9, 102190.7, 102137.7, 102060, 101965.9, 
    101861.3,
  100727.3, 101417.5, 102310.8, 102485.1, 102476.1, 102378.8, 102342.1, 
    102313.4, 102275.6, 102241, 102200.1, 102151.9, 102076.4, 101984.7, 
    101880.7,
  100444.1, 100231.7, 101147.3, 102435.5, 102499.9, 102417.4, 102348.8, 
    102327.4, 102291, 102251.5, 102204.4, 102157.1, 102086.2, 101998.7, 
    101896.7,
  100360.4, 99673.36, 99621.41, 101425.9, 102509.2, 102462.1, 102371.9, 
    102340.4, 102301.2, 102262.7, 102217.8, 102165.9, 102100.2, 102017.3, 
    101919.9,
  100617.7, 99852.57, 100293.6, 100800.5, 102442, 102494.5, 102408.3, 
    102354.3, 102319, 102278.4, 102228.8, 102175.3, 102112.3, 102036.3, 
    101944.2,
  99356.31, 99188.57, 100543.7, 100903.1, 101534.1, 102500.5, 102449.1, 
    102372.3, 102332.8, 102291.6, 102243, 102191.4, 102127.7, 102058.9, 
    101973.6,
  99395.66, 97862.38, 97709.78, 98941.26, 100709, 101503.4, 102522.2, 
    102426.5, 102338.1, 102311.8, 102254.1, 102207.9, 102144, 102078.4, 
    102000.6,
  102058.6, 102106.1, 102140.5, 102163.5, 102178.9, 102163.2, 102176.5, 
    102216.1, 102260.1, 102319.8, 102390.1, 102452, 102513.8, 102579.6, 
    102652.4,
  100634.7, 102098.5, 102169.2, 102188.8, 102207.3, 102196.3, 102213.8, 
    102262.6, 102301, 102358.4, 102442.1, 102520.5, 102600.9, 102663.7, 
    102715.4,
  100770.1, 101823.8, 102196.5, 102216.4, 102227.2, 102215.2, 102243.1, 
    102290.8, 102336.1, 102411, 102496.2, 102570.1, 102643.1, 102703.7, 
    102770.1,
  100457.4, 101766.8, 102195.3, 102220.4, 102237.3, 102245, 102271.8, 
    102323.3, 102367.8, 102452.7, 102535, 102621.1, 102686.4, 102754.3, 
    102816.8,
  100451.9, 101133.1, 102047.1, 102240.8, 102259.7, 102265.2, 102296.5, 
    102346.3, 102396.2, 102480.6, 102561.7, 102652.3, 102721.9, 102789.7, 
    102847.9,
  100145, 99945.53, 100854.6, 102173.4, 102274.2, 102286.2, 102318.4, 
    102363.5, 102409.4, 102498.6, 102577.3, 102677, 102747.9, 102815.9, 
    102870.8,
  100077.8, 99395.75, 99368.02, 101150.7, 102287.4, 102313.4, 102332.7, 
    102371.6, 102421.8, 102509.3, 102587.8, 102684.8, 102763.4, 102833.5, 
    102883.8,
  100319.6, 99565.45, 100025.1, 100540.5, 102207.8, 102328.5, 102345.1, 
    102373, 102426.8, 102511.6, 102593.7, 102687.6, 102772.1, 102833.2, 
    102885.8,
  99076.3, 98913.8, 100253.1, 100641.8, 101318.8, 102315.2, 102357.5, 
    102368.4, 102430, 102508.5, 102594.8, 102681.9, 102766.6, 102834.1, 
    102888.1,
  99133.86, 97624.18, 97462.28, 98666.17, 100489.5, 101242.1, 102374, 
    102373.2, 102412.3, 102503.4, 102585.5, 102673.3, 102755.3, 102828.3, 
    102876.2,
  101520.7, 101510.1, 101502.8, 101484.9, 101454.6, 101402, 101374.1, 
    101351.3, 101331, 101330.6, 101352.7, 101384.6, 101409, 101451.6, 101503.2,
  100148.9, 101571.9, 101577.7, 101536.1, 101481.3, 101432.8, 101405.9, 
    101387.6, 101391, 101402.4, 101407.1, 101414.7, 101453.4, 101515.6, 
    101603.8,
  100304.8, 101304, 101614.2, 101587.1, 101545.7, 101491.5, 101446.1, 
    101421.4, 101411.9, 101409, 101429, 101479.9, 101524.9, 101575.3, 101672.3,
  100023, 101270, 101645.6, 101635.6, 101594.1, 101541.1, 101497.5, 101478.3, 
    101482.5, 101469.9, 101505.9, 101534.8, 101575.7, 101653.5, 101753.2,
  100055.8, 100689.7, 101540.2, 101688.7, 101654.2, 101603.9, 101563.4, 
    101536.8, 101526, 101512.4, 101549.9, 101573.8, 101639.9, 101721.6, 
    101829.5,
  99804.92, 99550.8, 100386.4, 101649.2, 101694.8, 101650.9, 101607.4, 
    101586.3, 101565.2, 101568.6, 101600.6, 101637.9, 101701.9, 101803.5, 
    101916.7,
  99740.93, 99025.8, 98918.59, 100656.3, 101714.5, 101691.4, 101643.1, 
    101616.8, 101603.6, 101613.9, 101650.7, 101702.9, 101783.2, 101876.8, 
    101992.6,
  100033.2, 99223.16, 99598.77, 100065.2, 101646.7, 101710, 101664.7, 
    101651.1, 101655.5, 101669.2, 101716.2, 101776.6, 101849.9, 101948.3, 
    102063.7,
  98841.42, 98603.93, 99864.59, 100203, 100782.3, 101719.3, 101717.9, 
    101703.6, 101713, 101734.1, 101784.7, 101844.2, 101915.7, 102008.2, 
    102121.6,
  98924.09, 97375.74, 97157.99, 98281.26, 99993.72, 100756.5, 101783.4, 
    101778.8, 101757.3, 101803.6, 101838.2, 101902.7, 101972.4, 102064.5, 
    102181.2,
  101256.5, 101089.8, 100928.4, 100753.1, 100584.8, 100420.1, 100275.6, 
    100119, 99980.58, 99835.16, 99724.14, 99610.83, 99522.17, 99450.35, 
    99414.16,
  99943.82, 101215.9, 101099.2, 100930.6, 100754.3, 100566.1, 100407.6, 
    100265.9, 100129.4, 99991.38, 99879.69, 99775.27, 99671.43, 99602.85, 
    99562.49,
  100188.6, 101076.2, 101266.3, 101102, 100932.1, 100742.2, 100568.3, 
    100416.5, 100282.1, 100154.6, 100037.3, 99937.77, 99846.82, 99785.69, 
    99744.71,
  100008.9, 101148.8, 101405.1, 101260.1, 101103.7, 100921.5, 100749.3, 
    100593.8, 100451.4, 100324.4, 100208.6, 100114.8, 100030.1, 99963.68, 
    99916.41,
  100123.3, 100655.6, 101390.6, 101412.1, 101269.4, 101099.9, 100937.6, 
    100776.8, 100639.8, 100509.1, 100398, 100296.4, 100212.4, 100144.8, 
    100109.3,
  99936.76, 99594.29, 100334.6, 101497.7, 101433.6, 101272.9, 101124.1, 
    100975.2, 100832.2, 100701.5, 100590.1, 100488, 100404.7, 100338, 100303.8,
  99924.7, 99130.7, 98929.62, 100616.3, 101562, 101449.3, 101288, 101150.4, 
    101013.1, 100893.5, 100780.8, 100674.6, 100596.4, 100537.8, 100495.6,
  100276.3, 99408.82, 99674.23, 100105.8, 101596.8, 101595.6, 101441.7, 
    101327.3, 101191.3, 101078.1, 100962.9, 100863.8, 100793.8, 100730.7, 
    100678,
  99102.23, 98827.44, 100017.7, 100328.1, 100813.1, 101675.8, 101560.8, 
    101447.7, 101335.7, 101239.3, 101123.6, 101043.2, 100970.7, 100903.2, 
    100849.3,
  99199.59, 97601.77, 97333.16, 98448.48, 100062.9, 100787.6, 101710.7, 
    101633.5, 101454.9, 101383.9, 101272, 101206.2, 101117.9, 101053.9, 
    101007.8,
  101845.6, 101710.5, 101594, 101438.8, 101297.5, 101151.4, 101011.3, 
    100848.5, 100677.7, 100500.4, 100380.5, 100247, 100141.4, 100029.9, 
    99898.23,
  100483.3, 101791, 101720.3, 101586.5, 101432.1, 101262, 101120.1, 100995.9, 
    100863.1, 100719.6, 100562.5, 100422.6, 100288.2, 100176.4, 100072.1,
  100679.1, 101615.4, 101840.8, 101726.2, 101589.3, 101423.9, 101281.1, 
    101145.5, 101015.2, 100872.4, 100746.5, 100620.5, 100503.2, 100374.8, 
    100262.4,
  100447.1, 101650.4, 101939.1, 101848.6, 101716.3, 101563.7, 101410.9, 
    101280.2, 101161.4, 101042.5, 100923.9, 100803, 100689.3, 100578.5, 
    100474.2,
  100514.8, 101088.2, 101883.9, 101959.5, 101843.1, 101702.1, 101560.9, 
    101423.2, 101300.3, 101189.5, 101083.8, 100981.2, 100880.1, 100780.7, 
    100686.3,
  100292.6, 99980.25, 100794, 102003.8, 101965.3, 101832.5, 101699.9, 
    101570.6, 101447.9, 101336.2, 101234.9, 101141.5, 101051.4, 100964.4, 
    100878.1,
  100255.5, 99488.45, 99321.7, 101062.1, 102068.6, 101968.8, 101834.5, 
    101712.7, 101591.5, 101486.4, 101380.7, 101289.3, 101207.1, 101130.9, 
    101056.2,
  100576.9, 99741.57, 100053.6, 100514.9, 102073.9, 102087.2, 101967.8, 
    101861.9, 101739.5, 101637.5, 101535.9, 101446.2, 101363.2, 101288.7, 
    101219.4,
  99363.96, 99119.67, 100373.5, 100709.1, 101252.9, 102155.3, 102073.5, 
    101969.6, 101875.6, 101780.6, 101682.5, 101598.4, 101516.9, 101445.5, 
    101382.3,
  99435.57, 97833.73, 97626.41, 98774.57, 100471.2, 101227, 102215.2, 
    102126.5, 101974.6, 101917.9, 101811.1, 101738.9, 101658.3, 101593.9, 
    101530.4,
  102346.2, 102159.8, 101986.8, 101788.6, 101653.9, 101544.1, 101497.1, 
    101436.1, 101383.7, 101320.5, 101305.6, 101293.8, 101307.7, 101297.5, 
    101269,
  100950.4, 102193, 102064.7, 101902.5, 101736.4, 101603.4, 101521.3, 
    101460.8, 101406.7, 101373.6, 101340, 101307.7, 101292.5, 101267.3, 
    101289.8,
  101133.5, 102020, 102188.3, 102043.2, 101870.7, 101708.1, 101604.2, 
    101534.1, 101470.4, 101423.5, 101392.9, 101378.5, 101360.8, 101334.4, 
    101303.4,
  100880.8, 102070.7, 102304.7, 102182.7, 102018.5, 101860.2, 101731.3, 
    101643.6, 101574.3, 101523, 101485.6, 101458, 101431.1, 101409.9, 101392,
  100931.5, 101504.4, 102267.5, 102310.1, 102179.4, 102022.1, 101883.8, 
    101781.5, 101701.3, 101641.9, 101590, 101562.2, 101536.3, 101512.3, 
    101488.2,
  100696.9, 100374, 101170.1, 102352.5, 102312.3, 102172.3, 102043.8, 
    101936.4, 101845.7, 101778.6, 101719.3, 101675.4, 101639.5, 101609.1, 
    101585.7,
  100654.5, 99846.93, 99677.93, 101406.1, 102408.2, 102297.2, 102168.8, 
    102064.5, 101973.7, 101898.7, 101836, 101786.1, 101746.8, 101714.2, 
    101683.4,
  100968.4, 100085.5, 100390.7, 100833.8, 102400.1, 102403.8, 102289.7, 
    102187.2, 102094.4, 102015.8, 101950.2, 101895.8, 101850.4, 101812, 
    101779.7,
  99710.84, 99447.17, 100706.6, 101008.4, 101552, 102449.4, 102371.4, 
    102265.8, 102183.2, 102109.7, 102041.1, 101988.3, 101937.3, 101900.2, 
    101865.6,
  99771.07, 98131.66, 97913.96, 99059.62, 100767, 101521.3, 102497.5, 
    102402.6, 102260.4, 102214.1, 102131.1, 102084.7, 102028.8, 101987.4, 
    101953.8,
  103089.6, 103006.9, 102899.5, 102786.7, 102697, 102616.9, 102577.7, 
    102520.1, 102476.9, 102450.4, 102425.5, 102390.5, 102352.7, 102311.6, 
    102265.6,
  101595.6, 102941.8, 102864.3, 102737.1, 102610, 102542, 102492.9, 102450.9, 
    102413.6, 102398.8, 102377.1, 102351.3, 102324, 102301.6, 102270.2,
  101671.2, 102591.5, 102828.4, 102690.5, 102538.4, 102452.1, 102405.5, 
    102364.3, 102333, 102323.9, 102309.2, 102290.6, 102274.9, 102259.1, 
    102242.1,
  101360.3, 102515.2, 102778.8, 102650.6, 102449.1, 102353.1, 102299.4, 
    102260.7, 102236.2, 102227.8, 102221, 102220.2, 102212.9, 102210, 102200.8,
  101328.6, 101869.5, 102600.6, 102629.9, 102409.6, 102257.1, 102210.5, 
    102171.6, 102153.9, 102150.9, 102148.7, 102150.8, 102151.8, 102152.3, 
    102153.5,
  101055.4, 100685.4, 101433.4, 102565.9, 102428.2, 102229.6, 102170.6, 
    102130.9, 102112.2, 102103, 102110.2, 102119.9, 102123.6, 102123.7, 
    102121.4,
  100999.1, 100139.9, 99924.03, 101585.9, 102475.7, 102270.4, 102198.4, 
    102161.5, 102130, 102113, 102103, 102106.4, 102114.3, 102122.5, 102120,
  101342.9, 100390.9, 100640.6, 101007, 102516.1, 102385.8, 102282.9, 
    102234.8, 102192.4, 102164.5, 102141.5, 102144.2, 102145.3, 102145.1, 
    102141.6,
  100137.6, 99827.02, 101035.3, 101227.6, 101730.5, 102526.8, 102432, 
    102362.5, 102311.1, 102264.2, 102217.6, 102196.1, 102182.9, 102176.6, 
    102169.8,
  100244.1, 98548.08, 98274.05, 99365.3, 101027.6, 101700, 102601.6, 
    102508.7, 102394.9, 102363.4, 102303.3, 102275, 102239.1, 102222.5, 
    102205.3,
  102904.1, 102860.8, 102812.7, 102740.2, 102664.4, 102574.6, 102501.4, 
    102432.7, 102362.1, 102299.4, 102245.2, 102194.8, 102145.7, 102108.3, 
    102073.1,
  101527.3, 102916.7, 102903.1, 102831.6, 102745, 102650.7, 102569.3, 
    102509.2, 102444.1, 102384.1, 102334.2, 102288.7, 102242.6, 102203.6, 
    102169.5,
  101680.1, 102679.8, 102970.6, 102901, 102814.5, 102700, 102620, 102558.1, 
    102499.5, 102448.5, 102407.4, 102364.9, 102324.6, 102289.5, 102258.6,
  101437.2, 102684.5, 103014.8, 102959.8, 102861.5, 102738, 102649, 102580.3, 
    102523.5, 102484.2, 102452.9, 102425.1, 102398.4, 102375.3, 102353.3,
  101459.3, 102071, 102891.7, 102990.6, 102898, 102759, 102656.4, 102584.6, 
    102529.4, 102484.5, 102451.6, 102433.6, 102421, 102409.7, 102407.8,
  101206.7, 100908.7, 101736.7, 102947.9, 102930.1, 102762.6, 102649.7, 
    102564.1, 102505.8, 102462.7, 102436.3, 102418.9, 102400.4, 102393.9, 
    102387.4,
  101155.2, 100372.2, 100200.9, 101922.5, 102932.6, 102782.1, 102622.6, 
    102543.5, 102479.9, 102434.4, 102404.1, 102391.1, 102385.1, 102382.8, 
    102377.2,
  101469.3, 100591.8, 100898.9, 101312.1, 102876.7, 102802.3, 102612.8, 
    102528.2, 102456.5, 102416, 102385.1, 102379.1, 102377.5, 102387.1, 
    102366.7,
  100235, 99975.78, 101219.2, 101451.5, 101984.5, 102808.9, 102621, 102507.5, 
    102439, 102407.3, 102375.9, 102367.2, 102359.6, 102356.7, 102363,
  100313, 98656.27, 98425.5, 99545.61, 101199.1, 101900.9, 102708.3, 
    102548.2, 102438.8, 102426.2, 102397.5, 102389.1, 102376, 102374.9, 
    102367.1,
  102429.2, 102378, 102324.7, 102250, 102165.8, 102064, 101969, 101876, 
    101760.5, 101643.5, 101533.2, 101424.2, 101317.9, 101222.1, 101130.1,
  101078, 102447.5, 102444.8, 102375.5, 102293, 102196.2, 102098.7, 102009.8, 
    101915.1, 101809.7, 101703.2, 101600.3, 101498.4, 101402.5, 101317.2,
  101246.3, 102245, 102555, 102491, 102418, 102325.2, 102225.5, 102136.4, 
    102046.7, 101952, 101856.4, 101761.3, 101667.5, 101575.5, 101488.8,
  101043.6, 102287.3, 102643.7, 102594.1, 102520.5, 102434.3, 102341.8, 
    102256.4, 102168, 102080.9, 101992.5, 101908.1, 101821, 101737.8, 101659.1,
  101117.3, 101733.3, 102576.1, 102691.6, 102630.4, 102541.8, 102451.7, 
    102366, 102280.9, 102200.1, 102120.3, 102040, 101962.7, 101888.2, 101816.1,
  100900, 100630, 101469.3, 102710, 102734.2, 102646.5, 102560.2, 102469.8, 
    102386.9, 102304.1, 102227.5, 102154.2, 102084.6, 102014.6, 101948.5,
  100878.8, 100136.5, 100012.5, 101751.4, 102806.6, 102754.4, 102662.5, 
    102570.9, 102483.9, 102398.4, 102322.4, 102250.7, 102185.8, 102121.6, 
    102059.9,
  101212.9, 100378.5, 100734.9, 101206.7, 102808.9, 102837, 102747.8, 102663, 
    102569.4, 102483.6, 102402.2, 102332.7, 102267.2, 102211.8, 102152.1,
  99997.76, 99777.48, 101052.3, 101378.4, 101974.3, 102890.5, 102833.9, 
    102729.9, 102636.8, 102552.3, 102467.5, 102398.9, 102333.5, 102278.5, 
    102221.9,
  100079, 98480.45, 98295.85, 99458.68, 101173.4, 101941.5, 102909.2, 
    102837.8, 102689.2, 102609, 102518, 102450.3, 102384.7, 102325.2, 102272,
  102025, 102054.8, 102049.1, 102019.1, 101979.5, 101927.5, 101877.6, 
    101836.4, 101791.6, 101743.9, 101702.3, 101661.5, 101622.9, 101586.8, 
    101554.6,
  100676.6, 102090.4, 102160.5, 102139.8, 102111.6, 102066.9, 102012.1, 
    101970.4, 101927.4, 101883.3, 101837, 101794.1, 101753.2, 101714.3, 
    101679.6,
  100853, 101886.7, 102257.2, 102241.6, 102221.2, 102181.7, 102131.8, 102089, 
    102046.8, 102004.3, 101960, 101914.3, 101871, 101827.4, 101788.5,
  100634.1, 101909, 102329.5, 102331.9, 102312.6, 102279.1, 102234.2, 
    102190.3, 102150, 102109.9, 102068.7, 102024.5, 101981.9, 101938.3, 
    101895.8,
  100685.1, 101336.8, 102231.2, 102412.5, 102403.1, 102373.1, 102333.8, 
    102287.6, 102249.4, 102211.2, 102169.8, 102125.5, 102082.9, 102037.7, 
    101995.1,
  100438.2, 100226.2, 101094.8, 102389.2, 102480, 102451.8, 102416.7, 
    102376.1, 102337.8, 102300.1, 102258.4, 102215, 102170.2, 102125.2, 
    102081.5,
  100412.5, 99724.98, 99658.16, 101414.3, 102521.8, 102526.9, 102491.7, 
    102455.3, 102417.6, 102380.5, 102339.6, 102295.5, 102250.1, 102203.8, 
    102159.1,
  100693.8, 99923.27, 100351.3, 100857.5, 102486.2, 102578.6, 102551.8, 
    102523.7, 102487, 102453.5, 102411.7, 102372.2, 102325.1, 102278, 102231.5,
  99492.53, 99302.61, 100611.7, 100982, 101618.4, 102600.1, 102615.7, 
    102581.5, 102545.9, 102518.5, 102474.1, 102436.7, 102394.9, 102346.6, 
    102298.2,
  99553.02, 98023.95, 97853.73, 99034.38, 100806.5, 101578.2, 102655.1, 
    102644.4, 102594.3, 102575.7, 102533.7, 102497.2, 102456.3, 102412.9, 
    102363.8,
  102354.2, 102339.6, 102334.1, 102304.1, 102280.5, 102247.5, 102231.1, 
    102197.4, 102155.3, 102108.8, 102059.9, 102007.2, 101946.6, 101886.9, 
    101824.4,
  100899.7, 102301.1, 102368.9, 102351.7, 102330.9, 102303, 102276.1, 
    102255.1, 102219.2, 102175.9, 102132.7, 102089.2, 102042, 101989.6, 101937,
  101003.5, 102031.4, 102412.4, 102394.4, 102376.3, 102345.5, 102316.6, 
    102296.2, 102274.6, 102243.8, 102207.7, 102168.5, 102124.9, 102080.2, 
    102032.2,
  100708.6, 101986.8, 102419.5, 102425.2, 102417.8, 102393.9, 102371.8, 
    102348.7, 102325.4, 102304.3, 102279.1, 102250.8, 102217.3, 102178.9, 
    102139.8,
  100691.9, 101362.3, 102275.2, 102467.7, 102466.8, 102446, 102429, 102410.5, 
    102390.6, 102369.8, 102349, 102326.3, 102302.4, 102272.4, 102239.5,
  100401.8, 100200.5, 101088.6, 102401.6, 102496.1, 102486.1, 102475, 
    102460.1, 102449.9, 102437.8, 102421.4, 102402.3, 102382, 102357.7, 
    102331.3,
  100334.4, 99665.55, 99620.98, 101382.7, 102500.9, 102521, 102511.2, 
    102504.8, 102499.9, 102495.3, 102485.6, 102472, 102457, 102438.2, 102416.2,
  100584.2, 99833.24, 100275.8, 100784.5, 102415.4, 102517, 102517.3, 
    102522.6, 102527.8, 102530.4, 102531.5, 102528.2, 102521, 102509.8, 
    102493.9,
  99366.7, 99199.22, 100512.4, 100879.9, 101518.6, 102498, 102536.8, 
    102531.1, 102545.7, 102563.1, 102575.7, 102580.7, 102578.7, 102571.8, 
    102559.7,
  99415.58, 97921.19, 97759.67, 98945.58, 100713.8, 101468.4, 102538.5, 
    102534.1, 102553.3, 102591.1, 102612, 102625.4, 102627.7, 102625, 102617.6,
  102013.7, 102079.4, 102125.5, 102148.4, 102166.3, 102199.3, 102250.7, 
    102304, 102343.9, 102404.9, 102454.2, 102508, 102560.9, 102600.4, 102637.7,
  100571.8, 102033, 102126.9, 102160, 102181.1, 102198.2, 102239.4, 102295.1, 
    102336.6, 102391, 102444.1, 102508.7, 102561.7, 102615.1, 102657.4,
  100687.1, 101737.7, 102141.8, 102171.3, 102190.8, 102210.8, 102242.3, 
    102290.4, 102340.9, 102395.9, 102447.5, 102511.1, 102554.4, 102607.8, 
    102658,
  100378.6, 101686.2, 102133.9, 102175.4, 102211.8, 102229.3, 102257, 
    102297.6, 102344.8, 102396.7, 102454.5, 102517.3, 102567.9, 102620.6, 
    102663.5,
  100383.7, 101065, 101986.4, 102204.3, 102229, 102253.9, 102276.8, 102318.2, 
    102367.6, 102417, 102464.3, 102509.2, 102565.9, 102627.3, 102672.3,
  100104.3, 99915.95, 100811, 102137.8, 102246, 102273.6, 102295, 102335.3, 
    102383.9, 102430.9, 102482.7, 102533.6, 102581.8, 102629.1, 102668.6,
  100056.9, 99398.09, 99369.78, 101136.2, 102254.1, 102295.5, 102314.9, 
    102358.4, 102408, 102453.6, 102508.4, 102559.7, 102606.7, 102649.4, 
    102685.8,
  100320.5, 99577.23, 100035.7, 100548.5, 102175.2, 102301.2, 102325.9, 
    102374.8, 102423.8, 102469.2, 102533.1, 102587.5, 102633.2, 102674, 102710,
  99122.48, 98962.04, 100282.8, 100664.9, 101301.8, 102298.3, 102354.9, 
    102393.9, 102439.8, 102492.1, 102561.6, 102616.9, 102661.7, 102708.5, 
    102743.2,
  99193.68, 97711.25, 97540.78, 98731.95, 100499.5, 101274.1, 102374.8, 
    102416.8, 102442.9, 102512.9, 102585.2, 102642.9, 102685.9, 102733.5, 
    102768,
  101730.5, 101728.4, 101708.3, 101680.2, 101624.3, 101577.2, 101546, 
    101533.2, 101522.2, 101519.8, 101534.3, 101559.2, 101597.4, 101659.1, 
    101735.9,
  100305.8, 101710.7, 101768.6, 101751.5, 101713.9, 101669.4, 101639.6, 
    101629.7, 101621.7, 101621.2, 101636.7, 101670.2, 101703.7, 101763.8, 
    101836.2,
  100441.9, 101441.3, 101810.4, 101817.9, 101795, 101757.4, 101733.4, 
    101719.4, 101718.3, 101723.9, 101742, 101764.1, 101810.8, 101867.1, 
    101936.6,
  100173.7, 101419.6, 101843.9, 101855.2, 101869.2, 101846.2, 101830, 
    101816.9, 101817.6, 101830.4, 101834.5, 101863.9, 101917.6, 101971.1, 
    102030.6,
  100195.9, 100835.6, 101736.2, 101920.2, 101928.6, 101932.2, 101924.5, 
    101908, 101917.1, 101912.4, 101918.7, 101956.2, 102004, 102050.7, 102118,
  99942.22, 99736.03, 100602.3, 101895.9, 101988.3, 101990.3, 102000.2, 
    101989.2, 101994.7, 101978.9, 102002.9, 102033.5, 102084.3, 102134.7, 
    102200.4,
  99885.39, 99213.76, 99157.86, 100911.6, 102023.2, 102039.1, 102043.3, 
    102043.6, 102046.5, 102046.3, 102078.7, 102110.1, 102154, 102211.2, 
    102275.9,
  100172.9, 99415.84, 99838.45, 100340.6, 101958.6, 102070.7, 102082.7, 
    102089.8, 102093.8, 102108.4, 102140.7, 102178.4, 102220.8, 102276.6, 
    102338.8,
  98980.43, 98804.01, 100105.7, 100489.3, 101094.8, 102070.6, 102115, 
    102119.1, 102141.7, 102165.1, 102196.9, 102236.5, 102278.5, 102334.5, 
    102396.4,
  99049.92, 97561.98, 97404.7, 98572.8, 100299.3, 101092.5, 102154.7, 
    102173.7, 102168.5, 102210, 102239.5, 102289.4, 102330.4, 102388.7, 
    102446.2 ;

 sftlf =
  0.1986115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9611561, 0.1583273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7949425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7552791, 0.2484612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.9872221, 0.4156101, 0.04560489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.8345782, 0.2958934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.7792858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9990003, 0.3505592, 0.06537855, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.8140894, 0.2409153, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.9453563, 0.02902743, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  1.522432, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  122.465, 2.830728, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  113.0215, 29.31339, 0.004701966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  140.0874, 33.71546, 1.141547, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  141.9684, 87.21121, 14.52402, 0.1304746, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  165.7051, 185.2302, 111.1391, 5.227489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  172.6293, 232.1111, 238.8028, 89.74486, 0.6524738, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  149.5705, 217.5222, 183.4477, 142.7244, 6.651272, 0.2006134, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  253.9191, 270.7406, 160.8987, 135.4378, 83.93595, 3.422685, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  248.2018, 381.5977, 396.3867, 296.0411, 147.8827, 85.51294, 0.2661929, 0, 
    0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
