netcdf atmos_static_scalar_3.ck {
dimensions:
        lat = 6 ;
        lon = 7 ;
variables:
        float ck(lat, lon) ;
                ck:long_name = "vertical coordinate sigma value" ;
                ck:wrong_units = "wrong_unit" ;
                ck:missing_value = 1.e+20f ;
                ck:_FillValue = 1.e+20f ;
                ck:cell_methods = "time: point" ;
        float lat(lat) ;
        float lon(lon) ;
}
