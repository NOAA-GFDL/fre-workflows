netcdf atmos_daily.00010101-00010701.pr.tile4 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pr(time, grid_yt, grid_xt) ;
		pr:_FillValue = 1.e+20f ;
		pr:missing_value = 1.e+20f ;
		pr:units = "kg m-2 s-1" ;
		pr:long_name = "Precipitation" ;
		pr:cell_methods = "time: mean" ;
		pr:cell_measures = "area: area" ;
		pr:time_avg_info = "average_T1,average_T2,average_DT" ;
		pr:standard_name = "precipitation_flux" ;
		pr:interp_method = "conserve_order1" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:03 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile4.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile4.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.2466774, 0.6143242, 0.0668168, 0.2301621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.4924844, 0.2132108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.600569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1560082, 0,
  1, 1, 0.7132517, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02739768, 0,
  0.6230268, 0.6280472, 0.3043983, 0.08344039, 0, 0.3148882, 0.01188002, 0, 
    0, 0, 0, 0.08803581, 0, 0, 0,
  0, 0, 0, 0, 0.01144353, 0.8597386, 0.8205094, 0.5086318, 0.1258651, 
    0.08909279, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.291879, 0.6933324, 1, 0.9996726, 0.6666086, 0.08008575, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.611689, 0.7180831, 0.4623523, 0.2838529, 0.02767258, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0.002817577, 0.8915156, 0.5654301, 0.7485356, 0.3018697, 0, 0, 0, 
    0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pr =
  0.0001081887, 0.0001046199, 9.371072e-05, 9.009951e-05, 6.60707e-05, 
    4.940007e-05, 3.847138e-05, 3.621463e-05, 3.682214e-05, 3.690074e-05, 
    3.986833e-05, 3.571063e-05, 3.583044e-05, 4.657832e-05, 5.890123e-05,
  4.987934e-05, 5.482241e-05, 9.410775e-05, 8.321281e-05, 8.031804e-05, 
    9.022694e-05, 6.515281e-05, 5.162975e-05, 4.994209e-05, 4.669286e-05, 
    4.983995e-05, 4.948492e-05, 4.806573e-05, 5.790297e-05, 5.853715e-05,
  7.56838e-06, 1.6238e-05, 4.50459e-05, 7.434549e-05, 9.553545e-05, 
    9.163446e-05, 6.768306e-05, 5.44998e-05, 5.466418e-05, 6.1426e-05, 
    5.601239e-05, 5.968355e-05, 5.775705e-05, 6.561811e-05, 5.066306e-05,
  2.909376e-06, 5.48241e-06, 1.724562e-05, 7.097729e-05, 8.998905e-05, 
    0.0001040128, 8.405208e-05, 6.109393e-05, 6.208275e-05, 5.911403e-05, 
    6.137331e-05, 7.105203e-05, 7.492761e-05, 3.834488e-05, 3.693477e-05,
  1.842976e-06, 2.364439e-06, 1.47786e-05, 4.074825e-05, 9.817413e-05, 
    9.218635e-05, 0.0001049237, 8.320224e-05, 7.491779e-05, 6.226785e-05, 
    7.310425e-05, 7.182464e-05, 6.858942e-05, 4.993409e-05, 2.653822e-05,
  1.293556e-06, 1.862521e-06, 9.137445e-06, 5.036361e-05, 0.000105821, 
    9.89527e-05, 9.766006e-05, 8.05848e-05, 7.655469e-05, 7.210183e-05, 
    7.317578e-05, 7.036392e-05, 6.087621e-05, 5.116963e-05, 4.027776e-05,
  1.056584e-05, 1.934623e-06, 3.745846e-06, 3.837343e-05, 8.770591e-05, 
    7.528581e-05, 4.967919e-05, 5.202192e-05, 7.198821e-05, 9.114671e-05, 
    7.991046e-05, 6.878994e-05, 5.872474e-05, 4.689097e-05, 4.336357e-05,
  8.078097e-05, 2.034503e-05, 5.443358e-06, 2.580868e-05, 6.501624e-05, 
    4.168592e-05, 3.362558e-05, 3.841462e-05, 2.797147e-05, 3.967705e-05, 
    6.455577e-05, 6.080607e-05, 5.173051e-05, 5.525977e-05, 4.130483e-05,
  7.551413e-05, 4.845995e-05, 2.82344e-05, 3.36774e-05, 5.371876e-05, 
    3.240984e-05, 2.528738e-05, 2.06042e-05, 4.359015e-05, 4.869903e-05, 
    7.458976e-05, 6.191876e-05, 5.287956e-05, 4.148383e-05, 3.132792e-05,
  5.33877e-05, 6.797175e-05, 6.268861e-05, 5.733494e-05, 2.213962e-05, 
    2.364228e-05, 2.393479e-05, 3.513321e-05, 4.185243e-05, 5.332784e-05, 
    9.052843e-05, 5.061817e-05, 5.515912e-05, 3.383628e-05, 1.538476e-05,
  6.19086e-05, 7.623342e-05, 9.725763e-05, 9.01113e-05, 7.422398e-05, 
    5.710942e-05, 4.105728e-05, 3.50083e-05, 3.269596e-05, 3.614208e-05, 
    4.173234e-05, 3.634201e-05, 3.539267e-05, 3.435712e-05, 3.128286e-05,
  2.768214e-05, 1.520281e-05, 6.2919e-05, 5.418114e-05, 6.762816e-05, 
    7.570634e-05, 6.143469e-05, 5.772229e-05, 5.374067e-05, 5.219562e-05, 
    5.124656e-05, 5.115907e-05, 4.474784e-05, 3.672285e-05, 3.066327e-05,
  2.054709e-06, 2.143797e-06, 3.870922e-06, 3.042281e-05, 5.609522e-05, 
    6.400555e-05, 7.287179e-05, 7.057461e-05, 6.642245e-05, 5.728686e-05, 
    5.747522e-05, 5.17421e-05, 4.680967e-05, 3.941726e-05, 3.288936e-05,
  8.046947e-07, 2.527014e-07, 2.113754e-07, 3.064773e-05, 5.871015e-05, 
    6.879577e-05, 8.162745e-05, 8.303524e-05, 6.39537e-05, 6.348942e-05, 
    5.652135e-05, 5.367989e-05, 5.332137e-05, 3.31204e-05, 2.669217e-05,
  4.199175e-08, 3.933046e-09, 2.607958e-09, 5.544284e-06, 4.533696e-05, 
    7.33718e-05, 9.018301e-05, 8.321107e-05, 8.191516e-05, 6.727116e-05, 
    5.456734e-05, 5.622636e-05, 5.07971e-05, 3.727661e-05, 2.524979e-05,
  5.242643e-06, 3.664774e-07, 8.931105e-09, 7.332627e-08, 2.509861e-05, 
    3.935056e-05, 8.768945e-05, 0.0001333407, 0.0001158185, 9.315531e-05, 
    7.304626e-05, 4.661037e-05, 4.27021e-05, 3.945728e-05, 2.254153e-05,
  0.0001142527, 4.050995e-05, 5.882413e-06, 8.223711e-06, 3.120413e-05, 
    2.142259e-05, 1.758706e-05, 4.88179e-05, 9.661146e-05, 9.998478e-05, 
    8.667274e-05, 5.59441e-05, 3.755172e-05, 3.153017e-05, 2.291335e-05,
  0.0001297857, 0.0001452138, 0.0001046097, 4.827668e-05, 4.423091e-05, 
    2.849734e-05, 1.846821e-05, 2.50042e-05, 2.152049e-05, 3.419825e-05, 
    7.311474e-05, 6.456079e-05, 4.214905e-05, 2.73432e-05, 2.452721e-05,
  9.438135e-05, 0.0001240353, 0.0001298871, 0.0001038156, 7.622728e-05, 
    2.675907e-05, 2.367906e-05, 1.552786e-05, 1.776565e-05, 4.286503e-05, 
    5.81549e-05, 5.732382e-05, 4.121761e-05, 3.177472e-05, 3.849793e-05,
  5.017021e-05, 0.0001380442, 0.0001237723, 0.0001258186, 3.494634e-05, 
    5.568919e-05, 2.602825e-05, 1.50436e-05, 2.917192e-05, 3.979429e-05, 
    4.725177e-05, 5.176826e-05, 5.279855e-05, 5.655211e-05, 4.49255e-05,
  9.695924e-05, 0.0001104152, 9.851658e-05, 8.705661e-05, 5.346555e-05, 
    3.769237e-05, 1.761873e-05, 1.341237e-05, 1.537383e-05, 1.624354e-05, 
    1.742226e-05, 1.391143e-05, 1.748035e-05, 1.630413e-05, 1.751021e-05,
  3.313391e-05, 3.471445e-05, 8.644143e-05, 6.194854e-05, 6.477227e-05, 
    5.016969e-05, 3.208449e-05, 2.398571e-05, 2.554665e-05, 2.728755e-05, 
    2.544242e-05, 2.098294e-05, 2.289754e-05, 2.31071e-05, 1.951423e-05,
  2.253203e-06, 1.482635e-06, 4.932245e-06, 5.320023e-05, 6.27407e-05, 
    5.926103e-05, 5.880563e-05, 4.109895e-05, 3.277069e-05, 3.612941e-05, 
    3.189865e-05, 3.071457e-05, 2.964105e-05, 2.759834e-05, 2.222759e-05,
  8.694671e-07, 3.013561e-07, 2.584212e-06, 6.526131e-05, 6.553462e-05, 
    8.008001e-05, 6.360105e-05, 5.808516e-05, 4.937742e-05, 3.918365e-05, 
    4.047218e-05, 3.664603e-05, 3.876885e-05, 2.915126e-05, 2.514454e-05,
  1.29614e-08, 1.10661e-08, 8.123907e-08, 2.342487e-05, 6.451963e-05, 
    7.785743e-05, 8.905622e-05, 7.13713e-05, 5.850521e-05, 4.483488e-05, 
    4.169114e-05, 4.162334e-05, 4.156671e-05, 3.812187e-05, 2.886861e-05,
  1.576278e-09, 1.391011e-10, 1.079013e-09, 2.620069e-06, 6.633205e-05, 
    6.744601e-05, 0.0001208271, 0.0001323364, 9.392916e-05, 7.183531e-05, 
    4.952112e-05, 3.586359e-05, 3.712146e-05, 4.083784e-05, 3.52698e-05,
  9.337986e-06, 2.438005e-06, 7.435661e-07, 1.089914e-05, 7.479318e-05, 
    2.267024e-05, 2.28732e-05, 5.501109e-05, 0.0001175446, 0.0001008885, 
    7.010444e-05, 4.45928e-05, 3.731213e-05, 3.733282e-05, 3.450702e-05,
  0.0001138595, 8.942238e-05, 5.093779e-05, 3.469657e-05, 3.86472e-05, 
    4.823213e-05, 9.422049e-06, 8.885201e-06, 7.055105e-06, 6.044259e-05, 
    8.213941e-05, 6.589363e-05, 4.393212e-05, 3.329589e-05, 3.010188e-05,
  0.0001558934, 0.0001910911, 0.0001674285, 0.000100139, 6.534166e-05, 
    1.702666e-05, 7.076177e-06, 4.755364e-06, 2.182895e-05, 5.786885e-05, 
    7.756504e-05, 7.385719e-05, 5.438983e-05, 3.884154e-05, 2.878707e-05,
  0.0001182956, 0.0002316035, 0.0002700094, 0.0001725414, 1.865295e-05, 
    1.045054e-05, 7.552684e-06, 7.484231e-07, 2.133613e-05, 4.762943e-05, 
    7.125107e-05, 7.857964e-05, 6.110306e-05, 4.262465e-05, 2.870365e-05,
  4.835209e-05, 5.512598e-05, 4.501999e-05, 4.025838e-05, 1.836375e-05, 
    5.645114e-06, 6.237479e-07, 5.341152e-08, 2.520194e-07, 2.649142e-07, 
    6.645549e-07, 2.0913e-07, 1.855244e-06, 1.453941e-06, 3.811131e-06,
  2.856451e-05, 1.774111e-05, 4.165974e-05, 3.656094e-05, 4.633835e-05, 
    2.433059e-05, 8.791043e-06, 5.715992e-06, 3.609e-06, 3.063813e-06, 
    3.493202e-06, 3.396828e-06, 4.226015e-06, 5.082513e-06, 3.339839e-06,
  9.957741e-07, 9.030647e-07, 8.30863e-06, 2.670736e-05, 5.145426e-05, 
    4.178049e-05, 2.554506e-05, 1.760913e-05, 1.070749e-05, 9.328085e-06, 
    7.590605e-06, 7.7586e-06, 8.05849e-06, 6.165393e-06, 5.019914e-06,
  4.712912e-07, 1.312288e-06, 5.023805e-06, 4.588331e-05, 5.986817e-05, 
    5.662856e-05, 3.939988e-05, 2.691871e-05, 2.038276e-05, 1.879379e-05, 
    1.528446e-05, 1.197499e-05, 1.138573e-05, 6.775026e-06, 4.950035e-06,
  1.724196e-08, 5.796159e-08, 1.281765e-06, 3.862169e-05, 5.482327e-05, 
    7.722836e-05, 6.858558e-05, 3.84976e-05, 3.018336e-05, 2.016285e-05, 
    1.859915e-05, 1.389735e-05, 1.531886e-05, 1.120504e-05, 7.656578e-06,
  2.090442e-06, 5.649768e-07, 3.83019e-07, 2.136474e-05, 5.731799e-05, 
    8.216895e-05, 9.324803e-05, 8.02001e-05, 5.206357e-05, 3.327663e-05, 
    2.158638e-05, 1.220396e-05, 1.65486e-05, 1.205847e-05, 1.105002e-05,
  2.227027e-05, 1.563727e-05, 2.127687e-05, 2.858906e-05, 8.085123e-05, 
    4.506882e-05, 1.870537e-05, 6.514618e-05, 6.36227e-05, 4.700926e-05, 
    3.031432e-05, 1.896259e-05, 1.598849e-05, 1.315548e-05, 1.051044e-05,
  7.030096e-05, 5.494997e-05, 4.405811e-05, 4.206846e-05, 7.082957e-05, 
    4.207128e-05, 2.450839e-05, 1.630733e-05, 2.052989e-05, 3.152203e-05, 
    3.937591e-05, 2.536389e-05, 1.707366e-05, 1.284536e-05, 9.600179e-06,
  8.806628e-05, 6.547993e-05, 5.905114e-05, 6.215295e-05, 8.801477e-05, 
    5.493924e-05, 3.016119e-05, 9.283421e-06, 2.890395e-05, 4.947146e-05, 
    4.216602e-05, 3.338415e-05, 1.804047e-05, 1.487419e-05, 8.508345e-06,
  9.426704e-05, 7.881511e-05, 7.431541e-05, 8.490574e-05, 1.605101e-05, 
    8.038238e-05, 1.83672e-05, 8.323074e-06, 3.723108e-05, 4.541453e-05, 
    4.175647e-05, 3.42399e-05, 2.753579e-05, 1.227181e-05, 7.978203e-06,
  8.350616e-06, 4.241687e-06, 1.875142e-06, 1.754978e-07, 1.645523e-08, 
    9.521338e-10, 8.568528e-10, 8.746421e-12, 1.370245e-10, 3.52197e-09, 
    2.848236e-08, 5.671527e-08, 1.692588e-08, 3.376299e-09, 2.796605e-08,
  4.26588e-06, 1.529134e-06, 5.112552e-06, 1.507659e-06, 6.565701e-07, 
    4.607277e-09, 5.383096e-10, 2.332399e-09, 1.060102e-07, 1.374728e-07, 
    4.796892e-07, 2.165051e-07, 9.044951e-08, 3.279466e-08, 4.932739e-07,
  3.93895e-06, 5.803189e-07, 2.13739e-06, 3.980908e-06, 4.400091e-06, 
    1.489197e-06, 1.280886e-07, 2.586734e-07, 9.016298e-07, 3.301707e-06, 
    2.957676e-06, 1.81037e-06, 3.398321e-07, 1.91839e-07, 3.08326e-07,
  1.603621e-05, 1.805802e-06, 9.552743e-07, 1.057838e-05, 1.034559e-05, 
    8.692678e-06, 4.747569e-06, 5.05614e-06, 1.097208e-05, 1.695255e-05, 
    1.734584e-05, 9.681201e-06, 1.57908e-06, 7.513511e-07, 6.675891e-07,
  1.250641e-05, 4.418159e-06, 5.096892e-07, 1.400311e-05, 1.777382e-05, 
    1.958409e-05, 1.698169e-05, 1.265523e-05, 1.180435e-05, 1.515557e-05, 
    2.050748e-05, 1.846734e-05, 7.544983e-06, 8.270432e-07, 5.852154e-07,
  1.211787e-05, 3.552238e-06, 3.223987e-06, 2.598573e-05, 2.917047e-05, 
    1.448807e-05, 2.848848e-05, 2.701661e-05, 2.199588e-05, 2.490423e-05, 
    2.488062e-05, 1.50131e-05, 7.202776e-06, 1.666604e-06, 9.393622e-07,
  1.178019e-05, 9.630288e-06, 2.574026e-05, 4.371449e-05, 2.760912e-05, 
    5.103736e-06, 6.441116e-06, 1.256258e-05, 2.236681e-05, 2.309287e-05, 
    2.949606e-05, 1.910782e-05, 7.782653e-06, 2.086342e-06, 1.073644e-06,
  2.50117e-05, 2.908463e-05, 4.047026e-05, 5.928424e-05, 1.726874e-05, 
    1.039497e-05, 2.941587e-06, 1.516213e-06, 7.383416e-06, 2.02355e-05, 
    3.131499e-05, 2.233696e-05, 9.386952e-06, 2.683334e-06, 1.522367e-06,
  3.444437e-05, 4.513363e-05, 7.298973e-05, 2.728016e-05, 3.710764e-05, 
    1.134103e-05, 3.538021e-06, 1.346275e-06, 1.482509e-05, 2.90798e-05, 
    3.409637e-05, 2.665604e-05, 1.130552e-05, 2.925282e-06, 4.69274e-07,
  3.805689e-05, 6.734397e-05, 7.36742e-05, 2.47627e-05, 2.520447e-06, 
    1.62899e-05, 3.453637e-06, 1.945032e-06, 2.267259e-05, 3.0344e-05, 
    3.367823e-05, 3.170122e-05, 1.348189e-05, 1.830131e-06, 1.02321e-07,
  1.189693e-05, 3.06836e-06, 1.508878e-08, 5.062942e-08, 1.747423e-07, 
    2.321002e-07, 1.215583e-07, 5.534458e-09, 1.052536e-10, 3.09731e-11, 
    2.032338e-11, 7.681747e-09, 1.91874e-07, 7.957831e-10, 6.800303e-26,
  1.06047e-05, 1.146427e-06, 2.00832e-07, 4.822062e-07, 5.26732e-07, 
    3.346466e-07, 1.366555e-07, 6.516424e-08, 7.999247e-10, 8.986778e-11, 
    3.6751e-08, 4.983618e-07, 8.043025e-08, 7.685949e-10, 1.937014e-13,
  5.54538e-06, 6.350758e-07, 6.756197e-08, 4.991999e-07, 3.373016e-06, 
    2.019835e-06, 3.812156e-07, 4.044322e-07, 8.299026e-08, 1.174725e-07, 
    1.761859e-07, 1.051627e-06, 9.000151e-08, 1.252881e-09, 5.531245e-27,
  6.644514e-06, 1.13059e-06, 2.965374e-08, 2.337513e-06, 5.837026e-06, 
    6.614755e-06, 2.631185e-06, 1.599021e-06, 1.349236e-06, 8.917996e-07, 
    2.832182e-06, 3.193913e-06, 2.475747e-06, 6.718426e-09, 2.403404e-17,
  1.938607e-06, 2.391818e-07, 2.551829e-08, 3.107415e-06, 1.225043e-05, 
    1.630962e-05, 1.108622e-05, 4.743729e-06, 4.271872e-06, 4.086766e-06, 
    8.429278e-06, 7.728451e-06, 3.077193e-06, 1.013848e-08, 2.051193e-13,
  4.813867e-06, 1.85367e-07, 5.575251e-07, 6.165802e-06, 2.406086e-05, 
    1.344423e-05, 2.72455e-05, 1.764378e-05, 1.354059e-05, 6.95922e-06, 
    1.197072e-05, 9.464067e-06, 3.085337e-06, 9.611212e-08, 1.380521e-11,
  5.892364e-06, 3.652116e-06, 7.926224e-06, 2.826231e-05, 4.667333e-05, 
    1.71484e-05, 6.199233e-06, 7.39881e-06, 9.292059e-06, 7.856447e-06, 
    1.304334e-05, 1.188549e-05, 4.455158e-06, 1.121131e-06, 5.949923e-09,
  4.292595e-05, 2.714091e-05, 3.084104e-05, 4.917071e-05, 5.071326e-05, 
    1.468504e-05, 1.076451e-05, 8.36459e-06, 1.099284e-05, 8.60631e-06, 
    1.935057e-05, 2.10056e-05, 6.987654e-06, 1.555072e-06, 4.800114e-08,
  4.467983e-05, 4.679031e-05, 6.322422e-05, 5.4893e-05, 4.827749e-05, 
    5.256978e-05, 1.214924e-05, 6.811296e-07, 7.477484e-06, 2.036314e-05, 
    2.625107e-05, 2.779343e-05, 1.155221e-05, 2.030254e-06, 6.312977e-08,
  4.51853e-05, 7.309857e-05, 6.249135e-05, 7.94107e-05, 4.937665e-05, 
    6.947071e-05, 1.891657e-05, 7.099025e-06, 2.122818e-05, 2.814653e-05, 
    3.773181e-05, 3.639615e-05, 1.444561e-05, 2.174841e-06, 1.747347e-07,
  4.647643e-05, 3.401129e-05, 1.439661e-05, 7.187381e-06, 1.614427e-06, 
    4.866603e-09, 3.436205e-09, 1.101655e-07, 9.266977e-07, 1.692374e-05, 
    1.135563e-05, 2.887472e-07, 3.819988e-11, 4.90666e-13, 2.36874e-16,
  4.472907e-05, 2.766011e-05, 8.398682e-06, 5.511713e-06, 1.260929e-05, 
    8.946997e-06, 2.041283e-08, 2.61308e-07, 1.879491e-06, 5.897418e-06, 
    1.167849e-05, 8.986493e-07, 2.34051e-12, 7.670923e-14, 6.201524e-14,
  2.673433e-05, 1.647359e-05, 7.294012e-06, 5.381772e-06, 1.515088e-05, 
    1.237757e-05, 2.272993e-06, 3.261979e-07, 2.87433e-06, 7.265038e-06, 
    7.187546e-06, 1.235431e-06, 2.715314e-10, 5.97372e-14, 5.652341e-22,
  1.391976e-05, 1.032147e-05, 1.014277e-05, 1.453813e-05, 1.263641e-05, 
    3.527014e-05, 7.195576e-06, 2.376189e-06, 6.334973e-06, 1.39921e-05, 
    1.149833e-05, 3.672977e-06, 1.247219e-09, 8.850176e-13, 4.291738e-22,
  3.865687e-06, 7.862782e-06, 2.558804e-05, 1.920251e-05, 3.068912e-05, 
    7.389062e-05, 3.742301e-05, 6.441294e-06, 9.993637e-06, 1.760291e-05, 
    1.911334e-05, 8.271071e-06, 1.38275e-08, 3.348655e-14, 2.796386e-12,
  1.145597e-05, 7.121519e-06, 3.320833e-05, 4.948027e-05, 6.970882e-05, 
    7.485284e-05, 0.0001112447, 3.271703e-05, 1.338648e-05, 2.051545e-05, 
    2.551561e-05, 1.596175e-05, 2.356777e-09, 1.563609e-12, 2.506685e-22,
  1.182081e-05, 1.024428e-05, 5.076387e-05, 9.68875e-05, 0.0001085163, 
    6.200591e-05, 3.834756e-05, 4.382244e-05, 2.651725e-05, 3.17949e-05, 
    3.021226e-05, 1.799973e-05, 1.378939e-08, 2.908015e-10, 5.199613e-12,
  3.227401e-05, 3.723303e-05, 7.862377e-05, 0.0001197415, 0.00010256, 
    5.657054e-05, 5.211473e-05, 2.526677e-05, 1.642508e-05, 2.389627e-05, 
    3.069004e-05, 1.982849e-05, 3.397201e-07, 6.135004e-08, 2.52445e-10,
  5.024327e-05, 5.140251e-05, 7.792582e-05, 0.0001244909, 9.159661e-05, 
    4.16662e-05, 2.847583e-05, 3.486791e-05, 2.410974e-05, 3.385497e-05, 
    4.282812e-05, 1.939537e-05, 4.744767e-06, 4.203745e-08, 2.471546e-11,
  5.793768e-05, 4.709847e-05, 7.628701e-05, 0.00013145, 6.786543e-05, 
    3.88107e-05, 4.802473e-05, 3.922664e-05, 3.970885e-05, 3.671336e-05, 
    4.835651e-05, 3.22758e-05, 7.989985e-06, 7.869093e-07, 4.7437e-09,
  9.975016e-07, 8.393675e-08, 1.293669e-07, 1.909893e-07, 1.781379e-07, 
    1.47386e-06, 1.38745e-05, 2.34959e-05, 1.530837e-05, 1.498783e-05, 
    6.93366e-06, 1.704417e-06, 4.669075e-08, 1.328911e-08, 2.14237e-08,
  3.417507e-07, 5.440623e-08, 5.731262e-08, 9.571445e-08, 9.938034e-08, 
    2.498434e-07, 7.402482e-07, 4.432419e-06, 6.122461e-06, 7.065801e-06, 
    6.134368e-06, 2.358832e-06, 9.926977e-09, 3.260722e-09, 2.154077e-09,
  3.812116e-07, 1.765182e-08, 7.937879e-08, 5.077944e-08, 5.19399e-08, 
    4.528991e-08, 2.662854e-07, 3.747144e-07, 7.650145e-06, 1.314657e-05, 
    9.251772e-06, 7.156042e-06, 8.851364e-08, 5.060555e-09, 1.359962e-08,
  7.16749e-07, 3.335611e-08, 9.439233e-08, 1.423362e-07, 9.716804e-07, 
    3.682289e-07, 4.374537e-08, 9.013767e-08, 1.688031e-06, 6.031799e-06, 
    1.125357e-05, 1.045294e-05, 3.938907e-07, 1.301355e-08, 1.722353e-08,
  2.620673e-08, 7.814135e-09, 2.246126e-09, 1.176084e-07, 8.550804e-07, 
    9.222928e-07, 5.239475e-08, 3.750909e-08, 3.5548e-08, 1.919369e-06, 
    6.901125e-06, 2.038754e-05, 1.007134e-06, 3.101719e-09, 2.147529e-08,
  9.237838e-08, 3.071227e-07, 3.092002e-08, 4.451864e-08, 1.042714e-07, 
    6.579753e-07, 7.040582e-07, 1.033472e-07, 6.631345e-09, 2.27269e-07, 
    5.692244e-06, 2.049074e-05, 1.383682e-06, 9.794233e-09, 2.907518e-08,
  2.562646e-07, 6.804969e-08, 1.626041e-07, 4.975059e-08, 4.454312e-07, 
    3.106457e-07, 1.320835e-08, 4.278493e-08, 1.152417e-08, 4.749837e-08, 
    3.711366e-06, 2.280291e-05, 1.933118e-06, 3.921104e-09, 2.907873e-08,
  8.271459e-06, 2.264823e-06, 2.393664e-07, 2.30263e-07, 1.693188e-06, 
    1.200124e-06, 8.448487e-08, 3.436785e-07, 3.752716e-08, 1.332349e-07, 
    4.878445e-06, 2.059035e-05, 7.435848e-06, 1.172837e-09, 9.247391e-09,
  1.421897e-05, 4.025313e-06, 8.562503e-07, 1.372589e-06, 6.863138e-06, 
    5.192423e-07, 6.95398e-09, 4.677599e-09, 1.371293e-08, 1.48805e-07, 
    4.95657e-06, 2.45221e-05, 1.253116e-05, 1.224904e-09, 5.645657e-09,
  1.73814e-05, 3.906725e-06, 3.281343e-06, 4.565846e-06, 1.74854e-06, 
    1.609406e-06, 2.605141e-08, 7.286727e-09, 4.749438e-09, 6.824847e-08, 
    3.727829e-06, 2.792771e-05, 2.482173e-05, 4.290158e-08, 1.649336e-08,
  9.753566e-05, 0.0001824442, 0.0003116418, 0.000347156, 0.0004142713, 
    0.0005588787, 0.0007497658, 0.0008814128, 0.0008495693, 0.0005450568, 
    0.0004395757, 0.0004576397, 0.0006797097, 0.000881867, 0.0007631222,
  9.717862e-05, 0.0001559756, 0.0002455424, 0.0002904611, 0.0003232239, 
    0.0003991344, 0.0005931235, 0.0007884299, 0.0008258156, 0.0006052993, 
    0.00060676, 0.000544978, 0.0007919423, 0.001013444, 0.00104457,
  4.098446e-05, 0.000102623, 0.0001557858, 0.0002239244, 0.0002467315, 
    0.0002883144, 0.0004609117, 0.0006550145, 0.0008548964, 0.0009738731, 
    0.0008524971, 0.0006309946, 0.0006866516, 0.00103486, 0.001121089,
  2.026147e-05, 6.192043e-05, 8.641554e-05, 0.0001594328, 0.0001758903, 
    0.0001851487, 0.0003001077, 0.0005331088, 0.0009186133, 0.00103485, 
    0.0007499, 0.000580939, 0.0005842844, 0.0007778447, 0.0008975292,
  6.892524e-06, 3.080796e-05, 3.62741e-05, 9.001361e-05, 0.0001138033, 
    0.0001034458, 0.0001749693, 0.0003383945, 0.0006908757, 0.0007388876, 
    0.0005401403, 0.0003533591, 0.0002892775, 0.0003710574, 0.0004873943,
  3.465832e-06, 7.517797e-06, 1.340323e-05, 3.646447e-05, 5.249749e-05, 
    4.389478e-05, 5.834559e-05, 0.0001449542, 0.0003173531, 0.0003669916, 
    0.0002721544, 0.0001388577, 9.442364e-05, 7.660547e-05, 0.0001373235,
  1.237851e-07, 2.207291e-06, 4.061195e-06, 9.379102e-06, 2.028942e-05, 
    2.549235e-05, 6.263635e-06, 1.077348e-05, 8.353364e-05, 0.000145237, 
    0.0001277556, 7.304853e-05, 3.101014e-05, 1.597953e-05, 1.782445e-05,
  9.548097e-07, 2.76473e-07, 1.515511e-06, 3.03312e-06, 7.123107e-06, 
    1.219895e-05, 4.950852e-05, 0.000130563, 0.0001066672, 9.377596e-05, 
    7.38698e-05, 3.272961e-05, 1.699078e-05, 1.186828e-05, 1.031762e-05,
  1.565653e-06, 1.416599e-07, 9.609749e-07, 3.576207e-07, 1.836416e-06, 
    2.075347e-05, 3.365929e-05, 0.0001314688, 0.0001588295, 0.000138438, 
    8.40658e-05, 3.486526e-05, 1.371482e-05, 1.019083e-05, 9.764975e-06,
  3.707755e-06, 4.861286e-08, 6.485578e-07, 1.693908e-07, 4.325567e-07, 
    3.102139e-06, 1.1163e-05, 3.731599e-05, 0.0001098789, 0.0001781629, 
    8.477592e-05, 4.39355e-05, 1.775905e-05, 9.815324e-06, 7.804753e-06,
  0.0005644531, 0.0005999646, 0.0004159408, 0.0002631785, 0.0001145523, 
    2.55625e-05, 1.058878e-05, 1.162394e-05, 1.668977e-05, 2.19693e-05, 
    1.720887e-05, 1.056524e-05, 9.100212e-06, 6.14608e-06, 3.40664e-06,
  0.000543915, 0.0005338993, 0.0005451309, 0.0003404232, 0.0001464353, 
    3.481123e-05, 1.088571e-05, 1.207163e-05, 1.774793e-05, 2.457888e-05, 
    3.709035e-05, 2.18132e-05, 1.146323e-05, 5.75e-06, 3.465703e-06,
  0.0003844195, 0.0005301629, 0.0005752204, 0.000445604, 0.0002135762, 
    7.713764e-05, 6.256809e-05, 0.0001167462, 0.0001505622, 0.0001742884, 
    0.0001246029, 7.701341e-05, 5.961345e-05, 9.677782e-05, 0.0001156806,
  0.0006245378, 0.0009142709, 0.0008748299, 0.0006560569, 0.0003888241, 
    0.0003575484, 0.0004460682, 0.0004280577, 0.0002985213, 0.0001527089, 
    7.881254e-05, 0.00010598, 0.0002466163, 0.0004234535, 0.0004098688,
  0.0009818668, 0.001610375, 0.001417744, 0.001247135, 0.001004018, 
    0.0007780853, 0.0005663615, 0.0003110382, 0.0002143212, 0.0001674484, 
    0.0001548162, 0.0002600768, 0.0005339509, 0.0007028258, 0.0006959653,
  0.001415387, 0.00139743, 0.001540411, 0.001232636, 0.0007925376, 
    0.0003451966, 0.0002209512, 0.0002230796, 0.0002380283, 0.0002420065, 
    0.0002831909, 0.0004228483, 0.0006438391, 0.0007404127, 0.0008153407,
  0.001068482, 0.001187983, 0.001055417, 0.0004729429, 9.564048e-05, 
    6.86514e-05, 3.041526e-05, 4.670055e-05, 0.0001318331, 0.0002499247, 
    0.0003421098, 0.0004613143, 0.000628292, 0.0007273646, 0.0007894045,
  0.000662385, 0.0008228495, 0.000602155, 0.00027729, 4.96276e-05, 
    9.335294e-05, 0.0002230118, 0.0003504878, 0.0003698519, 0.0003797512, 
    0.0004595659, 0.0004842116, 0.0005407823, 0.0006248986, 0.0006781837,
  0.0004762841, 0.0006441596, 0.0004518977, 0.000180148, 0.0002526475, 
    0.0003704048, 0.0005546716, 0.0007804373, 0.0007671732, 0.0006883983, 
    0.0005179457, 0.0004564986, 0.0004415207, 0.0004418095, 0.0005207983,
  0.0002879444, 0.0004503635, 0.0003300597, 0.0001457256, 0.0001703914, 
    0.0002855639, 0.0007468352, 0.0008440068, 0.0009505532, 0.0007587889, 
    0.0004478939, 0.0003175647, 0.0002363859, 0.0002378345, 0.000311356,
  3.03834e-05, 5.310642e-05, 6.281819e-05, 5.768153e-05, 4.666533e-05, 
    3.564675e-05, 3.053524e-05, 4.850873e-05, 4.426167e-05, 3.206457e-05, 
    2.643877e-05, 3.001903e-05, 3.39989e-05, 2.705382e-05, 1.409394e-05,
  8.589594e-06, 1.900768e-05, 2.726897e-05, 3.206736e-05, 5.088198e-05, 
    5.102334e-05, 4.244351e-05, 3.81251e-05, 4.881856e-05, 4.257614e-05, 
    3.673405e-05, 3.975216e-05, 3.803817e-05, 2.718702e-05, 1.279767e-05,
  9.070781e-06, 7.275713e-06, 7.504122e-06, 1.231597e-05, 3.759408e-05, 
    5.894903e-05, 6.613827e-05, 6.375879e-05, 5.857366e-05, 5.245351e-05, 
    4.765923e-05, 4.253921e-05, 3.538469e-05, 2.703088e-05, 1.404855e-05,
  4.100274e-05, 3.101249e-05, 9.162056e-06, 1.443088e-05, 3.316477e-05, 
    5.019623e-05, 5.61626e-05, 6.321008e-05, 6.111046e-05, 5.907515e-05, 
    5.03949e-05, 4.920793e-05, 4.110007e-05, 1.594338e-05, 1.364748e-05,
  0.0001495327, 0.000118533, 5.120762e-05, 2.793493e-05, 3.43475e-05, 
    4.958733e-05, 5.93868e-05, 6.311731e-05, 6.619644e-05, 5.61835e-05, 
    4.891849e-05, 3.886403e-05, 3.341332e-05, 2.169994e-05, 1.669219e-05,
  0.0003758459, 0.0002308713, 0.0001311479, 6.200188e-05, 4.158589e-05, 
    4.584304e-05, 5.67204e-05, 5.50735e-05, 6.0669e-05, 5.757591e-05, 
    4.393943e-05, 2.628726e-05, 3.388234e-05, 2.403606e-05, 1.445851e-05,
  0.0003881477, 0.0002526218, 0.0001418759, 5.72106e-05, 3.950913e-05, 
    4.846515e-05, 3.671945e-05, 5.208908e-05, 4.402103e-05, 3.774082e-05, 
    3.348885e-05, 3.093592e-05, 2.651431e-05, 1.678933e-05, 1.365736e-05,
  0.000354466, 0.0002857706, 0.0001620463, 8.219843e-05, 5.543416e-05, 
    6.340355e-05, 5.651554e-05, 4.367315e-05, 2.674948e-05, 1.931974e-05, 
    2.799133e-05, 2.964512e-05, 1.976064e-05, 1.833242e-05, 1.408651e-05,
  0.0004600985, 0.0004349741, 0.0003092188, 0.000210829, 0.0002507624, 
    0.0001982588, 0.0001156833, 2.518313e-05, 2.203334e-05, 3.516179e-05, 
    2.924698e-05, 2.892754e-05, 2.406236e-05, 2.047877e-05, 1.286337e-05,
  0.0005288279, 0.0004630972, 0.0003370371, 0.0002520929, 0.0002710838, 
    0.0003449528, 0.0003658024, 0.0001345091, 0.0001649674, 0.0001402265, 
    0.0001006907, 0.0001410191, 5.239965e-05, 4.190493e-05, 2.895388e-05,
  2.122744e-07, 8.410648e-07, 4.97436e-07, 2.051588e-09, 2.489415e-08, 
    3.279952e-08, 5.157307e-08, 3.264063e-07, 5.121421e-07, 4.893199e-07, 
    2.619034e-07, 8.729634e-07, 2.837354e-06, 4.206253e-06, 3.78162e-06,
  2.127498e-06, 4.180558e-06, 1.453969e-06, 2.288655e-08, 5.74145e-07, 
    5.803166e-07, 3.862592e-07, 8.120912e-07, 4.073066e-07, 9.020895e-07, 
    2.230934e-06, 1.989486e-06, 3.38765e-06, 4.078692e-06, 2.310808e-06,
  1.582415e-05, 6.798149e-06, 2.131005e-06, 6.041833e-06, 4.921813e-06, 
    2.069488e-06, 3.619919e-06, 2.536692e-06, 2.630788e-06, 3.875688e-06, 
    5.896643e-06, 4.577901e-06, 8.18889e-06, 5.570773e-06, 6.358659e-06,
  2.426996e-05, 1.736721e-05, 3.190295e-06, 1.778147e-05, 1.297375e-05, 
    7.342039e-06, 5.899168e-06, 6.990629e-06, 7.974981e-06, 9.532071e-06, 
    9.23714e-06, 8.295061e-06, 1.009234e-05, 7.986493e-06, 7.799134e-06,
  9.475942e-06, 1.163421e-05, 1.851481e-05, 2.303096e-05, 2.595011e-05, 
    2.038111e-05, 1.642416e-05, 8.91016e-06, 1.149332e-05, 1.187168e-05, 
    1.48286e-05, 1.557012e-05, 1.638836e-05, 1.143664e-05, 6.367713e-06,
  9.27774e-06, 1.321031e-05, 1.518719e-05, 3.154239e-05, 4.321263e-05, 
    2.865534e-05, 2.919012e-05, 2.338026e-05, 1.830123e-05, 1.57186e-05, 
    1.447464e-05, 1.224069e-05, 1.378927e-05, 1.198572e-05, 7.187587e-06,
  3.020737e-05, 1.232664e-05, 2.36052e-05, 5.135558e-05, 7.124221e-05, 
    1.181864e-05, 4.817623e-06, 1.770221e-05, 1.829507e-05, 1.422427e-05, 
    1.278152e-05, 1.318642e-05, 1.179134e-05, 1.0664e-05, 8.555121e-06,
  6.93714e-05, 4.659852e-05, 5.761384e-05, 7.60539e-05, 8.051129e-05, 
    4.364568e-05, 1.355344e-05, 8.735276e-06, 8.189513e-06, 7.28474e-06, 
    1.468436e-05, 1.448454e-05, 1.276349e-05, 1.363194e-05, 1.217752e-05,
  3.042981e-05, 4.467179e-05, 7.271588e-05, 0.0001024534, 0.0001583559, 
    6.802049e-05, 4.618955e-05, 1.104288e-05, 1.323136e-05, 1.752028e-05, 
    1.983989e-05, 1.620695e-05, 1.479157e-05, 1.297917e-05, 1.333379e-05,
  1.962465e-05, 4.240709e-05, 7.231311e-05, 9.928788e-05, 8.161125e-05, 
    7.995354e-05, 4.782496e-05, 3.033636e-05, 3.30062e-05, 2.505324e-05, 
    2.451218e-05, 1.716927e-05, 1.543979e-05, 1.609288e-05, 1.587057e-05,
  1.454711e-09, 7.120111e-11, 1.954335e-11, 3.598152e-11, 2.239704e-11, 
    4.815394e-12, 2.172517e-12, 7.482155e-11, 1.11894e-10, 1.117854e-10, 
    3.598652e-10, 2.730145e-08, 3.116336e-09, 3.108123e-08, 9.9122e-09,
  1.457774e-08, 1.662436e-08, 1.210485e-09, 2.516812e-11, 2.518847e-12, 
    1.602578e-13, 6.575253e-13, 2.622789e-12, 2.402731e-09, 5.222998e-09, 
    8.185832e-08, 1.291714e-07, 5.305575e-08, 1.684897e-07, 6.49929e-08,
  5.86789e-07, 1.421404e-07, 1.759255e-08, 2.259386e-09, 1.749496e-12, 
    2.539522e-12, 1.313091e-12, 1.454605e-12, 1.152875e-07, 2.04375e-08, 
    3.100922e-09, 4.601293e-07, 9.947254e-07, 2.495592e-07, 3.031666e-07,
  4.717519e-07, 5.250713e-07, 3.627355e-08, 1.189498e-07, 2.608176e-08, 
    1.596155e-07, 2.662761e-07, 4.769598e-07, 4.327619e-08, 1.123975e-07, 
    1.033175e-07, 7.420845e-07, 1.693907e-06, 3.99822e-07, 1.206738e-07,
  7.346847e-07, 6.818588e-07, 1.288936e-07, 3.435663e-07, 1.476821e-06, 
    2.317924e-06, 1.26156e-06, 2.068021e-07, 2.726551e-08, 9.131754e-08, 
    8.050314e-07, 1.036346e-06, 7.047687e-07, 4.511173e-07, 7.122683e-07,
  1.335032e-06, 5.22993e-07, 8.652372e-08, 1.817534e-07, 5.449075e-06, 
    2.175624e-06, 4.6141e-06, 3.970169e-06, 2.751982e-06, 2.499915e-06, 
    5.142483e-06, 2.273405e-06, 1.150091e-06, 2.627493e-06, 4.357785e-07,
  2.290397e-05, 5.924038e-06, 4.480887e-06, 9.876842e-06, 1.827004e-05, 
    8.77566e-06, 3.169987e-06, 2.130401e-06, 3.356566e-06, 3.087919e-06, 
    4.289465e-06, 2.504789e-06, 1.977272e-06, 2.933229e-06, 2.146892e-06,
  2.22799e-05, 4.821749e-05, 4.370018e-05, 4.594567e-05, 3.781278e-05, 
    2.38973e-05, 1.995086e-05, 1.319332e-05, 2.594868e-06, 2.761852e-07, 
    4.13284e-06, 4.539948e-06, 2.376365e-06, 2.553033e-06, 1.85692e-06,
  2.887649e-05, 3.028112e-05, 6.004564e-05, 6.796604e-05, 7.844667e-05, 
    3.350213e-05, 2.147102e-05, 2.818688e-06, 9.84853e-07, 4.237888e-06, 
    7.223876e-06, 7.1524e-06, 5.155586e-06, 2.463903e-06, 2.597002e-06,
  2.302281e-05, 3.915787e-05, 6.468694e-05, 7.670515e-05, 4.100386e-05, 
    5.377835e-05, 2.739995e-05, 1.920432e-05, 1.876308e-05, 1.265719e-05, 
    1.302626e-05, 9.167364e-06, 6.529864e-06, 6.478246e-06, 4.85517e-06,
  3.355199e-08, 5.569781e-08, 1.749633e-07, 2.849362e-07, 3.817432e-07, 
    2.667648e-07, 1.312489e-07, 3.502138e-08, 4.074842e-08, 6.277136e-07, 
    1.474795e-06, 2.201952e-06, 2.605085e-06, 8.782621e-06, 2.162668e-05,
  7.459321e-08, 8.993763e-08, 3.760848e-08, 1.011972e-07, 2.621793e-07, 
    1.810158e-07, 7.20157e-08, 1.218053e-08, 1.394717e-09, 1.254274e-09, 
    1.300731e-08, 5.114368e-07, 2.025598e-06, 5.713342e-06, 9.479854e-06,
  3.247396e-08, 4.973514e-08, 3.413163e-08, 6.305912e-08, 1.574729e-07, 
    2.113809e-07, 6.369007e-08, 9.354332e-09, 2.305251e-08, 3.281932e-08, 
    1.483327e-08, 4.098955e-09, 4.782897e-07, 1.977745e-06, 2.163282e-06,
  4.666219e-08, 1.902752e-08, 7.449267e-09, 1.197768e-08, 4.397502e-08, 
    1.235712e-07, 1.788861e-07, 2.330582e-08, 1.635752e-08, 2.753633e-08, 
    6.454416e-09, 1.363907e-10, 1.451236e-07, 5.276256e-07, 4.769133e-07,
  8.178739e-08, 2.170961e-08, 2.158303e-09, 1.881642e-08, 1.045814e-08, 
    5.013138e-08, 1.271453e-07, 5.683192e-08, 3.353635e-08, 1.198263e-07, 
    9.472726e-08, 1.842436e-07, 1.876027e-07, 1.152598e-07, 8.242782e-08,
  2.758269e-07, 3.201361e-07, 8.759057e-09, 1.150838e-08, 3.448543e-09, 
    1.292528e-08, 2.603374e-08, 3.510088e-09, 4.792484e-08, 6.273672e-08, 
    4.10151e-07, 1.405325e-06, 1.004248e-06, 5.658289e-07, 1.492645e-08,
  1.261553e-06, 1.896832e-06, 9.060982e-07, 1.429141e-06, 9.218553e-07, 
    4.191215e-10, 1.192994e-09, 4.761561e-10, 4.491715e-10, 4.452644e-08, 
    1.309902e-07, 6.701307e-07, 4.045206e-06, 1.238564e-06, 9.606768e-09,
  7.632507e-06, 1.269606e-05, 1.776997e-05, 1.422654e-05, 3.615223e-06, 
    9.362123e-08, 1.441204e-08, 1.736161e-08, 2.28582e-11, 9.857215e-10, 
    4.310129e-07, 9.932513e-07, 3.866006e-06, 1.024717e-06, 6.686359e-07,
  1.341545e-05, 2.737062e-05, 3.165657e-05, 2.764329e-05, 3.637803e-05, 
    6.023433e-07, 1.240279e-08, 4.96788e-11, 4.41301e-09, 1.03905e-10, 
    4.484401e-08, 5.490743e-07, 2.214325e-06, 8.582503e-07, 5.415455e-07,
  2.033662e-05, 4.694391e-05, 4.275507e-05, 4.053915e-05, 2.10704e-05, 
    1.058423e-05, 1.128867e-06, 1.302408e-07, 1.77033e-07, 8.134732e-08, 
    1.83175e-07, 3.20945e-07, 7.72477e-07, 4.111274e-07, 2.367997e-06,
  0.0001883411, 0.0001723533, 0.0001435833, 9.489965e-05, 6.864218e-05, 
    6.616501e-05, 8.938572e-05, 0.0001347382, 0.0001890509, 0.0002345877, 
    0.0002459899, 0.0002321388, 0.000222421, 0.0002790197, 0.0003196051,
  0.0001901775, 0.0002123547, 0.0002171542, 0.0001641145, 0.0001463241, 
    0.0001300129, 0.0001358781, 0.0001456396, 0.0001973605, 0.0002484284, 
    0.0002755804, 0.0002463316, 0.0002420089, 0.0003173178, 0.0003450139,
  0.0001580165, 0.000194933, 0.0002201682, 0.0002204939, 0.0002199517, 
    0.0001977566, 0.0001813707, 0.0001716983, 0.000201857, 0.000255471, 
    0.0002879158, 0.000282212, 0.0002579605, 0.0003089588, 0.000313777,
  0.0001192151, 0.0001746174, 0.0001692276, 0.0002267623, 0.0002423647, 
    0.0002262294, 0.0002064442, 0.0002252756, 0.0002289749, 0.0002673835, 
    0.0002908784, 0.0002891016, 0.0002631954, 0.000306761, 0.0003141493,
  0.0001184864, 0.0001500003, 0.0001474468, 0.0001880949, 0.0002137769, 
    0.0002225159, 0.0002227176, 0.0002346951, 0.0002591414, 0.000289524, 
    0.0003008028, 0.0002914328, 0.0002935329, 0.0002893462, 0.0002919777,
  0.0001668456, 0.0001319362, 0.0001465939, 0.0001672624, 0.0001850824, 
    0.0001999733, 0.0002114683, 0.0002345409, 0.0002663542, 0.0003004431, 
    0.0003033994, 0.0002855214, 0.0003007848, 0.0002941965, 0.0002522142,
  9.139508e-05, 0.0001302824, 0.000142469, 0.0001503526, 0.0001689833, 
    0.0001541653, 0.0001696756, 0.0002113138, 0.0002487785, 0.0002864654, 
    0.0002821402, 0.0002745666, 0.0002836987, 0.0002943385, 0.0002529978,
  2.978744e-05, 7.309848e-05, 0.0001276608, 0.0001405578, 0.0001405269, 
    0.0001664953, 0.0001836603, 0.0002005228, 0.0002598042, 0.0002800404, 
    0.0002713612, 0.0002397974, 0.0002354812, 0.0002625502, 0.0002454514,
  1.185325e-05, 2.956405e-05, 7.040406e-05, 6.878563e-05, 0.0001352839, 
    0.0001645404, 0.000190411, 0.0002363307, 0.0002560254, 0.0002773251, 
    0.0002556429, 0.0002035028, 0.0001777258, 0.0002161008, 0.0002166364,
  8.317102e-06, 1.08081e-05, 2.28288e-05, 1.635668e-05, 7.500294e-05, 
    0.0001017576, 0.0001557563, 0.0002637788, 0.0002912965, 0.000287412, 
    0.0002609, 0.0001916298, 0.0001586708, 0.0001849195, 0.0001885979,
  0.0001104604, 0.000142642, 0.0001389716, 0.0001167151, 0.0001033445, 
    4.968952e-05, 2.948864e-05, 1.793543e-05, 1.167234e-05, 5.187586e-06, 
    3.660546e-07, 6.79087e-07, 7.723431e-07, 1.186151e-06, 9.646119e-07,
  0.000101573, 9.448264e-05, 0.000152294, 0.0001139615, 0.0001098458, 
    8.016864e-05, 4.367275e-05, 2.729846e-05, 1.803712e-05, 7.514627e-06, 
    1.348453e-06, 1.735909e-06, 1.691373e-06, 1.175918e-06, 7.992056e-07,
  4.689653e-05, 3.57344e-05, 7.790122e-05, 0.0001294554, 0.0001392707, 
    0.000101077, 6.991401e-05, 3.903859e-05, 2.476009e-05, 6.709222e-06, 
    5.119159e-06, 3.2209e-06, 2.957067e-06, 3.594564e-06, 1.610188e-06,
  4.935279e-05, 2.439867e-05, 3.96107e-05, 0.0001321618, 0.000120855, 
    0.0001084933, 8.84363e-05, 5.632616e-05, 2.874555e-05, 1.456585e-05, 
    1.011281e-05, 6.492266e-06, 4.432512e-06, 3.527764e-06, 2.680595e-06,
  1.974646e-05, 7.028887e-06, 2.911137e-05, 0.0001083583, 0.0001290947, 
    0.0001218104, 9.718558e-05, 6.770252e-05, 4.083604e-05, 2.593139e-05, 
    1.922869e-05, 1.262684e-05, 1.030025e-05, 5.048417e-06, 4.565927e-06,
  3.189903e-05, 2.405898e-05, 3.317694e-05, 7.909895e-05, 0.0001324997, 
    0.0001141685, 0.0001411189, 9.785991e-05, 7.036716e-05, 5.96594e-05, 
    2.889955e-05, 1.511763e-05, 1.203329e-05, 9.411507e-06, 5.043927e-06,
  8.100648e-05, 5.292022e-05, 7.358558e-05, 9.948372e-05, 0.0001454121, 
    6.41031e-05, 5.753131e-05, 0.0001191408, 9.951564e-05, 7.231237e-05, 
    5.235123e-05, 2.664307e-05, 1.580743e-05, 1.526126e-05, 9.116463e-06,
  0.0001875994, 0.0001676804, 0.0001636576, 0.0001699495, 0.0001649768, 
    0.0001303465, 5.399491e-05, 5.556368e-05, 8.56985e-05, 7.413603e-05, 
    5.980902e-05, 3.496156e-05, 2.001943e-05, 1.937166e-05, 1.481204e-05,
  0.0001689307, 0.0001962021, 0.0002294044, 0.000230213, 0.0002298062, 
    0.0001040777, 9.132244e-05, 7.061319e-05, 6.48679e-05, 6.163229e-05, 
    5.7673e-05, 6.030922e-05, 2.355581e-05, 2.204707e-05, 2.025985e-05,
  0.000137107, 0.0001729866, 0.00022789, 0.0002204182, 0.0001646391, 
    0.0001998107, 0.0001505048, 0.000105247, 7.86274e-05, 6.345497e-05, 
    5.795782e-05, 5.411956e-05, 6.034541e-05, 2.819122e-05, 2.641945e-05,
  4.836934e-05, 5.561973e-05, 5.888485e-05, 5.673816e-05, 4.457131e-05, 
    3.226759e-05, 2.305911e-05, 1.28271e-05, 7.172619e-06, 5.017963e-06, 
    3.942131e-07, 6.639094e-07, 2.618289e-06, 6.628097e-06, 9.246719e-06,
  4.044103e-05, 2.511457e-05, 4.456825e-05, 4.956541e-05, 4.592454e-05, 
    2.315745e-05, 1.752801e-05, 1.006077e-05, 4.709484e-06, 8.972418e-07, 
    4.194486e-07, 2.831033e-06, 9.502943e-06, 1.238804e-05, 1.276805e-05,
  1.58869e-05, 7.3803e-06, 1.874337e-05, 3.342707e-05, 3.634572e-05, 
    3.646032e-05, 7.472371e-06, 6.378107e-06, 2.447847e-06, 1.500265e-06, 
    9.750099e-07, 1.48115e-06, 6.707403e-06, 2.632299e-05, 1.773045e-05,
  3.927915e-06, 7.745091e-07, 9.102437e-07, 1.021992e-05, 2.724688e-05, 
    3.647524e-05, 1.971263e-05, 1.306366e-05, 9.959114e-06, 4.878852e-06, 
    4.280836e-06, 1.004714e-05, 1.024499e-05, 1.277556e-05, 1.66819e-05,
  3.402806e-07, 4.697419e-08, 1.470164e-07, 2.982405e-06, 2.623619e-05, 
    3.57972e-05, 2.895278e-05, 2.614515e-05, 2.42204e-05, 2.108758e-05, 
    1.693309e-05, 2.2465e-05, 2.92096e-05, 1.674655e-05, 1.420205e-05,
  3.741734e-06, 1.463914e-07, 5.073491e-08, 2.112019e-06, 3.485263e-05, 
    4.503803e-05, 4.938204e-05, 4.526637e-05, 4.472592e-05, 4.141944e-05, 
    3.170779e-05, 2.724829e-05, 3.935424e-05, 3.128343e-05, 1.603179e-05,
  3.629354e-05, 7.135188e-06, 2.90158e-06, 1.399327e-05, 5.26409e-05, 
    6.182869e-05, 3.929001e-05, 5.6477e-05, 4.376614e-05, 5.42305e-05, 
    5.892562e-05, 3.005498e-05, 3.239578e-05, 2.812931e-05, 2.472983e-05,
  0.0001157218, 6.58961e-05, 4.679286e-05, 6.063775e-05, 7.405003e-05, 
    7.754221e-05, 5.207862e-05, 4.643533e-05, 2.859836e-05, 5.502256e-06, 
    6.472833e-05, 5.892229e-05, 4.862127e-05, 3.342827e-05, 2.31266e-05,
  0.0001337016, 0.0001307414, 9.791473e-05, 0.0001318911, 8.962185e-05, 
    8.110543e-05, 5.416615e-05, 1.993459e-05, 6.322297e-06, 4.284824e-06, 
    5.50557e-05, 6.446628e-05, 5.671247e-05, 5.346335e-05, 3.558835e-05,
  7.53244e-05, 0.000116779, 0.0001755016, 0.0001838515, 0.0001204234, 
    0.0001000002, 4.518341e-05, 2.431873e-05, 1.892006e-05, 2.531518e-05, 
    5.08258e-05, 6.190947e-05, 6.569071e-05, 5.47244e-05, 4.2368e-05,
  1.13805e-05, 1.278107e-05, 1.367747e-05, 1.323365e-05, 9.198039e-06, 
    4.772246e-06, 2.457058e-06, 1.233942e-07, 2.194936e-07, 7.199296e-08, 
    2.942153e-07, 1.85877e-06, 1.584014e-05, 1.363579e-05, 1.342771e-05,
  4.357711e-06, 5.185224e-06, 7.014838e-06, 1.074527e-05, 9.153013e-06, 
    2.191599e-06, 2.248813e-07, 2.548169e-07, 3.972146e-07, 2.634907e-07, 
    2.626512e-06, 7.423644e-06, 1.745327e-05, 1.473957e-05, 1.168617e-05,
  3.139941e-07, 1.80674e-07, 2.488085e-07, 4.865497e-06, 1.237616e-05, 
    1.359424e-05, 7.275891e-06, 2.549109e-06, 3.330026e-06, 2.07832e-06, 
    4.994766e-06, 4.287962e-06, 1.158724e-05, 1.196955e-05, 7.521786e-06,
  3.42044e-09, 3.032075e-09, 2.867157e-09, 4.100969e-07, 7.619658e-06, 
    1.949626e-05, 1.089544e-05, 1.758959e-05, 1.732425e-05, 1.713344e-06, 
    5.994169e-06, 1.959014e-05, 2.595237e-05, 1.033008e-05, 7.591115e-06,
  6.172742e-10, 3.29e-11, 1.296541e-11, 2.189412e-09, 2.891644e-06, 
    1.64418e-05, 1.481856e-05, 2.21766e-05, 2.588106e-05, 2.665657e-05, 
    2.978517e-05, 2.624138e-05, 2.917012e-05, 2.189726e-05, 1.639235e-05,
  2.126947e-06, 3.135191e-09, 4.667977e-12, 1.891531e-12, 7.557722e-07, 
    3.95392e-06, 1.996001e-05, 1.904382e-05, 2.737325e-05, 2.877858e-05, 
    3.03137e-05, 2.495055e-05, 2.425692e-05, 2.563303e-05, 2.210642e-05,
  6.601821e-06, 2.207742e-06, 1.549628e-06, 1.300428e-06, 6.040166e-07, 
    1.685855e-06, 3.179924e-06, 1.315874e-05, 1.496316e-05, 2.279583e-05, 
    2.861402e-05, 2.757152e-05, 2.883628e-05, 2.90598e-05, 2.251183e-05,
  5.147477e-05, 3.977394e-05, 2.664464e-05, 2.123908e-05, 1.368466e-05, 
    6.51375e-06, 1.394204e-06, 8.704064e-07, 9.737006e-07, 4.847073e-06, 
    2.171322e-05, 2.867557e-05, 3.296824e-05, 2.797842e-05, 1.962712e-05,
  5.741107e-05, 6.764478e-05, 6.761606e-05, 7.478656e-05, 6.496364e-05, 
    9.990519e-06, 2.481054e-06, 3.946529e-07, 9.319692e-07, 3.11766e-06, 
    1.384611e-05, 2.403761e-05, 2.893566e-05, 2.497416e-05, 1.743624e-05,
  3.611513e-05, 6.142934e-05, 8.213007e-05, 0.0001014213, 4.509809e-05, 
    2.891764e-05, 1.43469e-05, 1.361047e-06, 5.347152e-06, 7.019532e-06, 
    1.332422e-05, 2.206685e-05, 3.272308e-05, 2.458983e-05, 1.744831e-05,
  1.624783e-05, 1.742888e-05, 1.459924e-05, 6.37914e-06, 4.105726e-07, 
    6.397372e-09, 3.763831e-10, 1.461367e-10, 1.38799e-07, 1.466227e-07, 
    9.910807e-07, 3.030261e-06, 6.469217e-06, 7.983588e-06, 6.054984e-06,
  3.852852e-06, 6.555086e-07, 1.348144e-05, 9.244832e-06, 8.303158e-06, 
    9.693414e-07, 1.486422e-07, 8.653574e-08, 2.78475e-07, 2.447219e-06, 
    3.620682e-06, 5.218234e-06, 8.984921e-06, 6.088527e-06, 6.45524e-06,
  4.561432e-06, 2.306469e-06, 3.516796e-07, 9.735882e-06, 1.431607e-05, 
    8.462032e-06, 3.214859e-06, 1.890088e-06, 2.904463e-06, 4.372942e-06, 
    7.946458e-06, 1.118284e-05, 1.133091e-05, 8.76456e-06, 7.841076e-06,
  7.574112e-06, 3.664069e-06, 2.831831e-07, 1.788938e-05, 2.239837e-05, 
    1.927642e-05, 1.353822e-05, 1.487974e-05, 1.184733e-05, 1.231403e-05, 
    1.362755e-05, 1.42522e-05, 1.371531e-05, 8.819276e-06, 9.559119e-06,
  4.59169e-06, 3.668021e-06, 1.055787e-06, 1.816311e-05, 2.705782e-05, 
    3.182104e-05, 2.523105e-05, 2.376287e-05, 2.057005e-05, 2.146199e-05, 
    1.857863e-05, 2.026998e-05, 1.550048e-05, 1.232754e-05, 1.157715e-05,
  1.180611e-05, 7.0105e-06, 6.059474e-06, 1.753318e-05, 2.929499e-05, 
    1.663348e-05, 2.851691e-05, 2.739685e-05, 2.513072e-05, 2.881973e-05, 
    2.337801e-05, 1.649813e-05, 1.463125e-05, 1.632716e-05, 1.319267e-05,
  1.20026e-05, 1.311149e-05, 2.266976e-05, 4.236726e-05, 3.608079e-05, 
    4.291776e-06, 3.745829e-07, 1.038039e-05, 1.699931e-05, 1.912065e-05, 
    2.178666e-05, 1.887811e-05, 1.796751e-05, 1.762196e-05, 1.320414e-05,
  2.694192e-05, 2.408247e-05, 2.499529e-05, 4.666338e-05, 3.63032e-05, 
    2.4434e-05, 1.422818e-05, 8.415966e-06, 2.255382e-06, 1.111621e-05, 
    1.584474e-05, 1.786143e-05, 1.936518e-05, 1.809164e-05, 1.474512e-05,
  3.778307e-05, 3.779528e-05, 5.593531e-05, 4.578951e-05, 5.964286e-05, 
    2.876204e-05, 1.070553e-05, 6.489795e-06, 1.328822e-05, 2.084756e-05, 
    1.95199e-05, 2.055186e-05, 1.691902e-05, 1.635805e-05, 1.318623e-05,
  4.183383e-05, 5.082777e-05, 6.059113e-05, 2.577707e-05, 3.227045e-05, 
    2.270508e-05, 1.457828e-05, 1.053307e-05, 2.690231e-05, 2.174506e-05, 
    2.257015e-05, 2.000101e-05, 1.770777e-05, 1.444581e-05, 1.07131e-05,
  4.208287e-05, 3.686226e-05, 3.590416e-05, 2.484374e-05, 7.95391e-06, 
    9.065766e-07, 1.99832e-08, 6.528827e-09, 8.516477e-11, 1.916563e-13, 
    1.705194e-25, 5.698356e-10, 5.062887e-08, 2.660009e-07, 1.241079e-07,
  3.70694e-05, 1.605931e-05, 2.89003e-05, 2.370362e-05, 2.08382e-05, 
    3.761983e-06, 5.180612e-08, 4.046033e-08, 1.848182e-08, 2.806361e-10, 
    5.440195e-18, 1.527714e-07, 1.657802e-07, 2.534188e-07, 4.530708e-07,
  1.66717e-05, 1.160308e-05, 1.013381e-05, 2.36316e-05, 2.993047e-05, 
    1.730963e-05, 5.450529e-06, 1.3129e-06, 1.096329e-07, 2.137516e-07, 
    2.719271e-07, 1.298948e-06, 4.504735e-07, 5.413487e-07, 9.379063e-07,
  1.054332e-05, 2.625912e-06, 3.094894e-06, 2.927275e-05, 3.545982e-05, 
    2.953319e-05, 2.526526e-05, 1.371848e-05, 3.500105e-06, 3.380279e-06, 
    3.97001e-06, 3.538056e-06, 3.376503e-06, 1.182491e-06, 1.403069e-06,
  1.344813e-07, 8.339401e-07, 2.227e-06, 2.365736e-05, 4.025599e-05, 
    4.649653e-05, 3.17555e-05, 2.807472e-05, 2.014807e-05, 1.998239e-05, 
    1.133139e-05, 1.393371e-05, 8.494053e-06, 2.588377e-06, 2.492356e-06,
  5.216194e-06, 5.314562e-06, 4.988046e-06, 2.003704e-05, 4.005498e-05, 
    2.899314e-05, 3.367742e-05, 4.403637e-05, 3.848525e-05, 3.70632e-05, 
    3.839755e-05, 1.907387e-05, 1.564702e-05, 7.606255e-06, 3.767745e-06,
  2.084786e-05, 1.764066e-05, 2.509987e-05, 4.296415e-05, 5.972114e-05, 
    2.100362e-05, 1.018569e-05, 1.610263e-05, 3.034116e-05, 3.265448e-05, 
    5.117295e-05, 3.230712e-05, 1.869959e-05, 1.023601e-05, 7.554572e-06,
  0.0001144211, 7.516541e-05, 6.881393e-05, 7.545666e-05, 7.770184e-05, 
    4.179553e-05, 1.701837e-05, 9.022328e-06, 6.295477e-06, 1.228193e-05, 
    4.476487e-05, 4.049786e-05, 2.199827e-05, 1.548743e-05, 1.525346e-05,
  0.0001365022, 0.0001278744, 0.0001253362, 0.0001263858, 0.0001347442, 
    2.981348e-05, 2.010404e-05, 4.75359e-06, 9.659207e-06, 2.433879e-05, 
    4.772737e-05, 4.113365e-05, 2.853452e-05, 1.792582e-05, 1.804481e-05,
  0.0001200872, 0.0001252383, 0.0001331362, 0.0001333975, 1.50973e-05, 
    3.943366e-05, 3.574725e-05, 1.203282e-05, 2.706164e-05, 3.512343e-05, 
    5.327518e-05, 4.544612e-05, 3.035415e-05, 2.004006e-05, 2.134674e-05,
  2.994099e-05, 2.568687e-05, 2.280843e-05, 1.98591e-05, 2.8999e-06, 
    4.119551e-07, 1.730217e-09, 7.159048e-10, 2.308453e-09, 1.149017e-08, 
    1.688537e-06, 5.649827e-06, 3.20923e-06, 6.809973e-07, 4.251813e-08,
  1.884439e-05, 1.666015e-05, 1.733499e-05, 1.574523e-05, 1.115462e-05, 
    2.849431e-06, 2.536373e-07, 4.482434e-09, 1.347506e-07, 6.241606e-07, 
    4.120212e-06, 5.276328e-06, 3.712929e-06, 1.13726e-06, 5.20305e-09,
  8.076184e-06, 1.012874e-05, 1.950654e-05, 2.183564e-05, 2.967852e-05, 
    2.82145e-05, 1.125894e-05, 3.915751e-06, 2.552258e-06, 6.883941e-06, 
    7.844829e-06, 9.42419e-06, 4.795475e-06, 2.123656e-06, 4.798637e-09,
  1.789571e-06, 4.470788e-06, 1.403359e-05, 3.615431e-05, 4.867609e-05, 
    6.010027e-05, 6.78622e-05, 3.033723e-05, 1.470579e-05, 1.669682e-05, 
    2.017831e-05, 1.518402e-05, 5.089857e-06, 8.134984e-08, 2.570252e-09,
  1.807022e-07, 9.679176e-07, 8.782401e-06, 3.189741e-05, 6.38398e-05, 
    7.29262e-05, 6.683711e-05, 9.293074e-05, 5.763339e-05, 3.912687e-05, 
    3.199628e-05, 1.639074e-05, 5.326296e-06, 3.960318e-07, 2.38325e-07,
  1.510985e-07, 1.732419e-07, 5.378453e-06, 2.055001e-05, 5.512902e-05, 
    7.359104e-05, 9.236034e-05, 8.213778e-05, 7.802272e-05, 6.877738e-05, 
    4.92928e-05, 1.38354e-05, 5.887005e-06, 1.057589e-06, 2.698988e-07,
  1.852885e-06, 2.386082e-07, 3.500768e-06, 1.209835e-05, 4.17162e-05, 
    5.173345e-05, 4.602186e-05, 6.075392e-05, 6.449453e-05, 7.487081e-05, 
    6.311292e-05, 2.592791e-05, 1.151515e-05, 4.076094e-06, 1.62394e-06,
  4.385841e-05, 2.196502e-05, 1.443704e-05, 1.59989e-05, 2.918256e-05, 
    3.783788e-05, 3.218995e-05, 4.56888e-05, 4.186152e-05, 4.230484e-05, 
    4.940246e-05, 2.713512e-05, 1.423619e-05, 6.738722e-06, 5.111011e-06,
  5.857354e-05, 5.835582e-05, 5.911952e-05, 3.398906e-05, 3.893117e-05, 
    1.656658e-05, 1.749343e-05, 2.47914e-05, 5.512392e-05, 5.243445e-05, 
    5.291086e-05, 3.761894e-05, 2.332269e-05, 1.411665e-05, 1.109287e-05,
  5.699428e-05, 6.478175e-05, 7.574667e-05, 7.346788e-05, 1.420982e-05, 
    9.211558e-06, 1.192956e-05, 2.470659e-05, 2.90801e-05, 3.324775e-05, 
    5.006767e-05, 3.940324e-05, 2.948765e-05, 2.348037e-05, 1.425889e-05,
  4.866382e-05, 6.077504e-05, 8.387803e-05, 8.871555e-05, 6.246792e-05, 
    2.303719e-05, 6.539263e-06, 9.607596e-07, 2.867412e-08, 3.270264e-08, 
    2.542945e-08, 2.604277e-07, 1.325976e-06, 1.189212e-06, 2.157045e-06,
  2.531846e-05, 1.06916e-05, 3.49154e-05, 2.782753e-05, 5.170258e-05, 
    4.466759e-05, 1.640516e-05, 1.267819e-06, 2.780087e-07, 3.954175e-08, 
    9.530663e-08, 2.617776e-06, 2.842374e-06, 2.704672e-06, 2.947469e-06,
  1.712533e-06, 7.043012e-07, 3.461132e-06, 1.933248e-05, 4.245627e-05, 
    6.582289e-05, 5.162854e-05, 1.663537e-05, 5.363965e-06, 8.249196e-07, 
    1.491772e-06, 5.144732e-06, 6.071608e-06, 4.48003e-06, 4.372522e-06,
  1.549274e-07, 1.614925e-08, 4.671485e-08, 1.017378e-05, 4.402203e-05, 
    5.874953e-05, 8.571721e-05, 6.378589e-05, 3.802852e-05, 1.342299e-05, 
    5.125099e-06, 1.200357e-05, 1.446385e-05, 6.615213e-06, 7.379723e-06,
  1.05898e-07, 5.323647e-09, 1.383439e-09, 2.919707e-06, 3.771428e-05, 
    6.478439e-05, 6.397601e-05, 9.661741e-05, 7.284255e-05, 4.583303e-05, 
    2.006432e-05, 2.354642e-05, 2.435828e-05, 1.359886e-05, 1.24436e-05,
  3.336697e-07, 3.581726e-08, 1.656355e-08, 2.029065e-06, 2.63401e-05, 
    4.662081e-05, 6.122188e-05, 6.70741e-05, 8.62161e-05, 9.155463e-05, 
    6.32486e-05, 4.739988e-05, 3.30329e-05, 2.670093e-05, 1.401805e-05,
  2.013231e-05, 6.64141e-06, 7.081996e-06, 1.411984e-05, 3.889806e-05, 
    2.093559e-05, 1.538171e-05, 1.900534e-05, 3.71407e-05, 3.990652e-05, 
    8.58282e-05, 8.375746e-05, 6.480291e-05, 3.325166e-05, 1.970119e-05,
  9.010557e-05, 7.27101e-05, 5.757503e-05, 6.373625e-05, 6.537096e-05, 
    4.8267e-05, 1.248486e-05, 6.314243e-06, 5.254896e-06, 2.014514e-05, 
    5.586212e-05, 0.0001103926, 9.039846e-05, 5.475157e-05, 2.65041e-05,
  7.41057e-05, 0.0001014204, 0.0001251167, 0.0001390846, 0.0001011681, 
    3.841352e-05, 3.884535e-05, 2.309767e-05, 3.367378e-05, 4.641854e-05, 
    6.234446e-05, 0.0001264302, 0.0001013322, 6.088855e-05, 3.885525e-05,
  5.95084e-05, 6.775446e-05, 0.0001201031, 0.0001921498, 7.081099e-05, 
    5.870263e-05, 4.339673e-05, 5.310532e-05, 9.740371e-05, 7.883531e-05, 
    0.0001000234, 0.0001171667, 0.0001090041, 7.965004e-05, 4.807357e-05,
  4.085889e-05, 4.135105e-05, 7.082915e-05, 5.112936e-05, 2.586796e-05, 
    1.354158e-05, 3.180347e-06, 3.575919e-07, 4.59909e-07, 7.809164e-07, 
    2.47157e-06, 4.108776e-06, 1.155327e-05, 2.106657e-05, 2.245494e-05,
  1.560452e-05, 1.021495e-05, 2.254516e-05, 3.312869e-05, 3.858832e-05, 
    2.338545e-05, 1.191088e-05, 3.040791e-06, 5.689254e-07, 5.050563e-06, 
    6.961642e-06, 1.575724e-05, 2.084112e-05, 2.220865e-05, 2.099719e-05,
  1.657447e-06, 7.896524e-07, 1.301744e-06, 1.958097e-05, 4.387189e-05, 
    4.591639e-05, 2.787987e-05, 1.695028e-05, 1.003814e-05, 1.584928e-05, 
    2.334228e-05, 1.691239e-05, 1.914874e-05, 1.093493e-05, 1.024481e-05,
  4.490704e-08, 1.582196e-08, 3.656153e-08, 1.443075e-05, 3.697525e-05, 
    5.748394e-05, 4.596726e-05, 4.050766e-05, 3.45652e-05, 2.945779e-05, 
    2.833053e-05, 2.762043e-05, 2.267481e-05, 1.374021e-05, 1.211414e-05,
  2.163727e-08, 3.542288e-09, 2.954111e-08, 6.607729e-07, 2.894594e-05, 
    4.621928e-05, 4.72363e-05, 6.336279e-05, 5.952082e-05, 5.702391e-05, 
    3.989682e-05, 3.493985e-05, 3.000346e-05, 1.801181e-05, 1.276938e-05,
  5.0122e-07, 7.771185e-09, 1.459841e-07, 5.115153e-07, 1.050005e-05, 
    2.659944e-05, 3.971578e-05, 4.312275e-05, 5.651218e-05, 6.135127e-05, 
    5.703076e-05, 3.912981e-05, 3.576078e-05, 2.330669e-05, 1.643195e-05,
  1.400912e-05, 4.218809e-06, 2.265142e-06, 6.181618e-06, 1.668708e-05, 
    1.054774e-05, 3.943552e-06, 8.856352e-06, 1.543078e-05, 3.66203e-05, 
    5.272344e-05, 4.59874e-05, 3.403366e-05, 2.479426e-05, 1.940381e-05,
  7.021156e-05, 5.020709e-05, 4.269806e-05, 3.643509e-05, 3.364317e-05, 
    1.580368e-05, 2.316135e-06, 6.933668e-07, 8.654398e-07, 2.080575e-06, 
    1.664988e-05, 3.603497e-05, 4.35767e-05, 3.178079e-05, 2.231874e-05,
  8.421107e-05, 9.203158e-05, 8.934891e-05, 7.594622e-05, 7.29188e-05, 
    2.085267e-05, 5.836531e-06, 5.735862e-07, 8.596812e-07, 4.149883e-06, 
    1.24569e-05, 2.849368e-05, 3.289741e-05, 3.292176e-05, 2.583355e-05,
  7.250296e-05, 8.360673e-05, 0.0001057856, 0.0001173987, 2.864024e-05, 
    3.946032e-05, 1.710509e-05, 6.075704e-06, 1.342576e-05, 1.420806e-05, 
    1.774688e-05, 1.830975e-05, 2.494072e-05, 2.953771e-05, 2.828768e-05,
  3.573151e-05, 3.405432e-05, 6.777507e-05, 4.35162e-05, 1.504539e-05, 
    3.358985e-06, 8.061242e-07, 5.029209e-08, 3.412386e-08, 3.094568e-09, 
    4.636887e-08, 5.421453e-08, 1.0949e-07, 8.157463e-07, 1.881266e-06,
  5.999187e-06, 6.304564e-06, 1.43189e-05, 3.953475e-05, 2.902196e-05, 
    1.418773e-05, 3.160848e-06, 4.656869e-07, 6.188595e-07, 3.575688e-07, 
    6.735883e-07, 2.710786e-07, 3.346066e-07, 1.194247e-06, 3.334651e-06,
  2.294857e-07, 3.689657e-07, 6.729329e-06, 2.052623e-05, 5.234137e-05, 
    4.086899e-05, 2.040712e-05, 1.017727e-05, 3.423206e-06, 3.936532e-06, 
    1.972028e-06, 2.117446e-06, 1.987024e-06, 1.53304e-06, 3.911392e-06,
  6.709039e-09, 1.10844e-08, 1.050619e-06, 2.285445e-05, 6.299923e-05, 
    7.672222e-05, 4.740816e-05, 3.213051e-05, 1.384404e-05, 8.765482e-06, 
    5.968937e-06, 4.269877e-06, 5.31271e-06, 1.537079e-06, 2.153281e-06,
  9.324658e-09, 1.244217e-09, 1.458838e-07, 6.279261e-06, 5.132643e-05, 
    8.776729e-05, 9.70229e-05, 7.999587e-05, 4.531293e-05, 3.12045e-05, 
    1.397328e-05, 8.630102e-06, 8.989735e-06, 8.311002e-06, 6.036395e-06,
  1.281345e-06, 2.495939e-09, 1.070256e-07, 1.784319e-06, 3.195583e-05, 
    6.020999e-05, 7.311776e-05, 9.973486e-05, 9.473626e-05, 6.258516e-05, 
    3.600712e-05, 1.631817e-05, 9.995377e-06, 1.032347e-05, 1.112414e-05,
  2.159885e-05, 3.709104e-06, 5.269108e-06, 1.327137e-05, 3.823507e-05, 
    2.786251e-05, 2.477681e-05, 2.798889e-05, 4.101492e-05, 5.861062e-05, 
    5.9504e-05, 3.241167e-05, 1.403629e-05, 1.083482e-05, 1.113973e-05,
  8.876748e-05, 5.963711e-05, 4.946514e-05, 4.49247e-05, 4.487237e-05, 
    2.893289e-05, 6.142274e-06, 3.161544e-06, 4.772685e-06, 1.519511e-05, 
    3.963855e-05, 4.65763e-05, 2.789445e-05, 1.43653e-05, 1.448719e-05,
  9.273249e-05, 0.0001033346, 0.0001055776, 9.017731e-05, 7.917931e-05, 
    1.141544e-05, 1.024744e-05, 2.632932e-06, 6.87388e-06, 3.075779e-05, 
    4.015043e-05, 4.364952e-05, 4.293008e-05, 2.71218e-05, 1.636855e-05,
  7.016589e-05, 9.512855e-05, 0.0001291434, 0.0001303527, 1.57608e-05, 
    1.311832e-05, 1.087859e-05, 1.239263e-05, 1.983385e-05, 4.874144e-05, 
    4.622598e-05, 5.035842e-05, 4.824427e-05, 3.619998e-05, 2.540479e-05,
  1.967071e-05, 1.439839e-05, 9.694026e-06, 3.389308e-06, 5.737905e-07, 
    1.126843e-07, 1.532171e-07, 2.194703e-07, 4.285577e-07, 8.440729e-07, 
    3.718175e-06, 4.254202e-06, 4.201584e-06, 4.268528e-07, 3.010067e-07,
  1.471444e-05, 4.798724e-06, 1.339685e-05, 5.536009e-06, 1.931174e-06, 
    3.096196e-07, 1.141381e-07, 2.339706e-07, 5.264037e-07, 1.371086e-06, 
    3.579693e-06, 4.965298e-06, 4.741751e-06, 7.148017e-07, 6.458675e-07,
  2.269507e-05, 7.973373e-06, 2.143526e-06, 1.35814e-05, 8.699384e-06, 
    2.413771e-06, 1.25824e-06, 1.477071e-06, 1.139008e-06, 3.300675e-06, 
    4.706474e-06, 7.154688e-06, 5.330457e-06, 1.599167e-06, 7.52322e-07,
  2.962051e-05, 1.024824e-05, 3.937566e-06, 2.13262e-05, 1.809789e-05, 
    1.330051e-05, 4.961957e-06, 5.869967e-06, 4.041603e-06, 8.405992e-06, 
    8.922602e-06, 1.109516e-05, 5.435881e-06, 1.652307e-06, 5.850958e-07,
  2.12689e-05, 7.592468e-06, 8.490963e-06, 2.631155e-05, 3.416804e-05, 
    2.738737e-05, 1.923987e-05, 1.649988e-05, 1.564784e-05, 1.789802e-05, 
    1.882202e-05, 1.763743e-05, 1.112475e-05, 5.294843e-06, 1.291919e-06,
  2.112219e-05, 7.925691e-06, 1.301085e-05, 2.880068e-05, 3.800046e-05, 
    1.14754e-05, 2.355698e-05, 2.72695e-05, 2.191623e-05, 2.446126e-05, 
    2.708698e-05, 1.887424e-05, 1.633417e-05, 9.60241e-06, 3.300236e-06,
  3.674742e-05, 1.322612e-05, 3.107513e-05, 4.564699e-05, 2.523665e-05, 
    6.728176e-06, 1.09254e-06, 1.547701e-06, 1.367285e-05, 1.767889e-05, 
    2.654102e-05, 1.708879e-05, 1.40226e-05, 9.64732e-06, 3.403849e-06,
  0.0001002273, 5.330753e-05, 5.76569e-05, 6.355564e-05, 2.261669e-05, 
    7.396937e-06, 3.404458e-06, 3.090969e-06, 8.317899e-07, 1.321752e-05, 
    2.249467e-05, 1.975599e-05, 1.203892e-05, 7.244061e-06, 2.92921e-06,
  0.000128677, 0.0001022795, 9.077917e-05, 5.934937e-05, 5.489002e-05, 
    1.944578e-05, 1.563445e-06, 2.130957e-06, 1.836427e-05, 2.979056e-05, 
    3.031075e-05, 2.667093e-05, 1.345989e-05, 6.47422e-06, 1.292034e-06,
  0.0001290178, 0.0001229741, 0.0001341765, 9.172549e-05, 4.105925e-05, 
    2.722044e-05, 5.153155e-06, 9.609915e-06, 3.512936e-05, 3.595607e-05, 
    3.174924e-05, 2.492871e-05, 1.303361e-05, 4.748152e-06, 7.814834e-07,
  2.559307e-05, 2.728631e-05, 3.311188e-05, 3.034947e-05, 1.884367e-05, 
    1.16151e-05, 3.42736e-06, 2.513203e-06, 8.413723e-07, 3.661869e-07, 
    1.005979e-06, 4.036777e-06, 1.036414e-05, 2.17872e-05, 1.674461e-05,
  9.834846e-06, 5.552212e-06, 1.187164e-05, 2.013079e-05, 1.778634e-05, 
    1.468311e-05, 4.713514e-06, 2.059554e-06, 7.644458e-07, 2.269401e-06, 
    5.514391e-06, 8.68875e-06, 7.80112e-06, 1.319411e-05, 1.171709e-05,
  1.771981e-06, 1.153826e-06, 1.436563e-06, 3.625739e-06, 1.033595e-05, 
    1.355417e-05, 7.775137e-06, 4.650887e-06, 3.804928e-06, 5.482641e-06, 
    6.721606e-06, 8.708086e-06, 1.152602e-05, 1.147778e-05, 6.747787e-06,
  6.011597e-07, 6.573788e-07, 5.68915e-07, 1.824611e-06, 1.30183e-05, 
    1.462328e-05, 1.132017e-05, 5.785019e-06, 1.42222e-05, 1.45403e-05, 
    1.026687e-05, 1.373142e-05, 1.296302e-05, 8.127541e-06, 6.404855e-06,
  1.776849e-07, 3.068541e-07, 3.169845e-07, 4.021101e-07, 6.15295e-06, 
    1.331803e-05, 1.278003e-05, 6.073693e-06, 1.702524e-05, 2.292388e-05, 
    1.954615e-05, 1.433799e-05, 1.078786e-05, 1.245067e-05, 1.204131e-05,
  3.384535e-06, 8.391018e-07, 3.862181e-07, 1.829683e-06, 2.297328e-06, 
    1.128383e-05, 1.236482e-05, 1.274547e-05, 5.528872e-06, 1.268748e-05, 
    1.355029e-05, 1.044555e-05, 1.243104e-05, 1.394626e-05, 9.407192e-06,
  4.118318e-05, 1.810208e-05, 1.387659e-05, 1.125529e-05, 8.190094e-06, 
    7.546871e-06, 2.195104e-06, 1.620615e-06, 2.847813e-06, 4.175195e-06, 
    6.149213e-06, 6.379099e-06, 1.153172e-05, 1.42988e-05, 9.598495e-06,
  7.948343e-05, 6.758457e-05, 6.118661e-05, 4.356944e-05, 3.035117e-05, 
    1.519054e-05, 1.498776e-06, 2.320746e-07, 1.638241e-07, 4.820353e-07, 
    5.591314e-06, 6.614068e-06, 9.848791e-06, 1.321768e-05, 1.159052e-05,
  8.277925e-05, 7.814189e-05, 8.786395e-05, 8.875454e-05, 4.607904e-05, 
    1.224236e-05, 2.81245e-06, 7.67317e-08, 2.018817e-07, 2.187198e-06, 
    6.199599e-06, 7.252853e-06, 1.011689e-05, 1.658814e-05, 1.232329e-05,
  8.121724e-05, 7.837719e-05, 0.0001057458, 0.0001154256, 2.987551e-05, 
    2.330978e-05, 1.209313e-05, 1.172053e-06, 4.98933e-06, 7.851087e-06, 
    8.152846e-06, 9.692872e-06, 1.271953e-05, 1.464421e-05, 1.386117e-05,
  0.0001006221, 0.0001376197, 0.0001903951, 0.0002479115, 0.0002733829, 
    0.0002794374, 0.0002306229, 0.0001402859, 6.344575e-05, 3.150512e-05, 
    2.181221e-05, 2.265617e-05, 2.033812e-05, 1.68629e-05, 1.351364e-05,
  7.224547e-05, 0.0001050889, 0.0001508407, 0.0001977513, 0.0002423189, 
    0.0002973499, 0.0003080576, 0.0002124946, 9.711093e-05, 5.230651e-05, 
    2.7688e-05, 2.45116e-05, 1.830366e-05, 1.964996e-05, 1.416208e-05,
  3.9739e-05, 8.129383e-05, 0.0001200499, 0.0001611887, 0.0001700393, 
    0.0002124188, 0.0002677353, 0.0002313813, 0.0001222222, 6.117806e-05, 
    2.959512e-05, 1.72233e-05, 1.600259e-05, 4.921762e-06, 5.487385e-06,
  2.436866e-05, 5.555399e-05, 8.547887e-05, 0.0001184131, 0.0001102895, 
    7.280982e-05, 0.0001238361, 0.0001626801, 0.0001051581, 4.874068e-05, 
    1.639611e-05, 1.131696e-05, 2.177163e-06, 1.443707e-06, 3.774893e-06,
  1.26426e-05, 3.288621e-05, 6.161177e-05, 8.338687e-05, 7.599483e-05, 
    1.658189e-05, 1.998368e-05, 5.950893e-05, 5.338951e-05, 2.103199e-05, 
    1.115077e-05, 6.455788e-06, 4.670054e-06, 2.926109e-06, 3.863648e-06,
  6.556157e-06, 1.810061e-05, 4.199219e-05, 5.985547e-05, 6.60548e-05, 
    2.445894e-05, 8.370237e-06, 1.777501e-05, 2.43271e-05, 7.757914e-06, 
    7.690287e-07, 5.55555e-07, 1.323172e-06, 1.94115e-06, 1.724338e-06,
  1.403626e-05, 2.122345e-05, 3.475082e-05, 4.782206e-05, 4.179812e-05, 
    2.99789e-05, 1.800528e-05, 8.947057e-06, 1.044659e-05, 4.5756e-06, 
    7.383778e-07, 8.593126e-08, 2.946267e-07, 1.574189e-07, 5.826124e-07,
  1.861424e-05, 1.958908e-05, 2.763589e-05, 3.652727e-05, 2.415512e-05, 
    2.329628e-05, 2.213968e-05, 1.848335e-05, 1.221146e-05, 2.567966e-06, 
    1.224282e-06, 9.699497e-07, 2.514842e-07, 2.317163e-07, 5.378975e-07,
  2.154022e-05, 2.321155e-05, 2.675817e-05, 2.924944e-05, 1.911203e-05, 
    9.512954e-06, 1.02285e-05, 1.066404e-05, 9.061774e-06, 3.787647e-06, 
    3.240659e-06, 1.699586e-06, 2.445409e-07, 3.089163e-07, 1.162106e-06,
  2.427155e-05, 2.559785e-05, 2.98447e-05, 2.715364e-05, 1.319038e-05, 
    6.752466e-06, 4.064162e-06, 4.758646e-06, 5.298203e-06, 2.040185e-06, 
    4.182081e-06, 6.275752e-06, 1.943162e-06, 2.721858e-06, 4.467415e-06,
  0.000100668, 0.0001596486, 0.000185972, 0.0003204641, 0.0002716001, 
    0.0002324252, 0.0001589696, 0.0001069008, 8.229331e-05, 6.329013e-05, 
    7.549808e-05, 0.0002436861, 0.0002007228, 0.0001525193, 4.328826e-05,
  9.50194e-05, 0.0001625198, 0.000285749, 0.0004063529, 0.0004241893, 
    0.0004106208, 0.0002945306, 0.0001628765, 0.0001145948, 9.387059e-05, 
    0.0001457258, 0.0001933882, 0.0002095915, 0.00014381, 7.683691e-05,
  8.43052e-05, 0.0001771167, 0.000325392, 0.0004438033, 0.000519321, 
    0.0005599409, 0.000438011, 0.0002139096, 0.0001288145, 0.0001394905, 
    0.0001946075, 0.0002682952, 0.0002081959, 0.0001100673, 0.000126565,
  8.000684e-05, 0.0001752582, 0.0002952435, 0.0004055393, 0.0005623512, 
    0.000619596, 0.0005283316, 0.0002945398, 0.000155164, 0.0001849597, 
    0.000217978, 0.0002749257, 0.0002018526, 0.0001118487, 0.000110236,
  6.329209e-05, 0.0001528854, 0.0003351764, 0.0004094083, 0.0006260871, 
    0.0006368148, 0.0005972408, 0.0003334952, 0.0001940972, 0.0002615548, 
    0.0002356697, 0.0002467472, 0.0001723439, 0.0001220417, 0.0001205198,
  5.198934e-05, 0.0001592041, 0.0002996353, 0.0005130109, 0.0006533907, 
    0.0006542168, 0.000604048, 0.0003486207, 0.0002445508, 0.0002534449, 
    0.000240224, 0.0002204843, 0.0001623544, 0.0001245945, 0.0001167411,
  3.461926e-05, 0.0001080139, 0.000218668, 0.0004626076, 0.000599184, 
    0.0007340083, 0.0005682, 0.000316157, 0.0002916155, 0.0002848693, 
    0.000234099, 0.000189251, 0.0001670607, 0.0001278243, 9.460707e-05,
  2.045734e-05, 6.457461e-05, 0.0001737949, 0.0004029364, 0.0006127139, 
    0.0008302211, 0.0006382787, 0.0003863707, 0.0003538982, 0.0002897864, 
    0.0002029055, 0.0001600915, 0.0001673405, 0.0001215018, 6.875777e-05,
  1.519462e-05, 4.072416e-05, 0.0001332577, 0.000279977, 0.0006379863, 
    0.0008205582, 0.0008012531, 0.0005587447, 0.0002918079, 0.0002597681, 
    0.0001634681, 0.0001299628, 0.0001483957, 0.0001043196, 3.495261e-05,
  9.86646e-06, 2.40208e-05, 9.122359e-05, 0.0002776018, 0.0005969711, 
    0.0006601919, 0.00088184, 0.0008969121, 0.000556563, 0.0002830049, 
    0.0001224735, 9.66782e-05, 0.0001043032, 6.075683e-05, 1.281681e-05,
  1.16529e-05, 1.503091e-05, 2.421404e-05, 3.587454e-05, 2.071647e-05, 
    1.573355e-05, 1.069717e-05, 4.565798e-06, 4.259207e-06, 7.210302e-06, 
    8.161665e-06, 7.992542e-06, 2.920026e-06, 3.072992e-06, 1.798789e-06,
  7.925651e-06, 1.714125e-05, 1.230372e-05, 2.788909e-05, 4.088215e-05, 
    3.544312e-05, 1.84715e-05, 1.485187e-05, 1.105456e-05, 1.003774e-05, 
    9.504336e-06, 8.096506e-06, 2.3297e-06, 6.461734e-06, 3.352801e-06,
  2.488372e-06, 1.21187e-05, 1.7582e-05, 1.677396e-05, 4.221783e-05, 
    6.712991e-05, 5.001025e-05, 2.798428e-05, 2.373887e-05, 1.946287e-05, 
    1.534617e-05, 7.02807e-06, 4.423421e-06, 6.737743e-06, 3.561871e-06,
  2.470561e-06, 1.007211e-05, 1.926182e-05, 1.590467e-05, 3.109688e-05, 
    4.97654e-05, 3.753191e-05, 3.692424e-05, 3.025742e-05, 1.558102e-05, 
    1.275144e-05, 3.842961e-06, 1.590628e-06, 4.495841e-06, 1.426104e-06,
  3.149364e-06, 5.491622e-06, 2.527586e-05, 2.131279e-05, 3.51023e-05, 
    2.918973e-05, 2.535066e-05, 2.564233e-05, 2.95117e-05, 1.896128e-05, 
    8.160583e-06, 5.249184e-06, 1.009679e-06, 1.516333e-06, 1.338109e-06,
  1.84364e-05, 1.413926e-05, 1.403109e-05, 3.322591e-05, 5.205085e-05, 
    1.43351e-05, 1.688231e-05, 1.480565e-05, 1.287325e-05, 1.286167e-05, 
    6.522209e-06, 9.738784e-07, 3.392301e-07, 3.111225e-07, 1.321326e-06,
  2.306172e-05, 1.200854e-05, 1.67746e-05, 5.458252e-05, 5.107949e-05, 
    1.448074e-05, 1.451249e-06, 2.345897e-06, 2.646099e-06, 3.232183e-06, 
    5.007232e-06, 1.469655e-06, 2.394121e-07, 2.585993e-08, 1.533841e-05,
  9.776541e-06, 1.670197e-05, 1.509235e-05, 8.379888e-05, 2.058409e-05, 
    2.85209e-05, 1.937748e-05, 8.176731e-06, 2.323712e-06, 1.277764e-07, 
    3.150287e-06, 1.27214e-06, 1.419712e-07, 4.26567e-06, 3.687483e-05,
  7.007397e-06, 1.097185e-05, 1.549177e-05, 7.31273e-05, 8.738785e-05, 
    4.49407e-05, 2.867756e-05, 1.980988e-05, 1.728448e-05, 7.651312e-06, 
    4.714087e-06, 1.742839e-06, 2.788405e-06, 2.611678e-05, 6.299953e-05,
  7.109836e-06, 8.281448e-06, 1.149232e-05, 4.461708e-05, 9.1707e-05, 
    6.498162e-05, 3.245692e-05, 2.392173e-05, 4.66262e-05, 2.719196e-05, 
    1.052558e-05, 5.656557e-06, 2.234975e-05, 5.350054e-05, 6.991687e-05,
  3.400501e-06, 2.226081e-06, 6.985495e-06, 1.416431e-05, 1.028693e-05, 
    1.081681e-05, 1.136587e-05, 1.746937e-05, 4.545744e-05, 9.068378e-05, 
    0.0001378002, 0.0001657724, 0.0001571317, 0.0001132063, 5.675152e-05,
  3.21436e-06, 2.111644e-06, 2.808739e-06, 6.429843e-06, 1.263789e-05, 
    2.811272e-05, 2.776744e-05, 2.894722e-05, 5.110536e-05, 9.46307e-05, 
    0.0001217677, 0.0001432019, 0.0001308379, 6.794247e-05, 1.970387e-05,
  2.020804e-06, 1.471052e-06, 6.925928e-07, 1.165352e-06, 6.195565e-06, 
    3.199666e-05, 6.640179e-05, 0.0001099396, 0.0001525104, 0.0001312701, 
    0.0001147489, 0.0001234617, 0.0001082885, 4.114335e-05, 3.031807e-06,
  1.929701e-06, 9.377968e-07, 4.428099e-07, 8.481897e-07, 6.046258e-06, 
    2.10075e-05, 6.232151e-05, 0.000171865, 0.0002657879, 0.0002431595, 
    0.0001747367, 0.0001369184, 9.310458e-05, 2.416992e-05, 1.924848e-06,
  3.961761e-07, 3.454319e-07, 3.984969e-07, 6.904204e-08, 2.707354e-06, 
    1.144914e-05, 3.035649e-05, 7.618078e-05, 0.0001586798, 0.0001834522, 
    0.0001490088, 9.594663e-05, 6.097191e-05, 2.545937e-05, 2.808064e-06,
  1.865755e-06, 1.229391e-06, 2.115859e-07, 3.324985e-07, 4.444349e-06, 
    1.538982e-06, 6.906178e-06, 9.506242e-06, 2.600051e-05, 4.766043e-05, 
    4.449053e-05, 3.336063e-05, 2.726528e-05, 1.588886e-05, 4.577817e-06,
  3.358967e-06, 3.438182e-06, 2.947409e-06, 4.322796e-06, 4.117313e-06, 
    1.807373e-06, 2.675906e-07, 3.142902e-07, 4.048265e-07, 1.604374e-06, 
    9.861597e-06, 6.822675e-06, 3.152355e-06, 8.039973e-06, 4.625696e-06,
  8.515118e-06, 7.187954e-06, 1.099484e-05, 1.494382e-05, 7.871085e-06, 
    5.436389e-06, 1.518873e-06, 5.245005e-07, 1.258571e-08, 2.183144e-07, 
    4.301833e-07, 2.333386e-06, 1.038153e-06, 5.079929e-06, 1.29055e-06,
  8.559526e-06, 9.180398e-06, 1.819264e-05, 2.889614e-05, 7.650487e-06, 
    3.280994e-06, 2.138054e-07, 2.002368e-07, 1.076243e-06, 2.062273e-06, 
    5.53927e-06, 8.36958e-06, 6.520281e-06, 6.554232e-06, 1.937196e-06,
  1.230517e-05, 1.048426e-05, 1.708139e-05, 2.210517e-05, 2.50298e-06, 
    3.071651e-06, 5.96568e-07, 1.682314e-07, 2.308836e-06, 1.548426e-06, 
    5.834906e-06, 7.809402e-06, 7.578298e-06, 7.942565e-06, 3.878505e-06,
  6.177772e-06, 4.619433e-06, 6.99884e-06, 5.640024e-06, 3.75984e-06, 
    3.167349e-06, 6.956041e-06, 9.763527e-06, 1.384446e-05, 7.434652e-06, 
    1.167259e-05, 2.878338e-05, 4.928451e-05, 8.937596e-05, 0.0001043659,
  3.985437e-06, 2.085133e-06, 2.168792e-06, 2.323169e-06, 3.445492e-06, 
    1.111877e-05, 2.177086e-05, 2.486139e-05, 2.923255e-05, 2.178252e-05, 
    2.29869e-05, 3.407553e-05, 7.273688e-05, 0.0001319071, 0.0001395164,
  2.284333e-06, 1.417287e-06, 1.188679e-06, 2.990723e-06, 6.093057e-06, 
    1.776479e-05, 4.847994e-05, 7.043214e-05, 6.963025e-05, 4.362515e-05, 
    3.222343e-05, 4.014666e-05, 8.24499e-05, 0.000145012, 0.0001495707,
  2.20473e-06, 2.312871e-06, 1.319393e-06, 4.402011e-07, 2.711693e-06, 
    1.825277e-05, 6.678888e-05, 0.000106274, 0.0001054447, 7.738926e-05, 
    5.380999e-05, 6.29291e-05, 0.0001063758, 0.0001545059, 0.0001439899,
  2.137905e-06, 1.844202e-06, 1.733433e-06, 4.708351e-07, 1.535306e-06, 
    9.873424e-06, 6.304505e-05, 0.0001133746, 0.0001535132, 0.0001751332, 
    0.0001328988, 0.0001243784, 0.0001593849, 0.0001692244, 0.000131426,
  2.073905e-06, 1.717702e-06, 9.477935e-07, 1.562308e-06, 3.799527e-06, 
    5.437396e-06, 4.240733e-05, 7.494392e-05, 0.000149877, 0.0002160838, 
    0.0002155253, 0.0001879704, 0.0002058651, 0.0001753382, 0.0001213762,
  4.222047e-05, 9.70507e-06, 2.856239e-06, 3.610477e-06, 8.570463e-06, 
    2.236796e-06, 1.730766e-05, 3.671963e-05, 8.086926e-05, 0.0001873293, 
    0.0002096934, 0.0001817251, 0.0001779217, 0.000150827, 0.0001032185,
  5.422295e-05, 7.35721e-05, 4.51812e-05, 2.238049e-05, 1.249236e-05, 
    4.424017e-06, 1.483549e-05, 3.354127e-05, 7.693974e-05, 0.0001604586, 
    0.0001955082, 0.0001653966, 0.0001321642, 0.0001051226, 7.706625e-05,
  3.719287e-05, 9.7431e-05, 0.0001346703, 5.336387e-05, 3.073196e-05, 
    3.506173e-06, 1.00117e-05, 2.78122e-05, 0.0001213507, 0.0001656029, 
    0.0001800614, 0.0001525493, 0.0001188983, 8.272654e-05, 5.875901e-05,
  1.431405e-05, 4.543039e-05, 0.0001072637, 6.615013e-05, 7.970787e-06, 
    8.010079e-06, 6.519847e-06, 3.314681e-05, 0.0001197593, 0.0001597139, 
    0.0001589301, 0.0001439572, 0.0001083623, 8.355493e-05, 5.038958e-05,
  4.118653e-06, 4.608681e-06, 1.460327e-06, 1.329179e-07, 6.437287e-10, 
    5.867955e-09, 1.663733e-09, 8.876934e-10, 5.031966e-10, 1.984817e-10, 
    1.425138e-06, 1.589391e-05, 2.30417e-05, 2.000445e-05, 1.322496e-05,
  1.236148e-06, 6.258043e-07, 3.916168e-06, 4.916319e-07, 8.172795e-08, 
    1.826915e-07, 1.269165e-08, 4.431911e-09, 1.773911e-09, 2.437075e-09, 
    4.615546e-07, 1.428202e-05, 1.694027e-05, 1.939343e-05, 1.004703e-05,
  6.478911e-06, 2.35221e-06, 3.10138e-07, 3.967883e-06, 2.176423e-06, 
    3.527672e-07, 7.730145e-07, 5.324214e-07, 8.107106e-08, 3.621904e-07, 
    3.036918e-06, 1.102047e-05, 1.301872e-05, 9.354513e-06, 9.147007e-06,
  8.203049e-06, 4.108359e-06, 8.501284e-07, 9.299016e-06, 9.438593e-06, 
    4.085846e-06, 2.131612e-06, 6.695977e-07, 4.440995e-07, 6.661957e-07, 
    4.59523e-06, 7.116813e-06, 7.009703e-06, 4.21611e-06, 3.901173e-06,
  4.028825e-06, 2.055795e-06, 1.098982e-06, 4.641578e-06, 6.948022e-06, 
    9.486714e-06, 7.086363e-06, 2.402711e-06, 1.644825e-06, 1.668907e-06, 
    6.239565e-06, 3.240895e-06, 3.110964e-07, 4.222637e-06, 4.691175e-06,
  2.055449e-06, 1.907128e-06, 1.884254e-06, 4.099374e-06, 6.422951e-06, 
    8.978915e-07, 5.418312e-06, 6.919202e-06, 2.493111e-06, 5.819533e-07, 
    8.105144e-07, 1.377371e-06, 5.131091e-07, 4.549417e-07, 5.363632e-08,
  1.985378e-05, 5.404678e-06, 3.362544e-06, 7.51405e-06, 5.866954e-06, 
    1.368231e-07, 1.249967e-07, 2.414015e-08, 9.258922e-08, 3.148335e-07, 
    9.66382e-07, 9.941084e-07, 5.440289e-07, 4.66668e-07, 1.228318e-07,
  4.654053e-05, 5.564381e-05, 4.892268e-05, 9.795482e-06, 3.481726e-06, 
    1.989405e-07, 4.384819e-08, 2.64441e-08, 1.055247e-09, 1.184037e-08, 
    3.377787e-08, 1.83831e-07, 1.333583e-07, 3.056108e-09, 6.740275e-12,
  5.896587e-05, 6.392987e-05, 0.0001263754, 4.708789e-05, 3.002765e-05, 
    2.701783e-07, 4.489812e-09, 6.646086e-10, 6.548785e-11, 1.021963e-10, 
    2.73057e-11, 3.858873e-10, 3.194902e-10, 2.838346e-16, 0,
  4.252274e-05, 5.171029e-05, 0.0001403987, 8.977853e-05, 5.994761e-06, 
    5.802171e-07, 7.231496e-07, 8.006521e-09, 1.162078e-07, 1.953422e-08, 
    2.889728e-28, 1.155353e-08, 2.87746e-10, 2.564223e-15, 2.238604e-14,
  3.379502e-06, 2.235702e-05, 6.483584e-05, 0.0001266056, 0.0002387871, 
    0.0003107872, 0.0003309632, 0.0002606673, 0.000113937, 5.785934e-05, 
    5.697541e-05, 5.148596e-05, 3.863745e-05, 1.471579e-05, 5.145817e-06,
  2.356609e-06, 5.473986e-06, 3.734558e-05, 0.0001204955, 0.0001631589, 
    0.0002442859, 0.0003994335, 0.0003896047, 0.0003079351, 0.0001106824, 
    2.748074e-05, 2.781258e-05, 1.910875e-05, 9.210599e-06, 3.491094e-06,
  2.075845e-06, 2.642353e-06, 1.657007e-05, 0.0001033763, 0.0001250216, 
    0.0001537052, 0.0002961108, 0.0004106353, 0.0003167777, 9.525527e-05, 
    2.142236e-05, 1.847834e-05, 1.203668e-05, 5.841194e-06, 1.59468e-06,
  2.056215e-06, 1.970133e-06, 5.535126e-06, 3.597926e-05, 0.0001003374, 
    9.425855e-05, 0.0001261973, 0.0003305355, 0.0003044326, 9.137742e-05, 
    1.253066e-05, 8.668629e-07, 1.055447e-06, 4.776551e-07, 1.216394e-06,
  1.334451e-06, 1.352685e-06, 2.22857e-06, 9.392294e-06, 5.81063e-05, 
    4.448938e-05, 2.842127e-05, 0.0001578637, 0.0002385378, 0.0001039396, 
    6.980767e-06, 4.835171e-07, 6.029049e-08, 6.727965e-07, 4.069506e-07,
  8.850777e-07, 8.885787e-07, 1.147792e-06, 8.826632e-07, 2.591779e-05, 
    6.752535e-05, 1.751796e-05, 3.781947e-05, 0.0001320471, 7.008518e-05, 
    5.466507e-06, 4.535338e-07, 1.39788e-08, 6.099178e-07, 4.703416e-07,
  6.361392e-07, 6.583703e-07, 5.905648e-07, 1.081738e-06, 3.424433e-06, 
    5.110867e-05, 3.551864e-05, 7.617623e-06, 4.850772e-05, 3.551929e-05, 
    7.940133e-06, 3.414103e-07, 4.251345e-08, 5.460321e-07, 7.749688e-07,
  7.946835e-06, 1.559847e-06, 2.019569e-06, 2.447107e-06, 2.651337e-06, 
    2.565815e-05, 3.436625e-05, 9.212884e-06, 1.63462e-05, 2.017994e-05, 
    8.522207e-06, 9.848123e-07, 5.463188e-07, 6.035666e-07, 6.344715e-08,
  1.533279e-05, 6.358233e-06, 6.210732e-06, 3.71642e-06, 7.428745e-06, 
    8.277777e-06, 1.729994e-05, 3.01582e-06, 6.97741e-06, 1.093423e-05, 
    5.010268e-06, 4.982539e-07, 2.656719e-07, 1.877317e-08, 3.720981e-08,
  2.316281e-05, 1.292328e-05, 1.746301e-05, 9.293572e-06, 2.099965e-06, 
    2.533958e-06, 1.114978e-05, 3.557398e-06, 2.838479e-06, 4.877322e-06, 
    3.078529e-06, 7.880469e-07, 1.587324e-07, 5.526647e-08, 1.352894e-07,
  7.688255e-07, 1.090577e-06, 3.889626e-06, 1.884628e-05, 3.731665e-05, 
    2.579739e-05, 1.893185e-05, 2.031781e-05, 1.632933e-05, 1.058527e-05, 
    4.681878e-05, 5.455614e-05, 4.736773e-05, 5.223074e-05, 1.90193e-05,
  1.64114e-06, 1.099745e-06, 3.008315e-06, 2.034229e-05, 6.024128e-05, 
    6.721867e-05, 7.469946e-05, 6.694715e-05, 8.657831e-05, 6.114251e-05, 
    5.449213e-05, 5.514892e-05, 3.833595e-05, 3.833513e-05, 2.139093e-05,
  1.872009e-06, 1.186193e-06, 2.200524e-06, 1.530466e-05, 7.042111e-05, 
    0.0001110434, 0.0001389173, 0.0001517031, 0.0001464878, 8.451509e-05, 
    7.534189e-05, 6.716149e-05, 3.48412e-05, 3.769882e-05, 2.113179e-05,
  1.71484e-06, 1.292202e-06, 1.459699e-06, 6.808547e-06, 5.808799e-05, 
    0.0001234398, 0.0001534386, 0.000260044, 0.0002196429, 0.0001700536, 
    0.000105017, 7.477823e-05, 5.854606e-05, 4.607758e-05, 1.475837e-05,
  8.149102e-07, 1.052186e-06, 1.188896e-06, 2.411197e-06, 4.295884e-05, 
    8.605489e-05, 0.0001556997, 0.000323603, 0.0003355898, 0.0002462517, 
    7.18041e-05, 4.420647e-05, 4.923715e-05, 2.669112e-05, 2.764941e-05,
  3.01933e-07, 7.616669e-07, 1.061299e-06, 1.780316e-07, 2.982492e-05, 
    0.000101942, 0.0001099716, 0.0002132939, 0.000457057, 0.0003806778, 
    0.0001799902, 5.459222e-05, 6.578951e-05, 4.595848e-05, 2.181547e-05,
  1.167807e-05, 7.013974e-06, 3.295927e-06, 9.957463e-07, 1.967589e-05, 
    8.554694e-05, 0.0001482388, 0.0001179167, 0.0003231716, 0.0004307696, 
    0.0002632583, 8.732657e-05, 4.463188e-05, 4.966751e-05, 2.548285e-05,
  1.75062e-05, 1.023198e-05, 1.437921e-05, 5.899576e-06, 4.814243e-06, 
    6.351952e-05, 0.0001389809, 0.0001326248, 0.0002435446, 0.0004738081, 
    0.0003795589, 0.0001556756, 4.592538e-05, 3.92691e-05, 3.031729e-05,
  1.391112e-05, 1.259827e-05, 1.655287e-05, 1.376681e-05, 9.116502e-06, 
    2.492383e-05, 0.0001052455, 0.0001082301, 0.0002088569, 0.000448425, 
    0.0004339426, 0.0002449176, 7.154881e-05, 3.603899e-05, 3.270813e-05,
  1.773602e-05, 1.869822e-05, 1.748593e-05, 2.172717e-05, 5.396995e-06, 
    1.197542e-05, 6.611557e-05, 9.548375e-05, 0.0001547264, 0.0003371346, 
    0.0004398465, 0.0003283305, 0.0001374601, 3.667103e-05, 1.917907e-05,
  2.511627e-06, 2.485093e-06, 9.794328e-06, 1.866047e-05, 3.466286e-05, 
    7.955451e-05, 0.0001075897, 9.134632e-05, 5.6467e-05, 2.204571e-05, 
    1.496818e-05, 5.78482e-06, 4.646171e-06, 3.329643e-06, 8.958527e-07,
  4.244432e-07, 8.740309e-07, 3.300052e-06, 1.239622e-05, 1.558959e-05, 
    5.769339e-05, 9.576123e-05, 9.740709e-05, 9.589985e-05, 9.161362e-05, 
    4.204853e-05, 1.592738e-05, 6.299032e-06, 1.659879e-06, 1.048184e-06,
  2.962693e-07, 5.081558e-07, 1.202403e-06, 5.527062e-06, 7.67983e-06, 
    3.255108e-05, 7.537872e-05, 8.810844e-05, 0.0001060474, 0.000129224, 
    8.533239e-05, 2.70423e-05, 8.518417e-06, 2.993069e-06, 3.6766e-07,
  3.329748e-07, 3.425667e-07, 6.232584e-07, 2.300193e-06, 3.688657e-06, 
    1.500195e-05, 3.906382e-05, 6.182124e-05, 7.889236e-05, 0.0001136078, 
    0.0001095092, 4.795519e-05, 1.295006e-05, 5.60544e-06, 1.900913e-06,
  1.070649e-07, 1.96492e-07, 4.602838e-07, 9.859384e-07, 8.402061e-07, 
    3.535741e-06, 1.174025e-05, 2.58449e-05, 3.665423e-05, 6.206065e-05, 
    8.546812e-05, 5.355498e-05, 2.102863e-05, 6.042289e-06, 5.077376e-06,
  2.12998e-07, 1.281244e-07, 4.684447e-07, 6.103336e-07, 5.882565e-07, 
    9.652507e-07, 1.511404e-06, 6.427721e-06, 1.229585e-05, 1.656491e-05, 
    4.624112e-05, 3.788601e-05, 2.282253e-05, 7.728316e-06, 8.577812e-06,
  1.675374e-05, 8.214612e-06, 4.348101e-06, 7.325846e-07, 5.593069e-07, 
    3.199905e-06, 3.459923e-06, 3.132307e-06, 1.10742e-05, 1.271735e-05, 
    2.99371e-05, 3.137541e-05, 2.154366e-05, 1.30268e-05, 5.226865e-06,
  4.293755e-05, 3.022736e-05, 2.874742e-05, 5.333374e-06, 5.358704e-06, 
    2.025924e-06, 3.696732e-06, 4.488882e-06, 9.057263e-06, 1.03345e-05, 
    2.785404e-05, 3.491531e-05, 2.248402e-05, 1.24674e-05, 6.645404e-06,
  4.004575e-05, 4.582206e-05, 4.598443e-05, 2.927594e-05, 1.657025e-05, 
    1.625373e-06, 1.254912e-06, 2.527565e-07, 2.365866e-06, 1.67453e-05, 
    2.87415e-05, 3.884153e-05, 2.14616e-05, 1.303462e-05, 7.393957e-06,
  3.841832e-05, 5.072984e-05, 6.157967e-05, 5.428667e-05, 8.035856e-06, 
    5.166801e-06, 1.410947e-06, 8.804937e-08, 9.394128e-07, 1.138235e-05, 
    2.301587e-05, 3.438769e-05, 2.723146e-05, 1.211524e-05, 3.168235e-06,
  2.732377e-06, 8.769665e-07, 4.153497e-06, 4.802122e-06, 2.943562e-06, 
    3.646971e-06, 1.507787e-05, 5.321926e-05, 8.523683e-05, 7.012864e-05, 
    5.411057e-05, 6.322531e-05, 5.250525e-05, 1.817338e-05, 3.880737e-07,
  2.223931e-07, 5.143747e-07, 7.826587e-07, 1.207209e-06, 2.998005e-06, 
    1.096678e-06, 9.749128e-06, 3.692162e-05, 6.727657e-05, 8.155207e-05, 
    8.477999e-05, 7.468819e-05, 6.0602e-05, 1.796718e-05, 2.889854e-07,
  1.197033e-07, 2.932189e-07, 4.368007e-07, 6.820168e-07, 1.61559e-06, 
    5.038803e-07, 6.889129e-06, 3.244249e-05, 5.395693e-05, 8.357113e-05, 
    0.0001060579, 8.758288e-05, 5.944619e-05, 2.243185e-05, 7.644912e-07,
  4.999687e-08, 1.448236e-07, 2.1217e-07, 5.551457e-07, 8.90463e-07, 
    2.582829e-07, 5.24521e-06, 3.024164e-05, 5.349678e-05, 7.356353e-05, 
    0.0001042702, 9.933749e-05, 6.05809e-05, 2.317194e-05, 2.695423e-06,
  6.514528e-09, 3.550904e-08, 1.346703e-07, 3.951551e-07, 5.238663e-07, 
    5.339647e-08, 1.966777e-06, 1.172571e-05, 3.647846e-05, 5.539603e-05, 
    9.90074e-05, 0.0001080436, 5.96234e-05, 3.051584e-05, 6.268218e-06,
  8.124122e-07, 4.500608e-09, 5.106615e-08, 2.846702e-07, 3.045259e-07, 
    7.954474e-07, 1.201042e-07, 2.706375e-06, 2.117331e-05, 5.162718e-05, 
    8.369261e-05, 0.0001071894, 5.396235e-05, 3.438729e-05, 1.1939e-05,
  1.074398e-05, 8.015657e-06, 7.312335e-06, 5.779023e-06, 8.645151e-06, 
    1.03506e-06, 1.622477e-06, 3.901378e-06, 2.110444e-05, 4.900411e-05, 
    7.681768e-05, 0.0001211314, 7.455078e-05, 3.726695e-05, 1.38084e-05,
  2.770068e-05, 2.444695e-05, 2.401541e-05, 1.885531e-05, 9.244421e-06, 
    1.837643e-06, 1.800069e-06, 6.548723e-06, 2.379591e-05, 4.449316e-05, 
    8.658085e-05, 0.0001186092, 8.371623e-05, 3.816961e-05, 1.652028e-05,
  3.331561e-05, 3.596533e-05, 3.916126e-05, 4.092746e-05, 1.198751e-05, 
    1.776684e-06, 5.277465e-07, 5.826669e-08, 8.069812e-06, 6.040922e-05, 
    8.835705e-05, 0.0001172554, 9.445044e-05, 4.308041e-05, 1.911774e-05,
  3.269145e-05, 3.845129e-05, 4.678149e-05, 4.148904e-05, 4.437091e-06, 
    5.122014e-06, 4.530661e-07, 1.144236e-07, 4.978026e-06, 2.916521e-05, 
    6.742519e-05, 0.0001070778, 9.493472e-05, 5.094621e-05, 2.26286e-05,
  2.006221e-06, 2.564165e-06, 2.493549e-06, 5.585133e-06, 4.588626e-05, 
    0.0001197389, 0.0002223603, 0.0002573204, 0.0002011347, 0.0001671453, 
    0.000121627, 9.896096e-05, 8.702982e-05, 1.284349e-05, 4.667165e-07,
  1.322728e-06, 1.574999e-06, 3.165138e-06, 3.714676e-06, 2.024323e-05, 
    6.959086e-05, 0.0001797175, 0.000247366, 0.0001983376, 0.0002132611, 
    0.0002265612, 0.0002056279, 9.851246e-05, 1.113839e-05, 6.855988e-08,
  9.956816e-07, 1.277889e-06, 2.070029e-06, 7.856029e-07, 8.816834e-06, 
    3.758598e-05, 0.0001287539, 0.0002482476, 0.0001977745, 0.0002009867, 
    0.0003075721, 0.0001728092, 0.0001029203, 1.6446e-05, 2.561348e-07,
  8.348701e-07, 1.051425e-06, 1.564271e-06, 3.749187e-07, 2.167306e-06, 
    2.233717e-05, 8.663131e-05, 0.0002271447, 0.0002192053, 0.0001813158, 
    0.0002900904, 0.0002339044, 9.30526e-05, 1.688486e-05, 8.826269e-08,
  4.311612e-07, 5.25592e-07, 1.22874e-06, 4.142088e-07, 4.749657e-07, 
    2.957289e-06, 4.48701e-05, 0.0001805436, 0.0002280426, 0.0001656166, 
    0.0002541151, 0.0002257815, 7.821867e-05, 1.745094e-05, 1.173358e-06,
  1.983213e-07, 3.110901e-07, 7.611227e-07, 3.83852e-07, 2.941704e-07, 
    3.659996e-06, 2.058692e-05, 0.0001127806, 0.0002194059, 0.0001909753, 
    0.0002567804, 0.0002302732, 5.630292e-05, 1.451119e-05, 3.849612e-06,
  1.480745e-06, 1.143831e-06, 6.119615e-07, 4.277314e-07, 1.186496e-06, 
    6.598247e-06, 2.467638e-05, 7.639515e-05, 0.0001569646, 0.0002190566, 
    0.0002855995, 0.000237042, 7.221223e-05, 1.851893e-05, 5.057233e-06,
  1.163537e-05, 7.581693e-06, 7.789905e-06, 2.616435e-06, 3.400593e-08, 
    5.420854e-06, 2.257476e-05, 8.042112e-05, 0.0001634601, 0.0002149759, 
    0.0002998363, 0.000268254, 8.817372e-05, 2.317718e-05, 6.078569e-06,
  2.04272e-05, 2.113438e-05, 1.743911e-05, 9.750165e-06, 4.118728e-06, 
    3.428123e-06, 9.489559e-06, 1.003548e-05, 9.664301e-05, 0.0001891955, 
    0.0002834283, 0.0002658216, 0.0001022488, 2.274485e-05, 6.284605e-06,
  2.07957e-05, 2.809345e-05, 3.168044e-05, 2.188988e-05, 4.747119e-06, 
    3.288177e-06, 6.437503e-06, 5.286831e-06, 4.30816e-05, 0.000107212, 
    0.000241444, 0.0002864897, 0.0001265351, 3.579792e-05, 7.80998e-06,
  3.708802e-06, 2.372364e-06, 1.672959e-06, 1.885152e-06, 2.946167e-05, 
    0.0001100161, 0.000229841, 0.0002834913, 0.0002895715, 0.0001998837, 
    8.314045e-05, 8.591365e-05, 6.266088e-05, 3.450547e-05, 2.018263e-05,
  1.403783e-06, 1.077759e-06, 1.531275e-06, 7.654361e-07, 9.436518e-06, 
    8.026583e-05, 0.0001889452, 0.0002845468, 0.0002939761, 0.000220855, 
    0.000119556, 9.396443e-05, 0.0001020204, 3.99762e-05, 2.038401e-05,
  1.014409e-06, 7.656552e-07, 1.163249e-06, 1.391685e-06, 4.606134e-06, 
    4.281279e-05, 0.0001455734, 0.0002447142, 0.0002704378, 0.0002130122, 
    0.0001390269, 9.211947e-05, 9.639865e-05, 4.425695e-05, 2.640094e-05,
  8.18721e-07, 5.284041e-07, 1.089637e-06, 4.492923e-07, 6.164659e-07, 
    3.000732e-05, 0.00010424, 0.0002074923, 0.0002387739, 0.0001744872, 
    0.0001301942, 9.242498e-05, 9.086238e-05, 3.437962e-05, 2.765581e-05,
  5.786083e-07, 4.016648e-07, 1.243092e-06, 8.067141e-07, 5.237578e-07, 
    2.168548e-05, 8.37428e-05, 0.0001828438, 0.0002185869, 0.0001548735, 
    0.0001162023, 0.0001206457, 0.0001103983, 3.792485e-05, 1.852287e-05,
  3.178858e-06, 3.65781e-07, 1.025906e-06, 1.266898e-06, 3.490837e-06, 
    4.833073e-06, 4.776699e-05, 0.0001808706, 0.0002260348, 0.0001820879, 
    0.0001222299, 0.0001575405, 0.0002195492, 6.879932e-05, 2.044901e-05,
  3.456965e-05, 3.327455e-05, 2.306574e-05, 1.043517e-05, 1.504968e-05, 
    2.097321e-05, 8.019317e-05, 0.0001737011, 0.0002072385, 0.0002484877, 
    0.000170579, 0.0001748636, 0.0002171188, 0.0001417189, 4.224536e-05,
  3.992994e-05, 3.153911e-05, 3.211546e-05, 2.37549e-05, 1.361123e-05, 
    2.138038e-05, 0.000102234, 0.0002069245, 0.0002495713, 0.0002651241, 
    0.0002742911, 0.0002222064, 0.0002060068, 9.9221e-05, 6.193186e-05,
  4.550035e-05, 3.481135e-05, 2.931022e-05, 3.512182e-05, 2.041859e-05, 
    1.288933e-05, 5.684857e-05, 7.006856e-05, 0.0002531268, 0.0003048521, 
    0.0003331467, 0.000304739, 0.0002722903, 0.0001597218, 5.974308e-05,
  4.87163e-05, 4.178943e-05, 3.150327e-05, 3.660798e-05, 8.579619e-06, 
    1.537022e-05, 4.301985e-05, 6.190779e-05, 0.0002324839, 0.000275997, 
    0.0003282702, 0.0003776466, 0.0003647217, 0.0002576293, 9.920444e-05,
  2.095234e-05, 1.933375e-05, 3.282702e-05, 3.340316e-05, 2.723484e-05, 
    1.299304e-05, 4.908375e-06, 4.317522e-06, 1.059724e-05, 9.014428e-06, 
    2.231201e-05, 3.991266e-05, 5.469966e-05, 5.749058e-05, 5.98611e-05,
  5.083095e-06, 2.857145e-06, 1.092047e-05, 1.621387e-05, 2.584721e-05, 
    3.090229e-05, 1.377773e-05, 1.348533e-05, 1.367789e-05, 1.824028e-05, 
    3.261367e-05, 5.562169e-05, 7.04738e-05, 5.360051e-05, 4.593573e-05,
  1.336896e-07, 8.389251e-08, 1.807196e-07, 2.462911e-06, 2.201373e-05, 
    3.558133e-05, 3.667568e-05, 1.997229e-05, 2.963314e-05, 4.239141e-05, 
    5.89507e-05, 7.06534e-05, 7.267853e-05, 5.989466e-05, 4.31773e-05,
  7.725828e-10, 4.713849e-10, 6.784815e-10, 6.898981e-07, 1.243942e-05, 
    3.158192e-05, 4.631178e-05, 3.172778e-05, 4.361733e-05, 5.022905e-05, 
    6.628223e-05, 7.543188e-05, 7.60874e-05, 4.477302e-05, 4.797265e-05,
  6.194109e-10, 3.638886e-13, 6.940075e-27, 8.040789e-10, 4.381925e-06, 
    2.843642e-05, 4.684832e-05, 3.814499e-05, 4.633171e-05, 5.673382e-05, 
    6.206311e-05, 6.090626e-05, 5.623237e-05, 5.075704e-05, 5.050468e-05,
  2.980755e-06, 2.045658e-07, 3.105996e-09, 3.803396e-11, 2.146898e-06, 
    1.286183e-05, 3.458653e-05, 3.907351e-05, 4.740571e-05, 5.325971e-05, 
    5.518636e-05, 3.589213e-05, 3.884531e-05, 4.907402e-05, 4.607921e-05,
  2.990671e-05, 2.022827e-05, 2.084397e-05, 2.046067e-05, 2.997497e-05, 
    7.169375e-06, 1.069263e-06, 4.360133e-06, 1.940647e-05, 2.738896e-05, 
    3.84634e-05, 4.068858e-05, 4.403439e-05, 4.129382e-05, 4.202969e-05,
  6.348902e-05, 6.085313e-05, 6.41981e-05, 6.852285e-05, 6.750367e-05, 
    2.784958e-05, 5.266299e-06, 2.40238e-06, 5.195217e-07, 6.06579e-07, 
    1.499258e-05, 3.269378e-05, 3.602046e-05, 4.170957e-05, 4.561375e-05,
  5.741399e-05, 6.902166e-05, 7.399641e-05, 9.464892e-05, 7.6169e-05, 
    2.189351e-05, 1.947437e-05, 5.334881e-06, 8.428807e-06, 1.533606e-05, 
    3.098124e-05, 3.510189e-05, 3.729544e-05, 4.116453e-05, 4.054258e-05,
  5.615974e-05, 6.527992e-05, 7.165154e-05, 8.715159e-05, 3.646637e-05, 
    3.704369e-05, 2.098974e-05, 2.579839e-05, 3.478516e-05, 3.609096e-05, 
    3.434869e-05, 3.74181e-05, 4.439581e-05, 4.026953e-05, 3.854552e-05,
  2.181685e-06, 1.698521e-06, 2.774414e-06, 7.052423e-06, 2.655458e-06, 
    2.167103e-06, 9.374377e-06, 3.081878e-05, 5.52032e-05, 7.361249e-05, 
    6.449454e-05, 5.110994e-05, 3.958428e-05, 2.728444e-05, 1.992304e-05,
  5.367242e-07, 5.536338e-07, 7.006338e-07, 1.743534e-06, 1.862609e-06, 
    4.972013e-07, 1.669331e-06, 5.770865e-06, 2.700904e-05, 3.962078e-05, 
    5.284898e-05, 5.357966e-05, 4.113332e-05, 2.726199e-05, 1.335973e-05,
  3.069511e-07, 5.23531e-07, 4.811111e-07, 4.603577e-07, 1.933358e-06, 
    2.149579e-06, 1.070453e-06, 4.542683e-06, 1.034558e-05, 2.412886e-05, 
    5.150615e-05, 5.523254e-05, 2.758553e-05, 1.390377e-05, 4.202544e-06,
  7.987326e-08, 3.476331e-07, 4.278943e-07, 3.584294e-07, 4.987591e-07, 
    1.484897e-06, 1.584111e-06, 5.579014e-06, 1.298087e-05, 2.506483e-05, 
    3.618079e-05, 3.9075e-05, 2.560361e-05, 8.972109e-06, 6.079789e-06,
  1.384663e-08, 6.983392e-08, 2.202625e-07, 2.766464e-07, 2.857797e-07, 
    9.872265e-07, 2.588487e-06, 4.401286e-06, 1.067986e-05, 2.177965e-05, 
    2.170903e-05, 1.919821e-05, 2.163835e-05, 1.196433e-05, 1.010509e-05,
  1.130007e-06, 1.22495e-08, 4.162022e-08, 1.284165e-07, 2.023339e-07, 
    8.729205e-07, 2.456173e-06, 3.216413e-06, 1.695085e-06, 4.384342e-06, 
    7.424083e-06, 1.357542e-05, 1.476021e-05, 8.055706e-06, 4.378735e-06,
  2.156477e-06, 1.987313e-07, 1.398447e-08, 7.055143e-07, 1.801289e-06, 
    1.993104e-06, 5.278887e-07, 4.283739e-07, 1.010064e-06, 3.978075e-07, 
    2.724585e-06, 1.181896e-05, 5.227738e-06, 3.558735e-06, 3.103884e-06,
  1.79848e-05, 1.515013e-05, 1.299885e-05, 1.051459e-05, 8.678808e-06, 
    3.849596e-06, 1.383243e-06, 2.383635e-07, 1.031297e-07, 2.5161e-08, 
    1.695122e-08, 1.684908e-07, 8.086485e-07, 3.625226e-06, 2.872008e-06,
  2.756629e-05, 3.002762e-05, 3.095534e-05, 2.937184e-05, 2.995714e-05, 
    2.940764e-06, 9.038026e-07, 1.445343e-07, 1.412217e-07, 1.326212e-06, 
    1.011917e-06, 1.156393e-07, 5.028348e-07, 3.244944e-06, 2.756484e-06,
  3.339924e-05, 3.992247e-05, 4.292904e-05, 5.005924e-05, 1.377379e-05, 
    8.685682e-06, 9.681799e-06, 2.095584e-06, 7.244194e-06, 6.286746e-06, 
    5.356288e-06, 3.190074e-06, 1.365072e-06, 3.500349e-06, 1.40887e-06,
  5.558623e-05, 6.593363e-05, 9.302707e-05, 0.0001221568, 0.0001877574, 
    0.0002908547, 0.0004326394, 0.0005236684, 0.0004899654, 0.000286979, 
    0.0001364031, 9.110948e-05, 3.345512e-05, 1.398999e-05, 5.916565e-06,
  4.659839e-05, 4.759235e-05, 8.836266e-05, 9.676405e-05, 0.0001566213, 
    0.0002365995, 0.0004012288, 0.0005781351, 0.000576013, 0.0003874618, 
    0.0002399969, 9.996406e-05, 3.653772e-05, 1.628106e-05, 4.953667e-06,
  3.840165e-05, 5.319197e-05, 7.881343e-05, 8.602785e-05, 0.0001185074, 
    0.0001942674, 0.0003591401, 0.0005420356, 0.0007001603, 0.0007779583, 
    0.0003158634, 0.000131127, 3.413233e-05, 1.576682e-05, 8.719505e-06,
  3.006973e-05, 5.252353e-05, 6.780846e-05, 7.517554e-05, 8.823999e-05, 
    0.0001497674, 0.0002920679, 0.0004290423, 0.0005786005, 0.0006267718, 
    0.0003980857, 0.0001310053, 3.332721e-05, 1.228374e-05, 8.500954e-06,
  1.864479e-05, 3.97379e-05, 6.455935e-05, 4.973483e-05, 5.067634e-05, 
    0.0001027386, 0.0002619824, 0.0003754546, 0.0005016999, 0.0005959665, 
    0.0004289248, 0.000139946, 3.33542e-05, 1.497945e-05, 5.620137e-06,
  1.366534e-05, 3.49945e-05, 2.878177e-05, 2.667499e-05, 3.574865e-05, 
    7.556444e-05, 0.0001807483, 0.0003405518, 0.0003861151, 0.0004430086, 
    0.0002876459, 9.757514e-05, 2.431183e-05, 8.600618e-06, 1.971346e-06,
  5.92277e-06, 1.255925e-05, 9.289944e-06, 1.237731e-05, 1.001465e-05, 
    9.298411e-05, 0.0001212962, 0.000171149, 0.0003462321, 0.0003680948, 
    0.0002862177, 6.973454e-05, 1.803542e-05, 8.008867e-06, 3.249056e-06,
  3.10311e-06, 5.993683e-06, 3.298469e-06, 3.926472e-06, 9.666302e-06, 
    5.669692e-05, 0.0001410992, 0.0001859381, 0.0002263039, 0.0002757965, 
    0.0002076714, 6.077224e-05, 1.391815e-05, 1.057133e-05, 7.142407e-06,
  2.701875e-06, 4.528156e-06, 5.201915e-06, 1.550785e-06, 1.227124e-05, 
    3.003483e-05, 9.22372e-05, 0.000138844, 0.0001315428, 0.0001426939, 
    0.000128196, 4.360927e-05, 1.264152e-05, 8.023893e-06, 7.362245e-06,
  1.895145e-06, 4.181412e-06, 7.964911e-06, 6.210765e-06, 5.680628e-06, 
    1.122886e-05, 5.273402e-05, 9.544149e-05, 0.0001042775, 8.701123e-05, 
    5.537914e-05, 2.618487e-05, 1.03354e-05, 6.04567e-06, 8.012964e-06,
  9.891633e-06, 8.110485e-06, 1.476918e-05, 2.067319e-05, 2.559465e-05, 
    1.525445e-05, 1.18138e-05, 2.64209e-05, 5.037077e-05, 4.531828e-05, 
    4.875369e-05, 6.25048e-05, 7.090039e-05, 7.672572e-05, 5.756584e-05,
  1.115893e-05, 4.761403e-06, 1.589182e-05, 2.689765e-05, 3.424218e-05, 
    3.981257e-05, 3.442622e-05, 2.660299e-05, 4.139107e-05, 5.479985e-05, 
    5.720745e-05, 7.79007e-05, 9.54214e-05, 8.97978e-05, 7.018235e-05,
  1.305271e-05, 9.879844e-06, 1.816831e-05, 3.154603e-05, 5.134532e-05, 
    4.967527e-05, 4.499031e-05, 3.111029e-05, 3.965259e-05, 5.429724e-05, 
    7.720557e-05, 9.908532e-05, 0.0001106113, 9.736143e-05, 8.359752e-05,
  1.900202e-05, 2.37562e-05, 2.391048e-05, 4.31954e-05, 5.987449e-05, 
    5.374082e-05, 4.377469e-05, 2.545408e-05, 2.683792e-05, 5.462688e-05, 
    0.0001326925, 0.0001302217, 0.0001079641, 8.326738e-05, 7.624168e-05,
  1.702067e-05, 3.244346e-05, 4.268263e-05, 5.481858e-05, 8.327152e-05, 
    6.620284e-05, 4.841164e-05, 2.901819e-05, 2.334846e-05, 4.76286e-05, 
    0.0001110064, 0.0001987036, 0.0001117011, 0.0001016828, 9.615353e-05,
  5.412856e-05, 5.296019e-05, 4.201268e-05, 6.178863e-05, 0.0001182585, 
    6.50825e-05, 3.971243e-05, 4.772509e-05, 4.678029e-05, 7.456674e-05, 
    9.995479e-05, 0.0001363155, 0.0001236942, 8.789767e-05, 7.832042e-05,
  5.183527e-05, 5.18862e-05, 4.345535e-05, 6.742604e-05, 0.0001416466, 
    0.0001009901, 3.44457e-05, 7.433444e-05, 0.0001187423, 0.0001565279, 
    0.0001662696, 0.0001412453, 0.0001134428, 9.012588e-05, 8.664733e-05,
  2.227049e-05, 4.131576e-05, 5.123717e-05, 6.230902e-05, 0.0001059271, 
    0.0001498373, 0.000165095, 0.0001872081, 0.0002514005, 0.0002875233, 
    0.0002582478, 0.0001235804, 7.348912e-05, 7.785171e-05, 8.873662e-05,
  2.00075e-05, 3.348645e-05, 5.188549e-05, 3.89206e-05, 0.0001059183, 
    0.0001803646, 0.0001608188, 0.0002665094, 0.0002965464, 0.0004015022, 
    0.0003950195, 0.0001720399, 5.957189e-05, 5.807673e-05, 7.137842e-05,
  1.526994e-05, 2.424659e-05, 4.323476e-05, 4.917179e-05, 9.849274e-05, 
    0.0001406338, 0.0001478562, 0.0002472821, 0.0002470034, 0.0004153432, 
    0.0004823992, 0.0002507663, 5.852007e-05, 4.266664e-05, 5.951298e-05,
  8.512065e-06, 4.987527e-06, 7.800731e-06, 1.060299e-05, 1.331625e-05, 
    9.254363e-06, 1.041887e-05, 1.078052e-05, 1.466639e-05, 1.410993e-05, 
    2.072214e-05, 3.654648e-05, 4.420838e-05, 2.602853e-05, 2.463824e-05,
  1.550913e-06, 8.843617e-07, 5.420745e-06, 6.250022e-06, 1.140608e-05, 
    2.676535e-05, 2.619675e-05, 1.889507e-05, 2.02461e-05, 2.141672e-05, 
    3.324538e-05, 6.112816e-05, 5.966998e-05, 3.346913e-05, 2.70028e-05,
  3.630696e-07, 1.379137e-07, 2.879516e-07, 2.560855e-06, 1.021144e-05, 
    2.047796e-05, 3.021603e-05, 3.458448e-05, 3.931484e-05, 4.044898e-05, 
    4.989066e-05, 6.855933e-05, 6.557763e-05, 3.421942e-05, 2.881637e-05,
  1.174562e-06, 2.251317e-07, 3.144603e-08, 4.28095e-06, 7.945035e-06, 
    1.528968e-05, 3.223001e-05, 4.537238e-05, 4.329479e-05, 4.72388e-05, 
    5.641866e-05, 6.492508e-05, 6.365902e-05, 2.848162e-05, 2.990334e-05,
  4.765599e-07, 1.779919e-07, 2.678248e-07, 1.9472e-06, 4.619275e-06, 
    1.228036e-05, 3.549224e-05, 5.059858e-05, 4.903935e-05, 5.510663e-05, 
    6.711065e-05, 6.997499e-05, 6.300733e-05, 3.334584e-05, 3.954825e-05,
  7.18973e-07, 2.247534e-07, 4.794475e-08, 4.057822e-07, 3.457246e-06, 
    6.852295e-06, 2.726691e-05, 3.779105e-05, 4.243185e-05, 4.916647e-05, 
    5.742996e-05, 6.309627e-05, 5.978409e-05, 4.441146e-05, 5.726404e-05,
  9.408039e-06, 7.271884e-06, 5.426148e-06, 6.96444e-06, 9.377723e-06, 
    6.847324e-06, 5.377276e-06, 3.645345e-06, 8.122088e-06, 2.041725e-05, 
    3.184367e-05, 4.803546e-05, 5.619519e-05, 5.251973e-05, 7.925495e-05,
  2.644765e-05, 2.529617e-05, 2.22385e-05, 2.263259e-05, 1.877462e-05, 
    1.090722e-05, 6.303528e-06, 6.989013e-07, 5.58113e-08, 3.892803e-08, 
    9.205737e-06, 3.292611e-05, 5.003568e-05, 6.258426e-05, 9.901365e-05,
  3.676386e-05, 3.188637e-05, 2.948557e-05, 2.73883e-05, 3.027177e-05, 
    6.359756e-06, 3.709212e-06, 1.415753e-06, 1.43877e-06, 3.142032e-06, 
    1.195046e-05, 2.993166e-05, 5.483456e-05, 7.86817e-05, 0.0001146398,
  4.034704e-05, 4.264397e-05, 3.161607e-05, 3.394166e-05, 5.67984e-06, 
    5.749412e-06, 3.99609e-06, 6.71504e-06, 2.199271e-05, 1.670752e-05, 
    1.495535e-05, 2.952894e-05, 7.249325e-05, 9.762361e-05, 0.0001354235,
  1.884782e-05, 1.460508e-05, 1.439684e-05, 1.568539e-05, 5.92472e-06, 
    3.806404e-07, 1.576685e-06, 1.049228e-07, 5.66519e-07, 2.055181e-07, 
    2.991964e-07, 1.373651e-05, 2.152298e-05, 1.848058e-05, 6.350275e-06,
  1.327586e-05, 6.317132e-06, 1.471161e-05, 1.061143e-05, 1.288384e-05, 
    6.837274e-06, 3.605394e-06, 2.910592e-06, 3.490714e-06, 1.355099e-07, 
    2.328484e-06, 2.10199e-05, 2.303282e-05, 1.372859e-05, 4.613081e-06,
  9.48936e-06, 5.160254e-06, 3.86019e-06, 9.448658e-06, 1.643483e-05, 
    1.272996e-05, 1.050013e-05, 6.538543e-06, 7.402145e-06, 4.584026e-06, 
    8.526336e-06, 1.515534e-05, 1.526292e-05, 7.575899e-06, 6.126653e-07,
  1.324587e-05, 3.681837e-06, 1.43968e-06, 1.508623e-05, 1.9974e-05, 
    1.939941e-05, 2.17431e-05, 1.904493e-05, 1.404313e-05, 8.838111e-06, 
    3.889254e-06, 1.513081e-05, 8.49068e-06, 2.993258e-07, 1.701703e-07,
  2.269104e-06, 6.994923e-07, 1.62158e-06, 9.62528e-06, 1.788735e-05, 
    2.482784e-05, 2.849672e-05, 3.216351e-05, 2.633951e-05, 1.576756e-05, 
    1.336754e-05, 7.761584e-06, 4.118362e-06, 1.131243e-06, 2.550848e-07,
  1.345823e-05, 7.801007e-06, 4.932698e-06, 9.643548e-06, 1.285775e-05, 
    1.304993e-05, 3.221868e-05, 4.083582e-05, 3.477206e-05, 2.674249e-05, 
    1.304877e-05, 7.352181e-06, 1.840771e-06, 1.330659e-06, 5.963195e-07,
  2.191744e-05, 1.49737e-05, 1.282718e-05, 1.061815e-05, 1.589809e-05, 
    5.625463e-06, 1.227705e-06, 5.41286e-06, 1.511189e-05, 2.032441e-05, 
    1.387775e-05, 7.74662e-06, 2.861676e-06, 1.05771e-06, 7.077632e-07,
  5.687706e-05, 3.662978e-05, 3.218247e-05, 1.86541e-05, 1.786056e-05, 
    1.188173e-05, 4.459868e-06, 2.732541e-06, 3.314116e-07, 4.414358e-06, 
    1.062413e-05, 7.645946e-06, 4.188981e-06, 2.026967e-06, 1.198682e-06,
  7.403351e-05, 6.517173e-05, 6.277156e-05, 3.728874e-05, 5.059341e-05, 
    1.529576e-05, 9.160586e-06, 4.242309e-06, 7.205894e-06, 1.130151e-05, 
    8.747334e-06, 7.09428e-06, 4.260084e-06, 2.568841e-06, 1.844266e-06,
  7.664014e-05, 7.084844e-05, 7.217161e-05, 6.058796e-05, 1.359482e-05, 
    1.718958e-05, 5.807014e-06, 9.801827e-06, 1.834763e-05, 1.382066e-05, 
    7.930178e-06, 5.394333e-06, 3.749949e-06, 3.273763e-06, 1.950259e-06,
  1.829231e-05, 1.64352e-05, 1.624974e-05, 1.31972e-05, 4.684316e-06, 
    1.038227e-06, 3.984176e-09, 1.655997e-08, 8.060572e-08, 2.767521e-07, 
    2.590835e-07, 2.135351e-06, 3.686023e-05, 7.812821e-05, 5.222491e-05,
  1.059196e-05, 6.210212e-06, 1.407281e-05, 1.007673e-05, 6.733148e-06, 
    2.033435e-06, 2.306172e-07, 3.505435e-07, 1.356857e-07, 2.204071e-07, 
    6.222966e-07, 5.941333e-06, 3.000336e-05, 5.399131e-05, 4.265826e-05,
  7.220421e-06, 4.093957e-06, 4.115918e-06, 8.714856e-06, 1.16851e-05, 
    6.070201e-06, 6.694514e-06, 4.16932e-06, 1.017771e-06, 2.082792e-06, 
    9.271575e-06, 1.160525e-05, 2.066656e-05, 2.77755e-05, 2.564964e-05,
  6.026492e-06, 2.023234e-06, 1.004048e-06, 1.098663e-05, 1.358476e-05, 
    5.978242e-06, 4.587508e-06, 5.055467e-06, 5.298404e-06, 1.6528e-05, 
    1.733438e-05, 1.275753e-05, 1.273205e-05, 1.453476e-05, 1.774675e-05,
  8.09028e-07, 4.480639e-07, 5.814226e-07, 8.636236e-06, 1.495428e-05, 
    1.530888e-05, 1.077011e-05, 1.740692e-05, 1.117545e-05, 2.521983e-05, 
    2.807771e-05, 1.627514e-05, 1.224686e-05, 1.429641e-05, 1.361706e-05,
  1.714553e-08, 1.347134e-08, 1.792352e-07, 6.466047e-06, 1.618337e-05, 
    1.77434e-05, 1.398696e-05, 1.427468e-05, 2.52904e-05, 3.913486e-05, 
    4.028326e-05, 2.086945e-05, 1.129519e-05, 1.132536e-05, 1.121896e-05,
  1.124827e-06, 1.947418e-06, 9.282758e-06, 2.288102e-05, 3.61424e-05, 
    9.616287e-06, 4.666517e-06, 5.637024e-06, 9.650223e-06, 1.995303e-05, 
    4.090575e-05, 2.492851e-05, 1.5159e-05, 9.705765e-06, 8.638852e-06,
  5.787253e-05, 5.375983e-05, 4.945316e-05, 4.554784e-05, 3.49855e-05, 
    1.147057e-05, 2.859692e-06, 7.872006e-07, 8.741569e-07, 5.554218e-07, 
    8.27961e-06, 3.368839e-05, 1.976816e-05, 9.982079e-06, 9.034211e-06,
  7.767176e-05, 7.510817e-05, 7.093091e-05, 6.24579e-05, 4.469655e-05, 
    9.392164e-06, 3.693381e-06, 2.83366e-07, 1.19775e-07, 1.937151e-06, 
    7.711492e-06, 2.462523e-05, 1.926506e-05, 1.202153e-05, 9.438766e-06,
  6.733874e-05, 7.864086e-05, 8.061255e-05, 8.22867e-05, 1.300611e-05, 
    7.831364e-06, 3.136624e-06, 3.471451e-06, 1.407449e-06, 7.681468e-06, 
    7.064808e-06, 1.643343e-05, 2.486687e-05, 1.544348e-05, 9.978346e-06,
  1.598559e-05, 1.861608e-05, 1.54783e-05, 1.720292e-05, 2.232222e-05, 
    2.878971e-05, 3.260216e-05, 4.793732e-05, 6.848753e-05, 7.097435e-05, 
    4.182843e-05, 3.209843e-05, 4.549216e-05, 3.076046e-05, 1.3108e-05,
  9.822299e-06, 8.051143e-06, 9.142053e-06, 8.276952e-06, 1.825228e-05, 
    2.183712e-05, 2.779075e-05, 3.855187e-05, 5.4625e-05, 6.447441e-05, 
    5.05723e-05, 3.327473e-05, 2.775637e-05, 1.88712e-05, 7.325976e-06,
  6.946083e-06, 4.929891e-06, 7.712957e-06, 5.160023e-06, 9.521357e-06, 
    1.764672e-05, 2.593228e-05, 3.652057e-05, 4.856769e-05, 5.782599e-05, 
    5.16101e-05, 2.483767e-05, 6.168328e-06, 4.205458e-06, 7.310267e-06,
  5.734909e-06, 4.211097e-06, 5.668423e-06, 5.059094e-06, 3.538164e-06, 
    6.644294e-06, 1.368505e-05, 2.413007e-05, 3.869494e-05, 4.507152e-05, 
    3.901424e-05, 2.060586e-05, 2.09362e-06, 8.779478e-07, 3.118852e-06,
  3.710006e-06, 3.301917e-06, 3.467338e-06, 2.675087e-06, 2.262613e-06, 
    1.943395e-06, 2.693455e-06, 5.057581e-06, 1.501398e-05, 3.161924e-05, 
    2.841364e-05, 1.561963e-05, 2.676458e-06, 1.150557e-06, 1.50849e-06,
  2.23466e-06, 2.321069e-06, 2.367242e-06, 1.693033e-06, 1.156086e-06, 
    2.807047e-06, 3.856259e-07, 5.309404e-07, 1.72995e-06, 1.238831e-05, 
    1.024776e-05, 3.404548e-06, 6.983068e-06, 1.214935e-06, 1.240768e-06,
  1.486315e-06, 1.658145e-06, 1.999084e-06, 2.309145e-07, 1.477256e-06, 
    3.699157e-06, 1.672176e-06, 1.06717e-06, 2.47316e-07, 8.029195e-07, 
    7.895303e-06, 5.026289e-06, 6.548782e-06, 2.358771e-06, 1.205868e-06,
  1.143116e-05, 6.630245e-06, 5.764426e-06, 2.653504e-06, 2.575192e-06, 
    3.90956e-06, 1.919052e-06, 1.086513e-06, 7.265108e-07, 8.36633e-08, 
    5.572906e-07, 7.091179e-06, 6.80266e-06, 5.490554e-06, 4.868227e-06,
  1.808695e-05, 1.932092e-05, 2.058668e-05, 1.146918e-05, 1.586547e-05, 
    2.227557e-06, 1.031903e-06, 7.895425e-08, 1.029319e-07, 3.626359e-07, 
    1.545252e-07, 4.833691e-06, 7.007096e-06, 5.320344e-06, 5.065246e-06,
  2.125059e-05, 2.381861e-05, 2.498345e-05, 2.745976e-05, 8.749402e-06, 
    2.284845e-06, 1.817494e-06, 2.25545e-07, 6.408543e-08, 5.815989e-08, 
    2.294282e-06, 1.949227e-06, 7.941276e-06, 4.840299e-06, 5.099268e-06,
  1.340745e-05, 1.117725e-05, 1.420895e-05, 8.928035e-06, 6.288084e-06, 
    5.917789e-06, 7.075377e-06, 1.208931e-05, 3.245697e-05, 4.504793e-05, 
    8.259408e-05, 0.0001353013, 0.000161087, 9.621254e-05, 5.269471e-05,
  6.88996e-06, 4.596689e-06, 1.222839e-05, 1.407452e-05, 1.693484e-05, 
    1.948774e-05, 1.673481e-05, 1.379872e-05, 3.063982e-05, 6.475437e-05, 
    0.0001224837, 0.0001320465, 0.0001416274, 0.0001084785, 6.935617e-05,
  8.001958e-06, 3.302109e-06, 4.253516e-06, 1.615215e-05, 3.349363e-05, 
    4.477555e-05, 4.065671e-05, 3.440368e-05, 5.600429e-05, 9.484342e-05, 
    0.0001635951, 0.0001678599, 0.000153113, 0.0001154799, 8.12527e-05,
  5.500534e-06, 2.774514e-06, 6.069942e-06, 2.028671e-05, 5.649369e-05, 
    7.283185e-05, 8.003585e-05, 6.619e-05, 8.919272e-05, 0.0001280708, 
    0.0001818161, 0.0001974475, 0.0001737989, 0.0001213413, 7.835195e-05,
  3.859039e-06, 2.725604e-06, 7.21067e-06, 2.063872e-05, 5.449106e-05, 
    7.183802e-05, 8.783802e-05, 8.317043e-05, 0.0001036644, 0.0001380852, 
    0.0001742004, 0.0001893414, 0.000156569, 0.0001137733, 7.154381e-05,
  6.435288e-06, 4.446179e-06, 5.204764e-06, 2.239854e-05, 2.294498e-05, 
    1.247347e-05, 3.653087e-05, 6.874005e-05, 0.0001075621, 0.0001425002, 
    0.0001658827, 0.0001570395, 0.0001476719, 0.0001001877, 6.524631e-05,
  3.742775e-06, 4.099861e-06, 7.878571e-06, 1.769884e-05, 2.138479e-05, 
    6.758834e-06, 4.518167e-06, 1.473521e-05, 5.318803e-05, 0.0001191762, 
    0.0001525349, 0.0001498258, 0.0001298791, 9.387924e-05, 6.458646e-05,
  1.264387e-05, 1.272909e-05, 1.274285e-05, 1.752873e-05, 3.625902e-05, 
    7.026333e-06, 5.175551e-06, 1.995834e-05, 3.786233e-05, 9.593036e-05, 
    0.0001582942, 0.0001473424, 0.000118053, 8.839203e-05, 5.5772e-05,
  2.298276e-05, 1.800952e-05, 1.828646e-05, 2.674216e-05, 4.716196e-05, 
    5.693182e-06, 3.988137e-07, 5.156741e-07, 5.08408e-05, 0.0001196675, 
    0.000167137, 0.000163326, 0.0001209885, 7.764824e-05, 4.934573e-05,
  2.72107e-05, 2.307539e-05, 2.566643e-05, 3.416544e-05, 1.203746e-05, 
    6.106143e-06, 4.174879e-06, 2.61525e-06, 4.328795e-05, 9.594714e-05, 
    0.0001613963, 0.0001633887, 0.0001375844, 7.365461e-05, 4.267833e-05,
  1.741306e-11, 6.004573e-11, 7.731652e-11, 7.560013e-12, 3.724018e-09, 
    1.14923e-09, 7.276334e-09, 2.93671e-09, 1.054161e-09, 3.935588e-11, 
    1.91353e-10, 2.378981e-09, 3.056096e-06, 4.687848e-06, 6.46368e-06,
  3.635173e-12, 3.613505e-12, 2.360617e-12, 2.925473e-10, 4.757145e-08, 
    3.048169e-09, 1.956308e-09, 4.410621e-09, 2.104027e-09, 1.554593e-09, 
    2.291569e-09, 4.623489e-07, 7.142703e-06, 1.111419e-05, 4.830401e-06,
  2.423128e-11, 1.105821e-17, 8.43695e-27, 4.356327e-08, 1.303891e-07, 
    1.310474e-07, 1.105541e-07, 5.36806e-08, 1.923424e-08, 4.238455e-07, 
    7.11978e-07, 1.299643e-06, 3.762e-06, 5.1077e-06, 2.853774e-06,
  2.824409e-11, 2.071131e-26, 9.319699e-28, 5.376418e-09, 6.806768e-08, 
    8.565847e-07, 2.974865e-06, 3.738185e-06, 2.345254e-06, 1.604508e-06, 
    6.319618e-07, 1.751516e-06, 2.812571e-06, 2.129303e-06, 1.936936e-06,
  7.748666e-09, 5.291088e-11, 3.564e-27, 9.17541e-10, 1.633928e-08, 
    8.764461e-07, 7.105036e-06, 7.50858e-06, 8.000894e-06, 7.39127e-06, 
    5.751413e-06, 4.463588e-06, 2.853702e-06, 2.183164e-06, 1.532861e-06,
  3.308293e-09, 2.621925e-11, 1.136736e-27, 8.063453e-08, 8.209417e-08, 
    3.352555e-07, 3.981996e-06, 9.157473e-06, 1.131467e-05, 9.965954e-06, 
    8.17458e-06, 4.885791e-06, 2.522944e-06, 1.774914e-06, 1.418991e-06,
  4.152238e-08, 8.196382e-08, 1.325703e-07, 4.156895e-08, 4.775333e-07, 
    5.497648e-09, 3.366318e-08, 2.386988e-08, 1.596677e-06, 6.65516e-06, 
    1.024754e-05, 8.056868e-06, 5.092887e-06, 2.154693e-06, 9.776029e-07,
  7.489488e-06, 2.140206e-06, 1.308646e-06, 9.040336e-07, 6.615773e-07, 
    2.060089e-07, 1.395094e-07, 4.518411e-07, 6.788348e-09, 6.52848e-09, 
    4.539449e-06, 9.916538e-06, 8.84258e-06, 3.690165e-06, 1.523063e-06,
  2.584145e-05, 7.116714e-06, 4.352023e-06, 4.627929e-06, 6.770549e-06, 
    4.820254e-07, 6.730377e-09, 8.783131e-09, 1.422034e-07, 6.587373e-07, 
    5.274681e-06, 6.284741e-06, 8.643243e-06, 7.734808e-06, 2.902265e-06,
  3.372067e-05, 1.843708e-05, 1.439079e-05, 1.280194e-05, 5.010035e-06, 
    1.088029e-06, 7.552482e-07, 8.822341e-07, 1.205773e-06, 3.295856e-06, 
    5.094013e-06, 9.230815e-06, 9.543426e-06, 8.902077e-06, 5.032937e-06,
  1.387806e-07, 8.013887e-08, 3.108669e-07, 1.552436e-07, 6.531456e-08, 
    1.125612e-06, 1.125033e-05, 6.497453e-05, 0.0001408671, 0.0001352346, 
    0.0001129187, 7.133593e-05, 3.556838e-05, 6.341626e-06, 1.425821e-06,
  2.261853e-07, 1.107602e-07, 5.77195e-08, 3.09025e-07, 3.311506e-07, 
    6.959116e-08, 5.966117e-06, 2.637623e-05, 0.0001217929, 0.0001360264, 
    8.429876e-05, 3.894761e-05, 2.258421e-05, 4.441573e-06, 2.190925e-06,
  7.195242e-07, 1.809407e-07, 6.344287e-08, 1.272791e-07, 1.086599e-06, 
    4.831637e-06, 7.110077e-06, 2.804833e-05, 8.926092e-05, 0.0001185212, 
    8.855145e-05, 3.235274e-05, 8.262919e-06, 3.354591e-06, 1.318029e-06,
  1.712433e-06, 3.435653e-07, 8.539934e-08, 4.230856e-08, 8.066488e-07, 
    4.78898e-06, 5.48216e-06, 1.502858e-05, 5.501895e-05, 0.0001088036, 
    7.01486e-05, 2.241045e-05, 4.945575e-06, 1.00898e-06, 9.730142e-07,
  9.157962e-07, 3.424733e-07, 9.83808e-08, 3.669113e-08, 3.364401e-07, 
    9.515474e-07, 6.189243e-06, 1.601269e-05, 4.832894e-05, 8.328725e-05, 
    5.437034e-05, 8.668419e-06, 3.091052e-06, 3.140321e-07, 6.45414e-07,
  2.892021e-07, 2.323043e-07, 6.915322e-08, 2.151342e-08, 1.386471e-07, 
    3.509636e-07, 2.066626e-06, 1.585478e-05, 5.789642e-05, 9.708772e-05, 
    3.991535e-05, 3.331461e-06, 1.626977e-06, 6.693484e-07, 1.883469e-07,
  5.102474e-08, 2.44836e-07, 1.594547e-07, 5.303197e-07, 5.7241e-07, 
    1.176801e-07, 1.30031e-07, 3.627035e-06, 4.32569e-05, 0.0001110841, 
    4.048304e-05, 3.733833e-06, 1.629654e-06, 6.326383e-07, 6.392649e-10,
  1.053337e-07, 6.202606e-07, 7.000336e-07, 2.153576e-06, 1.04845e-06, 
    1.968451e-07, 4.834044e-08, 1.449948e-06, 1.520083e-05, 6.096817e-05, 
    3.298643e-05, 3.252574e-06, 1.083433e-06, 3.107252e-07, 5.098378e-10,
  3.077835e-06, 1.619996e-06, 1.101559e-05, 7.27049e-06, 1.021587e-05, 
    5.298756e-08, 1.330239e-08, 1.393878e-08, 2.11702e-05, 8.528192e-05, 
    3.655122e-05, 4.988709e-06, 4.478042e-07, 3.829148e-08, 2.033482e-11,
  1.032108e-05, 7.643011e-06, 9.104472e-06, 1.37944e-05, 1.298845e-06, 
    3.664008e-08, 8.754792e-09, 1.132768e-06, 3.985133e-05, 7.856503e-05, 
    3.792781e-05, 6.662357e-06, 5.833026e-08, 5.321718e-09, 4.523474e-12,
  1.426285e-05, 1.697669e-05, 2.24763e-05, 3.388929e-05, 5.467044e-05, 
    9.709639e-05, 0.0002100379, 0.0003448692, 0.0003421404, 0.0002332264, 
    0.0002403424, 0.000242127, 0.0002091188, 0.0001481717, 7.405162e-05,
  5.296057e-06, 3.200672e-06, 1.087957e-05, 2.709124e-05, 5.535626e-05, 
    7.596818e-05, 0.0001832949, 0.0003699787, 0.0004253148, 0.0003417288, 
    0.000267107, 0.0002569029, 0.0002839131, 0.0001927506, 8.08397e-05,
  1.156876e-06, 2.0134e-06, 4.263408e-06, 1.502282e-05, 3.991557e-05, 
    7.123232e-05, 0.0001603291, 0.000361861, 0.0005070686, 0.0004170369, 
    0.0003866296, 0.0003118666, 0.000327909, 0.0001896376, 8.748326e-05,
  1.018339e-06, 1.574869e-06, 3.217493e-06, 1.092117e-05, 3.090494e-05, 
    6.806753e-05, 0.0001233881, 0.0003370099, 0.0005191566, 0.0004917441, 
    0.0004537567, 0.0003502417, 0.0003457592, 0.000122154, 9.82709e-05,
  6.322639e-07, 1.0404e-06, 2.804771e-06, 7.641586e-06, 2.419612e-05, 
    5.973587e-05, 9.080485e-05, 0.0002524447, 0.0004765665, 0.0005015525, 
    0.0004884037, 0.0004219981, 0.0003107936, 0.0002233556, 8.185769e-05,
  4.159934e-07, 7.158492e-07, 2.092262e-06, 5.944728e-06, 2.120272e-05, 
    6.388444e-05, 7.882603e-05, 0.0001476913, 0.000376979, 0.0005294124, 
    0.0004446413, 0.0003761998, 0.0003101096, 0.0001808216, 7.384687e-05,
  1.203191e-06, 8.353352e-07, 2.287535e-06, 4.693193e-06, 2.181203e-05, 
    6.735428e-05, 9.409552e-05, 0.000156552, 0.0002424178, 0.0004926862, 
    0.0004722767, 0.000391842, 0.0002577201, 0.0001287228, 6.04436e-05,
  2.15382e-05, 7.286753e-06, 4.463863e-06, 6.972781e-06, 2.494904e-05, 
    6.425013e-05, 0.0001059905, 0.0001721564, 0.0003002171, 0.000455356, 
    0.000421875, 0.0004027346, 0.0002963224, 0.0001315212, 4.884268e-05,
  3.218112e-05, 1.717446e-05, 1.032525e-05, 1.301887e-05, 3.159839e-05, 
    4.398701e-05, 7.642149e-05, 0.000103065, 0.000281801, 0.0005660739, 
    0.0004948868, 0.0003748193, 0.0002715183, 9.590784e-05, 1.169693e-05,
  4.133514e-05, 2.0983e-05, 1.468171e-05, 1.910269e-05, 2.153138e-05, 
    3.676659e-05, 8.223801e-05, 0.0001039087, 0.0002843472, 0.0005910564, 
    0.0005181814, 0.0003236159, 0.0002016549, 4.706415e-05, 1.276419e-06,
  5.172771e-05, 6.220775e-05, 8.695615e-05, 8.782807e-05, 5.989947e-05, 
    3.393518e-05, 3.104463e-05, 2.648958e-05, 2.066908e-05, 1.695942e-05, 
    8.113684e-06, 1.438069e-05, 2.741401e-05, 2.68009e-05, 2.974934e-05,
  1.122373e-05, 1.498721e-05, 4.979026e-05, 5.919166e-05, 7.969352e-05, 
    5.803359e-05, 3.049025e-05, 2.810802e-05, 2.304664e-05, 1.592944e-05, 
    1.525009e-05, 1.433051e-05, 3.122619e-05, 4.241271e-05, 4.464157e-05,
  8.046563e-07, 2.631791e-06, 1.126348e-05, 4.636551e-05, 7.251049e-05, 
    7.174611e-05, 5.382827e-05, 3.440983e-05, 2.080086e-05, 1.435382e-05, 
    2.263471e-05, 2.424459e-05, 3.553788e-05, 5.838733e-05, 4.956575e-05,
  4.705022e-08, 4.946959e-07, 1.527708e-06, 4.912218e-05, 7.146287e-05, 
    8.196425e-05, 6.014842e-05, 4.256088e-05, 3.518347e-05, 4.543116e-05, 
    2.666146e-05, 3.465444e-05, 4.452492e-05, 4.439756e-05, 3.323244e-05,
  4.244514e-10, 2.93153e-08, 3.713696e-08, 2.203413e-05, 6.881528e-05, 
    7.655031e-05, 5.91535e-05, 6.209424e-05, 6.130229e-05, 5.098781e-05, 
    4.485362e-05, 4.17861e-05, 3.473738e-05, 3.477459e-05, 3.604652e-05,
  1.308624e-08, 7.634037e-10, 4.366887e-07, 1.640029e-05, 3.702735e-05, 
    3.61065e-05, 7.461917e-05, 7.262213e-05, 7.482606e-05, 7.798861e-05, 
    5.975577e-05, 4.042684e-05, 4.100649e-05, 3.094758e-05, 3.563788e-05,
  2.282449e-05, 1.395439e-05, 2.419064e-05, 3.095104e-05, 4.901819e-05, 
    9.67171e-06, 7.26492e-06, 2.755113e-05, 5.28352e-05, 6.208342e-05, 
    7.838021e-05, 6.370446e-05, 3.477677e-05, 2.857733e-05, 4.596056e-05,
  8.305231e-05, 7.331359e-05, 6.22844e-05, 5.184807e-05, 4.111856e-05, 
    1.644468e-05, 3.101757e-06, 1.974323e-06, 3.385361e-06, 1.288096e-05, 
    5.220555e-05, 6.453211e-05, 4.877429e-05, 4.165531e-05, 6.034068e-05,
  8.57739e-05, 9.938367e-05, 8.788518e-05, 7.649795e-05, 4.726478e-05, 
    6.722739e-06, 7.207277e-06, 5.691335e-06, 1.376105e-05, 2.685305e-05, 
    5.408668e-05, 7.019058e-05, 5.649732e-05, 6.158881e-05, 9.257975e-05,
  8.226412e-05, 0.0001019647, 0.0001130933, 9.804231e-05, 1.871082e-05, 
    1.192245e-05, 4.448818e-06, 1.438449e-05, 3.937255e-05, 4.919607e-05, 
    6.973216e-05, 7.596623e-05, 5.97879e-05, 0.0001011051, 0.0001224654,
  2.984582e-05, 3.166809e-05, 5.081999e-05, 4.846665e-05, 3.0249e-05, 
    1.247146e-05, 7.102687e-06, 4.289482e-06, 4.625016e-06, 3.30985e-07, 
    7.360496e-08, 1.944117e-07, 7.721432e-07, 4.15021e-06, 6.556432e-06,
  1.326908e-05, 7.713401e-06, 3.513947e-05, 3.312716e-05, 4.645675e-05, 
    3.288087e-05, 2.173049e-05, 1.060371e-05, 2.107095e-06, 3.107726e-07, 
    3.647274e-07, 1.574645e-07, 1.465581e-06, 5.830138e-06, 1.122196e-05,
  1.688607e-05, 9.883377e-06, 7.865518e-06, 3.341819e-05, 5.527934e-05, 
    5.044689e-05, 4.240618e-05, 2.54114e-05, 2.124803e-05, 1.158956e-05, 
    1.160596e-06, 1.62955e-06, 2.445122e-06, 8.624939e-06, 1.129646e-05,
  1.895747e-05, 9.892984e-06, 3.881894e-06, 4.320546e-05, 4.92184e-05, 
    6.021332e-05, 6.027563e-05, 4.315438e-05, 4.822795e-05, 4.409011e-05, 
    2.86176e-05, 8.125794e-06, 1.109955e-05, 1.248275e-05, 1.24535e-05,
  2.465548e-06, 8.532645e-06, 1.261051e-05, 3.771824e-05, 5.467286e-05, 
    6.445017e-05, 6.966684e-05, 6.527946e-05, 7.282188e-05, 7.179653e-05, 
    6.451763e-05, 2.902776e-05, 1.341783e-05, 7.615388e-06, 9.146505e-06,
  1.602268e-05, 2.015782e-05, 1.902603e-05, 3.227057e-05, 5.077913e-05, 
    4.781524e-05, 6.140766e-05, 8.03554e-05, 9.005584e-05, 9.57239e-05, 
    9.170853e-05, 5.444846e-05, 2.490752e-05, 6.654842e-06, 7.680625e-06,
  3.663751e-05, 3.232825e-05, 3.954353e-05, 4.54758e-05, 6.595939e-05, 
    1.723893e-05, 8.043391e-06, 2.957936e-05, 6.061594e-05, 7.372089e-05, 
    8.429132e-05, 7.925463e-05, 3.935506e-05, 4.529272e-06, 8.98703e-06,
  7.960959e-05, 7.213011e-05, 7.5744e-05, 7.482203e-05, 5.407105e-05, 
    2.203975e-05, 6.045084e-06, 2.233879e-06, 3.69742e-06, 1.25404e-05, 
    5.127529e-05, 7.383346e-05, 5.557484e-05, 7.211936e-06, 1.024348e-05,
  6.870614e-05, 8.30833e-05, 9.487029e-05, 0.0001042885, 8.312759e-05, 
    2.065554e-05, 1.225259e-05, 7.110611e-06, 1.322498e-05, 3.129386e-05, 
    4.752455e-05, 5.713989e-05, 5.409456e-05, 2.443245e-05, 8.527463e-06,
  6.037513e-05, 7.297879e-05, 9.110871e-05, 0.0001250542, 3.567547e-05, 
    2.989707e-05, 1.454037e-05, 1.761464e-05, 4.359317e-05, 5.076361e-05, 
    4.310448e-05, 4.3768e-05, 4.393066e-05, 3.215437e-05, 1.164649e-05,
  3.178622e-07, 3.625077e-07, 8.96455e-07, 1.806637e-06, 1.282045e-06, 
    4.649022e-07, 1.195122e-08, 6.532511e-10, 2.696997e-09, 5.659911e-08, 
    2.802973e-07, 8.21412e-06, 2.967047e-05, 3.364346e-05, 2.332141e-05,
  1.102589e-07, 4.387343e-08, 3.008057e-07, 1.643013e-06, 3.200037e-06, 
    1.916834e-06, 7.208862e-08, 2.02736e-07, 9.058788e-08, 7.74506e-07, 
    1.659919e-06, 1.842314e-05, 3.678432e-05, 2.749208e-05, 1.613944e-05,
  6.528695e-09, 5.005941e-09, 2.638502e-08, 6.98611e-07, 4.147545e-06, 
    4.507061e-06, 1.383935e-06, 7.460234e-08, 4.611128e-07, 2.415521e-06, 
    1.839229e-05, 3.102786e-05, 2.503713e-05, 1.292165e-05, 1.253938e-05,
  2.815429e-09, 2.876656e-09, 3.798577e-08, 1.671161e-06, 6.8853e-06, 
    8.442279e-06, 8.619545e-06, 4.868969e-06, 8.462479e-06, 1.759471e-05, 
    2.665491e-05, 2.294088e-05, 1.47335e-05, 1.576082e-05, 1.474273e-05,
  1.682553e-09, 1.087108e-09, 4.20145e-08, 2.329482e-06, 7.514777e-06, 
    1.196187e-05, 1.668422e-05, 1.540198e-05, 2.386136e-05, 3.619603e-05, 
    3.653347e-05, 3.227645e-05, 2.611139e-05, 2.180213e-05, 1.914705e-05,
  7.44182e-09, 2.977321e-10, 8.232151e-08, 3.395706e-06, 5.748882e-06, 
    7.467002e-06, 1.430922e-05, 1.930713e-05, 1.916748e-05, 2.545098e-05, 
    3.261976e-05, 2.370204e-05, 1.651752e-05, 1.832267e-05, 1.46389e-05,
  5.810072e-07, 8.409825e-08, 1.050514e-06, 2.920889e-06, 5.932159e-06, 
    2.194167e-06, 1.058798e-06, 2.098619e-06, 3.344566e-06, 5.240156e-06, 
    1.353801e-05, 1.712635e-05, 1.242765e-05, 1.329697e-05, 1.490015e-05,
  1.206462e-05, 8.126445e-06, 8.033449e-06, 7.775391e-06, 1.030408e-05, 
    4.500148e-06, 4.163797e-07, 9.742477e-08, 1.261636e-07, 1.205852e-07, 
    1.491034e-06, 4.013587e-06, 9.487864e-06, 5.754776e-06, 6.39967e-06,
  1.763063e-05, 1.612321e-05, 1.96039e-05, 1.897992e-05, 2.448859e-05, 
    3.404825e-06, 5.117035e-07, 3.321478e-08, 6.396748e-10, 1.940831e-07, 
    2.101138e-06, 5.023465e-06, 9.92844e-06, 1.738316e-05, 5.293e-06,
  2.2409e-05, 2.397109e-05, 2.91538e-05, 3.641059e-05, 1.46174e-05, 
    3.19667e-06, 2.625606e-06, 2.090379e-07, 9.703582e-07, 2.216304e-06, 
    3.558829e-06, 5.995934e-06, 7.615889e-06, 1.283251e-05, 1.173581e-05,
  7.232656e-06, 6.52235e-06, 6.53061e-06, 1.797851e-06, 9.48982e-08, 
    5.949528e-10, 1.323524e-11, 5.443848e-11, 1.182852e-10, 7.154606e-11, 
    4.476702e-11, 4.836243e-07, 2.822391e-06, 3.527941e-06, 2.021954e-06,
  1.135291e-06, 4.08456e-07, 4.700591e-06, 2.911118e-06, 2.658413e-06, 
    8.755318e-08, 1.010055e-08, 2.304153e-11, 3.690018e-11, 4.620642e-11, 
    5.875654e-08, 4.196208e-06, 7.202972e-06, 5.097088e-06, 1.115919e-06,
  2.318441e-07, 6.764191e-08, 1.678887e-07, 5.009784e-06, 8.256507e-06, 
    5.428494e-06, 1.515113e-06, 2.185423e-08, 4.338795e-10, 3.115955e-09, 
    1.310529e-06, 7.831166e-06, 1.092995e-05, 8.193049e-06, 1.491822e-06,
  1.225315e-06, 1.483945e-07, 3.780967e-09, 9.615094e-06, 1.432889e-05, 
    1.341754e-05, 7.986263e-06, 4.493021e-06, 9.737347e-07, 1.173167e-06, 
    5.472171e-06, 1.38024e-05, 1.786656e-05, 1.230838e-05, 3.61082e-06,
  1.026085e-06, 6.161089e-08, 1.170478e-09, 5.735409e-06, 2.198245e-05, 
    1.599936e-05, 2.40371e-05, 1.956366e-05, 1.328831e-05, 1.148271e-05, 
    1.690742e-05, 2.513047e-05, 2.135507e-05, 1.356425e-05, 5.342833e-06,
  1.775498e-06, 1.626211e-07, 1.36331e-08, 6.61865e-06, 1.806891e-05, 
    1.51878e-05, 3.210129e-05, 3.867301e-05, 3.223761e-05, 2.761133e-05, 
    3.382851e-05, 2.94488e-05, 2.457473e-05, 2.047102e-05, 1.26612e-05,
  1.255343e-06, 1.086358e-06, 3.380564e-06, 1.795264e-05, 2.647312e-05, 
    4.308833e-06, 5.945904e-06, 9.63785e-06, 1.688655e-05, 3.229071e-05, 
    4.018638e-05, 3.843444e-05, 2.750792e-05, 1.893734e-05, 1.293017e-05,
  2.05634e-05, 1.200382e-05, 1.480727e-05, 2.598464e-05, 1.927848e-05, 
    3.525883e-06, 3.50365e-06, 2.186915e-06, 2.577326e-06, 1.568814e-05, 
    3.914955e-05, 3.794216e-05, 2.948615e-05, 1.728748e-05, 1.622726e-05,
  3.82288e-05, 2.897387e-05, 3.897705e-05, 3.5684e-05, 2.628185e-05, 
    5.300847e-06, 9.733338e-07, 4.630647e-06, 1.753787e-05, 3.595176e-05, 
    4.069419e-05, 4.247726e-05, 3.152207e-05, 2.369421e-05, 1.308336e-05,
  4.3537e-05, 3.861107e-05, 5.929249e-05, 4.733816e-05, 2.367953e-05, 
    1.035493e-05, 5.681389e-06, 8.518751e-06, 3.450051e-05, 4.096506e-05, 
    4.854419e-05, 4.686522e-05, 3.649118e-05, 2.347046e-05, 1.864135e-05,
  3.515714e-08, 7.647794e-08, 1.589213e-06, 7.534904e-07, 9.319685e-10, 
    5.026705e-10, 2.116436e-11, 1.215455e-14, 1.144088e-11, 2.785353e-11, 
    6.289554e-13, 1.170749e-14, 2.545934e-09, 5.222353e-11, 3.830026e-09,
  2.017837e-07, 1.713416e-07, 1.179875e-06, 1.575424e-06, 1.336172e-06, 
    8.227083e-09, 7.939311e-09, 3.718512e-14, 9.180367e-14, 8.551721e-14, 
    1.725369e-15, 1.489968e-25, 1.148943e-08, 1.989788e-08, 3.588267e-09,
  7.495055e-07, 3.535667e-07, 3.142548e-07, 1.648525e-06, 7.199578e-06, 
    3.509414e-06, 1.324356e-06, 1.18148e-07, 1.510184e-09, 1.157903e-11, 
    6.159878e-13, 1.607731e-13, 4.445216e-08, 5.587813e-08, 4.962575e-11,
  1.111232e-06, 3.573842e-07, 2.066471e-07, 3.58117e-06, 1.27394e-05, 
    1.399295e-05, 1.55211e-05, 7.949922e-06, 1.018701e-06, 1.606418e-09, 
    3.666355e-10, 3.314957e-12, 2.742563e-08, 4.274946e-08, 3.436189e-09,
  1.04084e-07, 7.103916e-08, 2.626107e-08, 1.366955e-06, 7.983318e-06, 
    1.229437e-05, 3.064757e-05, 2.526423e-05, 1.770399e-05, 5.159802e-06, 
    3.971696e-08, 6.331534e-09, 2.247845e-09, 3.252147e-09, 2.151303e-10,
  3.699297e-09, 2.111164e-09, 7.351217e-10, 1.526557e-06, 4.17874e-06, 
    9.026504e-06, 2.006426e-05, 3.056323e-05, 3.86815e-05, 2.012809e-05, 
    8.037387e-06, 1.710861e-07, 1.312222e-07, 3.208055e-09, 5.738518e-11,
  7.967184e-08, 1.049976e-06, 1.22653e-06, 4.12252e-06, 4.855707e-06, 
    2.090318e-06, 1.878321e-07, 4.086462e-06, 1.149886e-05, 1.976655e-05, 
    1.332771e-05, 2.140612e-06, 8.833931e-07, 4.031128e-07, 6.929739e-08,
  1.106399e-05, 9.153558e-06, 8.389742e-06, 6.358567e-06, 7.762682e-06, 
    1.901758e-06, 1.099585e-06, 4.018047e-07, 2.375194e-07, 3.100627e-06, 
    1.837633e-05, 8.50868e-06, 2.671156e-06, 1.620818e-06, 1.866044e-07,
  2.361343e-05, 2.282938e-05, 2.304067e-05, 1.70881e-05, 2.909201e-05, 
    1.024454e-06, 2.340403e-07, 1.888065e-08, 2.355571e-07, 1.219054e-05, 
    1.921335e-05, 1.538355e-05, 6.135505e-06, 3.425786e-06, 3.169253e-07,
  2.711579e-05, 3.111528e-05, 4.02545e-05, 3.978399e-05, 8.824158e-06, 
    1.513276e-06, 6.023425e-07, 8.234703e-10, 4.953349e-06, 2.14406e-05, 
    1.921815e-05, 2.017632e-05, 1.110529e-05, 5.936067e-06, 2.650877e-07,
  5.648937e-06, 1.928815e-05, 4.851464e-05, 8.276069e-05, 8.341654e-05, 
    8.168854e-05, 8.125238e-05, 3.409215e-05, 8.957064e-07, 3.013586e-06, 
    4.413837e-06, 4.098102e-06, 1.869574e-06, 1.941952e-06, 4.923305e-06,
  4.868593e-06, 8.469674e-06, 2.801405e-05, 6.460524e-05, 8.888979e-05, 
    8.870552e-05, 6.537898e-05, 3.362595e-05, 8.254502e-06, 1.246371e-06, 
    6.930871e-06, 2.630016e-06, 1.638232e-06, 2.178586e-06, 1.629276e-06,
  3.487485e-06, 4.514718e-06, 7.907059e-06, 3.285417e-05, 6.939916e-05, 
    7.780355e-05, 4.741682e-05, 2.319214e-05, 1.898069e-05, 8.813259e-06, 
    2.807691e-06, 3.117526e-07, 1.384374e-07, 8.663453e-08, 8.871595e-07,
  2.36252e-06, 1.515185e-06, 1.029417e-06, 9.960696e-06, 4.196434e-05, 
    6.444203e-05, 3.083928e-05, 1.170076e-05, 9.968461e-06, 2.191758e-06, 
    2.385001e-07, 4.964704e-08, 1.415929e-09, 3.628413e-08, 1.731436e-07,
  1.510366e-06, 3.707209e-07, 1.754649e-07, 3.599437e-06, 1.710722e-05, 
    3.859717e-05, 3.24324e-05, 4.511094e-06, 3.517703e-06, 1.015765e-06, 
    5.260738e-08, 1.447691e-08, 7.644427e-10, 1.248198e-08, 8.06805e-08,
  4.862453e-07, 2.321399e-07, 5.722361e-08, 7.490618e-07, 6.247989e-06, 
    2.555138e-05, 3.071409e-05, 5.47976e-06, 1.486516e-06, 1.439781e-06, 
    3.28204e-07, 4.739459e-10, 6.539531e-10, 1.62533e-08, 4.92118e-08,
  1.09203e-09, 1.424542e-08, 3.642428e-08, 2.814974e-07, 9.156043e-07, 
    8.594528e-06, 1.571146e-05, 8.571394e-06, 9.589417e-07, 2.063113e-06, 
    1.349473e-06, 3.471113e-07, 1.86913e-07, 1.335028e-08, 1.20787e-08,
  5.031057e-09, 1.64415e-08, 2.568221e-07, 1.103381e-06, 2.453302e-06, 
    1.857228e-06, 4.134498e-06, 5.089949e-06, 1.173392e-06, 5.645587e-07, 
    3.574588e-06, 9.837255e-07, 6.271903e-07, 2.27003e-07, 2.612467e-08,
  1.455433e-06, 8.113427e-07, 6.986357e-07, 1.041676e-06, 9.76758e-06, 
    8.407275e-07, 3.915581e-07, 1.274627e-07, 2.966186e-07, 3.004659e-06, 
    5.276033e-06, 4.36723e-06, 9.379983e-07, 5.545268e-07, 3.984359e-08,
  4.419489e-06, 3.254754e-06, 3.069448e-06, 2.932739e-06, 2.136547e-06, 
    5.791417e-07, 2.721865e-06, 8.986908e-07, 6.495433e-06, 7.202962e-06, 
    7.840122e-06, 5.578714e-06, 1.420066e-06, 7.246685e-07, 1.572576e-07,
  2.279716e-05, 1.748029e-05, 1.589103e-05, 9.352789e-06, 5.516997e-06, 
    7.094951e-06, 1.505606e-05, 3.500136e-05, 4.043956e-05, 4.268655e-05, 
    6.759579e-05, 7.939598e-05, 3.998914e-05, 8.472254e-06, 1.610054e-06,
  4.101383e-05, 2.267134e-05, 1.498818e-05, 1.943715e-05, 1.824057e-05, 
    2.779781e-05, 4.451638e-05, 5.255634e-05, 4.657735e-05, 3.808526e-05, 
    7.925186e-05, 0.00011075, 4.533713e-05, 9.091485e-06, 2.620145e-07,
  5.23352e-05, 3.070349e-05, 2.67334e-05, 3.072275e-05, 3.058625e-05, 
    5.029837e-05, 7.562253e-05, 8.523351e-05, 0.000129269, 0.0001042657, 
    0.0001095651, 0.0001299621, 5.194938e-05, 9.672076e-06, 4.585129e-08,
  5.652912e-05, 3.019632e-05, 2.693286e-05, 4.08788e-05, 4.36634e-05, 
    6.138641e-05, 0.0001025648, 0.0001207129, 0.000124474, 0.0001058488, 
    0.000149255, 0.0001589282, 5.459281e-05, 5.741505e-06, 2.552458e-07,
  4.498152e-05, 2.281302e-05, 2.761989e-05, 4.25616e-05, 5.119636e-05, 
    6.637623e-05, 0.0001042779, 0.0001343534, 0.0001289603, 0.0001587341, 
    0.0001882514, 0.0001548132, 5.755459e-05, 1.044189e-05, 3.9675e-07,
  2.557549e-05, 1.722179e-05, 1.70273e-05, 4.505598e-05, 6.939243e-05, 
    8.369637e-05, 0.0001023352, 0.0001412585, 0.000128686, 0.0001752451, 
    0.000199907, 0.0001448718, 6.013829e-05, 6.674294e-06, 5.453908e-07,
  2.011249e-05, 2.971873e-05, 4.176633e-05, 6.101396e-05, 7.128032e-05, 
    8.288438e-05, 9.639272e-05, 8.915196e-05, 0.0001043373, 0.0001350636, 
    0.0002212875, 0.0001325476, 5.379811e-05, 9.677035e-06, 2.188707e-07,
  5.626365e-05, 7.525921e-05, 7.939481e-05, 7.730809e-05, 8.032031e-05, 
    5.52773e-05, 7.120331e-05, 9.610395e-05, 0.0001074405, 8.94583e-05, 
    0.0001662702, 0.0001324567, 4.000218e-05, 1.262306e-05, 4.413959e-07,
  4.567745e-05, 7.87264e-05, 0.0001095944, 7.470824e-05, 7.856359e-05, 
    5.370687e-05, 5.587002e-05, 3.395599e-05, 5.304758e-05, 7.423644e-05, 
    0.000184366, 0.0001201207, 3.620296e-05, 1.215755e-05, 3.047183e-07,
  2.527889e-05, 6.043021e-05, 0.000121727, 0.0001121205, 4.784448e-05, 
    4.961306e-05, 8.65477e-05, 6.285357e-05, 6.757546e-05, 7.164824e-05, 
    0.0001288782, 0.0001038737, 3.884e-05, 9.182693e-06, 1.604219e-07,
  6.36543e-06, 8.510234e-06, 9.435753e-06, 1.433271e-05, 9.978725e-06, 
    1.471757e-06, 2.993561e-06, 1.357443e-05, 1.814218e-05, 1.831623e-05, 
    3.024518e-05, 6.348289e-05, 9.969415e-05, 0.000105912, 8.984229e-05,
  1.629829e-06, 1.516437e-06, 3.633643e-06, 6.030774e-06, 6.742915e-06, 
    2.578907e-06, 6.324553e-06, 9.655877e-06, 1.446783e-05, 1.969221e-05, 
    3.863476e-05, 8.069526e-05, 9.316811e-05, 0.00010487, 8.418463e-05,
  1.804574e-07, 8.750506e-08, 9.963187e-08, 1.112432e-07, 3.714717e-06, 
    6.461397e-06, 3.11697e-06, 9.216986e-06, 1.349867e-05, 2.211445e-05, 
    4.544843e-05, 6.893373e-05, 8.792438e-05, 8.776195e-05, 6.652129e-05,
  2.408068e-09, 1.409114e-09, 6.628599e-10, 2.45347e-09, 1.756756e-06, 
    6.245763e-06, 2.893375e-06, 8.63173e-06, 1.407526e-05, 3.048046e-05, 
    5.094322e-05, 5.880682e-05, 7.811702e-05, 8.064357e-05, 5.881145e-05,
  1.41338e-11, 4.353165e-12, 2.500824e-12, 4.333139e-10, 2.588821e-07, 
    3.693413e-06, 3.469511e-06, 1.01121e-05, 1.288977e-05, 2.988258e-05, 
    3.354387e-05, 3.849584e-05, 4.967891e-05, 8.321254e-05, 6.151382e-05,
  1.00344e-08, 6.528819e-11, 1.320951e-10, 2.053984e-10, 1.815196e-07, 
    2.533139e-06, 4.865894e-06, 3.240034e-06, 6.427379e-06, 1.01895e-05, 
    1.721162e-05, 1.985499e-05, 3.360025e-05, 7.256301e-05, 5.812146e-05,
  5.64273e-06, 5.536761e-08, 8.807028e-07, 3.331088e-06, 4.573227e-06, 
    4.750756e-07, 8.014085e-08, 7.742321e-08, 2.994445e-08, 4.787562e-07, 
    4.863647e-06, 9.565049e-06, 2.409722e-05, 5.960981e-05, 5.207484e-05,
  4.492222e-05, 3.472218e-05, 2.785814e-05, 1.409737e-05, 9.134101e-06, 
    1.131677e-06, 6.661452e-08, 1.770008e-07, 5.033131e-09, 4.458239e-07, 
    1.140346e-06, 3.868797e-06, 1.783177e-05, 5.182252e-05, 4.831819e-05,
  4.718544e-05, 5.365727e-05, 5.731972e-05, 3.780988e-05, 2.685417e-05, 
    1.642573e-06, 2.438766e-07, 7.66667e-09, 8.981312e-10, 3.285092e-07, 
    6.988149e-07, 5.170764e-06, 1.935092e-05, 5.454353e-05, 4.394005e-05,
  5.251765e-05, 5.260493e-05, 7.034397e-05, 6.510695e-05, 1.140116e-05, 
    2.844022e-06, 9.701179e-07, 1.392108e-07, 1.882603e-07, 1.111567e-07, 
    3.867086e-07, 3.400377e-06, 2.092192e-05, 5.80581e-05, 4.156387e-05,
  4.362933e-06, 4.713658e-06, 6.631459e-06, 4.501785e-06, 2.512469e-07, 
    1.918601e-06, 4.404122e-06, 1.606597e-05, 3.007902e-05, 5.298714e-05, 
    7.647611e-05, 0.0001405392, 0.0001617848, 0.0001006584, 5.365321e-05,
  2.515781e-07, 2.628625e-07, 2.98381e-06, 4.434316e-06, 2.805935e-06, 
    1.085706e-06, 3.179871e-06, 1.651632e-05, 3.106975e-05, 5.240669e-05, 
    0.0001005236, 0.000163789, 0.0001527165, 7.636056e-05, 3.63311e-05,
  7.910399e-09, 7.91183e-09, 1.136406e-07, 1.956007e-06, 2.357232e-06, 
    1.285132e-06, 2.931753e-06, 1.011145e-05, 3.44462e-05, 6.019945e-05, 
    0.0001382949, 0.000151268, 0.0001099257, 5.476115e-05, 3.272608e-05,
  5.7311e-11, 8.700492e-11, 3.28783e-09, 1.176149e-06, 3.581267e-06, 
    6.250751e-06, 3.481453e-06, 1.037933e-05, 2.825504e-05, 6.506158e-05, 
    0.0001358049, 0.0001280743, 7.779056e-05, 3.460552e-05, 2.650841e-05,
  0, 1.123572e-26, 6.512758e-11, 4.591372e-08, 1.467994e-06, 1.944678e-06, 
    3.246552e-06, 8.646511e-06, 2.520189e-05, 5.5892e-05, 8.224427e-05, 
    5.747906e-05, 3.537491e-05, 2.488523e-05, 1.812121e-05,
  5.468789e-10, 1.76816e-27, 1.10741e-10, 1.227654e-09, 2.329987e-07, 
    7.414511e-07, 8.140314e-07, 8.04671e-06, 1.974104e-05, 2.717207e-05, 
    3.640183e-05, 2.575322e-05, 1.685706e-05, 2.119329e-05, 1.709913e-05,
  3.691009e-08, 1.698057e-09, 5.747139e-07, 5.345828e-07, 2.442327e-06, 
    4.029159e-07, 1.128512e-07, 9.512571e-08, 3.915739e-07, 5.326865e-06, 
    7.845279e-06, 6.640756e-06, 1.242898e-05, 1.903335e-05, 1.522216e-05,
  1.027308e-05, 8.930435e-06, 3.898341e-06, 3.555796e-06, 7.932461e-06, 
    2.812049e-06, 9.696247e-08, 3.331526e-08, 3.775379e-08, 9.573933e-09, 
    1.655224e-07, 4.26018e-06, 1.872107e-05, 2.08111e-05, 1.346585e-05,
  2.535875e-05, 2.743252e-05, 2.750265e-05, 2.471085e-05, 2.134013e-05, 
    3.498362e-06, 1.176871e-07, 5.691218e-09, 1.58046e-07, 1.962698e-06, 
    1.0267e-05, 2.233223e-05, 2.638035e-05, 1.384922e-05, 8.874689e-06,
  2.160774e-05, 3.597796e-05, 4.815489e-05, 4.645086e-05, 1.162902e-05, 
    7.590661e-06, 4.285797e-07, 3.303627e-09, 1.760777e-06, 5.404523e-06, 
    9.559586e-06, 1.14869e-05, 1.385398e-05, 9.396809e-06, 9.070842e-06,
  5.514996e-10, 1.231671e-07, 1.123704e-06, 1.550041e-06, 3.882022e-07, 
    5.218217e-07, 1.824721e-06, 1.337009e-05, 7.869365e-05, 0.0001486111, 
    0.0001833746, 0.0002254377, 0.0002455159, 0.0001909197, 0.0001384277,
  8.332233e-12, 2.525216e-09, 7.910038e-08, 1.136787e-06, 3.548762e-08, 
    1.101249e-06, 8.995504e-07, 4.402379e-06, 5.424456e-05, 0.0001076657, 
    0.0001706743, 0.0002234999, 0.0002298307, 0.0001960249, 0.0001114766,
  5.02454e-14, 3.476659e-11, 1.46014e-09, 6.080157e-08, 1.273226e-07, 
    4.488887e-07, 4.488544e-06, 1.304834e-05, 3.240849e-05, 9.099366e-05, 
    0.0001478237, 0.000206132, 0.0001889716, 0.0001656045, 9.982043e-05,
  8.410408e-17, 6.851252e-26, 1.156005e-10, 6.876703e-09, 8.93576e-07, 
    1.36426e-06, 4.856165e-06, 8.520601e-06, 3.15159e-05, 6.125836e-05, 
    0.0001004436, 0.0001353952, 0.0001610677, 0.0001424693, 0.0001006923,
  1.269514e-19, 7.001694e-27, 3.730762e-25, 1.382305e-09, 2.24975e-07, 
    1.956457e-06, 2.837985e-06, 8.722753e-06, 1.665182e-05, 3.019858e-05, 
    5.129655e-05, 6.217311e-05, 0.0001024266, 0.0001324094, 0.0001065503,
  4.58032e-10, 4.827312e-28, 2.197869e-26, 2.134109e-10, 1.118397e-08, 
    7.98742e-07, 2.022843e-06, 2.033381e-06, 7.543812e-06, 7.92178e-06, 
    1.326901e-05, 2.24514e-05, 5.188137e-05, 9.448459e-05, 0.0001064686,
  4.552794e-08, 5.981384e-10, 2.907517e-11, 5.506632e-12, 7.70736e-08, 
    3.139891e-07, 1.072435e-07, 1.01887e-07, 2.857371e-09, 1.877142e-07, 
    6.235476e-06, 1.267749e-05, 2.122286e-05, 4.780051e-05, 5.920977e-05,
  5.097229e-06, 3.180102e-06, 1.246557e-06, 1.085215e-06, 9.591874e-07, 
    6.367704e-07, 1.15517e-07, 1.206354e-07, 1.124197e-07, 8.430374e-10, 
    1.210906e-06, 5.372031e-06, 7.823115e-06, 2.311795e-05, 2.862999e-05,
  1.805954e-05, 1.885992e-05, 1.55637e-05, 1.306762e-05, 1.39306e-05, 
    8.012309e-07, 5.317603e-08, 1.845199e-09, 6.249941e-09, 7.824935e-07, 
    1.994089e-06, 1.966518e-06, 3.82737e-06, 9.787073e-06, 1.106842e-05,
  2.302396e-05, 2.675277e-05, 3.022866e-05, 3.432643e-05, 9.854587e-06, 
    4.836057e-06, 2.965314e-07, 1.061311e-09, 1.958907e-08, 3.650067e-07, 
    3.326224e-06, 2.101172e-06, 3.589025e-06, 6.326809e-06, 7.811701e-06,
  1.436922e-07, 1.682975e-07, 7.588805e-08, 1.945566e-08, 4.818178e-07, 
    7.008897e-07, 1.263186e-05, 5.321448e-05, 0.0001666873, 0.000233964, 
    0.0003052629, 0.0003734233, 0.0003953299, 0.0002291433, 9.68499e-05,
  8.464499e-10, 5.627025e-09, 5.566935e-08, 4.771501e-08, 4.432061e-08, 
    2.286048e-06, 8.885495e-06, 4.429169e-05, 0.0001508563, 0.0002194688, 
    0.0003003862, 0.000374578, 0.0004270432, 0.0003305555, 0.0001476357,
  2.192821e-12, 9.907506e-10, 1.481546e-08, 2.396493e-08, 7.014565e-09, 
    2.615314e-06, 1.447211e-05, 3.717811e-05, 0.000130475, 0.0002459368, 
    0.0002938477, 0.0003173129, 0.000398232, 0.0004040554, 0.0001751047,
  1.390013e-16, 1.650373e-10, 4.99174e-09, 1.270103e-08, 7.803023e-08, 
    2.651657e-06, 1.241757e-05, 4.176757e-05, 0.0001014551, 0.0002181047, 
    0.0002944783, 0.0003024896, 0.0003485982, 0.0004330011, 0.0002927366,
  1.079891e-09, 6.20594e-10, 2.02799e-09, 1.778189e-08, 2.977074e-07, 
    2.190201e-06, 5.065053e-06, 8.33376e-06, 4.861161e-05, 0.0001560725, 
    0.0002781036, 0.0003128446, 0.000315088, 0.0004751261, 0.0004216415,
  4.244571e-07, 4.27279e-07, 2.494163e-07, 1.869991e-06, 2.035277e-06, 
    2.718934e-09, 9.824993e-07, 7.375256e-07, 6.228465e-06, 9.411175e-05, 
    0.000285464, 0.0003714092, 0.0003571134, 0.0005488621, 0.0005790919,
  1.347466e-05, 9.095644e-06, 8.9748e-06, 5.719844e-06, 5.488477e-06, 
    9.929042e-07, 8.930891e-07, 1.233044e-06, 3.880131e-06, 7.414707e-05, 
    0.0002655756, 0.0003589713, 0.000344655, 0.0005859954, 0.000694536,
  1.675992e-05, 1.483962e-05, 1.626706e-05, 1.263072e-05, 4.128799e-06, 
    7.270012e-07, 1.28984e-06, 4.300451e-06, 1.445605e-05, 4.362065e-05, 
    0.0002021695, 0.000270282, 0.0002575786, 0.0005132837, 0.0007090769,
  2.134864e-05, 2.26437e-05, 2.281601e-05, 2.777563e-05, 1.2014e-05, 
    6.343381e-07, 5.675523e-07, 4.381674e-08, 1.11432e-05, 5.952843e-05, 
    0.0001436402, 0.0001845784, 0.0001619795, 0.0003757279, 0.0006265346,
  2.558451e-05, 2.689236e-05, 2.956632e-05, 3.594518e-05, 5.306721e-06, 
    3.833246e-06, 6.398886e-07, 7.496123e-09, 3.439542e-06, 3.366769e-05, 
    9.096561e-05, 0.0001267913, 9.227565e-05, 0.0002222425, 0.0004615302,
  6.177821e-08, 1.34735e-06, 1.73186e-06, 5.354254e-06, 5.187053e-06, 
    1.21574e-06, 3.435361e-08, 1.842505e-06, 1.439046e-05, 4.473669e-05, 
    8.609505e-05, 0.0001172888, 0.0001427114, 0.0001421239, 0.0001168168,
  1.194135e-10, 5.711953e-09, 4.8497e-07, 1.600249e-06, 3.810877e-06, 
    1.129061e-05, 8.302925e-06, 8.751291e-06, 1.210427e-05, 4.515366e-05, 
    0.0001020694, 0.0001564611, 0.0001912581, 0.0001430173, 0.0001076127,
  4.920048e-14, 2.707675e-11, 1.151935e-09, 1.979994e-07, 2.331758e-06, 
    1.299796e-05, 2.572721e-05, 3.076199e-05, 3.182091e-05, 5.911855e-05, 
    0.000104504, 0.0001595434, 0.0001675109, 0.000141978, 9.836695e-05,
  1.343439e-27, 5.577801e-12, 8.868955e-12, 3.985875e-10, 1.772169e-06, 
    1.487255e-05, 2.992996e-05, 4.907743e-05, 4.986401e-05, 5.563404e-05, 
    8.066074e-05, 0.0001173237, 0.0001272722, 8.910364e-05, 8.801385e-05,
  1.691573e-09, 1.065461e-08, 3.897317e-08, 9.532002e-07, 1.317414e-05, 
    1.962095e-05, 3.076519e-05, 4.143635e-05, 4.262535e-05, 3.999021e-05, 
    5.148231e-05, 7.152215e-05, 9.51226e-05, 0.0001016832, 8.251123e-05,
  6.195049e-07, 3.3541e-06, 6.18458e-06, 1.633664e-05, 2.073104e-05, 
    1.019601e-05, 7.29094e-06, 8.904612e-06, 9.512698e-06, 1.524619e-05, 
    4.948974e-05, 7.60155e-05, 0.0001115148, 0.0001274498, 8.30873e-05,
  3.805187e-06, 6.404679e-06, 1.384522e-05, 2.473504e-05, 1.720885e-05, 
    6.540882e-07, 4.23887e-08, 2.75312e-08, 1.504558e-07, 2.373152e-05, 
    8.040207e-05, 0.0001400037, 0.0001549177, 0.0001451647, 6.434492e-05,
  4.104455e-06, 8.42262e-06, 1.559769e-05, 2.778703e-05, 6.258887e-06, 
    8.234545e-07, 4.667324e-07, 5.42808e-07, 2.564024e-06, 2.601318e-05, 
    0.000122855, 0.0001812954, 0.0002001279, 0.0001629728, 6.430124e-05,
  2.006648e-06, 1.083562e-05, 1.77018e-05, 2.621332e-05, 6.299237e-06, 
    1.761101e-07, 1.433538e-07, 1.361729e-08, 1.104075e-05, 8.725332e-05, 
    0.0002063415, 0.0002408662, 0.0002329621, 0.0002085029, 9.684026e-05,
  2.565052e-06, 1.039892e-05, 1.800375e-05, 2.198611e-05, 6.892682e-06, 
    7.220878e-07, 2.495949e-07, 1.468522e-08, 1.691475e-05, 0.0001121183, 
    0.0002052985, 0.0002534676, 0.0002843845, 0.000238186, 0.0001778765,
  1.260697e-06, 2.600516e-07, 4.633459e-07, 9.642725e-09, 1.117281e-08, 
    8.832961e-09, 3.943049e-09, 1.156368e-09, 4.208323e-10, 5.047114e-09, 
    1.247608e-06, 5.262003e-06, 7.860317e-06, 1.268889e-06, 4.405663e-06,
  1.000657e-05, 1.829772e-06, 1.082884e-06, 3.272658e-07, 1.68237e-08, 
    2.223052e-07, 6.17731e-09, 1.062954e-08, 1.471616e-09, 2.746942e-08, 
    5.142076e-06, 7.132708e-06, 9.946969e-06, 1.343792e-05, 1.302151e-05,
  2.834655e-05, 1.706254e-05, 1.731211e-07, 6.150294e-07, 5.645794e-07, 
    6.9286e-07, 1.663244e-06, 6.430759e-07, 1.42174e-07, 1.944022e-07, 
    6.821404e-06, 8.540323e-06, 9.928727e-06, 1.984936e-05, 1.978463e-05,
  2.846112e-05, 2.24124e-05, 2.602881e-06, 2.112797e-06, 5.445018e-07, 
    1.235524e-06, 3.671927e-06, 6.422561e-06, 6.782846e-06, 9.046574e-06, 
    6.29305e-06, 9.268355e-06, 1.548389e-05, 1.634081e-05, 2.175285e-05,
  1.259614e-05, 1.424658e-05, 1.091086e-05, 2.333892e-06, 1.675308e-06, 
    1.806611e-06, 6.447209e-06, 1.019398e-05, 1.575754e-05, 1.877631e-05, 
    1.450583e-05, 1.104671e-05, 1.774452e-05, 1.438298e-05, 1.969069e-05,
  3.835197e-06, 8.077187e-06, 1.426081e-06, 2.021534e-06, 2.73407e-06, 
    4.14282e-06, 5.531046e-06, 6.365996e-06, 1.041877e-05, 1.705288e-05, 
    1.439996e-05, 1.255543e-05, 1.464536e-05, 1.584845e-05, 1.515173e-05,
  2.464547e-07, 1.623944e-06, 1.304661e-06, 1.120429e-06, 4.678628e-06, 
    1.546552e-06, 5.158259e-08, 1.316791e-07, 3.00246e-07, 5.503891e-06, 
    4.752067e-06, 1.07872e-05, 1.458736e-05, 2.396035e-05, 2.840846e-05,
  2.784694e-06, 1.84752e-06, 1.503253e-06, 2.252151e-06, 4.096818e-06, 
    2.197623e-06, 2.909276e-08, 3.237631e-09, 2.508897e-08, 5.02889e-08, 
    6.020358e-07, 8.005199e-06, 1.533507e-05, 3.219542e-05, 3.244786e-05,
  6.297424e-06, 2.222235e-06, 2.713567e-06, 4.14594e-06, 6.375074e-06, 
    1.96642e-06, 4.252048e-09, 8.927807e-10, 7.071965e-11, 1.642356e-06, 
    5.721448e-06, 1.569234e-05, 2.441856e-05, 2.745058e-05, 3.301167e-05,
  1.990156e-06, 3.009553e-06, 4.709633e-06, 5.183977e-06, 6.711685e-06, 
    1.52627e-06, 3.460413e-07, 9.894778e-09, 2.582484e-06, 1.802105e-05, 
    3.742619e-05, 3.578599e-05, 3.134707e-05, 4.20955e-05, 6.057353e-05,
  1.014218e-05, 9.339758e-06, 1.665011e-05, 1.500579e-05, 2.820713e-06, 
    3.785155e-08, 3.635547e-08, 2.009132e-07, 8.069068e-08, 7.237769e-07, 
    2.738413e-06, 5.05486e-06, 7.161e-06, 7.442628e-06, 4.207772e-06,
  1.187676e-06, 5.529131e-07, 6.186406e-06, 1.248507e-05, 1.755794e-05, 
    5.159924e-06, 1.679766e-07, 5.8014e-07, 2.71256e-07, 1.015907e-06, 
    4.220452e-06, 9.077919e-06, 1.370174e-05, 8.742712e-06, 4.432857e-06,
  3.254097e-06, 1.956978e-06, 3.658442e-07, 1.06503e-05, 4.091691e-05, 
    2.668098e-05, 9.918353e-06, 3.213096e-06, 1.391155e-06, 6.266977e-06, 
    8.804004e-06, 1.411632e-05, 1.699949e-05, 1.072697e-05, 6.11319e-06,
  2.934151e-06, 1.208508e-06, 1.603768e-06, 3.162276e-05, 5.43667e-05, 
    5.078859e-05, 3.643976e-05, 3.012322e-05, 1.16646e-05, 1.167869e-05, 
    1.246632e-05, 2.246446e-05, 2.289649e-05, 1.016635e-05, 6.624494e-06,
  3.234717e-07, 5.960791e-07, 4.833224e-06, 3.334622e-05, 5.095487e-05, 
    5.970875e-05, 5.98769e-05, 4.067855e-05, 2.913084e-05, 2.217828e-05, 
    1.831587e-05, 2.498864e-05, 2.434817e-05, 1.461914e-05, 7.621116e-06,
  3.714754e-07, 1.217765e-06, 7.424047e-06, 2.02484e-05, 4.17288e-05, 
    4.13879e-05, 5.176618e-05, 6.630535e-05, 4.971531e-05, 4.151663e-05, 
    3.070633e-05, 2.194613e-05, 2.302924e-05, 2.062382e-05, 1.208732e-05,
  4.100753e-06, 4.327658e-06, 1.733742e-05, 4.640928e-05, 5.135614e-05, 
    6.409807e-05, 3.596663e-05, 4.053919e-05, 4.065592e-05, 4.332773e-05, 
    4.250012e-05, 3.793129e-05, 3.48762e-05, 2.584971e-05, 1.474647e-05,
  4.564986e-05, 2.567258e-05, 3.449082e-05, 6.062577e-05, 8.579979e-05, 
    7.857549e-05, 5.887153e-05, 3.284023e-05, 9.844318e-06, 2.410947e-05, 
    4.3374e-05, 5.428232e-05, 4.790248e-05, 2.928986e-05, 1.311721e-05,
  5.83266e-05, 5.025103e-05, 5.234186e-05, 6.143453e-05, 0.0001402403, 
    8.180891e-05, 2.788581e-05, 1.469438e-05, 2.374814e-05, 4.161016e-05, 
    6.000681e-05, 6.565356e-05, 5.188618e-05, 2.818467e-05, 8.638274e-06,
  4.910002e-05, 6.516794e-05, 7.467237e-05, 8.196593e-05, 0.0001005593, 
    6.085515e-05, 4.99289e-05, 2.084919e-05, 3.675048e-05, 4.827426e-05, 
    7.702072e-05, 7.115019e-05, 4.501184e-05, 2.302873e-05, 6.892304e-06,
  1.444826e-08, 5.458712e-09, 1.612944e-09, 1.318536e-10, 6.474542e-12, 
    4.963406e-27, 0, 0, 0, 0, 0, 1.899253e-09, 2.61278e-07, 6.633024e-07, 
    3.674328e-07,
  1.87133e-08, 6.605764e-09, 3.228048e-09, 2.069091e-09, 1.179861e-10, 
    5.916256e-12, 6.563336e-14, 2.669875e-10, 4.956325e-12, 7.640716e-14, 
    1.312968e-10, 5.598217e-07, 8.618305e-07, 1.580461e-06, 2.666672e-07,
  1.31045e-06, 1.868067e-07, 4.109363e-09, 4.057678e-09, 1.521784e-09, 
    8.769538e-11, 7.669445e-09, 2.315345e-08, 4.662699e-08, 4.905429e-09, 
    2.289863e-07, 1.613489e-06, 1.910187e-06, 7.156518e-08, 6.132512e-07,
  3.404724e-06, 9.527243e-07, 1.070979e-08, 2.301141e-09, 9.754703e-10, 
    2.413953e-09, 9.521758e-09, 3.716231e-08, 5.749263e-08, 3.976355e-07, 
    7.933217e-06, 7.709757e-06, 4.433395e-06, 5.466606e-08, 6.740203e-07,
  2.672086e-06, 1.164685e-06, 1.39498e-08, 4.162346e-09, 2.593374e-09, 
    9.572866e-10, 6.586479e-08, 1.823087e-06, 2.365334e-06, 4.775482e-06, 
    1.073051e-05, 8.788962e-06, 7.354397e-06, 1.381093e-06, 9.037257e-08,
  2.504252e-06, 1.519828e-06, 1.648818e-08, 2.600963e-07, 3.763187e-08, 
    1.891972e-07, 2.198552e-08, 5.641112e-07, 6.690598e-07, 3.653258e-06, 
    1.165344e-05, 6.358648e-06, 5.375805e-06, 3.215117e-06, 1.387762e-07,
  2.977073e-06, 2.256432e-06, 7.545044e-07, 3.073917e-06, 1.934839e-06, 
    2.114213e-07, 3.562889e-08, 1.32558e-08, 2.053093e-08, 2.897243e-07, 
    7.506417e-06, 8.284505e-06, 1.063085e-05, 4.575028e-06, 3.809118e-07,
  1.290847e-05, 1.125342e-05, 8.757277e-06, 4.751899e-06, 2.684874e-06, 
    5.155363e-07, 2.880301e-07, 3.767875e-08, 3.385622e-08, 1.769746e-08, 
    5.329263e-08, 5.645943e-06, 9.602714e-06, 6.945893e-06, 1.600072e-06,
  2.359235e-05, 3.289079e-05, 3.377105e-05, 2.466554e-05, 1.193014e-05, 
    2.807297e-06, 1.92905e-07, 1.488304e-08, 6.273718e-10, 5.639089e-10, 
    4.23889e-07, 2.968638e-06, 5.451924e-06, 5.612915e-06, 2.743493e-06,
  2.221965e-05, 3.1125e-05, 4.230702e-05, 4.261132e-05, 1.753282e-05, 
    2.997115e-06, 1.318464e-06, 2.328126e-08, 5.158254e-09, 6.275752e-09, 
    4.291282e-07, 1.999183e-06, 2.106934e-06, 3.825196e-06, 2.315108e-06,
  1.056851e-07, 2.041674e-07, 1.477298e-08, 1.15084e-08, 1.412697e-08, 
    9.942911e-09, 6.39412e-09, 1.625487e-09, 4.163248e-09, 6.238423e-09, 
    1.222505e-08, 1.174261e-07, 1.144948e-06, 5.840062e-07, 4.704079e-09,
  4.338791e-07, 4.195736e-08, 3.846105e-08, 1.074532e-08, 1.594205e-08, 
    3.177604e-08, 4.156331e-09, 2.445166e-09, 1.268839e-09, 2.124811e-09, 
    3.602723e-08, 1.271327e-07, 5.869553e-07, 3.304589e-07, 2.581638e-09,
  3.659843e-08, 2.668271e-08, 3.261447e-08, 1.171153e-08, 1.787488e-08, 
    6.31659e-08, 5.299136e-08, 8.936394e-10, 7.955459e-10, 8.259656e-08, 
    4.897595e-08, 2.693898e-08, 9.668386e-08, 6.955304e-08, 3.06357e-09,
  2.70449e-08, 3.410903e-08, 2.003688e-08, 1.673656e-08, 9.3882e-08, 
    3.588072e-07, 3.458094e-07, 4.144537e-08, 1.43739e-07, 2.111166e-07, 
    1.382063e-07, 2.339467e-07, 1.634725e-07, 2.015021e-07, 4.992461e-08,
  7.470669e-09, 1.773298e-08, 2.692181e-08, 2.360152e-07, 1.147916e-06, 
    1.312529e-06, 2.744507e-06, 2.87339e-06, 2.338334e-06, 2.07153e-06, 
    8.807828e-07, 5.268199e-07, 5.595051e-07, 4.190998e-07, 3.025909e-08,
  2.878488e-09, 1.203114e-08, 2.145357e-08, 3.894005e-07, 3.46656e-06, 
    2.151276e-06, 4.069256e-06, 5.111289e-06, 6.59728e-06, 8.695702e-06, 
    3.9553e-06, 2.153714e-06, 2.076183e-06, 4.631725e-07, 2.401128e-07,
  7.014378e-08, 4.903861e-09, 4.171513e-07, 1.84846e-06, 5.469323e-06, 
    7.475209e-06, 6.87213e-07, 3.863732e-07, 1.679569e-06, 4.509304e-06, 
    9.29857e-06, 8.055199e-06, 6.896385e-06, 2.368041e-06, 4.960197e-07,
  5.312139e-06, 3.301752e-07, 6.984961e-07, 3.563521e-06, 2.240531e-05, 
    2.057786e-05, 5.374106e-06, 1.033205e-06, 5.379516e-07, 5.869478e-07, 
    1.171427e-05, 1.233202e-05, 9.019493e-06, 2.06562e-06, 1.440937e-06,
  1.0976e-05, 3.196551e-06, 1.934605e-06, 8.48741e-06, 4.526493e-05, 
    3.065984e-05, 7.782239e-06, 3.003785e-06, 2.191163e-06, 7.699514e-06, 
    1.67481e-05, 1.737131e-05, 1.293792e-05, 4.149155e-06, 1.280475e-06,
  1.131665e-05, 8.696025e-06, 4.025958e-06, 1.137995e-05, 2.966145e-05, 
    1.798732e-05, 2.423092e-05, 1.308808e-05, 1.580153e-05, 1.607801e-05, 
    1.630742e-05, 2.125893e-05, 1.532096e-05, 4.066047e-06, 1.45339e-06,
  3.872058e-10, 2.832056e-10, 2.563662e-10, 3.678927e-09, 4.789472e-09, 
    2.319921e-09, 2.560767e-10, 1.134703e-10, 1.447181e-10, 1.039086e-10, 
    8.934135e-11, 1.085199e-07, 1.802916e-06, 6.091067e-06, 9.064262e-06,
  2.631931e-10, 4.467363e-10, 2.920639e-10, 6.843917e-10, 3.756286e-09, 
    3.840893e-09, 4.732198e-09, 1.531805e-09, 1.744213e-10, 5.883539e-11, 
    1.277338e-10, 8.781495e-08, 1.533672e-06, 8.347547e-06, 1.162579e-05,
  7.393496e-09, 6.392201e-10, 3.711473e-10, 6.506902e-10, 1.520943e-09, 
    2.567025e-09, 4.656075e-08, 6.01982e-08, 2.299559e-09, 1.325504e-10, 
    1.806404e-07, 6.056255e-07, 1.069281e-06, 5.274481e-06, 1.495964e-05,
  7.506069e-07, 2.695278e-08, 4.503293e-10, 4.92729e-07, 7.927837e-07, 
    5.914408e-07, 3.077046e-07, 8.405486e-07, 4.992867e-07, 7.616875e-07, 
    1.754254e-06, 2.212369e-06, 1.863521e-06, 4.823612e-06, 8.923704e-06,
  2.014056e-07, 2.295036e-08, 4.94735e-10, 7.05279e-07, 1.518663e-06, 
    1.720741e-06, 2.683086e-06, 2.077073e-06, 2.533178e-06, 4.273464e-06, 
    4.780513e-06, 4.11542e-06, 3.228755e-06, 4.319719e-06, 1.127731e-05,
  5.774845e-06, 1.291753e-06, 8.417636e-07, 1.538063e-06, 2.420461e-06, 
    2.949535e-06, 4.123895e-06, 6.893954e-06, 6.92766e-06, 1.081795e-05, 
    1.058533e-05, 3.308534e-06, 3.73896e-06, 5.89272e-06, 1.427023e-05,
  7.937831e-06, 6.409791e-06, 4.308516e-06, 4.352113e-06, 3.74209e-06, 
    3.88705e-07, 6.917591e-09, 3.118032e-08, 1.785347e-06, 5.902817e-06, 
    9.886023e-06, 9.841944e-06, 8.293351e-06, 7.383053e-06, 1.267276e-05,
  3.596778e-05, 2.157141e-05, 1.908447e-05, 7.235445e-06, 4.89603e-06, 
    3.959686e-07, 3.118823e-08, 2.312928e-08, 2.105911e-08, 3.370247e-08, 
    5.982562e-06, 9.246201e-06, 1.126867e-05, 1.16052e-05, 1.434284e-05,
  2.559816e-05, 3.441181e-05, 4.45864e-05, 2.424467e-05, 2.226792e-05, 
    5.434874e-07, 1.073821e-08, 1.406836e-09, 2.027169e-09, 1.957457e-06, 
    5.826457e-06, 1.242542e-05, 1.213895e-05, 1.254993e-05, 1.364869e-05,
  2.658869e-05, 3.809684e-05, 5.338625e-05, 5.512504e-05, 7.379827e-06, 
    1.213041e-06, 1.08446e-06, 1.810668e-06, 3.894486e-06, 5.127372e-06, 
    7.080798e-06, 1.301528e-05, 1.26332e-05, 1.495468e-05, 1.514011e-05,
  1.58384e-07, 4.275984e-07, 1.243547e-08, 4.922314e-06, 3.088298e-05, 
    3.439948e-05, 1.043102e-05, 1.316488e-07, 5.167749e-09, 7.572484e-08, 
    1.784345e-07, 1.145137e-06, 1.482927e-07, 1.25329e-07, 4.650184e-11,
  3.009127e-08, 2.493667e-07, 2.547784e-09, 8.242989e-09, 1.02136e-06, 
    6.418792e-06, 9.216143e-06, 1.798518e-07, 8.939216e-09, 1.313286e-07, 
    1.303011e-06, 1.670071e-06, 5.961407e-08, 5.404701e-08, 3.333852e-10,
  3.387666e-09, 5.324831e-08, 1.643223e-07, 2.148835e-09, 5.100962e-09, 
    5.514657e-07, 3.93464e-06, 2.47952e-06, 3.814757e-07, 1.239004e-06, 
    3.163656e-06, 1.284483e-06, 1.275846e-06, 2.259064e-07, 1.014333e-08,
  4.841211e-10, 1.124347e-08, 3.939896e-08, 2.588009e-08, 1.525838e-09, 
    8.724006e-09, 6.432343e-07, 3.463086e-06, 1.744157e-06, 2.614292e-06, 
    1.773439e-06, 3.015035e-06, 2.094086e-06, 3.113281e-07, 1.93497e-07,
  6.392514e-11, 1.500141e-09, 1.313018e-08, 3.071713e-08, 8.823882e-10, 
    8.524074e-10, 9.622e-09, 6.843314e-07, 2.877845e-06, 4.368704e-06, 
    3.513232e-06, 3.183456e-06, 1.821199e-06, 8.170836e-07, 4.553166e-07,
  1.468577e-08, 2.557953e-10, 2.428962e-09, 3.538534e-08, 1.130146e-09, 
    5.613844e-10, 6.539597e-10, 1.808497e-07, 2.664329e-06, 3.580611e-06, 
    3.510524e-06, 1.593357e-06, 1.424906e-06, 7.543194e-07, 1.030632e-07,
  1.288081e-06, 4.387584e-08, 1.100049e-09, 1.70262e-08, 1.092621e-09, 
    1.11792e-08, 1.538465e-08, 1.746753e-08, 1.539021e-07, 2.406676e-06, 
    5.336787e-06, 5.990629e-06, 2.435144e-06, 1.414991e-06, 1.69847e-07,
  2.171263e-05, 1.194131e-05, 8.755382e-06, 2.249754e-06, 4.262454e-08, 
    9.487438e-09, 4.122626e-09, 5.518354e-09, 4.264934e-09, 1.800658e-08, 
    1.113581e-06, 2.639633e-06, 2.336231e-06, 1.109774e-06, 6.024684e-07,
  1.968286e-05, 2.258958e-05, 3.135241e-05, 2.448029e-05, 1.703091e-05, 
    4.413704e-07, 3.533158e-09, 6.376134e-10, 2.137278e-10, 3.655547e-07, 
    3.251844e-06, 4.72613e-06, 2.930386e-06, 1.007379e-06, 7.681963e-07,
  2.433838e-05, 3.407871e-05, 3.839881e-05, 4.941832e-05, 1.408351e-05, 
    1.563517e-06, 2.777575e-07, 1.672981e-08, 1.042518e-06, 2.672676e-06, 
    4.408905e-06, 6.149752e-06, 5.782527e-06, 1.44446e-06, 2.630731e-07,
  3.467738e-07, 1.803433e-07, 1.235443e-08, 1.145137e-05, 0.0001661829, 
    0.000435148, 0.0004001185, 0.0003309935, 0.0001327669, 5.379949e-05, 
    3.485457e-05, 2.237759e-05, 1.338941e-05, 5.468188e-06, 5.270264e-06,
  1.873295e-07, 3.59725e-07, 9.835708e-08, 2.233159e-07, 3.758728e-05, 
    0.0002619187, 0.0003734493, 0.0003313481, 0.0002352035, 0.0001446571, 
    5.706699e-05, 2.360981e-05, 9.774296e-06, 7.550711e-06, 9.050742e-06,
  1.165699e-07, 2.675707e-07, 1.462722e-07, 5.468344e-09, 8.824806e-06, 
    0.0001336699, 0.0002988932, 0.0002432344, 0.000251695, 0.0002408521, 
    0.0001108653, 3.087035e-05, 1.160373e-05, 7.735983e-06, 7.63887e-06,
  6.32721e-08, 1.983561e-07, 1.463603e-07, 1.096599e-08, 9.32413e-09, 
    4.930342e-05, 0.0001846316, 0.0001752749, 0.0002172089, 0.0002416263, 
    0.0001844986, 3.836145e-05, 9.824269e-06, 4.089289e-06, 6.732041e-06,
  1.270916e-08, 1.054297e-07, 1.793099e-07, 1.17857e-08, 7.035279e-09, 
    1.120361e-05, 8.603471e-05, 0.0001271413, 0.0001514355, 0.000288126, 
    0.000215461, 4.945436e-05, 1.416358e-05, 5.203925e-06, 3.254648e-06,
  7.90685e-09, 3.706403e-08, 4.578991e-08, 7.582347e-08, 9.094557e-09, 
    2.105149e-06, 5.277593e-05, 8.195268e-05, 7.450741e-05, 0.0002340988, 
    0.0002202736, 5.698471e-05, 1.831996e-05, 2.890212e-06, 5.039608e-07,
  6.92804e-07, 1.230008e-08, 6.149556e-09, 4.348908e-09, 1.283312e-08, 
    6.487973e-06, 3.620597e-05, 9.008848e-05, 5.412798e-05, 0.0001181496, 
    0.000195199, 7.965844e-05, 2.376818e-05, 3.143061e-06, 1.023328e-07,
  1.17895e-05, 6.174043e-06, 2.663036e-06, 3.410424e-08, 3.906202e-09, 
    2.950225e-06, 2.675877e-05, 7.265672e-05, 7.516686e-05, 7.064161e-05, 
    0.0001207193, 7.964041e-05, 3.183408e-05, 4.18131e-06, 3.138572e-08,
  1.065357e-05, 1.602552e-05, 2.269045e-05, 4.8212e-06, 2.209863e-06, 
    1.146493e-06, 7.68958e-06, 2.450022e-05, 4.108368e-05, 4.016531e-05, 
    4.572371e-05, 5.688428e-05, 1.994789e-05, 4.869831e-06, 4.491805e-08,
  1.317255e-05, 2.373767e-05, 2.961158e-05, 2.897797e-05, 4.323349e-06, 
    6.879994e-07, 3.680317e-06, 6.285708e-06, 1.197597e-05, 7.426361e-06, 
    9.661263e-06, 1.865015e-05, 1.189469e-05, 2.055917e-06, 2.003407e-07,
  1.316038e-11, 3.119315e-10, 1.188605e-10, 3.180328e-10, 2.237419e-07, 
    4.941221e-06, 1.299189e-05, 2.249661e-05, 1.993726e-05, 1.414994e-05, 
    1.615772e-05, 3.92062e-05, 6.310963e-05, 5.527405e-05, 4.08712e-05,
  9.676937e-12, 1.005429e-10, 3.541639e-10, 2.378878e-10, 7.816625e-09, 
    5.279744e-06, 1.888574e-05, 2.573603e-05, 3.122202e-05, 3.14183e-05, 
    5.238257e-05, 7.422615e-05, 7.9912e-05, 6.561048e-05, 3.676034e-05,
  1.338833e-11, 8.480289e-11, 3.204598e-10, 3.363191e-10, 1.584932e-10, 
    3.28841e-06, 2.1984e-05, 2.960621e-05, 3.111373e-05, 4.189783e-05, 
    7.050568e-05, 9.673417e-05, 8.873235e-05, 5.840284e-05, 3.333289e-05,
  4.134454e-11, 5.499546e-11, 2.146353e-10, 6.388449e-10, 4.086257e-10, 
    3.386394e-06, 2.436735e-05, 4.462069e-05, 3.900182e-05, 4.542137e-05, 
    7.24602e-05, 7.895978e-05, 8.159146e-05, 4.729345e-05, 3.673914e-05,
  6.512504e-11, 4.576544e-11, 2.399793e-10, 7.184274e-10, 6.766789e-10, 
    2.945657e-07, 1.724546e-05, 6.855799e-05, 6.133885e-05, 6.515623e-05, 
    9.379534e-05, 0.0001107863, 7.53623e-05, 5.868818e-05, 3.304363e-05,
  3.00679e-10, 3.707047e-11, 2.246545e-10, 3.602199e-09, 1.368027e-09, 
    1.915318e-07, 3.436213e-06, 5.296665e-05, 0.0001186863, 0.0001098297, 
    0.0001371575, 9.520832e-05, 6.988792e-05, 5.611463e-05, 3.49793e-05,
  5.27516e-07, 6.237992e-09, 1.84097e-08, 1.718562e-08, 1.728951e-09, 
    3.300281e-07, 9.217414e-06, 8.557725e-05, 0.0001133363, 0.000169625, 
    0.0002048482, 0.000136766, 8.250953e-05, 5.713857e-05, 3.920919e-05,
  1.027543e-05, 5.110573e-06, 2.351225e-06, 2.141119e-07, 7.919364e-08, 
    3.838652e-07, 1.247911e-05, 8.964155e-05, 0.0001503252, 0.0001970601, 
    0.0002754293, 0.0001569527, 8.775496e-05, 6.64141e-05, 4.553351e-05,
  1.524109e-05, 1.782716e-05, 1.392944e-05, 8.969029e-06, 6.421356e-06, 
    5.809896e-07, 3.868156e-06, 6.049974e-05, 0.0001214772, 0.0002030891, 
    0.0003187689, 0.0003046824, 0.0001258681, 7.626928e-05, 5.105437e-05,
  1.756212e-05, 2.231046e-05, 2.67005e-05, 2.239002e-05, 7.152923e-06, 
    1.244304e-06, 3.909166e-06, 4.26081e-05, 8.561998e-05, 0.0001385062, 
    0.0002450003, 0.0003265816, 0.0001778003, 7.997978e-05, 5.367854e-05,
  4.393502e-10, 8.532986e-11, 7.793115e-11, 4.531543e-12, 2.585969e-16, 
    5.667172e-12, 1.785841e-15, 2.192904e-14, 2.644595e-09, 2.051189e-08, 
    4.804976e-07, 1.289747e-05, 3.789263e-05, 5.236722e-05, 3.796518e-05,
  2.114319e-09, 4.384423e-10, 7.398753e-11, 5.864131e-11, 3.381061e-14, 
    1.005558e-15, 3.040074e-15, 1.494107e-14, 3.129462e-09, 1.554914e-08, 
    1.108988e-06, 1.237314e-05, 3.725738e-05, 3.244051e-05, 1.965857e-05,
  4.30117e-09, 1.115104e-09, 2.373797e-10, 5.780078e-11, 4.470962e-12, 
    1.163441e-12, 1.571094e-15, 8.095749e-10, 8.081348e-09, 8.930031e-08, 
    2.178702e-06, 1.785696e-05, 2.285273e-05, 2.374685e-05, 1.269486e-05,
  6.320414e-09, 2.577242e-09, 4.672747e-10, 7.379403e-11, 1.796093e-12, 
    4.175237e-11, 2.736686e-11, 9.047836e-10, 1.048873e-07, 6.010378e-07, 
    9.665995e-06, 1.221848e-05, 1.441412e-05, 9.620137e-06, 1.155949e-05,
  1.067777e-08, 3.126815e-09, 1.018741e-09, 1.349002e-10, 1.043056e-11, 
    2.362869e-09, 3.167436e-12, 3.578777e-08, 7.320567e-07, 3.773994e-06, 
    1.406777e-05, 9.912679e-06, 5.2527e-06, 1.104344e-05, 5.72031e-06,
  8.446904e-09, 3.658039e-09, 1.376255e-09, 1.977935e-10, 2.694832e-11, 
    6.641031e-11, 1.304788e-08, 1.863415e-07, 5.897808e-07, 4.931601e-06, 
    8.048879e-06, 3.06221e-06, 2.453179e-06, 2.720002e-06, 4.521294e-06,
  1.025987e-08, 2.857261e-09, 1.35093e-09, 6.739652e-10, 1.333906e-10, 
    4.021114e-12, 3.507448e-10, 5.566515e-09, 6.704724e-09, 5.117013e-07, 
    4.741782e-06, 3.636725e-06, 1.389573e-06, 9.198319e-07, 2.133324e-06,
  1.789395e-07, 4.730879e-08, 5.789069e-09, 6.013745e-10, 8.833742e-10, 
    9.71731e-11, 3.073705e-12, 1.070325e-11, 2.375044e-11, 2.896086e-08, 
    1.985492e-07, 1.726832e-07, 1.351667e-07, 1.324424e-07, 8.350031e-06,
  4.835067e-07, 2.586778e-07, 7.571767e-08, 5.232696e-09, 1.049702e-06, 
    5.011174e-09, 8.945903e-10, 1.91615e-17, 2.980075e-14, 6.143022e-10, 
    1.284055e-08, 2.766698e-08, 1.106836e-07, 1.21177e-06, 6.109765e-06,
  1.872369e-06, 1.518791e-06, 1.516222e-06, 1.176895e-06, 8.735764e-07, 
    3.649048e-08, 7.898231e-09, 2.202276e-12, 6.500668e-17, 9.676312e-10, 
    1.133178e-08, 1.729567e-08, 1.209416e-08, 5.331913e-07, 1.760379e-06,
  2.889149e-09, 2.220661e-08, 6.013693e-08, 8.804513e-08, 1.163408e-07, 
    8.48401e-08, 3.438346e-09, 2.3024e-09, 2.48666e-08, 4.805818e-06, 
    6.376702e-05, 0.0001363806, 0.0001052954, 2.240423e-05, 1.036906e-07,
  5.327556e-09, 5.748729e-09, 4.784202e-08, 8.258084e-08, 1.314187e-07, 
    8.28442e-08, 3.634498e-08, 1.416565e-08, 1.238292e-08, 5.565595e-06, 
    8.289474e-05, 0.0001431292, 6.664531e-05, 5.767186e-06, 2.198005e-08,
  9.69244e-08, 5.988467e-09, 3.569939e-08, 7.186716e-08, 1.94044e-07, 
    1.4662e-07, 6.278213e-08, 2.462401e-08, 5.048717e-09, 5.155364e-06, 
    8.524599e-05, 0.0001296605, 4.630198e-05, 2.371323e-06, 4.163315e-09,
  1.996244e-06, 3.902425e-07, 7.50995e-09, 4.154733e-08, 1.991159e-07, 
    2.534774e-07, 1.380883e-07, 4.200274e-08, 3.201803e-08, 3.785443e-06, 
    7.012185e-05, 9.389698e-05, 2.790275e-05, 1.009864e-06, 1.875778e-08,
  1.213207e-06, 4.886768e-07, 6.231053e-08, 6.95116e-09, 7.005524e-08, 
    5.351716e-08, 4.232705e-08, 5.758675e-08, 2.153552e-06, 4.06456e-06, 
    5.173386e-05, 5.788342e-05, 1.577264e-05, 4.511652e-07, 6.83177e-08,
  5.408404e-06, 1.493229e-06, 4.939149e-08, 4.027622e-09, 7.420405e-09, 
    7.86988e-09, 6.940978e-09, 1.842387e-06, 2.580541e-06, 4.715679e-06, 
    2.849049e-05, 3.301044e-05, 6.655295e-06, 1.270816e-07, 2.461641e-08,
  1.46639e-05, 1.29602e-05, 4.68201e-06, 1.471383e-06, 2.066184e-07, 
    3.04365e-08, 4.536779e-09, 6.094342e-07, 6.238952e-07, 1.807622e-06, 
    2.131698e-05, 2.327898e-05, 3.196461e-06, 1.36976e-07, 1.110013e-07,
  8.945484e-06, 7.767259e-06, 7.744926e-06, 4.477903e-06, 5.588755e-08, 
    1.652907e-07, 8.210272e-09, 2.64287e-08, 2.266778e-08, 2.09752e-07, 
    9.608388e-06, 1.765842e-05, 4.962464e-06, 1.063414e-07, 1.216576e-07,
  5.748304e-06, 4.944688e-06, 1.093839e-05, 2.265632e-05, 2.528847e-05, 
    1.588056e-06, 7.302526e-08, 6.056714e-08, 2.06722e-09, 2.546245e-06, 
    1.14447e-05, 1.669019e-05, 5.932648e-06, 5.901942e-08, 2.936959e-08,
  2.235745e-06, 4.851554e-06, 1.19737e-05, 3.199618e-05, 1.857871e-05, 
    4.715231e-06, 3.235102e-07, 2.971417e-08, 1.688736e-06, 3.655824e-06, 
    8.931327e-06, 1.521852e-05, 7.1395e-06, 5.370756e-07, 1.479933e-07,
  2.515657e-23, 2.401885e-11, 3.447248e-09, 7.155606e-09, 2.052405e-08, 
    1.588974e-07, 2.208519e-07, 3.70994e-08, 2.192343e-09, 5.428666e-10, 
    1.064536e-09, 2.039662e-05, 8.113735e-05, 7.769471e-05, 3.41317e-05,
  3.681845e-16, 2.68139e-10, 8.2454e-10, 2.744834e-09, 1.260441e-08, 
    8.769647e-08, 4.932397e-08, 6.980755e-08, 1.911718e-08, 3.295728e-09, 
    2.530836e-07, 4.336722e-05, 0.0001352712, 0.0001106581, 5.320991e-05,
  1.021366e-25, 1.798703e-11, 1.339089e-11, 1.916826e-09, 2.507054e-07, 
    1.057871e-06, 1.011925e-06, 6.825618e-07, 2.642675e-07, 5.919714e-09, 
    1.812289e-06, 6.029248e-05, 0.0001620568, 0.0001375179, 6.953823e-05,
  6.191474e-18, 3.20334e-14, 4.706802e-12, 2.138407e-09, 2.768934e-08, 
    6.558534e-07, 3.179114e-06, 2.896546e-06, 9.092566e-07, 1.892455e-07, 
    3.527998e-06, 7.417973e-05, 0.0001601915, 0.0001366634, 8.01239e-05,
  1.479084e-11, 4.28368e-10, 6.378208e-11, 1.424052e-09, 1.409561e-09, 
    1.282369e-07, 2.877908e-06, 3.806823e-06, 1.947707e-06, 1.11923e-06, 
    4.894505e-06, 7.469275e-05, 0.0001383709, 0.0001237741, 8.513974e-05,
  5.288321e-10, 9.144172e-07, 4.589435e-07, 4.076401e-07, 1.2276e-09, 
    2.402264e-09, 8.547959e-09, 1.588398e-06, 2.712909e-06, 3.209112e-06, 
    6.145875e-06, 7.35844e-05, 0.0001230853, 0.0001157236, 7.849149e-05,
  8.336001e-11, 1.31606e-06, 1.505043e-06, 1.082694e-06, 1.532548e-07, 
    5.914323e-08, 9.71126e-10, 3.77841e-09, 1.077502e-08, 1.135987e-08, 
    1.888947e-06, 5.085875e-05, 0.0001115665, 0.0001152758, 6.792563e-05,
  1.246536e-11, 4.791874e-10, 1.906849e-07, 2.520044e-06, 1.907186e-06, 
    3.835655e-07, 3.26892e-08, 6.123447e-09, 6.135135e-09, 7.31566e-09, 
    6.923875e-07, 2.663738e-05, 0.0001000231, 0.0001123073, 5.856966e-05,
  4.959975e-12, 9.688324e-12, 3.759716e-10, 3.514683e-06, 6.476444e-06, 
    1.058545e-06, 2.587828e-08, 3.913723e-09, 5.573729e-09, 6.187218e-09, 
    5.094992e-07, 1.295072e-05, 8.856503e-05, 0.0001237767, 6.170003e-05,
  2.421375e-11, 2.854294e-12, 6.287257e-11, 1.283605e-06, 8.815343e-06, 
    3.695803e-06, 4.861789e-07, 3.702566e-08, 3.222627e-07, 4.529251e-07, 
    2.199994e-07, 1.079765e-05, 7.341215e-05, 0.0001411475, 6.617482e-05,
  7.990173e-05, 9.900503e-05, 9.39555e-05, 7.242689e-05, 8.270823e-05, 
    9.621344e-05, 5.636574e-05, 1.592345e-07, 3.720699e-09, 1.301642e-09, 
    1.248373e-07, 3.753344e-06, 2.524075e-06, 1.096153e-06, 1.297919e-06,
  7.52223e-05, 8.906376e-05, 9.773466e-05, 8.829706e-05, 8.726716e-05, 
    9.829419e-05, 7.05419e-05, 1.186932e-06, 1.46146e-09, 7.069479e-08, 
    4.274318e-06, 4.091152e-06, 5.438638e-07, 6.133074e-07, 1.071129e-06,
  6.790848e-05, 8.457487e-05, 8.302324e-05, 8.944325e-05, 9.042528e-05, 
    9.598851e-05, 7.442669e-05, 8.51315e-06, 1.592268e-06, 5.621946e-06, 
    4.833047e-06, 2.783807e-06, 1.080915e-06, 8.032783e-07, 1.188178e-06,
  4.91953e-05, 5.952091e-05, 6.132577e-05, 7.96692e-05, 8.363745e-05, 
    9.099156e-05, 7.812669e-05, 2.218387e-05, 4.978122e-06, 5.13192e-06, 
    3.505211e-06, 3.046659e-06, 2.279957e-07, 1.091504e-06, 9.097794e-07,
  2.527403e-05, 3.145232e-05, 5.149584e-05, 6.482293e-05, 6.841529e-05, 
    8.929556e-05, 7.848936e-05, 3.608892e-05, 7.788791e-06, 4.410795e-06, 
    3.979137e-06, 1.71332e-06, 4.431582e-08, 5.390361e-07, 1.935527e-06,
  1.664197e-05, 2.288135e-05, 2.671196e-05, 4.531992e-05, 5.027961e-05, 
    7.445969e-05, 7.961417e-05, 4.319378e-05, 6.685941e-06, 5.010887e-06, 
    2.591881e-06, 1.097431e-06, 3.723449e-07, 2.920138e-07, 2.199333e-06,
  2.773876e-06, 2.237967e-05, 5.353654e-05, 5.456245e-05, 3.72947e-05, 
    6.672544e-05, 6.029314e-05, 2.875765e-05, 2.511214e-06, 1.18072e-06, 
    5.42754e-07, 4.643301e-07, 8.639193e-07, 2.695129e-06, 1.884401e-06,
  7.158261e-05, 8.535666e-05, 8.095039e-05, 6.649656e-05, 4.224783e-05, 
    2.727098e-05, 3.222217e-05, 1.857713e-05, 2.508757e-06, 1.213514e-06, 
    9.620329e-07, 5.403898e-07, 1.114249e-06, 1.480186e-06, 2.255448e-06,
  8.260334e-05, 0.0001051447, 0.0001072662, 7.149576e-05, 6.389913e-05, 
    3.088179e-05, 5.414504e-06, 2.750472e-07, 4.142715e-07, 1.266041e-06, 
    1.127694e-06, 1.127709e-06, 1.280651e-06, 7.142955e-07, 4.934841e-06,
  4.831149e-05, 7.761307e-05, 9.379701e-05, 6.969547e-05, 6.143976e-05, 
    4.03449e-05, 1.934265e-05, 2.834566e-07, 3.508751e-06, 4.322827e-06, 
    8.909605e-06, 6.884782e-06, 2.66108e-06, 1.886019e-06, 7.156136e-06,
  1.160755e-06, 8.62806e-07, 6.514603e-08, 2.069692e-07, 7.374469e-07, 
    1.122261e-05, 0.0001275235, 0.0001460659, 0.000128167, 0.0001275138, 
    0.0001372422, 0.0001593615, 0.0001282639, 9.945404e-05, 6.253514e-05,
  1.008967e-06, 8.450791e-07, 4.947433e-07, 9.619978e-08, 3.991574e-07, 
    5.759061e-06, 8.77507e-05, 0.000154926, 0.0001442576, 0.000161882, 
    0.0001963387, 0.0001931342, 0.0001511743, 0.0001111061, 7.369364e-05,
  1.374364e-06, 2.517226e-07, 2.083686e-07, 1.127904e-07, 3.780038e-07, 
    4.009446e-06, 6.624989e-05, 0.0001635207, 0.000174284, 0.0002034764, 
    0.0002317094, 0.0002162562, 0.000159795, 0.0001069237, 6.433162e-05,
  4.506256e-06, 3.662903e-07, 4.696444e-09, 2.408666e-06, 5.244419e-06, 
    7.441234e-06, 4.799917e-05, 0.0001688507, 0.0002025036, 0.0002072438, 
    0.0002329298, 0.0002213996, 0.0001572119, 9.806483e-05, 5.959443e-05,
  4.000395e-06, 2.384614e-06, 5.851622e-07, 7.716694e-06, 1.651027e-05, 
    1.576652e-05, 4.524081e-05, 0.0001493605, 0.0002062939, 0.0002060155, 
    0.0002302901, 0.000223582, 0.00015659, 9.830783e-05, 6.038584e-05,
  1.098529e-05, 7.607495e-06, 5.164268e-06, 4.55968e-06, 1.119697e-05, 
    9.453628e-06, 4.697163e-05, 0.0001664997, 0.0002059905, 0.0002214527, 
    0.000209601, 0.0001937271, 0.0001525041, 8.670636e-05, 6.120848e-05,
  1.220684e-05, 1.117334e-05, 9.95521e-06, 4.64075e-06, 9.221512e-06, 
    1.528932e-05, 5.027635e-05, 0.0001627366, 0.0002130056, 0.0001483438, 
    0.0001741729, 0.0001630367, 0.0001374189, 0.0001145498, 5.845048e-05,
  1.151761e-05, 7.42983e-06, 6.626578e-06, 1.043256e-05, 8.680288e-06, 
    2.129658e-05, 5.777091e-05, 0.0001465078, 0.0001910971, 9.175841e-05, 
    0.0001254359, 0.000138192, 0.0001398833, 0.0001055659, 5.600874e-05,
  1.740243e-05, 1.859653e-05, 1.877368e-05, 2.356111e-05, 3.438123e-05, 
    1.383331e-05, 1.659481e-05, 1.468703e-05, 7.185728e-05, 0.0001490029, 
    0.0001403213, 0.0001218919, 0.000121439, 0.0001226053, 3.763396e-05,
  2.738615e-05, 3.296262e-05, 3.41811e-05, 2.706642e-05, 3.089075e-05, 
    1.200014e-05, 2.957396e-05, 3.112022e-05, 0.0001252168, 0.0001857189, 
    0.0001736688, 0.0001448616, 0.0001469863, 0.0001406038, 3.117679e-05,
  3.07183e-08, 7.787297e-08, 2.81555e-07, 6.253236e-09, 3.441189e-08, 
    5.29303e-08, 1.794785e-08, 6.834133e-09, 4.216918e-09, 3.284784e-08, 
    4.703709e-07, 1.068632e-06, 1.205765e-05, 3.049441e-05, 2.748089e-05,
  1.334893e-06, 4.879479e-07, 2.817396e-07, 2.893806e-07, 9.885001e-08, 
    9.863258e-08, 7.801911e-08, 1.559277e-08, 3.214643e-08, 1.351618e-08, 
    8.600029e-07, 3.22272e-06, 2.192849e-05, 4.209559e-05, 3.640841e-05,
  4.079142e-06, 1.161782e-06, 2.080191e-08, 1.331859e-06, 2.109849e-06, 
    1.192541e-07, 2.978773e-08, 2.559039e-08, 1.731211e-08, 7.875327e-08, 
    1.767558e-06, 1.001677e-05, 3.452824e-05, 5.099986e-05, 3.810322e-05,
  9.808816e-06, 3.949935e-06, 1.270496e-07, 4.520839e-06, 7.56378e-06, 
    8.414054e-07, 5.228072e-07, 2.314209e-06, 3.508107e-07, 3.752668e-07, 
    6.018264e-06, 2.289798e-05, 4.570146e-05, 5.57854e-05, 4.12718e-05,
  5.70043e-06, 2.849503e-06, 3.521385e-07, 8.148734e-06, 7.565208e-06, 
    3.974645e-06, 2.213685e-06, 3.606237e-06, 2.464955e-06, 3.885678e-06, 
    1.209753e-05, 3.077432e-05, 5.063242e-05, 5.889926e-05, 5.211353e-05,
  4.253606e-06, 1.450471e-06, 2.008194e-06, 7.272356e-06, 5.483394e-06, 
    4.726885e-06, 3.944996e-06, 5.775116e-06, 3.633845e-06, 6.264342e-06, 
    2.039924e-05, 3.924253e-05, 4.72684e-05, 5.843019e-05, 5.800518e-05,
  5.012186e-07, 1.851852e-06, 4.837872e-06, 7.750895e-06, 4.00029e-06, 
    7.680826e-07, 6.114995e-08, 5.913711e-08, 2.498266e-07, 5.885941e-06, 
    2.707456e-05, 4.872038e-05, 4.81793e-05, 6.023602e-05, 6.056144e-05,
  3.056724e-06, 3.555257e-06, 6.361799e-06, 1.260289e-05, 3.482661e-06, 
    2.964489e-07, 5.970053e-08, 1.723689e-08, 2.86708e-09, 2.099e-06, 
    2.391334e-05, 5.141395e-05, 5.275589e-05, 7.065425e-05, 6.559415e-05,
  9.73082e-06, 5.902416e-06, 7.80707e-06, 9.494031e-06, 4.163393e-06, 
    9.927292e-08, 2.783966e-09, 1.828267e-08, 1.089459e-07, 2.649005e-06, 
    2.645768e-05, 6.037299e-05, 6.167075e-05, 8.925972e-05, 7.375453e-05,
  1.298354e-05, 6.860695e-06, 1.686533e-05, 3.9109e-06, 5.259223e-07, 
    4.161317e-07, 1.30422e-08, 2.08158e-08, 2.904063e-07, 4.471643e-06, 
    3.113777e-05, 6.542588e-05, 7.332391e-05, 0.0001042987, 8.82522e-05,
  3.990743e-06, 1.565155e-06, 2.578586e-06, 6.473103e-08, 2.060461e-08, 
    1.085339e-07, 1.712002e-07, 2.163532e-07, 1.582096e-07, 2.14299e-08, 
    6.581332e-10, 1.515789e-12, 1.927758e-10, 2.097973e-12, 9.13929e-24,
  1.412267e-06, 7.828446e-07, 5.007151e-07, 2.75376e-08, 1.441671e-08, 
    7.427705e-08, 9.36769e-08, 2.64987e-07, 1.569516e-07, 5.249685e-08, 
    1.204754e-09, 1.007859e-12, 2.895746e-11, 2.535563e-12, 2.148218e-18,
  5.470338e-06, 4.235246e-07, 1.225181e-07, 6.008266e-07, 4.831977e-07, 
    5.912462e-08, 6.542871e-08, 1.857333e-07, 9.00027e-08, 3.024179e-08, 
    7.369691e-09, 2.407448e-12, 7.477576e-09, 5.081283e-11, 2.974232e-24,
  7.754385e-07, 6.260436e-07, 1.788923e-08, 3.340248e-06, 1.778501e-06, 
    2.580367e-06, 2.196568e-06, 5.256002e-07, 1.9819e-07, 2.607335e-08, 
    1.670117e-08, 8.971011e-08, 3.194206e-08, 2.684211e-09, 1.743044e-14,
  6.308402e-07, 3.344794e-07, 3.622974e-08, 2.622477e-06, 2.870545e-06, 
    1.126871e-05, 1.19206e-05, 4.333604e-06, 1.635064e-06, 2.87051e-07, 
    7.468754e-08, 1.700525e-07, 1.426315e-07, 6.061624e-08, 2.478324e-10,
  3.714439e-06, 2.368117e-07, 7.487782e-10, 2.294082e-06, 5.177869e-06, 
    1.176733e-05, 2.183996e-05, 1.684296e-05, 7.156269e-06, 4.233517e-06, 
    9.852234e-07, 7.322225e-07, 1.09588e-07, 7.32149e-08, 2.620748e-10,
  4.677764e-06, 2.550226e-06, 5.16212e-06, 6.152791e-06, 1.542646e-05, 
    1.628028e-05, 1.150144e-05, 2.001806e-06, 3.652288e-06, 8.149007e-06, 
    4.78173e-06, 1.2781e-06, 2.403771e-08, 1.439726e-08, 2.891694e-10,
  1.676948e-05, 1.137604e-05, 1.243986e-05, 1.408017e-05, 2.397595e-05, 
    1.426976e-05, 1.250891e-05, 4.148374e-06, 2.876192e-06, 2.77993e-06, 
    8.135047e-06, 2.901592e-06, 6.036167e-07, 6.416356e-08, 1.186207e-09,
  2.293508e-05, 1.817253e-05, 1.837585e-05, 2.617197e-05, 6.894863e-05, 
    3.190364e-05, 7.816683e-06, 5.939996e-06, 9.614219e-06, 1.061233e-05, 
    1.11883e-05, 5.20694e-06, 3.169984e-06, 3.870967e-07, 2.148473e-08,
  2.551281e-05, 2.750738e-05, 2.583194e-05, 3.739461e-05, 5.165442e-05, 
    2.542758e-05, 1.763205e-05, 1.59722e-05, 2.112279e-05, 1.6426e-05, 
    1.286184e-05, 6.606557e-06, 4.597981e-06, 1.380563e-06, 8.00495e-08,
  6.874086e-06, 7.778014e-06, 1.625865e-05, 4.337023e-05, 0.0001347576, 
    0.0002782065, 0.0004039461, 0.0004816241, 0.0004817164, 0.0002895844, 
    1.191224e-05, 1.430307e-06, 3.772322e-07, 1.548861e-06, 1.792491e-06,
  3.837943e-06, 2.034821e-06, 1.040585e-05, 4.514029e-05, 0.00011017, 
    0.0002346767, 0.0003334992, 0.0004689313, 0.000477983, 0.0002651274, 
    1.336868e-05, 1.411049e-06, 9.230041e-07, 9.460879e-07, 7.079639e-07,
  5.028433e-06, 3.478428e-06, 6.609606e-06, 3.160526e-05, 8.775621e-05, 
    0.0001740977, 0.0002749712, 0.000367679, 0.0004255597, 0.0002563531, 
    2.118599e-05, 2.552398e-06, 7.704779e-07, 3.642592e-07, 2.379085e-07,
  3.960163e-06, 2.76689e-06, 2.906972e-06, 1.930877e-05, 5.669686e-05, 
    0.0001122425, 0.0001785467, 0.000213308, 0.0003127192, 0.000235017, 
    3.812669e-05, 2.838148e-06, 5.642596e-07, 1.500888e-07, 1.266907e-07,
  1.752927e-06, 9.731413e-07, 1.779249e-06, 1.20925e-05, 2.852099e-05, 
    5.286307e-05, 0.0001065261, 0.0001023323, 0.0001623842, 0.0001821329, 
    5.005146e-05, 7.888531e-06, 2.042276e-06, 5.654646e-07, 1.734849e-07,
  1.186688e-06, 3.514292e-07, 1.83868e-07, 4.734389e-06, 1.034292e-05, 
    2.297318e-05, 6.975188e-05, 8.735251e-05, 6.080875e-05, 0.0001181868, 
    4.546244e-05, 8.926273e-06, 3.34315e-06, 1.473349e-06, 4.397058e-07,
  1.345827e-06, 8.212962e-09, 1.943174e-07, 3.416421e-06, 4.617848e-06, 
    1.090669e-05, 3.762056e-05, 5.11839e-05, 2.167547e-05, 5.232278e-05, 
    3.958426e-05, 9.402179e-06, 5.990754e-06, 3.066376e-06, 1.496772e-06,
  6.938834e-06, 1.174297e-06, 1.546264e-06, 3.193885e-06, 4.147447e-06, 
    3.357565e-06, 2.778455e-05, 7.189801e-05, 3.327333e-05, 9.027024e-06, 
    1.961742e-05, 6.39069e-06, 8.502243e-06, 6.10709e-06, 3.696379e-06,
  1.56788e-05, 5.118236e-06, 4.973168e-06, 3.70316e-06, 7.827794e-06, 
    2.961193e-06, 2.159537e-06, 3.185474e-05, 3.510903e-05, 1.384496e-06, 
    6.549008e-06, 4.650287e-06, 3.85163e-06, 4.838066e-06, 4.375756e-06,
  2.268249e-05, 1.156458e-05, 8.494951e-06, 9.177012e-06, 3.209227e-06, 
    1.701214e-06, 1.793742e-06, 1.368542e-05, 3.113355e-05, 1.275304e-06, 
    3.342842e-07, 1.913079e-06, 2.35633e-06, 3.959359e-07, 3.037295e-06,
  8.373506e-10, 6.374135e-08, 4.484002e-07, 1.931907e-06, 8.487043e-06, 
    2.979133e-05, 3.669789e-05, 4.599763e-05, 5.773357e-05, 7.599705e-05, 
    5.902491e-05, 5.078368e-05, 0.0001516133, 0.00013614, 7.445648e-05,
  5.461776e-10, 7.571538e-10, 2.009518e-07, 1.555518e-06, 2.092038e-05, 
    6.260693e-05, 8.499423e-05, 0.0001656513, 0.0001958279, 0.000165065, 
    7.93179e-05, 9.89531e-05, 0.0001127996, 0.0001331438, 0.0001056451,
  3.689878e-10, 1.370208e-09, 5.747244e-08, 5.984402e-06, 4.39822e-05, 
    9.123144e-05, 0.0001211105, 0.0002806157, 0.0003566824, 0.000284615, 
    0.0002086889, 7.027918e-05, 0.0001116924, 0.0001469531, 0.0001248033,
  2.268261e-10, 5.666368e-09, 2.002703e-08, 8.092285e-06, 6.211866e-05, 
    0.0001029302, 0.0001353305, 0.0002742639, 0.0004825295, 0.0004541402, 
    0.0001820785, 7.411493e-05, 0.0001150038, 0.0001539328, 0.0001317236,
  4.822736e-10, 4.174145e-09, 1.358458e-08, 8.109615e-06, 6.63546e-05, 
    0.0001105059, 0.0001390308, 0.0002318953, 0.0005318869, 0.0005593466, 
    0.0003118437, 9.432103e-05, 0.000115846, 0.0001586918, 0.0001437108,
  4.537532e-08, 4.499556e-08, 1.925526e-08, 1.808053e-05, 8.473967e-05, 
    0.000101583, 0.0001536215, 0.0002456576, 0.0005192577, 0.0006121449, 
    0.0003715666, 0.0001014463, 9.489266e-05, 0.0001485435, 0.0001434564,
  4.480876e-06, 2.819159e-06, 3.337905e-07, 1.51932e-05, 9.059097e-05, 
    9.432552e-05, 0.0001338967, 0.0001967008, 0.0004245833, 0.0006264551, 
    0.0004303858, 0.0001148183, 7.921619e-05, 0.0001410163, 0.0001367263,
  3.331009e-06, 3.855886e-06, 1.961906e-06, 8.885438e-06, 7.930599e-05, 
    9.225982e-05, 0.0001529959, 0.000236438, 0.0003822353, 0.0006116214, 
    0.000504034, 0.0001718359, 6.989998e-05, 0.0001254836, 0.0001293417,
  4.20199e-06, 4.146067e-06, 2.816705e-06, 1.244922e-05, 6.303978e-05, 
    8.130291e-05, 0.0001256683, 0.0002363845, 0.0003684941, 0.00054467, 
    0.0005646339, 0.0002179783, 8.446038e-05, 0.000117254, 0.0001185175,
  4.600477e-06, 4.935132e-06, 4.155361e-06, 1.370301e-05, 4.456438e-05, 
    7.622101e-05, 0.000109445, 0.0001999953, 0.0002858963, 0.0004710799, 
    0.0005680522, 0.0003001647, 7.295683e-05, 0.0001351052, 0.0001059519,
  5.614599e-12, 6.02954e-13, 6.949515e-13, 1.110132e-13, 1.939015e-24, 
    1.402806e-16, 9.975798e-15, 7.879593e-18, 2.725905e-17, 5.560406e-11, 
    1.092002e-09, 1.878344e-10, 6.388715e-11, 2.581493e-07, 2.420175e-06,
  2.407764e-12, 2.090037e-17, 7.063157e-29, 2.007753e-27, 9.103464e-26, 
    3.321302e-17, 1.088298e-12, 6.148438e-17, 1.312601e-16, 4.328371e-13, 
    1.716546e-10, 3.410088e-10, 8.1153e-11, 1.338503e-07, 5.619098e-07,
  1.244678e-12, 7.818036e-28, 0, 2.007602e-29, 2.340269e-27, 1.432254e-25, 
    5.953447e-13, 1.127395e-12, 9.397068e-10, 7.13037e-11, 1.030847e-09, 
    1.43028e-10, 2.279791e-10, 1.496749e-09, 4.313768e-09,
  7.281035e-11, 6.400869e-27, 1.821962e-29, 0, 3.828826e-14, 2.425309e-10, 
    6.033908e-11, 2.259872e-09, 7.173652e-08, 1.828747e-07, 1.51042e-07, 
    6.540753e-11, 6.165523e-09, 8.178329e-10, 5.126728e-09,
  1.45041e-10, 1.760852e-12, 1.372857e-26, 7.68095e-11, 5.249782e-12, 
    1.846524e-07, 3.962232e-08, 9.912301e-08, 3.475637e-07, 2.014061e-07, 
    1.671951e-07, 2.104216e-09, 7.165164e-09, 1.011525e-09, 1.785183e-09,
  4.748229e-10, 4.016572e-11, 1.714678e-14, 1.523634e-11, 3.192226e-07, 
    2.978231e-07, 5.811969e-07, 1.58786e-07, 4.901784e-07, 6.723517e-07, 
    3.75274e-07, 2.844344e-08, 2.377335e-08, 9.107281e-10, 2.733453e-09,
  1.084657e-09, 7.229651e-10, 9.407043e-10, 5.391541e-09, 3.665784e-09, 
    2.030661e-07, 6.383729e-10, 7.797968e-09, 9.656235e-08, 1.808912e-08, 
    3.205935e-08, 5.49164e-09, 2.485048e-08, 1.886381e-09, 6.177667e-08,
  6.033675e-08, 1.998225e-07, 1.582366e-07, 3.324474e-09, 4.197486e-10, 
    1.475702e-08, 6.321212e-09, 2.451645e-10, 3.388131e-09, 2.173755e-10, 
    1.085689e-10, 8.273375e-11, 4.70433e-09, 3.558102e-08, 1.580784e-07,
  1.052371e-07, 1.641022e-07, 4.209288e-07, 3.81603e-07, 7.08765e-07, 
    1.354333e-07, 4.850578e-13, 1.363945e-08, 3.374697e-11, 2.626446e-12, 
    5.322542e-09, 3.074926e-08, 3.990015e-08, 2.678595e-08, 4.870857e-07,
  4.197923e-07, 7.439664e-07, 1.007205e-06, 7.501516e-07, 3.003846e-07, 
    5.161502e-08, 2.945491e-09, 7.072398e-16, 1.435967e-07, 5.13948e-07, 
    1.882212e-07, 5.398701e-08, 1.056595e-07, 2.181163e-07, 1.557378e-06,
  4.123711e-05, 4.011603e-05, 3.349323e-05, 2.06573e-05, 2.512849e-05, 
    3.423235e-05, 2.215815e-05, 5.690913e-06, 6.528585e-07, 1.369919e-06, 
    7.052355e-07, 4.031425e-07, 2.979926e-07, 2.339783e-07, 3.087958e-07,
  2.55396e-05, 3.061712e-05, 2.022706e-05, 7.039868e-06, 2.920115e-06, 
    6.452414e-06, 1.024219e-05, 4.172386e-06, 6.460012e-07, 1.313956e-06, 
    1.657314e-07, 8.92743e-08, 1.042474e-07, 5.803909e-07, 2.124792e-07,
  1.43283e-05, 1.959461e-05, 9.968941e-06, 2.304679e-06, 1.219733e-06, 
    3.828594e-07, 9.4431e-07, 2.038499e-06, 9.706388e-07, 1.84697e-06, 
    1.15615e-07, 8.421508e-08, 1.742412e-07, 4.025776e-07, 4.594361e-07,
  9.052882e-06, 1.046987e-05, 2.297877e-06, 1.358179e-06, 1.300007e-06, 
    3.378428e-07, 8.074505e-07, 8.143422e-07, 1.629433e-06, 1.92906e-06, 
    3.911562e-07, 1.747772e-08, 9.802913e-08, 8.743213e-08, 1.708219e-07,
  5.900239e-06, 6.191576e-06, 4.637929e-06, 1.56539e-06, 7.729518e-07, 
    6.371714e-07, 1.908516e-06, 1.384415e-06, 1.694453e-06, 9.905306e-07, 
    1.650522e-07, 5.007929e-09, 2.895892e-09, 1.429089e-08, 4.253584e-09,
  4.466926e-06, 5.933601e-06, 2.875373e-06, 2.990287e-06, 1.407128e-06, 
    5.090189e-07, 5.725836e-07, 1.817494e-06, 1.65591e-07, 8.482888e-07, 
    1.872707e-07, 2.34372e-08, 1.506882e-09, 3.04727e-09, 6.871567e-10,
  5.325043e-07, 2.914725e-06, 3.097916e-06, 2.811072e-06, 2.16131e-06, 
    7.718525e-07, 2.608716e-07, 7.915621e-08, 1.644173e-07, 3.243265e-07, 
    8.297277e-08, 1.018067e-07, 1.811905e-09, 9.00175e-10, 1.974832e-09,
  1.30011e-07, 7.064467e-07, 1.067745e-06, 1.211019e-06, 8.984879e-07, 
    5.49303e-07, 6.679874e-07, 7.098655e-07, 1.21283e-07, 1.615753e-08, 
    5.718922e-08, 8.036162e-08, 1.18549e-09, 1.603609e-09, 4.255077e-09,
  1.240374e-09, 2.860733e-09, 7.174264e-09, 1.735824e-08, 3.363479e-07, 
    1.675455e-07, 9.943766e-08, 2.468727e-08, 3.29076e-08, 3.309288e-09, 
    1.857807e-08, 1.675689e-08, 2.117725e-09, 4.517671e-09, 7.261382e-09,
  2.488178e-09, 1.41389e-09, 1.021012e-09, 5.139338e-09, 6.62411e-09, 
    1.122992e-08, 4.723399e-08, 6.404925e-09, 2.085606e-09, 1.440736e-09, 
    5.795214e-10, 6.680564e-10, 3.937272e-10, 8.31629e-11, 1.920513e-10,
  0.0001686022, 0.000235492, 0.000283989, 0.0002473209, 0.0001414832, 
    7.905412e-05, 2.963732e-05, 5.303784e-07, 6.357585e-08, 9.252317e-08, 
    1.874743e-07, 1.443293e-06, 5.849652e-06, 6.217131e-06, 2.900852e-06,
  0.0002101845, 0.0002993874, 0.0003566798, 0.0002967958, 0.0002021578, 
    0.0001132093, 5.528316e-05, 4.472938e-06, 4.333877e-07, 7.251241e-07, 
    1.461936e-06, 7.541898e-06, 1.11099e-05, 8.894116e-06, 7.715922e-06,
  0.0002410323, 0.0003660592, 0.0004073863, 0.0003465756, 0.0002513139, 
    0.0001680667, 6.957688e-05, 6.427123e-06, 1.141703e-06, 1.358643e-06, 
    9.588152e-06, 1.006883e-05, 1.13313e-05, 9.654274e-06, 5.951091e-06,
  0.0002097298, 0.0003377398, 0.000381686, 0.0003784327, 0.0002720438, 
    0.0001989157, 9.027788e-05, 1.352629e-05, 4.166047e-06, 1.045314e-05, 
    1.312508e-05, 1.15175e-05, 1.24729e-05, 8.303468e-06, 7.00051e-06,
  0.0001228473, 0.0002587283, 0.0003588995, 0.0003761421, 0.0003003662, 
    0.0002243248, 0.0001293977, 2.240448e-05, 1.437188e-05, 1.798928e-05, 
    1.315095e-05, 6.487568e-06, 7.38855e-06, 9.498699e-06, 4.830114e-06,
  0.000107351, 0.0001909719, 0.0002553695, 0.0003668124, 0.0003309058, 
    0.0002668813, 0.0001793297, 4.459721e-05, 1.065062e-05, 1.673615e-05, 
    9.590108e-06, 3.774841e-06, 5.640047e-06, 4.85459e-06, 3.53385e-06,
  6.754456e-05, 0.0001146502, 0.0002632958, 0.0003560208, 0.000291771, 
    0.0003336958, 0.0002172967, 6.221575e-05, 1.735231e-06, 7.287068e-06, 
    9.672161e-06, 4.658378e-06, 3.366452e-06, 3.700733e-06, 4.121682e-06,
  0.0002444054, 0.0002110149, 0.0002681322, 0.000332691, 0.0002741189, 
    0.000233349, 0.0002256626, 0.0001132844, 1.113635e-05, 4.285328e-06, 
    1.033437e-05, 6.627064e-06, 2.375287e-06, 2.726332e-06, 2.655837e-06,
  0.0003705067, 0.0002844318, 0.0001948438, 0.0002366401, 0.0003274529, 
    0.0002490369, 0.0001579756, 1.792798e-05, 1.233819e-05, 1.357962e-05, 
    1.724038e-05, 1.007447e-05, 2.195654e-06, 1.498943e-06, 8.799321e-07,
  0.000360149, 0.0002772471, 0.0001796411, 0.0001679821, 0.0002777123, 
    0.0002406865, 0.0002535612, 7.520193e-05, 2.213668e-05, 1.215638e-05, 
    1.22173e-05, 8.370664e-06, 2.602887e-06, 3.043744e-06, 2.652215e-06,
  0.0001847077, 0.0001677057, 0.0001155844, 8.750146e-05, 8.202284e-05, 
    1.835798e-05, 9.758278e-06, 1.107151e-06, 1.89097e-07, 5.294543e-07, 
    8.081816e-08, 9.467595e-08, 3.032084e-06, 4.217362e-06, 1.70833e-06,
  0.0001638386, 0.0001748412, 0.000158941, 0.0001067757, 0.00013389, 
    3.788012e-05, 6.469282e-06, 1.317034e-06, 5.400631e-07, 9.956785e-07, 
    4.321025e-07, 3.92594e-07, 3.513657e-06, 2.833783e-06, 1.328023e-06,
  0.0001187851, 0.0001679805, 0.0001850404, 0.0001393602, 0.0001765097, 
    0.0001038175, 1.978986e-05, 5.674491e-06, 1.612631e-06, 1.332067e-06, 
    3.240585e-07, 1.425873e-05, 5.505432e-06, 1.738454e-06, 8.776722e-07,
  5.327899e-05, 0.0001047361, 0.0001582082, 0.0001652682, 0.0002091612, 
    0.0001718699, 4.503945e-05, 1.798268e-05, 6.371317e-06, 2.313154e-06, 
    0.0001018535, 3.324309e-05, 4.500605e-06, 3.03975e-06, 3.094153e-06,
  6.606377e-06, 3.168632e-05, 8.501224e-05, 0.0001331969, 0.0002200597, 
    0.0002341158, 7.297573e-05, 4.156097e-05, 2.351048e-05, 0.0003257599, 
    5.361744e-05, 2.254283e-05, 2.242774e-06, 1.772954e-06, 8.099624e-07,
  7.576972e-06, 7.074226e-06, 5.0781e-06, 6.01908e-05, 0.0001727067, 
    0.0002810118, 0.0001362478, 7.806753e-05, 6.637246e-05, 0.0003689254, 
    0.0001222492, 5.054394e-06, 5.245946e-07, 3.282782e-07, 9.326133e-07,
  6.788889e-06, 6.467684e-06, 1.600215e-06, 6.200553e-06, 5.065274e-05, 
    0.0003230207, 0.0002231009, 0.000141003, 0.0001044307, 6.521655e-05, 
    4.350614e-05, 7.801702e-06, 8.102133e-07, 1.005366e-07, 1.223608e-06,
  3.737272e-06, 5.567896e-06, 1.68938e-06, 2.138797e-06, 4.07939e-06, 
    0.0002612315, 0.0003229387, 0.0002352459, 0.0002105644, 0.0001019809, 
    3.706028e-05, 8.372874e-06, 1.593696e-06, 3.612087e-07, 2.996197e-06,
  9.686222e-07, 1.703792e-06, 8.898448e-07, 2.26005e-06, 3.262498e-06, 
    0.0001337878, 0.0003178387, 0.0001978729, 3.220222e-05, 8.021221e-05, 
    5.228562e-05, 3.422004e-06, 2.040553e-06, 1.627917e-07, 3.661376e-06,
  3.271816e-07, 3.505569e-07, 6.250033e-07, 2.802281e-06, 2.047903e-06, 
    2.268122e-05, 0.0003247253, 0.0003316556, 0.0001213007, 7.65908e-05, 
    0.0001256774, 1.980037e-05, 2.990287e-06, 1.00477e-06, 4.456395e-06,
  5.627605e-07, 8.055674e-06, 0.0001224026, 0.000239421, 0.0001592491, 
    1.420419e-05, 8.231817e-06, 2.264146e-05, 2.61814e-05, 5.209456e-08, 
    3.15416e-08, 4.148339e-09, 1.658938e-07, 3.090229e-06, 6.564524e-06,
  1.604559e-06, 7.467024e-07, 6.979265e-05, 0.0002471882, 0.0002192613, 
    3.849325e-05, 9.520628e-06, 3.56767e-06, 8.829208e-07, 2.019935e-07, 
    1.382956e-07, 1.094493e-08, 1.749905e-06, 5.410134e-06, 8.352898e-06,
  3.674419e-05, 1.696367e-05, 2.992552e-05, 0.0002118966, 0.0002755319, 
    0.0001620038, 1.53746e-05, 4.155602e-06, 1.258147e-06, 3.168385e-07, 
    2.252879e-07, 6.231787e-07, 4.43547e-06, 8.381018e-06, 1.030047e-05,
  9.790889e-05, 8.046848e-05, 3.631931e-05, 0.000125069, 0.0003010715, 
    0.0002382278, 3.286541e-05, 2.245516e-05, 2.188378e-06, 1.216447e-06, 
    1.184034e-06, 9.262638e-07, 4.409728e-06, 9.229925e-06, 1.425593e-05,
  0.0001152315, 0.0001344572, 0.0001115882, 7.565205e-05, 0.000245512, 
    0.0002569564, 0.0001028705, 4.541258e-05, 1.405821e-05, 0.0001137399, 
    4.651961e-05, 1.723753e-06, 2.1021e-06, 8.505568e-06, 1.214972e-05,
  8.589062e-05, 0.0001315226, 0.0001720652, 0.0001141575, 0.0001890492, 
    0.0002647946, 0.0001916798, 6.923771e-05, 7.105062e-05, 0.0002535293, 
    7.872041e-05, 8.230075e-06, 7.533239e-06, 9.337266e-06, 1.073965e-05,
  2.475387e-05, 8.190026e-05, 0.0001715057, 0.0001865847, 0.0001755729, 
    0.0002883105, 0.0002140361, 0.0001230549, 0.0001155074, 3.188071e-05, 
    3.35668e-05, 1.396435e-05, 1.02821e-05, 1.038726e-05, 9.698922e-06,
  5.022197e-06, 3.884092e-05, 0.0001534521, 0.0002263302, 0.0001965393, 
    0.0002804947, 0.0002552398, 0.0002477256, 0.0002613044, 4.640091e-05, 
    1.192626e-05, 1.264335e-05, 1.22929e-05, 1.097475e-05, 9.658123e-06,
  5.370791e-07, 1.536276e-05, 0.0001182315, 0.00021509, 0.0002481652, 
    0.0002617957, 0.000245701, 0.0001469159, 0.0001063585, 4.89476e-05, 
    7.900715e-06, 1.008208e-05, 1.592662e-05, 1.02366e-05, 9.001229e-06,
  1.443571e-08, 6.964889e-06, 0.0001032147, 0.000207202, 0.0002412164, 
    0.0002249129, 0.0002118703, 0.0001915867, 0.0001749723, 8.878719e-05, 
    9.162072e-06, 1.020197e-05, 1.359522e-05, 9.433699e-06, 8.22614e-06,
  3.565968e-08, 8.884307e-08, 8.536986e-08, 3.126274e-06, 3.870897e-05, 
    8.718445e-05, 9.424709e-05, 0.0001312644, 8.470388e-05, 4.090906e-05, 
    4.776776e-05, 3.862624e-06, 5.217307e-06, 3.361554e-08, 4.327751e-07,
  2.718547e-08, 2.957194e-08, 3.865203e-08, 2.863277e-06, 1.118744e-05, 
    4.568319e-05, 5.018755e-05, 0.0001219613, 0.0001109779, 1.457193e-05, 
    1.876426e-05, 1.36258e-05, 3.164061e-05, 1.790872e-05, 1.852729e-06,
  4.875195e-08, 3.979347e-08, 1.841947e-07, 6.543789e-06, 1.241023e-05, 
    1.858554e-05, 2.954832e-05, 7.143514e-05, 0.0001181611, 3.769554e-05, 
    1.714961e-05, 1.990547e-05, 3.068788e-05, 1.585089e-05, 8.944735e-06,
  2.908604e-08, 2.273585e-08, 2.604924e-07, 1.739924e-05, 1.253337e-05, 
    4.589174e-06, 1.59653e-05, 2.459277e-05, 0.0001015818, 7.716401e-05, 
    3.261326e-05, 2.792457e-05, 1.951209e-05, 3.770198e-05, 1.457734e-05,
  1.605281e-08, 8.575181e-09, 2.802757e-07, 1.044836e-05, 1.899278e-05, 
    7.148092e-06, 6.734937e-06, 1.139829e-05, 6.223968e-05, 8.314179e-05, 
    4.376469e-05, 3.872381e-05, 1.656623e-05, 1.974118e-05, 1.791021e-05,
  5.850939e-08, 1.104973e-07, 2.456125e-07, 6.904983e-06, 3.38278e-05, 
    1.800282e-05, 1.149698e-05, 6.88415e-06, 3.255281e-05, 8.331466e-05, 
    5.369235e-05, 3.051828e-05, 1.283269e-05, 1.888161e-05, 2.229042e-05,
  2.78216e-08, 6.930038e-08, 3.96676e-07, 2.387212e-06, 4.820214e-05, 
    5.013566e-05, 2.893158e-05, 1.107462e-05, 1.946661e-05, 4.457687e-05, 
    4.58389e-05, 2.057584e-05, 1.359651e-05, 1.743138e-05, 2.069669e-05,
  2.333848e-08, 9.836937e-08, 3.661088e-07, 1.742025e-06, 2.317907e-05, 
    9.848981e-05, 8.091607e-05, 3.97922e-05, 3.177221e-05, 3.826024e-05, 
    4.554543e-05, 2.325563e-05, 1.405266e-05, 1.603282e-05, 2.06151e-05,
  1.045102e-08, 5.90139e-08, 1.344111e-07, 1.850863e-06, 1.601066e-05, 
    0.0001231068, 0.0001246563, 8.265445e-05, 4.846043e-05, 7.755162e-05, 
    8.705e-05, 4.138277e-05, 1.621673e-05, 1.407636e-05, 1.987537e-05,
  6.815593e-08, 9.811814e-08, 8.503662e-08, 7.544836e-07, 1.594145e-06, 
    0.0001104762, 0.0001925616, 0.0001405249, 0.00010787, 7.99976e-05, 
    0.0001059583, 7.054659e-05, 2.820309e-05, 1.513413e-05, 2.01171e-05,
  2.723039e-08, 2.594204e-08, 8.034603e-08, 4.260236e-06, 2.786751e-05, 
    9.499973e-05, 0.0002009588, 0.0002593605, 0.0001575507, 0.0001253833, 
    0.0001109722, 4.939007e-05, 1.560025e-05, 1.042775e-05, 3.48317e-05,
  3.294948e-09, 9.349583e-09, 2.44617e-08, 2.230794e-06, 1.438262e-05, 
    3.342782e-05, 8.364712e-05, 0.0001938109, 0.0001641684, 0.0001415814, 
    0.0001956044, 0.0001286842, 3.511556e-05, 1.671082e-05, 1.078905e-05,
  7.589316e-08, 1.243715e-07, 3.305351e-08, 2.327343e-06, 8.065246e-06, 
    1.598824e-05, 1.580024e-05, 9.001089e-05, 0.0001687332, 0.0001335895, 
    0.0002265871, 0.0002139666, 8.721539e-05, 1.871282e-05, 1.485617e-05,
  5.929314e-08, 5.448983e-08, 1.350321e-08, 7.534404e-07, 3.086303e-06, 
    6.084867e-06, 5.929917e-06, 2.645377e-05, 0.0001171946, 0.0001476084, 
    0.0002039766, 0.0002459994, 0.0001032259, 4.848833e-05, 2.067009e-05,
  4.337554e-08, 2.672994e-08, 4.260174e-10, 6.6516e-08, 4.025596e-07, 
    1.888887e-06, 3.10958e-06, 3.538604e-06, 6.978607e-05, 0.00014358, 
    0.0001883231, 0.0002478474, 0.0001868937, 3.511246e-05, 1.836583e-05,
  2.149757e-08, 3.769745e-09, 1.265447e-10, 6.231224e-09, 9.063834e-08, 
    3.410269e-07, 1.00979e-06, 1.827476e-06, 2.369583e-05, 0.0001197279, 
    0.0001935836, 0.0002475223, 0.0002423292, 0.0001026551, 2.608963e-05,
  2.723969e-12, 5.852927e-11, 9.592931e-10, 1.758716e-09, 1.674339e-08, 
    3.118194e-08, 6.494373e-07, 1.576453e-06, 3.376908e-06, 5.945643e-05, 
    0.0001612258, 0.0002354364, 0.0002759618, 0.0001835461, 4.537606e-05,
  7.135073e-10, 3.681258e-11, 1.368681e-08, 7.453902e-09, 7.355909e-10, 
    2.553897e-09, 3.526438e-07, 1.180803e-06, 1.346957e-06, 1.88807e-05, 
    9.490963e-05, 0.0001968071, 0.0002749359, 0.0002504258, 9.289926e-05,
  3.815152e-10, 1.053043e-08, 7.750006e-09, 2.25446e-08, 5.914653e-09, 
    8.308939e-09, 3.282376e-08, 2.583207e-07, 9.316461e-07, 7.151439e-06, 
    5.233656e-05, 0.0001449461, 0.0002381292, 0.0002724803, 0.0001592533,
  5.218464e-08, 2.750914e-08, 1.643661e-07, 1.493295e-08, 6.826378e-09, 
    3.033731e-09, 2.152497e-08, 2.451818e-07, 7.609735e-07, 5.030348e-06, 
    2.739636e-05, 8.682856e-05, 0.0001904002, 0.0002816012, 0.0002234802,
  7.879868e-07, 3.846705e-07, 2.138451e-07, 3.669016e-06, 3.186126e-05, 
    6.581203e-05, 0.0001224178, 0.0001879473, 0.0002398656, 0.0002476325, 
    0.000201038, 0.0001507628, 0.0001343437, 1.418141e-05, 8.067652e-07,
  1.765809e-06, 1.096838e-06, 4.55443e-07, 9.557037e-07, 2.024467e-05, 
    5.308663e-05, 0.000132614, 0.0002203472, 0.0002822773, 0.0002786816, 
    0.0002468278, 0.0002988617, 0.0001919774, 1.320802e-05, 1.991797e-06,
  2.871425e-06, 1.843021e-06, 4.854406e-07, 7.7609e-07, 1.054726e-05, 
    3.683978e-05, 0.0001417541, 0.0002541651, 0.0002878583, 0.0003057744, 
    0.000290023, 0.0002217862, 0.000215198, 2.989344e-05, 4.18352e-06,
  2.946331e-06, 2.255867e-06, 7.040085e-07, 6.522899e-07, 6.779571e-06, 
    1.147668e-05, 0.0001209239, 0.0002603814, 0.0003059082, 0.0003165406, 
    0.0003224068, 0.0002448319, 0.0001770442, 3.314221e-05, 7.813742e-06,
  2.044315e-06, 2.037817e-06, 1.06805e-06, 4.326786e-07, 3.873663e-06, 
    7.927659e-06, 8.807827e-05, 0.0002389451, 0.0003201604, 0.0003196166, 
    0.0003605732, 0.0004351693, 0.0001504558, 5.246534e-05, 1.039461e-05,
  7.406504e-07, 1.300995e-06, 8.628871e-07, 3.609934e-07, 2.880638e-06, 
    4.015814e-06, 5.583709e-05, 0.0002131686, 0.0002973655, 0.0003199276, 
    0.0003840414, 0.0003365201, 0.0001737032, 6.227288e-05, 9.133772e-06,
  1.81068e-08, 1.828067e-07, 6.326969e-07, 2.656871e-07, 7.68003e-07, 
    5.985419e-06, 3.929462e-05, 0.0001803466, 0.0002343668, 0.0002870205, 
    0.0004021466, 0.0004565408, 0.0002059961, 7.319105e-05, 1.73862e-05,
  3.725878e-10, 3.738899e-08, 1.043971e-07, 3.514668e-07, 1.837832e-07, 
    5.229859e-06, 5.691104e-05, 0.0001940219, 0.0002186747, 0.0002837245, 
    0.0004593358, 0.000555766, 0.0002840937, 7.853109e-05, 2.779718e-05,
  1.690297e-10, 8.531187e-09, 3.335809e-07, 4.184719e-07, 2.306319e-06, 
    5.850283e-06, 1.847501e-05, 8.556158e-05, 0.0002530738, 0.0002850198, 
    0.0004940861, 0.0006456291, 0.000390528, 9.586851e-05, 3.546842e-05,
  1.653415e-10, 1.843329e-07, 7.715814e-07, 3.003648e-07, 2.060163e-06, 
    4.69782e-06, 1.259107e-05, 3.519924e-05, 0.0001954067, 0.0002211276, 
    0.0004050553, 0.0006846936, 0.000514648, 0.000132445, 4.246253e-05,
  3.927393e-08, 1.912856e-08, 1.64159e-08, 5.476691e-08, 1.259568e-07, 
    2.110042e-05, 0.0001277401, 0.0004097336, 0.0005203206, 0.0003949379, 
    0.0003010473, 0.0002015119, 9.379887e-05, 8.585596e-07, 8.724075e-08,
  4.945801e-08, 4.841179e-08, 2.22855e-08, 1.816311e-08, 2.696401e-08, 
    5.470171e-07, 4.253673e-05, 0.0002001725, 0.0004324964, 0.0003749151, 
    0.0002882179, 0.0002073233, 5.01606e-05, 1.363979e-06, 2.384352e-07,
  6.5931e-08, 4.438878e-08, 2.843078e-08, 1.930226e-08, 1.693607e-08, 
    6.564222e-08, 8.166583e-06, 9.641548e-05, 0.0002942861, 0.0003256738, 
    0.0002429903, 0.0001902036, 0.0001023504, 7.509986e-06, 4.853036e-07,
  1.254225e-07, 1.000092e-07, 6.552268e-08, 4.425873e-08, 1.202825e-08, 
    1.012115e-08, 5.357403e-07, 4.24866e-05, 0.000168776, 0.0002445267, 
    0.00016661, 0.0001470511, 0.000131209, 5.395921e-05, 4.112891e-06,
  8.139045e-08, 1.319176e-07, 1.046255e-07, 6.43635e-08, 2.93404e-08, 
    1.138529e-08, 9.52739e-09, 9.361359e-06, 8.208343e-05, 0.0001561768, 
    0.000115379, 7.179757e-05, 0.0001058621, 7.946145e-05, 2.163497e-05,
  1.04573e-08, 9.307237e-08, 1.010507e-07, 8.925801e-08, 1.489471e-08, 
    2.259455e-09, 1.079258e-07, 7.769419e-07, 3.818654e-05, 9.123934e-05, 
    9.157933e-05, 3.391762e-05, 4.14986e-05, 6.59556e-05, 3.338468e-05,
  1.608045e-09, 2.991876e-08, 1.035232e-07, 5.662072e-08, 1.319743e-08, 
    1.960892e-09, 2.107151e-09, 4.072664e-09, 8.058865e-06, 4.606626e-05, 
    6.611436e-05, 4.155317e-05, 1.6658e-05, 2.91683e-05, 2.649215e-05,
  7.890319e-07, 1.330249e-08, 5.886788e-08, 3.074874e-08, 1.302323e-08, 
    3.971833e-09, 1.296888e-09, 5.904718e-09, 4.84193e-08, 2.251532e-05, 
    5.319158e-05, 6.057668e-05, 2.651046e-05, 9.498305e-06, 8.219098e-06,
  3.297177e-07, 5.268617e-07, 2.151312e-07, 2.372862e-08, 1.556174e-07, 
    2.498248e-09, 1.666096e-09, 6.025698e-09, 7.653284e-07, 1.735348e-05, 
    4.337851e-05, 6.961363e-05, 5.475343e-05, 1.251536e-05, 4.210596e-06,
  3.996848e-08, 4.842795e-08, 1.241174e-06, 7.535007e-07, 1.071585e-07, 
    1.333214e-08, 1.315993e-08, 1.034208e-08, 1.534845e-06, 1.693959e-05, 
    4.520893e-05, 6.33222e-05, 4.790809e-05, 1.813913e-05, 8.446571e-06,
  7.413134e-08, 1.50917e-07, 1.244649e-06, 2.947479e-06, 1.494664e-05, 
    0.0001060958, 0.0002065939, 0.0003413509, 0.0005454223, 0.0006654588, 
    0.0006389356, 0.0005174767, 0.0005785606, 0.0001210635, 2.001379e-05,
  7.721421e-08, 4.4419e-08, 1.487285e-07, 1.622166e-06, 3.247648e-06, 
    2.189462e-05, 0.0001342158, 0.000241468, 0.0004936582, 0.0007081018, 
    0.0007842288, 0.0007516205, 0.0006450524, 0.0002253324, 1.519705e-05,
  4.299234e-09, 8.354948e-08, 5.234389e-08, 2.932451e-07, 1.490118e-06, 
    3.085778e-06, 5.748633e-05, 0.0001607185, 0.0003459839, 0.0006893239, 
    0.00077881, 0.0007933951, 0.0006162187, 0.0005073649, 3.748036e-05,
  2.239503e-07, 1.44256e-07, 4.242747e-08, 2.26237e-08, 1.492194e-07, 
    1.145565e-06, 8.661737e-06, 7.561314e-05, 0.0002017805, 0.0005781397, 
    0.0007276452, 0.0006914075, 0.0006852908, 0.0003801695, 8.821409e-05,
  1.768228e-07, 1.402636e-07, 2.78822e-08, 3.963672e-08, 2.66428e-09, 
    3.76343e-08, 1.962787e-06, 1.495018e-05, 0.000119169, 0.0002990388, 
    0.0006465964, 0.0005464426, 0.0005712623, 0.0006214762, 0.0002804142,
  5.442647e-09, 1.216497e-08, 8.225513e-09, 2.974347e-08, 2.067186e-09, 
    1.510535e-11, 1.319462e-07, 2.608798e-06, 2.132029e-05, 8.85396e-05, 
    0.0004451818, 0.0004860348, 0.0005152213, 0.0006256034, 0.000487275,
  1.718323e-13, 5.365025e-11, 1.054928e-09, 3.811369e-08, 3.041847e-09, 
    5.596991e-11, 5.302347e-10, 8.172283e-07, 1.385004e-06, 2.119229e-05, 
    0.0001558065, 0.0004683771, 0.000459642, 0.0005708449, 0.0005980305,
  8.022067e-14, 3.104372e-12, 1.288972e-10, 2.137396e-08, 8.476945e-09, 
    3.585249e-10, 5.141426e-08, 6.949957e-07, 7.228372e-07, 2.948807e-07, 
    2.725321e-05, 0.0003227452, 0.0004855027, 0.0005465859, 0.0006442949,
  4.925451e-13, 5.931106e-13, 1.926937e-11, 5.085025e-09, 2.320774e-07, 
    3.828407e-08, 2.181352e-11, 2.075693e-08, 3.022234e-08, 1.805399e-07, 
    1.217305e-05, 0.0001173471, 0.0004512481, 0.0005184421, 0.0006416901,
  3.268562e-12, 1.999426e-12, 8.059775e-12, 3.244114e-08, 3.512178e-08, 
    3.558133e-09, 1.237424e-10, 8.843468e-09, 5.910224e-09, 3.485831e-08, 
    5.569116e-07, 2.731292e-05, 0.0002978696, 0.0005343628, 0.0006432272,
  5.515339e-07, 7.620833e-07, 3.791428e-06, 3.688365e-06, 1.38709e-05, 
    5.749794e-05, 7.227154e-05, 4.847281e-05, 4.717395e-05, 4.082616e-05, 
    7.262953e-05, 0.0001036101, 8.994425e-05, 3.636971e-05, 1.509078e-05,
  6.330249e-07, 3.366562e-07, 1.017025e-06, 2.152434e-06, 5.158917e-06, 
    2.691681e-05, 8.613923e-05, 7.596082e-05, 6.417438e-05, 7.010361e-05, 
    0.0001212176, 0.0001808231, 0.0001421328, 4.858786e-05, 5.503223e-06,
  4.126566e-07, 2.731564e-07, 2.500981e-07, 1.202577e-06, 2.696536e-06, 
    1.066142e-05, 6.698277e-05, 8.647026e-05, 8.343308e-05, 0.0001204794, 
    0.000211, 0.0002669138, 0.0001949775, 8.078526e-05, 6.946085e-06,
  2.586827e-07, 3.67331e-07, 2.872106e-07, 6.271007e-07, 2.35888e-06, 
    3.073894e-06, 2.68385e-05, 9.000266e-05, 0.0001051488, 0.0001718919, 
    0.0002788508, 0.0003215449, 0.0002304302, 9.018192e-05, 1.108029e-05,
  1.568371e-07, 3.643225e-07, 4.627422e-07, 5.122217e-07, 6.549342e-07, 
    2.232919e-06, 1.084692e-05, 7.122044e-05, 0.0001413849, 0.0002111048, 
    0.0003152605, 0.0003732415, 0.0002634563, 9.266174e-05, 1.765765e-05,
  2.118681e-07, 3.350353e-07, 4.381874e-07, 4.401564e-07, 3.420477e-07, 
    4.44286e-07, 1.063823e-05, 5.337698e-05, 0.000156486, 0.0002474053, 
    0.0003848129, 0.0004494449, 0.0003221859, 0.0001022426, 1.557547e-05,
  3.05646e-07, 4.827816e-07, 3.562787e-07, 8.417373e-07, 2.161581e-07, 
    7.194953e-08, 6.418252e-06, 4.455193e-05, 9.759486e-05, 0.0002430518, 
    0.0004172509, 0.0005364611, 0.0004033362, 0.0001385096, 2.6965e-05,
  2.123392e-08, 2.556262e-07, 2.145366e-07, 9.592706e-07, 1.29327e-07, 
    4.060816e-08, 6.919803e-06, 6.607514e-05, 0.0001396063, 0.0002224822, 
    0.000423036, 0.0005772972, 0.0005086793, 0.0002249109, 5.859911e-05,
  2.33199e-08, 1.313459e-07, 4.024369e-07, 1.725953e-06, 2.462315e-07, 
    2.943698e-08, 4.291887e-07, 2.003127e-05, 0.000118478, 0.0002080565, 
    0.0003682993, 0.0005660171, 0.0005572475, 0.0002796861, 6.717132e-05,
  1.983217e-08, 1.146474e-07, 2.388327e-07, 1.674474e-07, 4.587729e-07, 
    1.830218e-08, 1.347075e-07, 9.349775e-06, 7.551075e-05, 0.0001660094, 
    0.0003189315, 0.0005790631, 0.0005714751, 0.0003515155, 7.981798e-05,
  7.053016e-09, 2.508843e-08, 2.583158e-08, 8.075583e-08, 1.440907e-07, 
    1.010401e-07, 6.832235e-08, 5.12947e-08, 2.227223e-07, 1.970976e-06, 
    5.328343e-05, 0.0001503143, 0.0002439745, 0.000253835, 0.0001388756,
  7.149501e-09, 7.844842e-10, 1.588031e-08, 8.833254e-08, 1.143471e-06, 
    1.584268e-06, 3.237268e-08, 8.013888e-08, 5.457727e-08, 1.024971e-06, 
    4.271639e-05, 0.0001469513, 0.0002260895, 0.0001938124, 0.0001029262,
  2.531029e-07, 7.146587e-08, 1.357469e-09, 2.185093e-09, 1.814751e-06, 
    3.027101e-06, 1.550651e-06, 1.477441e-06, 2.18319e-07, 3.75576e-06, 
    5.155307e-05, 0.0001399467, 0.0002055183, 0.0001651232, 8.204748e-05,
  2.683153e-06, 3.278738e-07, 5.612055e-07, 3.08877e-07, 9.419373e-07, 
    2.05712e-07, 2.864741e-06, 6.508637e-07, 3.140263e-06, 6.633404e-06, 
    3.169588e-05, 8.60253e-05, 0.0001463927, 0.0001302482, 6.995388e-05,
  2.055589e-06, 1.264958e-06, 3.44017e-06, 7.524645e-07, 8.820691e-07, 
    6.005624e-09, 1.269278e-07, 3.503549e-07, 2.151304e-07, 6.211954e-07, 
    6.421809e-06, 3.13299e-05, 8.481449e-05, 0.0001082201, 5.536619e-05,
  1.401717e-05, 3.053758e-06, 2.576157e-08, 4.752919e-09, 4.051551e-08, 
    5.477525e-11, 8.127341e-08, 3.124685e-07, 1.176305e-07, 4.616562e-08, 
    1.832082e-06, 1.139208e-05, 5.376665e-05, 8.138866e-05, 4.254622e-05,
  5.871314e-09, 4.213971e-08, 1.546038e-09, 2.036263e-08, 2.768966e-08, 
    2.72812e-10, 3.25774e-09, 3.002864e-07, 3.625877e-07, 8.005447e-08, 
    3.140386e-06, 2.342292e-05, 4.574273e-05, 5.594067e-05, 3.1443e-05,
  3.091227e-09, 2.051149e-09, 1.145737e-10, 7.087186e-10, 5.90003e-09, 
    3.366913e-09, 1.124485e-08, 2.593294e-07, 9.225708e-08, 5.273439e-08, 
    8.90858e-06, 2.450315e-05, 3.140168e-05, 2.499015e-05, 1.879968e-05,
  8.929185e-11, 2.010157e-10, 9.180105e-09, 7.135182e-08, 1.9313e-07, 
    1.916418e-08, 4.655554e-10, 9.466576e-09, 1.519764e-06, 7.126822e-06, 
    1.429617e-05, 1.633891e-05, 1.441965e-05, 1.213353e-05, 9.790137e-06,
  2.381738e-09, 2.573581e-09, 1.210257e-07, 3.245541e-08, 3.965325e-08, 
    3.324842e-08, 6.977293e-09, 9.077933e-09, 1.220027e-07, 4.925157e-06, 
    9.748797e-06, 1.429506e-05, 1.042436e-05, 8.99532e-06, 7.016155e-06,
  1.200533e-07, 1.632132e-07, 1.196965e-07, 3.230455e-07, 1.575924e-07, 
    2.180599e-08, 2.397949e-08, 4.015559e-06, 1.957972e-07, 2.010967e-06, 
    7.926505e-05, 0.0002258313, 0.000282293, 0.0002103158, 0.0001045638,
  3.374479e-08, 6.120776e-08, 5.215987e-08, 2.792638e-07, 7.076861e-07, 
    1.488782e-06, 1.374212e-06, 1.719556e-06, 1.154437e-07, 2.112547e-06, 
    0.0001121459, 0.0003220799, 0.0003256554, 0.000226413, 0.0001151587,
  1.550063e-06, 1.595028e-06, 6.025341e-08, 3.059893e-08, 1.592018e-06, 
    3.691346e-06, 6.115542e-06, 5.57407e-06, 1.610127e-06, 2.455949e-06, 
    0.000107101, 0.0003497085, 0.0003731929, 0.0002637234, 0.0001565679,
  2.075972e-05, 1.264416e-05, 4.090753e-06, 4.455836e-07, 1.503447e-06, 
    1.557879e-06, 5.320517e-06, 4.957744e-06, 4.139878e-06, 1.032897e-05, 
    8.176604e-05, 0.000306615, 0.0003573592, 0.0002897638, 0.0001983527,
  4.884257e-05, 4.441955e-05, 3.263886e-05, 5.248604e-06, 1.242093e-06, 
    1.534597e-06, 1.721582e-06, 1.108331e-06, 8.555318e-08, 1.881986e-05, 
    6.189966e-05, 0.0002321743, 0.0003455263, 0.0003222206, 0.0002954052,
  4.320537e-05, 3.949252e-05, 1.294519e-06, 7.406853e-06, 1.93776e-06, 
    2.337585e-08, 4.760027e-08, 1.346992e-07, 9.601347e-07, 1.532235e-05, 
    4.583004e-05, 0.0001718931, 0.0003560262, 0.0004122225, 0.0004189412,
  1.781117e-05, 1.258041e-05, 1.16976e-06, 1.881473e-07, 1.247392e-08, 
    7.087356e-07, 1.260992e-08, 6.727768e-08, 9.891426e-08, 4.899443e-06, 
    3.479418e-05, 0.0001277436, 0.0002924875, 0.0004183628, 0.0004894029,
  1.405949e-05, 8.817623e-06, 9.408561e-08, 1.820404e-07, 6.244986e-09, 
    4.978773e-07, 9.925843e-07, 4.274535e-08, 1.180625e-07, 5.041779e-06, 
    3.532648e-05, 9.14054e-05, 0.0001762883, 0.0002884481, 0.0003417567,
  7.685599e-06, 1.627747e-06, 1.484023e-09, 6.587436e-09, 1.383397e-06, 
    7.699779e-07, 1.208187e-09, 1.054465e-06, 1.135417e-05, 2.250742e-05, 
    4.478542e-05, 5.943705e-05, 7.213933e-05, 0.0001322154, 0.0001803897,
  1.005461e-05, 5.686315e-06, 1.13566e-07, 9.369234e-10, 2.453137e-06, 
    1.424196e-07, 4.886152e-07, 2.235436e-07, 1.224385e-05, 2.486497e-05, 
    3.690827e-05, 2.604677e-05, 3.554368e-05, 5.796841e-05, 8.973423e-05,
  2.154399e-07, 2.269555e-07, 1.749057e-07, 5.60845e-08, 5.052907e-09, 
    4.294143e-09, 4.719536e-09, 2.657896e-08, 1.92527e-07, 8.621788e-07, 
    5.200753e-06, 3.161349e-05, 8.281869e-05, 6.972533e-05, 4.956054e-05,
  3.097816e-08, 9.379725e-08, 1.549909e-07, 7.654785e-08, 6.234951e-09, 
    5.112526e-10, 5.538562e-09, 9.676955e-08, 1.868341e-08, 2.838531e-07, 
    1.353416e-05, 6.386155e-05, 0.000110208, 7.434979e-05, 4.729992e-05,
  1.589983e-08, 1.067072e-08, 4.59386e-08, 8.517413e-08, 2.067516e-08, 
    3.770409e-08, 1.831807e-07, 3.955025e-07, 5.519341e-07, 1.531307e-06, 
    2.921147e-05, 0.0001113733, 0.0001420271, 9.446083e-05, 6.203627e-05,
  4.398293e-06, 1.229935e-05, 1.552562e-08, 1.963895e-08, 2.273675e-08, 
    9.202509e-07, 1.186061e-06, 1.927854e-06, 1.978035e-06, 6.181794e-06, 
    3.358522e-05, 0.000125934, 0.00016642, 0.0001188013, 7.74588e-05,
  9.978067e-06, 1.318604e-05, 1.102888e-06, 9.23272e-10, 1.35048e-07, 
    3.128328e-07, 1.054047e-06, 5.191533e-07, 1.967175e-06, 1.11242e-05, 
    3.551477e-05, 0.0001245122, 0.0001884712, 0.0001485468, 9.997255e-05,
  2.170579e-05, 1.649075e-05, 1.436459e-06, 4.64141e-06, 8.188376e-07, 
    7.357402e-07, 1.400276e-09, 1.68033e-09, 6.840907e-09, 7.224594e-06, 
    2.951624e-05, 8.390204e-05, 0.0001537063, 0.0001481589, 0.000110916,
  2.032493e-09, 2.530279e-05, 1.147621e-05, 1.724058e-06, 1.319759e-06, 
    2.339454e-06, 2.735191e-09, 1.079774e-09, 1.283484e-08, 2.252129e-06, 
    2.560007e-05, 5.663404e-05, 7.77637e-05, 0.0001051356, 0.0001044833,
  1.430072e-06, 8.685011e-06, 1.302422e-05, 5.30428e-06, 1.593111e-06, 
    6.374494e-06, 5.556523e-06, 2.502888e-06, 1.753885e-06, 1.173225e-05, 
    5.211939e-05, 6.850022e-05, 5.440203e-05, 4.534254e-05, 8.096196e-05,
  9.951325e-06, 1.679729e-05, 1.049897e-05, 8.260186e-07, 1.730986e-05, 
    5.19681e-06, 8.504562e-07, 3.149595e-06, 5.63469e-05, 8.984199e-05, 
    0.000125021, 0.000122491, 6.736116e-05, 3.456253e-05, 5.086629e-05,
  1.534407e-05, 2.856842e-05, 1.226089e-05, 5.844965e-06, 1.657069e-05, 
    5.807673e-06, 2.368411e-06, 4.064969e-06, 3.563357e-05, 6.512543e-05, 
    0.000145631, 0.0001428329, 6.461496e-05, 3.497651e-05, 3.237315e-05,
  1.60068e-06, 1.380393e-06, 2.996383e-06, 6.407482e-06, 6.875963e-07, 
    5.05347e-09, 2.720323e-08, 4.593603e-08, 1.615995e-07, 6.608619e-07, 
    1.336829e-06, 1.383036e-05, 3.935025e-05, 3.368943e-05, 1.24648e-05,
  1.109192e-06, 1.381008e-06, 1.776612e-06, 6.503159e-06, 5.33832e-06, 
    2.327013e-07, 7.249358e-09, 3.353408e-08, 1.796088e-08, 1.039697e-06, 
    1.610499e-05, 4.378267e-05, 6.260907e-05, 3.414457e-05, 7.98906e-06,
  1.010343e-06, 4.624118e-07, 2.069799e-06, 5.297324e-06, 2.189551e-05, 
    8.788665e-06, 1.416581e-06, 4.219388e-07, 1.911018e-06, 9.654046e-06, 
    4.756394e-05, 9.082013e-05, 6.853484e-05, 3.540418e-05, 7.507116e-06,
  6.553915e-06, 1.035353e-05, 9.12113e-06, 2.018075e-05, 2.450927e-05, 
    1.064123e-05, 1.661449e-06, 3.627627e-07, 3.736853e-06, 2.831929e-05, 
    9.215459e-05, 0.0001233199, 9.822297e-05, 4.623718e-05, 5.446473e-06,
  1.117988e-05, 1.152626e-05, 1.850221e-05, 4.911787e-06, 9.970663e-06, 
    1.147234e-06, 6.111765e-08, 5.005822e-09, 4.586503e-06, 3.316686e-05, 
    6.027391e-05, 0.000147256, 0.0001082504, 4.424057e-05, 6.892372e-06,
  2.480278e-05, 2.445122e-05, 1.373431e-05, 3.474946e-06, 5.107385e-06, 
    5.349087e-07, 4.712463e-08, 5.551729e-09, 1.894367e-05, 3.33461e-05, 
    0.000101478, 0.000158116, 0.0001123844, 3.626985e-05, 2.702402e-06,
  6.324696e-05, 9.280157e-05, 8.064376e-05, 5.69274e-06, 5.569706e-07, 
    2.584509e-07, 2.258789e-07, 3.455994e-06, 2.058875e-06, 8.287435e-06, 
    9.018686e-05, 0.0001988244, 0.0001450642, 2.195891e-05, 5.696186e-07,
  5.948278e-05, 0.0001140394, 4.639482e-05, 1.798389e-06, 8.523593e-08, 
    5.502878e-07, 9.523392e-07, 6.764841e-07, 6.775153e-06, 6.955362e-06, 
    6.908813e-05, 0.0002303103, 0.000134586, 3.215286e-05, 7.528163e-07,
  6.719717e-06, 2.038598e-05, 1.828828e-05, 1.776622e-07, 2.205372e-06, 
    1.85999e-06, 4.027124e-07, 5.150232e-06, 1.700522e-05, 5.370786e-05, 
    0.0001399917, 0.0003179222, 0.0001680062, 3.287557e-05, 2.488427e-06,
  3.003502e-08, 1.546512e-07, 8.88276e-07, 3.8607e-07, 8.63844e-06, 
    2.369664e-06, 1.213688e-06, 1.419069e-05, 6.849129e-06, 7.287237e-05, 
    0.000168785, 0.0004310844, 0.0002330915, 3.526199e-05, 7.537725e-06,
  4.874622e-08, 6.865658e-08, 3.489009e-08, 3.513009e-09, 1.059102e-07, 
    2.285049e-08, 1.906989e-08, 2.740236e-08, 1.606065e-07, 1.542174e-05, 
    0.0001016495, 0.0001915323, 0.0003026251, 0.0003559319, 0.0004355269,
  8.856588e-09, 3.990971e-08, 2.417046e-08, 8.296534e-09, 1.216901e-07, 
    6.739891e-07, 1.613852e-07, 5.68168e-08, 4.635339e-08, 3.214269e-06, 
    7.002808e-05, 0.0001803151, 0.0002794462, 0.0002874566, 0.0002831425,
  1.610782e-05, 3.704605e-06, 5.574591e-09, 7.933349e-08, 2.089756e-06, 
    4.939164e-06, 3.192541e-06, 1.563457e-06, 7.814677e-07, 4.154993e-06, 
    4.36134e-05, 0.0001522804, 0.0002586633, 0.0002539708, 0.000187466,
  3.78029e-05, 1.79681e-05, 1.45563e-07, 4.743103e-08, 6.448874e-06, 
    9.135277e-06, 8.76608e-06, 6.066794e-06, 3.247513e-06, 8.124615e-06, 
    1.848159e-05, 0.0001052322, 0.0002270376, 0.0002431385, 0.0001497081,
  3.971977e-05, 2.755914e-05, 6.749372e-06, 5.429835e-09, 4.070796e-06, 
    3.686948e-06, 6.563297e-06, 7.735293e-06, 6.184162e-06, 1.119936e-05, 
    9.580114e-06, 5.49927e-05, 0.0001718553, 0.0002536614, 0.0001532511,
  4.860063e-05, 2.788771e-05, 1.362043e-08, 3.949451e-07, 3.868102e-06, 
    3.343833e-06, 8.96558e-07, 2.875217e-06, 3.441048e-06, 8.458132e-06, 
    6.995773e-06, 2.013802e-05, 0.0001169403, 0.000196791, 0.0001579198,
  3.685535e-05, 1.385614e-05, 1.278957e-05, 7.422305e-06, 4.267284e-06, 
    3.276554e-06, 1.635865e-06, 1.300906e-08, 2.685789e-07, 2.073599e-06, 
    3.918526e-06, 8.910529e-06, 6.819842e-05, 0.0001322899, 0.0001330397,
  2.66591e-05, 3.511661e-05, 3.358311e-05, 1.460059e-05, 6.93622e-06, 
    1.350178e-05, 1.889459e-05, 1.380358e-05, 9.175213e-06, 2.192669e-06, 
    6.663842e-06, 3.785463e-05, 7.537148e-05, 8.844839e-05, 0.0001065671,
  4.112232e-05, 7.036451e-05, 3.602489e-05, 1.741703e-05, 3.373252e-05, 
    7.867377e-06, 2.827039e-05, 5.491137e-05, 7.298701e-05, 2.973416e-05, 
    2.71046e-05, 4.944671e-05, 7.766087e-05, 8.414076e-05, 8.235216e-05,
  1.535842e-05, 3.265481e-05, 5.021824e-05, 2.188284e-05, 3.287448e-05, 
    3.499393e-05, 9.60351e-05, 0.000217957, 0.0001674824, 8.22627e-05, 
    6.98353e-05, 9.309974e-05, 0.0001017416, 5.404505e-05, 5.396951e-05,
  2.482804e-07, 7.700858e-08, 4.364722e-08, 2.691606e-07, 6.709119e-08, 
    1.692209e-08, 2.396954e-08, 2.194054e-08, 9.015829e-08, 6.318855e-06, 
    2.601056e-05, 7.542946e-05, 0.0001473967, 0.0001147427, 5.828795e-05,
  2.127856e-07, 5.966305e-08, 1.400285e-08, 6.106083e-07, 1.066642e-07, 
    1.954667e-07, 9.768856e-07, 2.152069e-08, 2.793173e-08, 2.757848e-06, 
    3.424167e-05, 9.478362e-05, 0.0001120259, 0.0001002293, 5.967782e-05,
  1.948382e-07, 2.816344e-07, 1.242988e-07, 8.927499e-07, 7.114937e-08, 
    1.956647e-08, 3.332847e-06, 3.215049e-06, 8.795637e-08, 1.722025e-06, 
    2.8632e-05, 8.606743e-05, 0.0001150572, 0.0001283254, 9.176171e-05,
  4.037319e-07, 5.58833e-07, 9.311098e-08, 1.841773e-06, 2.049149e-08, 
    1.348468e-07, 6.870191e-06, 7.064019e-06, 1.294631e-06, 9.069488e-06, 
    2.090909e-05, 6.688063e-05, 0.0001407655, 0.0001946674, 0.0001482683,
  1.318188e-06, 1.517901e-06, 2.77014e-07, 3.003772e-08, 1.100678e-07, 
    1.391726e-07, 5.170825e-06, 9.086771e-06, 3.188879e-06, 8.198209e-06, 
    1.442854e-05, 4.537035e-05, 0.0001383526, 0.0002649778, 0.000222359,
  5.160936e-06, 3.878773e-06, 5.027282e-08, 1.508994e-08, 4.496857e-07, 
    2.174226e-07, 7.159287e-08, 2.305298e-07, 4.640342e-06, 8.160296e-06, 
    1.059161e-05, 2.81725e-05, 0.0001193116, 0.0002892001, 0.0002922461,
  2.31287e-07, 1.358767e-07, 3.204503e-07, 1.819227e-07, 5.339933e-07, 
    1.707211e-06, 2.217239e-08, 2.643389e-09, 4.822851e-07, 4.717821e-06, 
    9.687542e-06, 2.210974e-05, 9.861829e-05, 0.0002743186, 0.0003491656,
  8.808446e-09, 1.367512e-08, 2.281789e-06, 1.06515e-06, 8.033359e-07, 
    4.112565e-06, 3.394373e-06, 8.61719e-07, 8.59785e-07, 7.944344e-06, 
    1.319881e-05, 2.062072e-05, 7.23649e-05, 0.0002443879, 0.0004096544,
  4.222636e-06, 3.697558e-06, 2.08607e-06, 1.518467e-06, 5.962433e-06, 
    2.491617e-06, 2.514183e-07, 1.660856e-06, 1.426367e-05, 1.905282e-05, 
    1.45868e-05, 1.744708e-05, 5.443015e-05, 0.0002029803, 0.0004210404,
  2.996496e-06, 2.788679e-06, 1.389524e-06, 2.803589e-07, 7.283775e-06, 
    3.683323e-06, 1.654969e-06, 2.530398e-08, 4.858494e-06, 1.291218e-05, 
    1.254246e-05, 1.785262e-05, 3.949043e-05, 0.0002010234, 0.000403911,
  2.124613e-07, 3.332068e-07, 3.277721e-07, 2.374546e-07, 1.416917e-07, 
    3.311682e-06, 1.369342e-05, 2.935156e-05, 6.406355e-05, 9.929037e-05, 
    8.092105e-05, 1.735803e-05, 1.011295e-05, 1.777526e-05, 8.549644e-06,
  6.944824e-07, 8.994241e-07, 1.805234e-07, 1.828725e-07, 6.549404e-08, 
    1.465542e-06, 1.075063e-05, 2.369602e-05, 4.268867e-05, 5.548557e-05, 
    3.188909e-05, 3.07877e-06, 3.957758e-06, 3.103528e-06, 1.021214e-06,
  4.173601e-06, 3.60836e-06, 4.421854e-07, 2.355088e-07, 1.233303e-07, 
    3.640582e-07, 5.45726e-06, 2.066172e-05, 4.848987e-05, 2.72568e-05, 
    1.370226e-05, 4.831225e-06, 1.017678e-06, 4.036729e-07, 1.494756e-08,
  9.121477e-06, 4.666018e-06, 1.247093e-07, 1.302231e-07, 1.176667e-07, 
    8.498329e-09, 6.067623e-06, 6.580135e-05, 6.786196e-05, 4.457865e-05, 
    1.33456e-05, 4.623754e-06, 2.977278e-06, 1.398063e-06, 5.097059e-08,
  3.162317e-06, 2.563249e-06, 2.058961e-07, 1.559839e-07, 5.04708e-08, 
    5.430138e-09, 2.309402e-07, 2.7528e-05, 4.487627e-05, 5.498671e-05, 
    2.50694e-05, 7.653619e-06, 4.694246e-06, 1.93201e-06, 5.67132e-07,
  9.304854e-08, 8.923598e-08, 1.253874e-07, 1.605977e-07, 7.293558e-08, 
    5.436463e-09, 5.89235e-10, 6.909051e-07, 8.750575e-06, 4.045774e-05, 
    3.27316e-05, 1.547477e-05, 7.284639e-06, 3.717978e-06, 1.487241e-06,
  2.409317e-09, 1.172647e-08, 1.166118e-07, 6.606489e-08, 4.439721e-08, 
    2.483372e-08, 6.781419e-10, 2.96788e-07, 1.155207e-07, 1.023807e-05, 
    2.957719e-05, 2.371125e-05, 9.736302e-06, 6.269743e-06, 2.965326e-06,
  5.520083e-10, 7.892488e-10, 5.057438e-09, 8.724006e-09, 1.097599e-08, 
    3.99126e-08, 2.023286e-09, 1.176357e-06, 1.989105e-06, 1.32789e-06, 
    1.81678e-05, 2.66609e-05, 1.290366e-05, 5.116888e-06, 4.910778e-06,
  4.357314e-11, 6.511468e-11, 4.27568e-10, 1.744887e-09, 6.454718e-09, 
    5.119265e-09, 3.968517e-09, 5.295076e-07, 4.865472e-07, 5.671496e-06, 
    1.765538e-05, 1.980034e-05, 1.178523e-05, 5.136006e-06, 6.658997e-06,
  8.529405e-13, 1.831662e-13, 9.63273e-11, 1.127012e-09, 2.446483e-07, 
    2.576631e-09, 5.754739e-09, 5.146364e-09, 1.285537e-06, 4.028965e-06, 
    9.711794e-06, 1.225519e-05, 7.022094e-06, 6.781928e-06, 5.763845e-06,
  8.713493e-07, 5.974895e-07, 3.414152e-06, 6.87815e-06, 1.334012e-05, 
    1.044014e-05, 2.265458e-05, 6.988805e-05, 0.0001459971, 0.0002654259, 
    0.0003132953, 0.0002634295, 0.0001940516, 0.000128248, 0.0001173983,
  5.147325e-07, 2.531115e-07, 4.739828e-07, 5.112058e-06, 3.154546e-05, 
    6.47094e-05, 7.151612e-05, 9.141063e-05, 0.0001950678, 0.0003292188, 
    0.0003782464, 0.0002723435, 0.0001745352, 0.0001002363, 0.0001426937,
  4.134809e-06, 8.109371e-07, 6.395426e-07, 6.355224e-06, 3.943929e-05, 
    0.000105175, 0.0001761487, 0.000150813, 0.0002789886, 0.0004035876, 
    0.0003992462, 0.0002991618, 0.0001421936, 0.0001337241, 0.000175438,
  1.389671e-05, 2.134764e-06, 1.228466e-06, 4.421174e-06, 3.573084e-05, 
    0.0001242102, 0.0002239522, 0.0002853964, 0.0004188716, 0.0004967491, 
    0.0004563199, 0.000341765, 0.0001647761, 0.0001645729, 0.0001983656,
  9.774028e-06, 1.967719e-06, 2.694737e-06, 1.491494e-05, 0.0001224455, 
    0.0003090769, 0.0004537493, 0.0005365803, 0.0006069884, 0.0006033579, 
    0.0004800188, 0.0002905988, 0.0002180422, 0.0002050512, 0.0002087365,
  6.480261e-06, 3.130917e-07, 6.636566e-06, 9.161129e-05, 0.0003001055, 
    0.0004397962, 0.0006072828, 0.0007418412, 0.0007227974, 0.000628889, 
    0.0005215543, 0.0003251307, 0.0002759872, 0.0002244053, 0.000217092,
  7.297136e-08, 6.193691e-07, 2.792477e-05, 0.0001691295, 0.0003399061, 
    0.000407523, 0.0004843521, 0.0005879863, 0.0007097208, 0.0006084518, 
    0.000477708, 0.0003356378, 0.0002839613, 0.0002414212, 0.0002138093,
  1.362039e-07, 4.064121e-06, 3.831317e-05, 0.000124707, 0.0002087811, 
    0.000285381, 0.0003477209, 0.0004446793, 0.0005537411, 0.0004873055, 
    0.0005018918, 0.0004065565, 0.0003056292, 0.0002615865, 0.0001978947,
  3.437795e-07, 8.557123e-06, 1.620786e-05, 3.719775e-05, 0.0001289372, 
    0.0002014945, 0.0002553272, 0.0003654353, 0.0004858402, 0.0005109312, 
    0.0005105933, 0.0004177626, 0.0003618416, 0.0002865157, 0.0002013365,
  5.106471e-07, 4.652877e-06, 4.727646e-06, 1.788953e-05, 0.0001095635, 
    0.0001614551, 0.0002316864, 0.0003901596, 0.0004768621, 0.0005397162, 
    0.0005455472, 0.000499549, 0.0003909718, 0.0002909528, 0.000212854,
  5.315265e-09, 4.484646e-08, 7.179138e-07, 2.554692e-06, 1.182767e-06, 
    1.101967e-09, 4.171224e-07, 7.37148e-07, 4.027259e-07, 4.912286e-07, 
    1.134957e-06, 1.381683e-06, 1.61953e-06, 1.111823e-06, 7.641148e-07,
  3.438625e-09, 2.332213e-07, 7.601327e-07, 1.917176e-06, 3.554733e-06, 
    1.191934e-06, 6.830928e-07, 1.028258e-06, 1.07403e-06, 4.971342e-07, 
    4.040247e-07, 1.424956e-06, 1.500602e-06, 3.862905e-07, 3.585267e-07,
  1.947114e-07, 7.736656e-07, 5.509752e-07, 7.03846e-07, 1.778793e-06, 
    3.873702e-06, 3.38927e-06, 2.75719e-06, 2.755337e-06, 1.41345e-06, 
    1.91262e-06, 2.007942e-06, 1.381463e-06, 8.08595e-07, 2.2268e-07,
  2.048757e-06, 1.623156e-06, 1.782833e-07, 6.257466e-07, 1.347537e-06, 
    3.620057e-06, 5.484817e-06, 5.69902e-06, 7.057614e-06, 5.91282e-06, 
    5.364661e-06, 2.721454e-06, 2.659749e-06, 7.362173e-07, 5.490987e-07,
  1.633557e-06, 3.631126e-06, 1.898112e-06, 2.807528e-09, 5.390869e-07, 
    2.913963e-06, 5.477618e-06, 7.114355e-06, 9.057578e-06, 1.041449e-05, 
    8.662835e-06, 3.12747e-06, 3.116959e-06, 1.695877e-06, 1.143787e-06,
  9.394061e-06, 2.957731e-06, 3.583398e-07, 1.264294e-06, 5.63746e-06, 
    6.92946e-06, 6.100211e-06, 5.814935e-06, 8.250357e-06, 1.28627e-05, 
    1.114687e-05, 2.853464e-06, 1.906021e-06, 1.178194e-06, 7.994553e-07,
  1.50188e-05, 1.728753e-05, 2.136682e-05, 2.733755e-05, 2.724639e-05, 
    1.473977e-05, 3.636844e-06, 1.239698e-06, 4.103045e-06, 6.872062e-06, 
    1.082755e-05, 7.894895e-06, 2.288026e-06, 1.014844e-06, 5.052714e-07,
  1.311976e-05, 1.881951e-05, 2.19943e-05, 2.745759e-05, 3.187875e-05, 
    3.643602e-05, 2.338285e-05, 1.146215e-05, 1.002996e-06, 1.870659e-07, 
    8.880277e-06, 6.425058e-06, 4.476363e-06, 1.463215e-06, 4.654295e-07,
  1.312815e-05, 1.867259e-05, 2.468963e-05, 2.953995e-05, 6.576622e-05, 
    4.57067e-05, 3.691386e-05, 2.097171e-05, 1.224328e-05, 7.061642e-06, 
    7.620394e-06, 1.536363e-05, 9.747033e-06, 2.683599e-06, 7.186269e-07,
  2.819408e-05, 2.785429e-05, 1.830583e-05, 5.499794e-05, 0.0001206984, 
    0.0001442298, 0.0001687802, 0.0001601156, 0.0001116181, 4.113352e-05, 
    1.62106e-05, 8.413737e-06, 4.122098e-06, 3.464063e-06, 2.503378e-06,
  8.645001e-10, 9.411152e-11, 1.021043e-08, 3.123698e-09, 1.188052e-10, 
    4.085558e-11, 2.769546e-12, 8.030156e-13, 2.085997e-13, 6.583657e-24, 
    1.355455e-23, 1.454672e-10, 4.271957e-11, 9.143533e-11, 1.705635e-07,
  9.003696e-09, 3.552888e-09, 1.473197e-10, 1.059828e-08, 7.039765e-08, 
    5.274961e-10, 3.925779e-12, 2.430416e-13, 2.707557e-24, 5.9227e-24, 
    4.958132e-24, 2.173065e-11, 9.925307e-11, 2.692715e-09, 7.549075e-08,
  1.078258e-06, 1.059801e-06, 4.589694e-08, 1.575589e-08, 2.085479e-07, 
    9.909103e-08, 2.171455e-08, 7.706685e-09, 4.163831e-09, 3.467167e-24, 
    4.546207e-24, 8.935424e-08, 2.611808e-10, 1.081358e-08, 9.324014e-09,
  1.989717e-06, 1.468149e-06, 1.320961e-08, 3.760258e-08, 8.654599e-08, 
    1.820989e-09, 1.463369e-07, 6.122183e-07, 1.642674e-06, 1.555142e-06, 
    1.912901e-06, 2.701564e-06, 6.925569e-07, 2.24388e-07, 1.040722e-07,
  6.240027e-07, 1.192435e-07, 1.853801e-09, 3.412512e-11, 9.194712e-11, 
    3.358292e-11, 4.267061e-09, 5.793128e-09, 5.810483e-07, 3.293455e-06, 
    4.730312e-06, 6.734322e-06, 4.295333e-06, 6.197742e-07, 4.027781e-07,
  3.453354e-08, 1.748335e-09, 1.77403e-11, 4.924992e-11, 2.076182e-09, 
    2.38673e-10, 1.689611e-10, 5.949428e-11, 1.1223e-06, 4.969161e-06, 
    9.327148e-06, 7.198146e-06, 4.880118e-06, 1.063132e-06, 1.952614e-07,
  2.273533e-08, 2.80727e-07, 4.349876e-07, 2.248654e-07, 1.05884e-07, 
    1.803017e-07, 3.551316e-10, 1.398946e-09, 4.982816e-10, 4.517192e-07, 
    5.540441e-06, 7.378522e-06, 7.315365e-06, 2.94919e-06, 6.960049e-07,
  1.980327e-07, 1.427495e-06, 3.624252e-06, 1.987544e-06, 2.909158e-06, 
    4.570752e-06, 3.409144e-06, 1.905674e-06, 7.814213e-09, 6.430506e-10, 
    1.070951e-06, 5.713857e-06, 6.920292e-06, 3.249347e-06, 7.837771e-07,
  1.085065e-07, 1.07327e-06, 3.942004e-06, 5.436852e-06, 2.670807e-05, 
    6.027664e-06, 1.444963e-06, 7.050447e-07, 7.408963e-07, 6.598475e-07, 
    3.576102e-07, 3.140147e-06, 4.164574e-06, 3.068696e-06, 1.508334e-06,
  2.732958e-06, 2.288872e-06, 3.972486e-06, 7.184542e-06, 2.132023e-05, 
    4.845801e-06, 9.659889e-06, 2.255135e-06, 7.031828e-06, 5.037808e-06, 
    2.608451e-06, 2.032141e-06, 3.117655e-06, 3.28341e-06, 2.291066e-06,
  3.780892e-06, 2.566476e-06, 2.414769e-06, 1.892971e-06, 8.693452e-07, 
    1.818757e-06, 1.784915e-06, 2.586576e-07, 7.871495e-10, 2.372824e-06, 
    1.699353e-05, 2.188242e-05, 6.15967e-06, 8.311261e-07, 3.334506e-09,
  6.538685e-06, 4.28307e-06, 2.884225e-06, 1.834904e-06, 1.829741e-06, 
    1.286982e-06, 1.828476e-06, 1.768093e-07, 3.173316e-09, 1.816327e-06, 
    1.019841e-05, 1.246559e-05, 2.896556e-06, 9.027593e-08, 5.901413e-11,
  1.129217e-05, 8.340339e-06, 2.468426e-06, 1.983489e-06, 8.319195e-07, 
    1.527489e-06, 1.067231e-06, 4.670449e-07, 1.160567e-08, 4.737823e-06, 
    1.382625e-05, 8.530416e-06, 2.577938e-07, 4.548735e-09, 5.720237e-08,
  1.761678e-05, 1.27273e-05, 2.25318e-06, 2.029869e-06, 1.480964e-06, 
    1.023245e-06, 1.313927e-06, 1.148083e-06, 2.991731e-06, 1.029489e-05, 
    1.272356e-05, 7.984237e-06, 1.416118e-07, 1.5854e-07, 2.162851e-07,
  7.541195e-06, 6.872162e-06, 4.635842e-06, 2.487937e-06, 2.921901e-06, 
    2.528651e-06, 1.167867e-05, 1.280839e-05, 1.191656e-05, 1.183226e-05, 
    1.128137e-05, 4.041075e-06, 1.411759e-07, 1.777139e-07, 5.710406e-08,
  6.126302e-06, 2.304136e-06, 1.25598e-06, 4.728586e-06, 5.983836e-06, 
    3.380975e-06, 6.935254e-06, 5.892213e-06, 5.557603e-06, 1.327241e-05, 
    7.373365e-06, 2.276412e-06, 7.824872e-07, 1.779786e-07, 7.953602e-08,
  1.037965e-07, 7.459064e-08, 4.211826e-06, 9.364209e-06, 6.639481e-06, 
    7.010365e-06, 1.148612e-06, 1.259201e-06, 3.207857e-06, 2.284721e-06, 
    6.720438e-06, 5.944661e-06, 2.112253e-06, 5.521176e-08, 3.842639e-09,
  6.762228e-07, 2.394223e-06, 1.252182e-05, 2.097341e-05, 9.83002e-06, 
    7.5136e-06, 7.604959e-06, 4.032036e-06, 1.577992e-07, 4.465853e-07, 
    6.659669e-06, 8.438498e-06, 5.986878e-06, 1.491461e-06, 1.006702e-08,
  4.372564e-06, 5.374583e-06, 2.292971e-05, 2.565448e-05, 5.000939e-05, 
    7.123013e-06, 1.366541e-06, 1.101717e-07, 2.655798e-08, 9.028296e-07, 
    8.72959e-06, 1.023284e-05, 5.378688e-06, 2.136031e-06, 7.925631e-07,
  1.259162e-05, 1.250343e-05, 2.643981e-05, 1.848172e-05, 2.051246e-05, 
    4.623717e-06, 1.945364e-06, 1.673903e-07, 1.6626e-06, 2.27801e-06, 
    8.368525e-06, 1.15347e-05, 4.686958e-06, 1.602598e-06, 1.127322e-06,
  1.241253e-09, 2.911544e-08, 3.493541e-08, 9.883786e-07, 3.83354e-05, 
    0.0001078164, 0.0001096839, 5.840686e-05, 7.290979e-05, 9.73444e-05, 
    0.0001618195, 0.000276593, 0.0002419814, 8.986145e-05, 3.222924e-05,
  5.248494e-10, 2.460821e-08, 2.676254e-08, 8.26976e-08, 8.822335e-06, 
    5.453296e-05, 0.0001032275, 6.653722e-05, 6.764349e-05, 0.0001133752, 
    0.0002134309, 0.0003118639, 0.0002774638, 8.463365e-05, 6.535884e-05,
  1.967585e-09, 3.945186e-08, 3.521113e-08, 2.035764e-08, 1.515405e-06, 
    2.575781e-05, 7.458831e-05, 7.741255e-05, 6.628118e-05, 0.0001466407, 
    0.000301021, 0.000406555, 0.0002884831, 0.0001167296, 6.866371e-05,
  1.363001e-08, 4.879299e-08, 2.563516e-08, 3.912324e-08, 5.434749e-08, 
    7.795569e-06, 4.597178e-05, 7.724274e-05, 7.528553e-05, 0.0001807851, 
    0.0003801609, 0.0004273777, 0.0003066749, 0.0001692372, 5.320783e-05,
  2.676456e-09, 1.325389e-08, 1.168628e-08, 3.684369e-08, 3.733506e-08, 
    2.553747e-06, 1.889744e-05, 6.288736e-05, 8.878233e-05, 0.0001995942, 
    0.000433018, 0.0004361589, 0.0002793513, 0.0001981395, 7.381442e-05,
  2.222646e-09, 1.282043e-10, 2.483818e-09, 7.471162e-08, 2.339033e-08, 
    3.323877e-07, 9.31212e-06, 4.025123e-05, 9.345066e-05, 0.0002243376, 
    0.0004771838, 0.0004264667, 0.0002515759, 0.0001730595, 0.0001083482,
  1.665765e-09, 2.146536e-09, 2.318928e-09, 8.619399e-08, 1.451677e-07, 
    2.611103e-05, 3.625214e-05, 5.932267e-05, 6.608458e-05, 0.0001750005, 
    0.0004795437, 0.0004017297, 0.0002155233, 0.0001611794, 0.0001143291,
  1.353825e-06, 3.265883e-07, 2.672458e-07, 3.84969e-07, 8.387986e-06, 
    1.733575e-05, 4.41361e-05, 5.725995e-05, 8.312226e-05, 0.0001066159, 
    0.0004762002, 0.0003632726, 0.0001877801, 0.0001411486, 0.0001317069,
  2.386069e-06, 1.035095e-06, 2.380665e-06, 5.810622e-06, 5.492901e-05, 
    2.012608e-05, 1.09251e-05, 2.822588e-06, 3.074464e-05, 0.0001662696, 
    0.0004083261, 0.0003505831, 0.0001690961, 0.0001289561, 0.0001122646,
  2.391913e-06, 1.726918e-06, 5.247647e-06, 1.546539e-05, 6.006179e-05, 
    1.928795e-05, 2.959934e-05, 2.397083e-05, 7.376862e-05, 0.0001917569, 
    0.0003958858, 0.0003299942, 0.0001500654, 0.0001288251, 0.0001023195,
  4.557196e-09, 6.450163e-10, 3.838457e-11, 2.472431e-11, 7.084448e-12, 
    3.033983e-11, 6.037646e-11, 7.167943e-12, 5.260251e-11, 1.041457e-08, 
    9.99161e-07, 1.140771e-06, 1.286535e-06, 1.360756e-06, 6.109386e-08,
  8.792704e-07, 1.745688e-08, 2.100967e-09, 1.461979e-10, 8.854328e-11, 
    5.244068e-11, 1.03595e-11, 7.01257e-11, 2.950145e-12, 1.265723e-09, 
    4.411176e-07, 1.252037e-06, 1.497069e-06, 7.120453e-07, 8.497539e-07,
  1.042618e-05, 1.59455e-06, 1.175616e-08, 2.841111e-09, 4.612581e-10, 
    4.624517e-11, 6.248234e-12, 2.689021e-11, 1.45546e-10, 2.379217e-07, 
    1.709307e-06, 2.179552e-06, 3.869544e-06, 1.345029e-06, 7.863144e-07,
  7.146296e-06, 3.147865e-06, 1.306159e-08, 6.95217e-09, 2.535754e-09, 
    4.787049e-10, 5.889142e-11, 9.307665e-12, 1.70835e-11, 1.803032e-07, 
    1.721272e-06, 4.076023e-06, 3.651073e-06, 2.281181e-06, 1.138861e-06,
  4.950431e-07, 1.375111e-06, 7.315331e-07, 4.996375e-09, 2.913612e-09, 
    1.087833e-09, 4.221962e-10, 5.773715e-11, 4.539192e-09, 1.338366e-06, 
    4.140539e-06, 4.978085e-06, 5.31665e-06, 2.760256e-06, 1.46117e-06,
  3.346499e-08, 1.143662e-07, 2.190175e-09, 2.476884e-09, 2.11256e-09, 
    1.005726e-09, 6.444998e-10, 1.163164e-10, 3.782539e-08, 1.206639e-06, 
    4.372717e-06, 6.750194e-06, 5.033864e-06, 2.730876e-06, 1.898406e-06,
  5.950496e-08, 3.670095e-09, 1.19023e-09, 1.36285e-09, 2.780945e-08, 
    1.365302e-08, 2.884311e-09, 3.880055e-10, 2.104108e-07, 1.329296e-06, 
    3.484019e-06, 6.863545e-06, 6.164505e-06, 2.801929e-06, 1.13472e-06,
  3.050971e-06, 7.843797e-07, 4.197424e-08, 2.030918e-08, 4.277036e-09, 
    1.022968e-08, 1.440282e-07, 1.852384e-07, 1.023497e-07, 1.402294e-08, 
    3.120821e-06, 9.489286e-06, 9.909138e-06, 3.924373e-06, 1.523387e-06,
  1.628798e-06, 1.77067e-06, 3.773479e-06, 2.208232e-06, 3.111038e-06, 
    7.859679e-08, 2.26775e-09, 1.204992e-08, 2.9153e-06, 8.333833e-06, 
    1.472932e-05, 1.903126e-05, 1.607266e-05, 5.967242e-06, 6.028884e-06,
  4.626702e-06, 3.991209e-06, 5.965108e-06, 7.622608e-06, 8.451071e-06, 
    7.290046e-08, 9.191187e-09, 1.795881e-07, 8.634105e-06, 2.584635e-05, 
    3.484362e-05, 2.675381e-05, 1.347714e-05, 1.016945e-05, 1.873805e-05,
  6.696996e-05, 7.315527e-05, 7.218814e-05, 2.600543e-05, 2.578211e-06, 
    9.585008e-07, 5.394504e-07, 7.148964e-07, 1.518665e-08, 6.986777e-08, 
    1.902094e-08, 3.132595e-08, 4.013383e-11, 1.098071e-10, 2.817897e-10,
  9.007435e-05, 5.998244e-05, 5.350226e-05, 2.578229e-05, 3.103831e-06, 
    7.074377e-07, 8.436845e-08, 5.038396e-08, 3.018383e-08, 9.294931e-08, 
    8.785481e-08, 1.397178e-08, 1.604589e-11, 1.252928e-10, 6.033395e-11,
  0.0001903306, 0.0001114412, 5.474881e-05, 1.550691e-05, 6.398484e-07, 
    4.138052e-07, 3.201521e-07, 1.030904e-08, 2.01754e-07, 6.465489e-07, 
    8.094961e-08, 1.599822e-08, 5.656239e-11, 4.845999e-12, 7.815113e-11,
  0.0001578212, 0.0001665595, 0.0001060838, 2.012173e-05, 6.161729e-07, 
    3.180006e-07, 5.059873e-07, 4.687026e-07, 3.781661e-06, 1.810907e-06, 
    2.404087e-07, 2.826228e-08, 4.295761e-10, 6.355478e-11, 1.217444e-11,
  7.740862e-05, 0.0001497184, 0.0001645625, 8.518976e-05, 1.599376e-05, 
    1.777425e-06, 4.395277e-06, 2.82978e-06, 7.234196e-06, 5.124268e-06, 
    7.82017e-07, 1.649334e-07, 3.834152e-10, 9.728576e-11, 1.001804e-10,
  2.083349e-05, 9.546642e-05, 0.0001748547, 0.0001424491, 6.717217e-05, 
    1.108566e-05, 1.189752e-06, 1.957434e-06, 4.19676e-06, 1.022643e-05, 
    2.346879e-06, 2.522996e-07, 2.209355e-10, 1.855405e-10, 1.057457e-10,
  9.451497e-07, 3.205496e-05, 0.0001151189, 0.0001477614, 7.703499e-05, 
    3.177539e-05, 2.848776e-06, 4.227184e-06, 4.202989e-06, 5.113019e-06, 
    2.58229e-06, 1.348345e-07, 4.281139e-11, 1.734363e-10, 2.822191e-11,
  7.028417e-10, 3.18449e-06, 5.010705e-05, 0.0001066473, 8.649187e-05, 
    2.51798e-05, 1.603371e-05, 9.713642e-06, 4.791093e-06, 7.53275e-06, 
    4.789329e-06, 1.527011e-07, 1.998242e-11, 1.676426e-11, 5.642969e-10,
  6.507555e-09, 7.279489e-08, 1.648569e-05, 5.701092e-05, 7.049643e-05, 
    3.359344e-05, 6.984884e-06, 4.041598e-07, 6.522734e-06, 1.366577e-05, 
    6.937639e-06, 2.748924e-07, 5.889694e-10, 9.709679e-13, 2.274829e-11,
  1.534273e-09, 7.679287e-09, 5.267264e-07, 2.551205e-05, 3.372705e-05, 
    2.772349e-05, 2.063449e-05, 6.938489e-06, 4.38735e-06, 4.961447e-06, 
    5.724145e-06, 1.749672e-06, 3.191555e-09, 1.612119e-11, 4.742833e-13,
  0.0002629536, 0.000327337, 0.0002796831, 8.43943e-05, 4.189324e-05, 
    3.749171e-05, 4.48276e-05, 6.802548e-05, 7.18156e-05, 3.649103e-05, 
    3.584658e-05, 4.108849e-05, 2.660202e-05, 1.207263e-05, 4.309739e-07,
  0.0002824061, 0.0003685328, 0.0003833401, 0.0002502867, 7.905001e-05, 
    4.970709e-05, 3.912603e-05, 5.376374e-05, 7.531778e-05, 4.818857e-05, 
    4.446344e-05, 5.466092e-05, 3.730725e-05, 1.217864e-05, 2.4209e-07,
  0.0003176738, 0.000417978, 0.0004759227, 0.0004332582, 0.0001609939, 
    7.894039e-05, 4.370039e-05, 4.244702e-05, 6.687126e-05, 6.292848e-05, 
    6.172029e-05, 5.106024e-05, 3.188171e-05, 7.79911e-06, 1.130485e-06,
  0.0003009436, 0.0004167696, 0.0005219222, 0.0005346392, 0.0002997324, 
    0.0001079614, 6.717224e-05, 4.078011e-05, 6.07717e-05, 8.86514e-05, 
    5.691646e-05, 5.44723e-05, 3.027012e-05, 3.751655e-06, 3.651476e-06,
  0.0002618244, 0.0003490006, 0.000523333, 0.0006117906, 0.0004075269, 
    0.0001692789, 9.70004e-05, 6.00628e-05, 7.700479e-05, 9.452184e-05, 
    5.856216e-05, 4.544654e-05, 2.49339e-05, 4.927118e-06, 3.327854e-06,
  0.0003050725, 0.0003419427, 0.0004785889, 0.0006511105, 0.0005296452, 
    0.0002675282, 0.0001398723, 9.769998e-05, 8.586414e-05, 9.448206e-05, 
    6.234678e-05, 3.696257e-05, 2.444526e-05, 2.880494e-06, 1.771341e-06,
  0.0001635013, 0.0003294996, 0.0004557154, 0.0006779462, 0.0006337779, 
    0.0003857867, 0.0002338757, 0.0001740792, 9.655831e-05, 6.572624e-05, 
    6.019131e-05, 4.101007e-05, 1.599405e-05, 2.733604e-06, 1.417745e-06,
  7.782454e-05, 0.0002147778, 0.0004768867, 0.0006947345, 0.0006448106, 
    0.0003537114, 0.0002737306, 0.0002168381, 0.0001140245, 4.902772e-05, 
    5.498938e-05, 4.144747e-05, 1.134286e-05, 3.067078e-06, 1.756707e-06,
  3.827189e-05, 0.0001323237, 0.0004136547, 0.0006527885, 0.0007020339, 
    0.0003913706, 0.0002182602, 8.78548e-05, 7.622453e-05, 9.696362e-05, 
    5.585236e-05, 3.670948e-05, 9.725995e-06, 3.186404e-06, 1.367572e-06,
  1.694112e-05, 7.937246e-05, 0.0003015854, 0.0006988994, 0.0006808973, 
    0.0004590794, 0.0003716787, 0.0002553029, 0.0002043094, 9.468588e-05, 
    6.104985e-05, 2.865944e-05, 7.671621e-06, 6.364461e-06, 1.305485e-06,
  1.375552e-09, 3.857336e-10, 5.621693e-08, 4.532421e-09, 1.711559e-07, 
    1.083329e-06, 1.293766e-06, 3.84967e-06, 3.922751e-06, 7.655061e-06, 
    2.404099e-05, 3.184579e-05, 2.918699e-05, 3.324045e-05, 3.0021e-05,
  1.601339e-08, 1.880717e-07, 1.50034e-09, 2.902858e-08, 3.955869e-07, 
    1.251423e-06, 9.952203e-07, 3.193496e-06, 4.107294e-06, 5.949633e-06, 
    2.265021e-05, 3.259339e-05, 3.637723e-05, 4.58327e-05, 4.021465e-05,
  2.212452e-05, 1.297233e-05, 9.517555e-07, 1.924575e-07, 2.250095e-06, 
    5.090574e-06, 3.616177e-06, 3.320699e-06, 3.770074e-06, 8.161214e-06, 
    2.829972e-05, 2.927877e-05, 3.966382e-05, 5.263146e-05, 3.915299e-05,
  4.181658e-05, 2.347077e-05, 6.088907e-06, 4.70946e-06, 6.901167e-06, 
    1.087802e-05, 8.885183e-06, 7.986576e-06, 6.440255e-06, 1.094272e-05, 
    2.860716e-05, 3.084864e-05, 3.908337e-05, 5.304227e-05, 3.914696e-05,
  3.385409e-05, 2.531761e-05, 3.051587e-05, 2.070989e-05, 2.34073e-05, 
    2.256512e-05, 1.774291e-05, 1.206272e-05, 8.48141e-06, 1.910539e-05, 
    4.080991e-05, 3.51989e-05, 4.314007e-05, 5.204102e-05, 3.89518e-05,
  3.304476e-05, 3.656974e-05, 4.324485e-05, 8.411804e-05, 7.500685e-05, 
    4.687485e-05, 3.620148e-05, 1.953499e-05, 1.416018e-05, 3.060081e-05, 
    4.244821e-05, 3.562337e-05, 4.153388e-05, 4.631421e-05, 3.573261e-05,
  1.452555e-05, 1.774864e-05, 2.360943e-05, 3.268692e-05, 6.307987e-05, 
    3.537617e-05, 8.32842e-06, 3.928235e-06, 1.440565e-05, 2.958464e-05, 
    4.29573e-05, 4.134233e-05, 5.143724e-05, 4.183823e-05, 3.5874e-05,
  3.225992e-06, 3.369299e-06, 5.183498e-06, 1.526392e-05, 2.121016e-05, 
    3.412059e-05, 1.926933e-05, 3.786713e-06, 1.593956e-06, 1.186744e-05, 
    4.206707e-05, 3.234372e-05, 5.678379e-05, 4.526097e-05, 3.33679e-05,
  1.020141e-06, 8.936487e-07, 1.621815e-06, 1.156213e-05, 2.673472e-05, 
    8.887187e-06, 1.003497e-05, 1.106774e-05, 1.057266e-05, 2.4885e-05, 
    3.22825e-05, 4.261149e-05, 5.517478e-05, 4.637694e-05, 3.113637e-05,
  6.720865e-08, 1.985623e-07, 3.616269e-07, 3.487149e-06, 1.955704e-05, 
    3.38362e-06, 6.332814e-06, 7.902796e-06, 2.763057e-05, 3.90908e-05, 
    5.125121e-05, 6.79093e-05, 6.256716e-05, 4.025126e-05, 3.383933e-05,
  2.414088e-11, 2.528812e-11, 4.769898e-07, 1.457688e-06, 2.104425e-07, 
    1.655348e-09, 7.920368e-10, 8.650724e-09, 9.14741e-09, 2.469269e-08, 
    4.08282e-08, 1.531946e-07, 7.114939e-06, 1.23927e-05, 1.738211e-05,
  1.683104e-10, 1.345553e-07, 6.923416e-11, 4.609846e-07, 1.010667e-06, 
    9.755222e-08, 1.605981e-07, 4.103608e-07, 5.929291e-09, 2.294644e-08, 
    1.290048e-07, 5.893305e-07, 3.235808e-06, 1.210939e-05, 1.380574e-05,
  4.886034e-06, 6.315417e-06, 4.169573e-07, 4.657636e-07, 3.105269e-06, 
    4.581795e-06, 1.999956e-06, 1.562105e-06, 1.524984e-06, 2.28009e-07, 
    5.735713e-07, 2.325194e-06, 1.263793e-05, 1.040462e-05, 6.426087e-06,
  2.447564e-05, 1.359925e-05, 5.406801e-06, 4.500208e-06, 1.388094e-05, 
    1.616008e-05, 1.342905e-05, 1.222355e-05, 8.224045e-06, 1.108584e-05, 
    1.45065e-05, 1.603765e-05, 1.356468e-05, 7.68373e-06, 7.463706e-06,
  2.567957e-05, 2.922189e-05, 9.149672e-06, 1.975432e-05, 3.545755e-05, 
    3.447182e-05, 3.21101e-05, 2.53259e-05, 2.05314e-05, 2.700731e-05, 
    1.959482e-05, 1.881256e-05, 1.736097e-05, 1.511167e-05, 9.306163e-06,
  2.390617e-05, 1.908122e-05, 3.108677e-05, 3.597607e-05, 5.246171e-05, 
    4.749025e-05, 4.084933e-05, 3.297162e-05, 2.933334e-05, 3.372751e-05, 
    3.162583e-05, 2.211122e-05, 1.962703e-05, 1.560274e-05, 1.270616e-05,
  8.082809e-06, 1.040067e-05, 2.474285e-05, 2.205219e-05, 4.200263e-05, 
    3.13687e-05, 1.67665e-05, 1.088538e-05, 1.280844e-05, 2.558881e-05, 
    3.591171e-05, 3.315726e-05, 2.607552e-05, 1.610975e-05, 1.345526e-05,
  2.802787e-06, 2.095107e-06, 1.10101e-05, 1.195841e-05, 1.007317e-05, 
    1.279001e-05, 2.152718e-05, 1.244403e-05, 3.146385e-06, 1.792629e-06, 
    1.851263e-05, 2.668038e-05, 2.243593e-05, 1.688276e-05, 1.503401e-05,
  4.146416e-06, 8.194816e-06, 7.614139e-06, 1.381208e-05, 2.23081e-05, 
    4.687465e-06, 4.34868e-06, 9.770801e-06, 2.585485e-05, 2.752752e-05, 
    2.680001e-05, 2.773044e-05, 2.282678e-05, 1.487731e-05, 1.148943e-05,
  7.249253e-06, 1.010455e-05, 1.291753e-05, 1.308503e-05, 1.59206e-05, 
    6.486097e-06, 4.025219e-06, 5.020914e-06, 3.959914e-05, 6.009463e-05, 
    6.388948e-05, 4.922907e-05, 2.963518e-05, 1.643533e-05, 1.041069e-05,
  3.859033e-08, 3.624533e-08, 1.603114e-06, 5.004043e-06, 3.066403e-06, 
    3.274206e-07, 5.320133e-07, 2.812907e-07, 1.420028e-08, 1.058399e-08, 
    1.319453e-07, 8.31868e-07, 4.80938e-06, 4.360377e-06, 8.457307e-07,
  9.39196e-08, 1.957368e-07, 2.239928e-08, 2.209464e-07, 2.584184e-06, 
    2.30214e-06, 5.161486e-07, 3.643086e-06, 1.853757e-06, 9.845794e-07, 
    2.723857e-06, 6.409212e-06, 1.079012e-05, 6.812829e-06, 1.92379e-06,
  1.657181e-06, 2.673791e-06, 1.167659e-07, 9.624441e-08, 4.139773e-06, 
    8.387896e-06, 6.177215e-06, 8.237802e-06, 5.575073e-06, 8.560658e-06, 
    1.139868e-05, 1.659614e-05, 1.294158e-05, 7.063428e-06, 3.017601e-06,
  4.107247e-06, 2.132236e-06, 1.866247e-06, 1.556892e-06, 7.770795e-06, 
    2.067481e-05, 3.261292e-05, 2.98514e-05, 2.728234e-05, 2.774402e-05, 
    2.189298e-05, 1.733285e-05, 1.416012e-05, 4.702809e-06, 2.968535e-06,
  6.891684e-07, 2.116964e-06, 2.035254e-06, 2.297603e-07, 2.493605e-06, 
    2.036335e-05, 4.095621e-05, 5.171639e-05, 5.268697e-05, 5.33893e-05, 
    4.982792e-05, 3.625207e-05, 2.162783e-05, 9.251067e-06, 2.7219e-06,
  5.80241e-07, 1.07689e-06, 2.74274e-08, 2.129325e-07, 1.934254e-06, 
    6.964876e-06, 1.295357e-05, 2.746616e-05, 4.102156e-05, 5.958773e-05, 
    6.695473e-05, 4.337548e-05, 2.371822e-05, 1.189108e-05, 4.431462e-06,
  6.23788e-09, 6.699956e-09, 5.487709e-07, 1.047487e-06, 1.994864e-06, 
    6.767195e-06, 3.814229e-06, 5.392579e-06, 7.551041e-06, 2.276326e-05, 
    4.899634e-05, 5.274948e-05, 3.606066e-05, 1.633226e-05, 5.987077e-06,
  1.321422e-08, 2.306771e-08, 2.143577e-07, 2.305295e-06, 2.217413e-06, 
    6.565112e-06, 1.259133e-05, 7.176554e-06, 2.381506e-06, 2.986473e-07, 
    1.895234e-05, 4.112109e-05, 3.640746e-05, 1.946082e-05, 9.21561e-06,
  1.018808e-08, 6.885752e-08, 3.870256e-08, 2.46115e-06, 9.690051e-06, 
    4.255406e-06, 7.156615e-07, 3.962986e-06, 3.618134e-05, 4.216662e-05, 
    4.447852e-05, 4.474313e-05, 3.169581e-05, 1.964529e-05, 9.229701e-06,
  2.208538e-09, 9.024176e-09, 4.620859e-07, 1.959171e-06, 8.745297e-06, 
    5.645571e-06, 7.050422e-06, 1.447703e-06, 3.929621e-05, 9.792556e-05, 
    0.0001764553, 0.0001031415, 3.029841e-05, 1.703015e-05, 1.023995e-05,
  2.636867e-08, 6.242567e-09, 5.2888e-07, 6.508923e-06, 3.779711e-06, 
    2.714124e-06, 3.4477e-08, 3.005058e-09, 1.310276e-10, 3.800809e-09, 
    4.064699e-08, 1.840188e-08, 5.119146e-07, 1.036383e-07, 2.058523e-09,
  3.2238e-08, 2.916779e-08, 6.86215e-09, 6.823484e-07, 1.611158e-06, 
    3.721348e-07, 3.615976e-08, 6.790782e-09, 1.880253e-10, 2.749687e-10, 
    8.086749e-09, 2.009503e-08, 1.638288e-07, 5.916667e-07, 2.098293e-08,
  3.959563e-06, 1.957755e-06, 5.54585e-09, 2.165117e-08, 8.413384e-07, 
    2.690591e-06, 1.917754e-07, 3.756294e-09, 2.161225e-10, 9.263215e-10, 
    1.787577e-08, 4.77331e-07, 5.300753e-07, 7.448974e-08, 1.95574e-08,
  1.557496e-05, 9.640959e-06, 3.893417e-07, 9.428333e-09, 1.069678e-06, 
    6.118571e-06, 5.51282e-06, 3.523885e-06, 1.571487e-06, 1.461699e-06, 
    1.874352e-06, 1.335368e-06, 7.317013e-07, 2.330968e-07, 1.376394e-08,
  1.648657e-05, 2.284687e-05, 5.187326e-06, 6.125558e-08, 1.274562e-06, 
    5.030911e-06, 1.320765e-05, 1.473682e-05, 1.760464e-05, 2.288656e-05, 
    1.310055e-05, 5.70084e-06, 3.678276e-06, 1.212619e-06, 3.664561e-07,
  1.702238e-05, 1.506689e-05, 1.39607e-06, 1.064776e-06, 2.512147e-06, 
    6.410843e-06, 8.343412e-06, 1.497619e-05, 1.867404e-05, 2.728654e-05, 
    2.373743e-05, 1.419235e-05, 5.733429e-06, 3.610652e-06, 6.783504e-07,
  1.343354e-07, 1.044625e-05, 4.660255e-06, 1.556246e-07, 5.862516e-07, 
    5.340706e-06, 6.247568e-07, 1.252225e-06, 4.840588e-06, 8.834912e-06, 
    1.564765e-05, 1.842595e-05, 1.094279e-05, 5.091505e-06, 1.727189e-06,
  1.435081e-08, 3.538336e-06, 6.253069e-06, 3.790047e-06, 1.231454e-06, 
    1.590565e-06, 3.489962e-06, 1.152928e-06, 2.106918e-09, 2.896087e-09, 
    6.261511e-06, 1.126007e-05, 1.022043e-05, 3.980969e-06, 1.13431e-06,
  7.757971e-09, 2.000083e-06, 4.549209e-07, 1.169231e-07, 3.173527e-06, 
    9.175635e-07, 5.463045e-08, 3.457421e-07, 1.79916e-06, 2.625391e-06, 
    4.32533e-06, 6.281206e-06, 8.250764e-06, 3.162214e-06, 1.859092e-06,
  3.075734e-09, 2.347235e-08, 6.122713e-08, 6.31595e-08, 2.039403e-06, 
    2.76308e-07, 2.107792e-06, 2.696306e-07, 9.528914e-06, 1.961018e-05, 
    1.651083e-05, 1.24228e-05, 6.097295e-06, 3.631099e-06, 2.263022e-06,
  1.370695e-10, 1.418143e-12, 4.52014e-13, 1.332717e-13, 5.022908e-27, 
    1.791832e-08, 1.779031e-08, 6.511651e-09, 1.214494e-09, 1.552874e-08, 
    7.679612e-08, 1.289714e-06, 4.629949e-06, 1.603495e-06, 7.798899e-07,
  1.885218e-09, 1.658649e-10, 7.036247e-12, 2.170839e-12, 4.730974e-14, 
    2.508446e-10, 1.214517e-08, 1.1618e-08, 3.972916e-09, 1.395117e-07, 
    1.701218e-07, 1.03993e-06, 3.097947e-06, 1.789622e-06, 1.124241e-07,
  1.733406e-08, 2.021438e-09, 1.653199e-10, 7.148136e-12, 5.189617e-14, 
    6.701158e-28, 2.823128e-09, 2.788546e-08, 1.42498e-09, 1.013707e-06, 
    1.716895e-06, 2.929021e-06, 2.407263e-06, 2.37822e-06, 3.071443e-07,
  6.47605e-07, 5.052564e-07, 2.904889e-10, 1.408879e-10, 2.687902e-12, 
    3.30692e-15, 4.621339e-08, 4.543412e-07, 1.036684e-06, 7.613503e-06, 
    7.791449e-06, 3.632919e-06, 2.50635e-06, 1.761153e-06, 7.044119e-07,
  6.999146e-07, 5.200855e-07, 6.366822e-08, 1.015214e-10, 4.661128e-11, 
    5.709536e-07, 7.091894e-07, 1.29005e-06, 4.339648e-06, 1.658614e-05, 
    2.072947e-05, 1.122094e-05, 4.024952e-06, 2.886831e-06, 2.195288e-06,
  2.525387e-08, 1.306891e-07, 7.468995e-09, 1.085063e-09, 3.542237e-11, 
    1.796997e-06, 7.581743e-07, 2.465181e-06, 3.063581e-06, 9.754252e-06, 
    2.152455e-05, 1.897948e-05, 9.732734e-06, 3.100859e-06, 2.388459e-06,
  3.196544e-08, 3.170018e-08, 1.505041e-08, 2.466158e-09, 1.683839e-07, 
    6.209687e-06, 3.867242e-06, 1.85027e-06, 2.56523e-06, 5.056051e-06, 
    1.157032e-05, 2.232562e-05, 1.888163e-05, 6.28255e-06, 2.061117e-06,
  6.420071e-08, 2.638503e-08, 5.291772e-08, 4.783759e-08, 2.97707e-06, 
    1.050049e-05, 1.337955e-05, 1.009025e-05, 1.659027e-06, 2.683744e-09, 
    7.508712e-06, 1.367713e-05, 2.189785e-05, 9.567561e-06, 2.503858e-06,
  7.184123e-08, 8.34113e-08, 2.774414e-07, 1.404892e-06, 2.997434e-05, 
    1.75006e-05, 1.747591e-06, 1.216205e-06, 2.16325e-06, 2.319145e-06, 
    2.978022e-06, 6.742361e-06, 1.449974e-05, 1.127081e-05, 3.704438e-06,
  6.466833e-08, 1.78203e-07, 6.980719e-08, 6.363563e-08, 1.845021e-05, 
    7.751652e-06, 3.418032e-06, 6.562708e-06, 3.186869e-06, 7.41656e-06, 
    1.063278e-05, 8.409993e-06, 7.642781e-06, 9.547006e-06, 5.525814e-06,
  3.987193e-08, 7.726021e-08, 1.130009e-07, 1.282832e-07, 2.128028e-07, 
    1.55141e-07, 9.551673e-08, 4.947258e-08, 3.365084e-08, 2.286054e-06, 
    1.45077e-05, 1.508508e-05, 1.913598e-05, 2.818884e-06, 2.821023e-07,
  7.881815e-09, 9.057094e-08, 6.585057e-08, 1.013908e-07, 6.535225e-08, 
    8.622023e-08, 6.556524e-08, 2.256566e-08, 1.771466e-08, 5.765717e-07, 
    7.161467e-06, 1.180126e-05, 1.366047e-05, 3.364148e-06, 4.649576e-07,
  2.439502e-10, 1.410802e-08, 2.370561e-08, 3.854823e-08, 3.264929e-08, 
    4.081985e-08, 4.703301e-08, 1.74675e-08, 1.653832e-08, 7.137538e-07, 
    2.208965e-06, 3.37503e-06, 7.742102e-06, 4.149476e-06, 5.966649e-07,
  1.839328e-10, 1.62837e-10, 1.042357e-09, 4.486532e-10, 4.16892e-09, 
    1.571535e-08, 1.896884e-08, 2.3497e-08, 1.905715e-08, 2.50091e-08, 
    1.24998e-08, 2.472909e-08, 1.792912e-07, 1.747592e-06, 7.277079e-07,
  1.85741e-09, 2.832791e-09, 8.997923e-11, 3.967488e-11, 1.347737e-10, 
    1.324165e-09, 7.003945e-09, 1.188053e-08, 6.713703e-09, 2.633073e-08, 
    9.098326e-09, 2.838134e-08, 1.00694e-08, 4.245528e-08, 5.963495e-07,
  2.516707e-08, 1.735811e-08, 1.007643e-08, 6.355687e-09, 1.644228e-10, 
    1.214264e-10, 1.857527e-09, 8.036013e-09, 5.384138e-09, 1.386128e-09, 
    5.983443e-09, 1.042917e-08, 2.666783e-08, 7.242924e-09, 4.802165e-08,
  2.576659e-08, 1.409372e-07, 4.540617e-08, 2.226045e-09, 1.500925e-09, 
    7.700326e-11, 1.848568e-10, 1.866563e-09, 3.83358e-09, 5.219149e-09, 
    1.212831e-09, 1.716938e-09, 1.00251e-08, 1.150784e-08, 3.412008e-09,
  2.898599e-08, 4.027599e-08, 1.539048e-07, 1.028834e-08, 2.986477e-10, 
    9.849611e-11, 5.930013e-11, 1.587713e-08, 7.662599e-10, 5.879668e-10, 
    6.201679e-10, 2.737633e-11, 3.789971e-10, 5.518625e-09, 2.194003e-08,
  1.741191e-08, 1.280967e-08, 2.090855e-07, 1.68432e-08, 5.52775e-10, 
    2.033782e-10, 1.374911e-10, 2.432321e-11, 1.290562e-12, 4.176332e-11, 
    9.0066e-11, 2.563853e-11, 1.122512e-09, 5.947944e-10, 2.164991e-08,
  4.424526e-09, 1.300574e-08, 1.054006e-08, 1.167271e-08, 9.46352e-09, 
    1.58833e-08, 1.884324e-09, 4.26956e-11, 2.530841e-12, 8.221283e-12, 
    2.426011e-11, 9.14274e-12, 6.927019e-11, 7.505462e-10, 2.365211e-08,
  1.498588e-06, 4.165647e-06, 1.759777e-05, 3.464757e-05, 3.512602e-05, 
    4.484007e-05, 9.269892e-05, 0.0001275773, 0.0001956761, 0.0002648847, 
    0.000291225, 0.0002868315, 0.0002803771, 0.0002680842, 0.0001979076,
  1.499333e-07, 8.412453e-07, 5.684032e-06, 1.251711e-05, 1.145394e-05, 
    7.381131e-06, 2.364221e-05, 6.599976e-05, 0.0001142588, 0.0001785899, 
    0.0002244504, 0.000234867, 0.00021551, 0.0002013469, 0.0001581416,
  7.029927e-08, 6.828812e-07, 5.593703e-07, 2.251026e-06, 2.968818e-06, 
    5.126975e-06, 6.607079e-06, 3.473609e-05, 6.54117e-05, 0.0001128906, 
    0.0001621675, 0.0002018345, 0.0001860157, 0.0001589769, 0.0001124825,
  9.75717e-08, 2.700106e-07, 1.351778e-07, 2.352011e-07, 7.146789e-07, 
    1.933736e-06, 3.686353e-06, 1.210393e-05, 2.11768e-05, 5.681117e-05, 
    9.621902e-05, 0.0001497194, 0.0001533454, 0.0001282835, 6.822059e-05,
  1.14921e-07, 8.558056e-08, 8.534532e-08, 6.729864e-08, 6.550351e-08, 
    1.850303e-07, 2.218889e-06, 3.50475e-06, 9.664501e-06, 1.709552e-05, 
    3.211913e-05, 6.458579e-05, 0.0001049203, 9.218919e-05, 3.959415e-05,
  1.077101e-07, 6.029493e-08, 1.329796e-08, 3.730373e-08, 6.404535e-08, 
    2.048304e-08, 4.875615e-07, 9.630338e-07, 4.821838e-06, 8.260711e-06, 
    9.649463e-06, 1.28531e-05, 2.047044e-05, 5.032965e-05, 3.369695e-05,
  1.031456e-07, 5.850651e-08, 1.198074e-08, 5.972327e-09, 7.67282e-09, 
    8.797834e-09, 7.459216e-08, 4.110961e-08, 7.572629e-07, 5.293141e-06, 
    6.661477e-06, 3.516068e-06, 3.016399e-06, 7.602658e-06, 1.120173e-05,
  6.455492e-08, 2.452301e-08, 8.641308e-09, 6.123288e-09, 6.624733e-09, 
    2.725673e-09, 1.028186e-08, 1.250732e-07, 3.224673e-06, 2.938019e-06, 
    3.674828e-06, 4.203657e-08, 2.458667e-07, 2.383356e-07, 3.55522e-07,
  3.041497e-08, 4.385111e-09, 5.033857e-09, 4.672855e-09, 9.640796e-09, 
    3.288992e-08, 3.019018e-08, 1.264118e-06, 1.380989e-06, 1.365283e-06, 
    1.529402e-06, 3.709723e-08, 1.181577e-07, 1.513452e-07, 1.301483e-07,
  8.211177e-09, 3.122725e-09, 2.592806e-09, 2.428599e-09, 9.952548e-09, 
    3.307052e-08, 1.596652e-06, 3.207372e-06, 8.271933e-06, 3.936455e-06, 
    1.625122e-06, 1.187131e-07, 6.273319e-07, 1.291545e-07, 1.685336e-07,
  8.84546e-05, 9.454269e-06, 1.997916e-05, 0.000177988, 0.000395689, 
    0.0006173447, 0.000621479, 0.0003714107, 0.0001317371, 6.367335e-05, 
    6.237531e-05, 8.824121e-05, 0.0001201771, 0.000127038, 0.0001115516,
  4.044519e-05, 2.398895e-05, 1.583338e-05, 0.0001318412, 0.0003811334, 
    0.000667438, 0.0007584492, 0.0005026834, 0.00021939, 0.0001163493, 
    9.856001e-05, 0.0001174108, 0.0001693387, 0.0002003243, 0.0001771079,
  6.941694e-05, 3.124048e-05, 2.609227e-05, 0.0001239235, 0.0003992605, 
    0.0006716773, 0.0008539619, 0.0006622829, 0.0003230795, 0.0001688515, 
    0.0001130808, 0.0001151894, 0.0001893552, 0.0002600163, 0.0002671944,
  6.285108e-05, 3.133906e-05, 2.078289e-05, 0.0001032238, 0.0003763756, 
    0.0006416475, 0.0008721757, 0.0007422638, 0.0004496283, 0.0002076187, 
    0.0001138928, 0.0001048142, 0.0001538395, 0.000279768, 0.0003356914,
  4.481409e-05, 1.953075e-05, 1.564176e-05, 9.105739e-05, 0.0003387103, 
    0.0005421619, 0.0007670287, 0.0007543484, 0.0005208175, 0.0002721492, 
    0.0001386943, 9.403878e-05, 0.0001154209, 0.0002325238, 0.0003422567,
  3.861419e-05, 1.224695e-05, 1.350818e-05, 0.0001137351, 0.0003747598, 
    0.0005364592, 0.0006227231, 0.0006373542, 0.0005493804, 0.0003375174, 
    0.000167179, 9.268933e-05, 9.60328e-05, 0.0001581566, 0.0003044317,
  1.825774e-05, 1.838339e-05, 3.350576e-05, 0.0001944128, 0.0005390811, 
    0.0007016247, 0.0005490906, 0.0003876715, 0.0004356362, 0.0003702547, 
    0.0001937028, 9.658878e-05, 7.192764e-05, 0.0001011291, 0.0002144881,
  2.089533e-05, 1.675945e-05, 6.243995e-05, 0.0003341486, 0.0007030753, 
    0.0008120388, 0.0006616186, 0.0004437374, 0.000417336, 0.0003565479, 
    0.0002236705, 0.0001088583, 5.985044e-05, 7.37522e-05, 0.0001423551,
  1.768034e-05, 1.661258e-05, 0.0001198968, 0.0004846736, 0.0007950716, 
    0.0009566936, 0.0006830281, 0.000427389, 0.0003390365, 0.0003329773, 
    0.0002330062, 0.0001308292, 7.051479e-05, 6.699358e-05, 0.000113225,
  8.928007e-06, 3.337877e-05, 0.0002690961, 0.0005788957, 0.0008031215, 
    0.0008275356, 0.0006789246, 0.0004636057, 0.0003417358, 0.0003015872, 
    0.0002080303, 0.0001178832, 7.226656e-05, 6.323419e-05, 0.000108019,
  2.420865e-09, 1.850009e-08, 3.449753e-09, 5.160294e-10, 2.60174e-10, 
    3.623752e-10, 3.633948e-10, 9.293156e-11, 9.32221e-10, 2.853668e-10, 
    2.428903e-10, 4.996679e-11, 1.574883e-09, 1.471443e-07, 2.550832e-06,
  2.079569e-08, 1.915967e-08, 2.603866e-08, 2.946607e-09, 7.092017e-09, 
    4.062486e-08, 7.700114e-10, 5.312526e-09, 1.402707e-10, 1.00889e-09, 
    1.36434e-09, 2.979345e-11, 1.79899e-10, 1.193862e-08, 7.923052e-07,
  1.345944e-07, 5.295874e-08, 2.781463e-08, 9.603309e-09, 2.031548e-09, 
    1.260983e-08, 3.921368e-07, 1.845753e-07, 2.098622e-08, 1.934252e-07, 
    2.727691e-07, 1.21848e-08, 1.750999e-08, 2.745069e-11, 1.33173e-07,
  1.694945e-07, 1.623129e-07, 6.48926e-08, 3.019079e-08, 5.440561e-09, 
    3.477378e-08, 2.81615e-07, 4.172194e-07, 2.59551e-07, 1.014881e-08, 
    2.131414e-07, 4.378438e-08, 2.179775e-10, 2.091507e-13, 2.648159e-08,
  1.165073e-07, 1.223842e-07, 6.208326e-08, 2.666165e-08, 2.037483e-08, 
    2.935635e-07, 2.246211e-07, 5.45664e-07, 3.120405e-07, 9.399462e-08, 
    1.73669e-08, 1.108174e-07, 4.77279e-10, 3.840028e-22, 1.060246e-09,
  4.724249e-08, 2.847267e-08, 3.718676e-08, 3.71043e-08, 2.035032e-07, 
    6.869287e-07, 9.580051e-07, 9.050422e-07, 2.494439e-07, 2.034569e-07, 
    5.455838e-11, 8.75312e-08, 3.484664e-08, 7.116143e-13, 1.819456e-09,
  7.103624e-09, 1.202931e-08, 1.887962e-08, 8.694771e-08, 5.847868e-07, 
    1.165071e-05, 1.434958e-06, 4.378538e-07, 6.949274e-11, 1.727021e-12, 
    4.693168e-11, 1.17924e-07, 4.500442e-08, 6.304554e-10, 1.626555e-15,
  1.157195e-07, 1.57134e-07, 2.25149e-07, 6.815415e-07, 4.622094e-06, 
    2.429165e-05, 1.486615e-05, 5.509937e-06, 3.307675e-08, 4.406083e-13, 
    5.985309e-12, 4.267099e-08, 1.107881e-07, 8.341119e-11, 1.70117e-15,
  2.526227e-06, 2.852205e-06, 3.1194e-06, 5.060848e-06, 4.135637e-05, 
    1.800534e-05, 1.68864e-06, 5.066341e-08, 3.30132e-08, 2.302122e-11, 
    9.069804e-11, 1.025436e-09, 7.922035e-11, 4.694466e-09, 2.501377e-16,
  1.006844e-05, 1.891965e-05, 4.55298e-05, 7.572023e-05, 9.409209e-05, 
    7.02855e-05, 2.564676e-05, 6.391875e-07, 1.270445e-06, 3.749469e-07, 
    1.395026e-07, 3.306532e-09, 5.046257e-10, 5.932983e-16, 6.725643e-17,
  2.946197e-05, 2.124922e-05, 1.775954e-06, 6.293469e-06, 1.649594e-05, 
    0.0001374627, 0.0002020375, 0.0003220496, 0.0005522202, 0.0006646617, 
    0.0005803456, 0.0003329227, 0.0001081759, 1.474879e-05, 1.817572e-06,
  1.086611e-05, 2.865946e-05, 4.858957e-06, 1.04013e-06, 1.020276e-05, 
    4.054767e-05, 0.0001588591, 0.0002193276, 0.0003895519, 0.0005666022, 
    0.0006077758, 0.0004638824, 0.0002011922, 4.130379e-05, 1.911867e-06,
  7.998457e-08, 6.497459e-06, 1.415616e-05, 1.298612e-06, 4.322164e-06, 
    1.366953e-05, 6.692202e-05, 0.0001795085, 0.0002590022, 0.0003968035, 
    0.0005003688, 0.000508846, 0.0003202754, 0.0001118281, 1.011022e-05,
  1.906013e-07, 1.136204e-07, 3.78628e-07, 1.638208e-07, 3.247112e-07, 
    7.972873e-06, 3.405703e-05, 0.0001076065, 0.0002107448, 0.0003064086, 
    0.0003852836, 0.0003879124, 0.0003204857, 0.0001629179, 2.486188e-05,
  1.189796e-07, 1.48214e-07, 1.059069e-07, 3.674632e-08, 3.501033e-08, 
    2.254265e-06, 1.03868e-05, 4.705787e-05, 0.0001297723, 0.0002407343, 
    0.0003001125, 0.0002814335, 0.0002116431, 0.0001473849, 4.556197e-05,
  6.965321e-08, 1.130672e-07, 9.678845e-08, 9.425288e-08, 2.336207e-08, 
    4.197461e-08, 5.749707e-06, 1.881405e-05, 6.393973e-05, 0.0001420813, 
    0.0002251882, 0.0002042515, 0.0001123677, 8.721971e-05, 4.400657e-05,
  5.216982e-09, 3.513879e-08, 6.488123e-08, 6.523238e-08, 5.436273e-08, 
    5.878771e-08, 4.210806e-07, 5.413809e-06, 2.000713e-05, 6.775914e-05, 
    0.0001567396, 0.0001810454, 7.11023e-05, 2.877015e-05, 1.760958e-05,
  4.764044e-10, 6.918025e-09, 3.037434e-08, 6.306139e-08, 7.810038e-08, 
    7.627397e-08, 3.148944e-08, 5.016399e-06, 1.319852e-05, 2.71317e-05, 
    8.748893e-05, 0.0001471065, 7.221643e-05, 1.239207e-05, 6.25611e-06,
  1.349338e-11, 6.936222e-10, 6.511704e-09, 3.799565e-08, 6.911071e-08, 
    6.630264e-08, 4.85931e-08, 1.578947e-08, 3.395179e-06, 1.096823e-05, 
    3.578894e-05, 0.0001018381, 6.99973e-05, 1.132711e-05, 4.649915e-06,
  2.405301e-11, 6.049793e-12, 3.017573e-10, 6.228562e-09, 4.644712e-08, 
    5.839201e-08, 5.134834e-08, 1.816914e-08, 1.11912e-08, 2.013038e-06, 
    8.509606e-06, 4.521277e-05, 6.427887e-05, 9.308204e-06, 2.185122e-06,
  3.246807e-07, 3.820106e-06, 3.82182e-05, 0.0002948206, 0.0006095217, 
    0.0009117587, 0.0008595541, 0.0005071966, 0.000212489, 0.0001120216, 
    7.747645e-05, 5.139329e-05, 6.998212e-05, 9.219259e-05, 9.171508e-05,
  9.534997e-08, 2.221249e-06, 1.052979e-05, 0.0001500613, 0.0004946885, 
    0.0007163944, 0.0009236324, 0.0008050368, 0.0004512319, 0.0003062582, 
    0.0001865315, 7.555448e-05, 8.278816e-05, 0.0001226391, 0.0001450044,
  2.637591e-06, 2.040097e-06, 1.909198e-06, 5.54513e-05, 0.0003684509, 
    0.0005852344, 0.0008226803, 0.0009038794, 0.0007505396, 0.0004835738, 
    0.0003270904, 0.0001517213, 9.992997e-05, 0.0001669678, 0.0001729029,
  2.710413e-06, 4.485522e-06, 1.954008e-07, 3.028617e-06, 0.0001941905, 
    0.0005038182, 0.0006450826, 0.0008677912, 0.0008504164, 0.0006570906, 
    0.0004366337, 0.0002319019, 0.000152548, 0.0002343776, 0.0002035522,
  1.280476e-07, 5.805729e-07, 1.76156e-07, 1.057692e-07, 7.111916e-05, 
    0.0003909732, 0.0005123925, 0.0006653545, 0.0008810443, 0.0008160625, 
    0.0005715906, 0.0003253569, 0.000272815, 0.0003219135, 0.000235991,
  3.510153e-07, 1.616832e-07, 1.118786e-07, 1.243568e-07, 3.451768e-06, 
    0.0002336634, 0.0004584681, 0.0005018268, 0.0007501775, 0.0008740691, 
    0.0007194151, 0.0004172866, 0.0003815225, 0.0004079277, 0.0002719626,
  1.248449e-06, 7.412522e-07, 7.616081e-08, 1.092266e-07, 1.2647e-07, 
    9.155926e-05, 0.0002712494, 0.0003390068, 0.0005405201, 0.0008658263, 
    0.0008347092, 0.0005561388, 0.0004303445, 0.0004330172, 0.0002848342,
  1.842378e-06, 8.258141e-07, 6.665206e-08, 9.354172e-08, 1.414881e-07, 
    6.797748e-06, 0.0002237635, 0.0004949839, 0.0005843159, 0.0007773219, 
    0.0009544563, 0.0007910582, 0.0005113795, 0.0003848982, 0.0002648848,
  3.882107e-06, 3.151779e-06, 1.626592e-06, 6.951597e-08, 8.605985e-08, 
    4.129941e-07, 4.698167e-05, 0.0002780234, 0.0004607854, 0.0006051087, 
    0.0009474885, 0.001061071, 0.0007320502, 0.0003934288, 0.0002719969,
  5.279878e-06, 3.618663e-06, 1.855645e-06, 3.894404e-08, 6.148046e-08, 
    9.275578e-08, 1.837544e-05, 0.0001309516, 0.0003204408, 0.000486739, 
    0.000729477, 0.001219037, 0.001009467, 0.0005296696, 0.0003159663,
  1.443246e-08, 4.144135e-08, 1.039849e-08, 2.688006e-09, 4.438205e-09, 
    3.813689e-09, 1.357231e-09, 3.758335e-10, 3.171336e-10, 2.547675e-08, 
    4.16877e-07, 1.52968e-06, 2.016491e-06, 2.016632e-06, 5.171499e-07,
  1.111072e-08, 4.308281e-09, 3.084448e-09, 2.600045e-07, 2.378789e-07, 
    9.159766e-08, 8.252823e-09, 1.929613e-09, 2.107144e-09, 1.194574e-06, 
    1.297574e-06, 2.371502e-06, 8.490088e-06, 4.88185e-06, 7.681583e-07,
  4.368793e-06, 7.356334e-06, 1.208847e-07, 9.250542e-07, 7.509294e-07, 
    1.920649e-06, 6.552949e-07, 1.719724e-07, 1.287367e-07, 1.971276e-06, 
    4.050675e-06, 1.355468e-05, 1.368018e-05, 1.535129e-05, 8.284382e-06,
  7.744196e-06, 9.560911e-06, 6.766145e-06, 4.977464e-06, 1.959976e-06, 
    3.780101e-06, 3.556423e-06, 4.837457e-06, 1.945957e-06, 3.192693e-06, 
    7.419234e-06, 1.576854e-05, 2.632271e-05, 8.936819e-06, 6.879344e-06,
  1.088398e-06, 7.187018e-06, 5.294661e-06, 2.60169e-06, 1.363696e-06, 
    1.296494e-06, 9.663387e-07, 6.736732e-07, 2.360801e-06, 5.235177e-06, 
    1.615245e-05, 1.523608e-05, 1.02209e-05, 1.257049e-05, 6.968411e-06,
  1.636609e-05, 1.087988e-05, 1.884501e-06, 1.692766e-06, 3.359832e-06, 
    1.671653e-06, 1.445856e-06, 6.039759e-07, 1.074032e-07, 6.208853e-06, 
    2.221947e-05, 1.817621e-05, 1.055718e-05, 7.583137e-06, 7.196521e-06,
  3.290876e-05, 2.482113e-05, 1.481707e-05, 8.443641e-06, 7.655067e-06, 
    3.387195e-07, 1.683417e-07, 2.189222e-08, 1.461361e-07, 1.054134e-05, 
    2.985456e-05, 2.978671e-05, 1.607608e-05, 9.378688e-06, 4.703585e-06,
  2.578934e-05, 3.341094e-05, 1.960758e-05, 2.26881e-05, 4.382568e-06, 
    1.80977e-06, 5.137388e-07, 1.077645e-06, 6.913511e-06, 1.084717e-05, 
    3.435364e-05, 4.579473e-05, 2.298495e-05, 1.327082e-05, 5.924654e-06,
  2.139345e-05, 2.948179e-05, 3.023177e-05, 3.515715e-05, 3.402228e-05, 
    4.673677e-06, 1.074407e-06, 2.584104e-07, 1.21832e-05, 2.015553e-05, 
    3.695176e-05, 5.150141e-05, 2.55795e-05, 1.254981e-05, 9.910782e-06,
  1.946118e-05, 2.710447e-05, 2.866232e-05, 2.634391e-05, 2.936372e-05, 
    1.928897e-05, 8.819191e-06, 4.288918e-06, 2.282172e-05, 3.415653e-05, 
    4.581203e-05, 5.878464e-05, 3.698731e-05, 1.352381e-05, 9.337921e-06,
  6.126892e-05, 6.220782e-05, 3.456406e-05, 7.190294e-06, 4.083848e-07, 
    9.797656e-08, 6.758076e-08, 1.723892e-08, 1.778649e-08, 2.028693e-06, 
    7.038176e-06, 1.302173e-05, 9.493486e-06, 8.21614e-07, 8.67163e-08,
  4.884229e-05, 3.69297e-05, 3.299263e-05, 1.084018e-05, 2.456303e-06, 
    8.993268e-07, 2.131971e-07, 4.418379e-08, 4.485891e-08, 6.7301e-07, 
    5.683819e-06, 1.106829e-05, 6.799385e-06, 2.407215e-06, 1.247693e-06,
  4.040981e-05, 2.356704e-05, 1.753255e-05, 1.068586e-05, 3.801735e-06, 
    1.083049e-06, 5.659343e-07, 6.224577e-07, 1.550177e-06, 1.194217e-06, 
    2.15072e-06, 4.818748e-06, 5.332721e-06, 2.295401e-06, 9.443844e-08,
  2.809319e-05, 1.471508e-05, 8.438227e-06, 5.80596e-06, 2.134543e-06, 
    5.058484e-06, 7.079276e-07, 4.604312e-07, 7.049897e-07, 7.107356e-07, 
    1.609203e-06, 7.405681e-07, 6.670481e-07, 2.937416e-07, 5.596937e-09,
  5.980241e-06, 4.708356e-06, 4.89884e-06, 3.066977e-06, 2.997713e-06, 
    3.423388e-06, 1.535138e-06, 2.214675e-07, 4.060211e-07, 1.625811e-06, 
    2.136485e-06, 3.107823e-07, 3.023282e-07, 7.30463e-08, 6.452768e-08,
  2.837943e-06, 5.09154e-06, 1.922635e-06, 3.045873e-06, 3.384438e-06, 
    1.666197e-06, 5.410037e-07, 3.117615e-07, 1.293142e-07, 1.400186e-06, 
    1.345443e-06, 1.383565e-07, 9.952356e-08, 4.81873e-07, 7.234497e-08,
  4.347775e-06, 5.830959e-06, 2.694656e-06, 7.909885e-06, 9.687468e-07, 
    6.082046e-07, 6.728634e-08, 6.157775e-09, 7.943956e-10, 2.65926e-08, 
    1.055271e-06, 9.332696e-07, 1.632591e-08, 1.397811e-06, 2.277678e-07,
  7.10927e-06, 8.463781e-06, 6.670979e-06, 5.749345e-06, 2.278872e-07, 
    2.056692e-07, 3.399645e-07, 3.501794e-07, 2.140784e-07, 1.78908e-08, 
    1.687186e-06, 5.701705e-07, 2.619612e-07, 7.295412e-07, 6.832209e-07,
  7.927331e-06, 7.988532e-06, 8.214795e-06, 3.445938e-06, 1.169743e-05, 
    6.155691e-07, 8.496261e-08, 4.74177e-07, 2.948531e-06, 3.227264e-06, 
    4.558273e-06, 4.730015e-06, 3.053161e-06, 8.761373e-07, 1.57471e-06,
  9.080702e-06, 7.857999e-06, 9.088941e-06, 4.165802e-06, 1.009443e-05, 
    4.200648e-06, 2.440072e-06, 5.123784e-07, 5.898629e-06, 4.92828e-06, 
    6.585256e-06, 2.036967e-06, 9.362116e-07, 2.77203e-06, 2.123472e-06,
  2.759526e-05, 4.682187e-05, 5.373355e-05, 4.440376e-05, 2.065562e-05, 
    1.352987e-05, 1.382928e-05, 1.203794e-05, 1.506061e-05, 7.583151e-05, 
    0.0001515352, 7.20124e-05, 1.366142e-05, 1.924073e-06, 2.275746e-06,
  3.620249e-05, 5.012611e-05, 6.707556e-05, 3.904905e-05, 1.430608e-05, 
    1.035551e-05, 1.421408e-05, 2.015988e-05, 3.343709e-05, 0.000151239, 
    0.0002021796, 6.933306e-05, 7.151952e-06, 1.629425e-06, 3.34105e-06,
  3.461208e-05, 5.287075e-05, 6.489002e-05, 3.458062e-05, 1.545963e-05, 
    8.138041e-06, 1.310872e-05, 2.093192e-05, 7.736326e-05, 0.0002090245, 
    0.0001822133, 4.575269e-05, 5.204606e-06, 2.057051e-06, 1.366782e-06,
  2.821456e-05, 3.596954e-05, 3.389976e-05, 2.55107e-05, 1.419635e-05, 
    7.357982e-06, 7.389351e-06, 2.015683e-05, 0.0001148805, 0.000219062, 
    0.0001313544, 2.471764e-05, 7.115785e-06, 5.762272e-07, 1.715602e-06,
  1.499717e-05, 2.193533e-05, 3.008947e-05, 1.880842e-05, 1.313842e-05, 
    6.082471e-06, 4.605992e-06, 1.701373e-05, 0.0001016871, 0.0001713047, 
    7.941991e-05, 7.496535e-06, 1.156498e-06, 1.47007e-06, 4.618505e-06,
  1.07863e-05, 1.783051e-05, 1.294277e-05, 1.215782e-05, 1.014836e-05, 
    7.075329e-06, 8.679101e-06, 1.365051e-05, 8.524752e-05, 0.0001079307, 
    3.376321e-05, 5.101888e-06, 2.946286e-06, 1.745012e-06, 1.639531e-06,
  5.843093e-06, 7.467724e-06, 7.01311e-06, 8.32414e-06, 7.707917e-06, 
    9.782954e-06, 1.105707e-05, 1.422469e-05, 4.559388e-05, 6.058113e-05, 
    2.478036e-05, 8.035042e-06, 1.509602e-06, 1.160056e-06, 8.421976e-07,
  3.654672e-06, 3.072452e-06, 5.133434e-06, 5.478339e-06, 6.313603e-06, 
    1.239924e-05, 1.910116e-05, 1.92179e-05, 3.167262e-05, 3.091011e-05, 
    1.446501e-05, 6.73507e-06, 1.813823e-06, 2.407939e-07, 2.111432e-06,
  3.146887e-06, 3.381415e-06, 3.037329e-06, 2.399398e-06, 1.651492e-05, 
    1.556661e-05, 1.423326e-05, 1.543602e-05, 3.308945e-05, 2.580977e-05, 
    9.447604e-06, 5.366308e-06, 7.901079e-07, 2.193321e-06, 1.45238e-06,
  5.643808e-06, 3.443819e-06, 4.281997e-06, 3.019024e-06, 8.957442e-06, 
    1.153601e-05, 3.29668e-05, 4.312763e-05, 4.905623e-05, 2.443696e-05, 
    1.345294e-05, 4.585153e-06, 3.675351e-06, 3.84199e-06, 1.77163e-06,
  7.26697e-06, 1.830075e-05, 1.322438e-05, 1.655396e-06, 5.519847e-07, 
    1.666789e-06, 2.107634e-05, 8.079129e-05, 0.0002406915, 0.0002610059, 
    0.0001722827, 5.646107e-05, 2.625365e-05, 2.420868e-06, 2.058682e-06,
  1.263531e-05, 1.32978e-05, 7.077829e-06, 1.02206e-06, 1.653253e-07, 
    2.268632e-06, 2.750555e-05, 9.892543e-05, 0.0002604635, 0.0003027167, 
    0.0001593382, 2.537858e-05, 4.785519e-06, 3.395511e-06, 3.491005e-06,
  1.691745e-05, 1.391634e-05, 5.553222e-06, 3.808409e-06, 5.71789e-06, 
    2.990591e-06, 3.770367e-05, 0.0001155095, 0.0002501862, 0.0003583805, 
    0.0001737079, 2.021523e-05, 4.352576e-06, 3.699241e-06, 3.277039e-06,
  1.872039e-05, 1.720893e-05, 3.452963e-06, 8.283859e-06, 1.681059e-05, 
    5.535655e-06, 5.281791e-05, 0.0001365224, 0.0002944068, 0.00047041, 
    0.0001912011, 1.433538e-05, 4.715834e-06, 2.316466e-06, 2.783307e-06,
  4.764596e-06, 5.012999e-06, 9.924062e-07, 9.721557e-06, 2.088898e-05, 
    2.768864e-05, 8.438202e-05, 0.0001873932, 0.0004165897, 0.0006096872, 
    0.0002210905, 1.057229e-05, 4.164527e-06, 4.015058e-06, 3.620278e-06,
  2.945795e-06, 5.751913e-07, 6.724009e-08, 2.545565e-06, 1.362126e-05, 
    5.241261e-05, 0.0001273814, 0.0002664984, 0.0005850584, 0.0006242035, 
    0.000133729, 4.239408e-06, 1.82271e-06, 2.969393e-06, 2.743429e-06,
  1.728336e-08, 1.179978e-08, 1.938071e-08, 1.936332e-07, 5.116749e-06, 
    0.0001175299, 0.0001791898, 0.0003191717, 0.0006110467, 0.0005232824, 
    6.149147e-05, 8.619581e-06, 2.160504e-06, 1.67954e-06, 6.728295e-07,
  9.431494e-08, 5.996088e-08, 2.118478e-08, 9.644583e-09, 2.93763e-06, 
    0.0001707167, 0.0002822127, 0.0004087508, 0.0005905843, 0.0003419764, 
    2.456503e-05, 6.279784e-06, 4.153639e-06, 4.376139e-06, 1.651435e-06,
  7.672119e-08, 1.801699e-07, 2.668328e-08, 8.096556e-09, 3.736704e-06, 
    0.0002389354, 0.0004427845, 0.0004956376, 0.0004871016, 0.0001916651, 
    2.06794e-05, 1.168206e-05, 9.070821e-06, 8.784339e-06, 3.523022e-06,
  5.150696e-07, 4.50027e-08, 1.443896e-07, 1.351153e-08, 5.766158e-06, 
    0.00024058, 0.0005000246, 0.0006143136, 0.0004691677, 0.0001605039, 
    2.638545e-05, 2.011584e-05, 1.316756e-05, 8.352868e-06, 6.674812e-06,
  1.571618e-07, 3.500863e-08, 3.419112e-09, 1.190531e-08, 2.042381e-06, 
    6.141353e-06, 2.575064e-06, 4.848841e-08, 6.008133e-07, 6.90362e-06, 
    4.192882e-05, 0.0003247512, 0.000599073, 0.0006585907, 0.0003673836,
  2.775848e-08, 5.617883e-06, 7.036998e-10, 9.369497e-09, 1.800551e-07, 
    6.005566e-07, 2.658824e-07, 5.292972e-07, 5.147787e-06, 3.765207e-05, 
    9.455859e-05, 0.0003074385, 0.0004924457, 0.0006068244, 0.0003505153,
  1.452029e-05, 1.232227e-05, 7.322321e-08, 1.58728e-08, 1.871282e-06, 
    5.458998e-07, 6.60587e-07, 2.39395e-06, 1.244514e-05, 5.800492e-05, 
    0.0001294539, 0.000303721, 0.0003964811, 0.0005327283, 0.0003051599,
  3.507629e-05, 4.226783e-05, 2.076385e-05, 2.304376e-06, 1.13829e-05, 
    3.929843e-06, 2.532692e-06, 7.806405e-06, 1.929878e-05, 6.270695e-05, 
    0.0001368753, 0.0002643525, 0.0003416608, 0.0004675235, 0.0002702585,
  4.582795e-05, 3.504059e-05, 2.789216e-05, 9.473763e-06, 2.730835e-05, 
    6.842296e-06, 5.266947e-06, 1.616027e-05, 2.454077e-05, 5.277219e-05, 
    0.0001154099, 0.0002143215, 0.000333027, 0.0004416007, 0.0002391532,
  2.316134e-05, 1.297983e-05, 7.997124e-07, 1.622889e-06, 2.544873e-05, 
    1.571785e-05, 6.584256e-06, 2.901833e-05, 4.461043e-05, 6.60084e-05, 
    8.776422e-05, 0.0001781814, 0.0003160327, 0.0004014608, 0.000226697,
  5.988091e-08, 3.757015e-08, 1.160118e-08, 2.913692e-07, 3.708411e-06, 
    4.115902e-05, 3.492438e-05, 5.178973e-05, 7.02685e-05, 8.669175e-05, 
    7.517759e-05, 0.0001431299, 0.0002752632, 0.0003971694, 0.0002162917,
  2.512208e-07, 6.769401e-08, 6.114157e-09, 6.380345e-10, 7.130666e-06, 
    7.641337e-05, 9.243011e-05, 9.407061e-05, 9.297818e-05, 0.000107537, 
    6.1149e-05, 0.0001200827, 0.0002353373, 0.0003708297, 0.0001754965,
  1.375056e-07, 2.704477e-07, 9.038778e-08, 6.924418e-08, 2.770728e-05, 
    0.0001026776, 0.0001221775, 8.570479e-05, 0.0001541041, 0.0001357006, 
    6.805555e-05, 9.542447e-05, 0.0002070854, 0.0003435558, 0.0001180675,
  6.472079e-08, 4.063349e-08, 1.876308e-06, 3.301448e-06, 8.342622e-05, 
    0.0002057906, 0.0002365765, 0.0002335917, 0.0002637806, 0.0001588099, 
    8.008664e-05, 8.461904e-05, 0.0002148832, 0.0003012411, 5.847547e-05,
  1.549802e-09, 3.578579e-10, 4.558786e-11, 8.935969e-12, 1.038321e-09, 
    2.143064e-07, 1.366822e-11, 2.047547e-10, 1.582568e-09, 5.963274e-10, 
    2.120558e-08, 2.257211e-05, 7.291668e-05, 7.811791e-05, 6.944401e-05,
  2.13024e-09, 1.584988e-08, 4.356258e-10, 2.418965e-12, 1.023917e-10, 
    6.509243e-09, 4.049312e-11, 2.852643e-11, 7.94375e-10, 1.165261e-10, 
    3.946878e-08, 3.850897e-05, 0.0001149475, 0.0001028891, 0.0001424949,
  7.440423e-09, 3.920253e-08, 1.374818e-09, 4.055847e-12, 2.78145e-13, 
    1.814077e-13, 1.517198e-12, 8.878473e-12, 1.830597e-10, 2.484202e-10, 
    8.247129e-07, 5.673386e-05, 0.0001335897, 0.000129029, 0.0001867975,
  3.660047e-09, 2.95373e-07, 3.546172e-08, 1.581566e-09, 6.196541e-12, 
    1.277134e-14, 1.297827e-12, 4.064129e-12, 5.250657e-12, 3.003283e-09, 
    8.041587e-07, 4.904377e-05, 0.0001567524, 0.0001584418, 0.0002247681,
  1.277253e-07, 5.257052e-09, 1.210629e-06, 1.44557e-10, 4.751393e-12, 
    1.043149e-12, 3.334291e-13, 4.374067e-12, 9.446802e-12, 7.80276e-09, 
    3.405097e-07, 3.941041e-05, 0.0001522539, 0.0001701012, 0.0002335905,
  2.966825e-06, 2.186336e-08, 1.031458e-09, 1.123591e-11, 5.620049e-12, 
    1.584716e-12, 2.025905e-22, 9.46638e-13, 9.898316e-13, 2.277261e-08, 
    4.69975e-08, 2.350554e-05, 0.0001581719, 0.0001754868, 0.000217059,
  6.126341e-08, 1.157438e-08, 1.67121e-08, 2.087456e-11, 4.50695e-11, 
    6.162789e-09, 1.164778e-13, 1.048661e-16, 2.23675e-12, 3.389468e-08, 
    2.659198e-08, 1.436883e-05, 0.0001747408, 0.0001764929, 0.0002123071,
  4.279033e-07, 3.732308e-07, 1.268461e-07, 4.408184e-10, 9.384329e-11, 
    4.726697e-08, 2.031128e-08, 7.521387e-08, 4.723516e-10, 3.618331e-08, 
    2.031199e-08, 1.520461e-05, 0.0001870002, 0.000184483, 0.0002355485,
  2.283839e-06, 2.887009e-06, 1.251081e-06, 7.475418e-08, 1.030004e-05, 
    1.972421e-07, 2.81187e-11, 4.028566e-10, 2.684926e-10, 9.219268e-09, 
    1.17732e-07, 2.041718e-05, 0.0001877913, 0.000216554, 0.0002727422,
  1.028978e-05, 2.340847e-06, 4.260922e-06, 1.66088e-06, 1.649987e-05, 
    2.043202e-06, 5.086212e-10, 3.76519e-14, 2.528951e-13, 9.182493e-11, 
    3.324788e-07, 1.553309e-05, 0.0001664017, 0.0002657645, 0.0003109048,
  0.0001359283, 0.0002826471, 0.0002601115, 9.677071e-05, 3.568063e-05, 
    1.164758e-05, 7.540878e-06, 3.142907e-06, 1.27974e-06, 1.695335e-06, 
    2.627241e-06, 3.225241e-06, 6.739789e-06, 4.879872e-06, 4.989524e-06,
  0.0002548499, 0.0003428459, 0.0003855037, 0.0001585522, 3.704561e-05, 
    5.600493e-06, 6.23799e-06, 2.344614e-06, 6.245679e-07, 3.180212e-06, 
    4.436379e-06, 5.631373e-06, 8.431846e-06, 6.280057e-06, 6.639802e-06,
  0.0002854244, 0.0004181013, 0.0004759961, 0.0002213078, 3.424574e-05, 
    2.144288e-06, 3.798371e-06, 2.986583e-06, 1.560821e-06, 5.313821e-06, 
    8.374761e-06, 6.77724e-06, 8.377543e-06, 8.267892e-06, 6.576757e-06,
  0.0002656668, 0.0003631218, 0.0004891343, 0.0002701083, 2.923833e-05, 
    2.485196e-07, 1.163368e-06, 1.160947e-06, 1.706818e-06, 6.912673e-06, 
    6.982293e-06, 6.825557e-06, 6.01924e-06, 7.766312e-06, 5.876519e-06,
  0.0001694997, 0.0002739066, 0.000445443, 0.0002863536, 3.192043e-05, 
    2.891903e-08, 2.29731e-07, 1.460742e-06, 2.50522e-06, 3.666255e-06, 
    5.856151e-06, 5.81069e-06, 3.478084e-06, 5.280344e-06, 5.60442e-06,
  9.310571e-05, 0.0002071317, 0.0003480031, 0.0002655271, 3.4391e-05, 
    2.392454e-08, 1.187579e-06, 6.50186e-07, 3.907847e-06, 3.626565e-06, 
    3.172819e-06, 2.309171e-06, 3.355961e-06, 2.53138e-06, 3.301159e-06,
  2.890338e-05, 0.0001980405, 0.0003397002, 0.0002377308, 3.02369e-05, 
    2.743392e-06, 3.144237e-06, 4.813709e-08, 3.47703e-07, 1.428416e-06, 
    1.640955e-06, 3.321105e-06, 2.427906e-06, 2.207116e-06, 1.981744e-06,
  9.575936e-05, 0.0002611736, 0.0003501204, 0.000232805, 2.674201e-05, 
    5.822939e-07, 1.826338e-06, 3.079212e-06, 1.042536e-06, 2.416171e-07, 
    1.801364e-06, 2.082591e-06, 2.674399e-06, 2.249705e-06, 3.31064e-06,
  0.0001518878, 0.000276962, 0.0003170221, 0.0001810832, 2.458845e-05, 
    1.242797e-06, 6.710324e-07, 1.102606e-07, 5.093443e-07, 2.264765e-07, 
    9.871421e-07, 5.029422e-07, 2.575655e-06, 2.854505e-06, 9.015866e-07,
  0.000153005, 0.0002459521, 0.0002967442, 0.0001299754, 4.962264e-06, 
    7.66966e-07, 3.504126e-06, 2.875322e-06, 1.412219e-07, 3.741281e-08, 
    1.265271e-07, 4.929602e-07, 1.770768e-06, 1.886131e-06, 4.573409e-07,
  9.142485e-07, 8.50682e-06, 4.145677e-05, 7.685877e-05, 0.000148411, 
    0.000250255, 0.0003428835, 0.0002976489, 0.0001298154, 3.706836e-05, 
    9.399904e-05, 6.106345e-05, 1.228785e-05, 2.926539e-06, 4.414369e-06,
  3.531759e-07, 1.267322e-05, 6.596634e-05, 0.0001563454, 0.0001799487, 
    0.0001714538, 0.0003083034, 0.0003531504, 0.0002226838, 4.595647e-05, 
    4.919248e-05, 5.62576e-05, 2.720279e-05, 8.166072e-06, 6.48682e-06,
  7.097314e-08, 2.442233e-05, 9.466246e-05, 0.0002598229, 0.0002346614, 
    0.0001123913, 0.0002357152, 0.0003809246, 0.0003059956, 0.0001117854, 
    4.326406e-05, 7.025865e-05, 3.976957e-05, 1.167305e-05, 7.456734e-06,
  5.652261e-08, 2.844505e-05, 0.0001204025, 0.0003147063, 0.0003148094, 
    0.0001083374, 0.0001500559, 0.00033897, 0.0003372129, 0.0001862927, 
    8.917403e-05, 9.933243e-05, 6.071438e-05, 2.248662e-05, 6.274856e-06,
  7.931868e-09, 1.73919e-05, 0.0001487037, 0.0003176383, 0.0004308255, 
    0.0001528688, 6.280265e-05, 0.0002825361, 0.0003505792, 0.0002790413, 
    9.543401e-05, 5.473579e-05, 6.848697e-05, 3.756835e-05, 3.023928e-06,
  1.455274e-08, 1.659357e-05, 0.0001755449, 0.0003423652, 0.0005447413, 
    0.0002179872, 5.402745e-05, 0.0002042627, 0.0003585631, 0.0003371105, 
    0.0001885987, 6.088047e-05, 6.510933e-05, 5.606459e-05, 1.340606e-06,
  8.574933e-09, 2.808552e-05, 0.0001890469, 0.0003567255, 0.0006093652, 
    0.0003168632, 7.745402e-05, 0.0001513311, 0.0003360295, 0.0003612021, 
    0.000233936, 7.855798e-05, 5.442167e-05, 6.295629e-05, 4.233667e-06,
  2.142053e-08, 5.078789e-05, 0.0002153197, 0.0003744538, 0.0005773124, 
    0.0002766918, 0.0001003105, 0.0001290113, 0.0002952871, 0.0003391942, 
    0.0002520179, 0.0001062734, 4.303468e-05, 6.430984e-05, 1.690248e-05,
  1.449714e-08, 6.269158e-05, 0.0002255359, 0.0003674503, 0.0005602675, 
    0.0002665134, 5.459501e-05, 1.787052e-05, 0.0001635982, 0.0002911917, 
    0.0002648095, 0.0001306882, 3.540942e-05, 6.594216e-05, 2.705629e-05,
  2.61957e-08, 7.611387e-05, 0.0002516706, 0.0004078555, 0.0005167491, 
    0.0002960198, 0.0001225626, 5.729292e-05, 0.0001566458, 0.0002786268, 
    0.0002527962, 0.00014603, 3.746459e-05, 5.467623e-05, 2.468076e-05,
  3.340606e-07, 1.955982e-07, 3.792666e-06, 7.481896e-06, 4.018341e-05, 
    8.708972e-05, 0.0001512735, 0.000183627, 0.0001135693, 0.0001193819, 
    0.0001989652, 5.406029e-05, 1.892443e-05, 9.390847e-06, 8.710213e-06,
  2.862172e-07, 9.300438e-08, 1.007448e-07, 2.917812e-06, 2.729497e-05, 
    6.005748e-05, 9.082069e-05, 0.000177447, 0.0001221059, 8.467039e-05, 
    0.0002352259, 0.0001147822, 2.669247e-05, 2.169413e-05, 8.99108e-06,
  2.514145e-07, 8.894713e-08, 6.699605e-09, 2.237246e-07, 6.721202e-06, 
    5.26125e-05, 5.924538e-05, 0.0001345846, 0.000138996, 6.785521e-05, 
    0.0001666667, 0.0001578723, 3.940269e-05, 3.324423e-05, 1.09865e-05,
  5.44751e-08, 2.601913e-08, 7.372414e-09, 1.43172e-08, 3.051648e-07, 
    2.881412e-05, 5.418296e-05, 7.892271e-05, 0.0001326788, 8.171163e-05, 
    8.948529e-05, 0.0001642724, 4.253148e-05, 4.284851e-05, 1.682108e-05,
  1.714499e-07, 1.469791e-07, 8.341038e-08, 1.618886e-08, 2.261694e-08, 
    8.891926e-06, 4.772448e-05, 5.744118e-05, 0.0001047242, 9.959731e-05, 
    5.647372e-05, 0.0001390313, 3.250243e-05, 3.573408e-05, 3.351629e-05,
  1.850754e-06, 2.251467e-06, 1.271072e-08, 3.891261e-08, 2.03785e-09, 
    6.1004e-07, 1.775579e-05, 4.513971e-05, 7.359259e-05, 9.328601e-05, 
    6.791673e-05, 0.0001235993, 4.420084e-05, 2.145904e-05, 4.415647e-05,
  5.879706e-09, 7.732314e-08, 6.507151e-08, 2.194378e-09, 7.892774e-10, 
    8.076281e-09, 9.877102e-06, 3.668049e-05, 5.64334e-05, 6.909355e-05, 
    6.227083e-05, 0.000100543, 7.312345e-05, 1.717194e-05, 4.48672e-05,
  3.990094e-10, 8.098512e-10, 5.674689e-09, 5.390595e-08, 1.991517e-09, 
    7.776509e-10, 1.210876e-06, 2.289988e-05, 4.454513e-05, 4.86876e-05, 
    3.26165e-05, 6.13138e-05, 0.0001082802, 2.940031e-05, 4.475472e-05,
  3.097894e-10, 1.583812e-09, 8.388788e-09, 9.599495e-09, 9.162928e-07, 
    1.569559e-09, 6.121149e-09, 4.200791e-06, 1.379453e-05, 2.299466e-05, 
    1.05935e-05, 1.265845e-05, 9.324884e-05, 5.277168e-05, 5.534035e-05,
  9.939136e-08, 2.646972e-08, 6.543737e-09, 2.573069e-08, 1.561743e-06, 
    3.441286e-09, 1.32947e-09, 7.991964e-07, 1.064769e-05, 5.118122e-06, 
    4.081103e-06, 1.393807e-06, 5.157233e-05, 6.168276e-05, 7.129657e-05,
  2.477381e-06, 1.012309e-05, 0.0001015264, 0.0001650818, 0.0002049634, 
    0.0002918278, 0.0003706866, 0.0003471372, 0.0002806196, 0.0001503835, 
    0.0001121394, 4.062546e-05, 2.553827e-06, 1.944718e-06, 3.467247e-06,
  3.148754e-06, 4.261739e-06, 6.193375e-05, 0.0001398607, 0.0001842079, 
    0.0002681824, 0.000428295, 0.0004543109, 0.0003449759, 0.0002221888, 
    0.0001819782, 0.0001286878, 1.571187e-05, 3.945438e-06, 5.013406e-06,
  6.043661e-06, 1.384182e-05, 2.882861e-05, 0.0001004048, 0.0001457049, 
    0.000216077, 0.0004165259, 0.0005325677, 0.0004235446, 0.0002636044, 
    0.0002483784, 0.0001827909, 4.472744e-05, 5.277378e-06, 4.238685e-06,
  1.312188e-05, 1.902764e-05, 1.37757e-05, 4.447035e-05, 0.0001289798, 
    0.0001811119, 0.0003536489, 0.0005615953, 0.0005123792, 0.0002934753, 
    0.0002671695, 0.0001886767, 5.082741e-05, 4.963807e-06, 5.745086e-06,
  8.951058e-06, 1.097501e-05, 1.080871e-05, 1.612656e-05, 0.0001194111, 
    0.0001946322, 0.0003255562, 0.0005737856, 0.0006159127, 0.0004045352, 
    0.0002483134, 0.0001547543, 3.695272e-05, 4.2439e-06, 4.033051e-06,
  7.349983e-06, 3.886239e-06, 8.016422e-06, 1.119344e-05, 0.0001040521, 
    0.0001983645, 0.0003414222, 0.0005850272, 0.0007626709, 0.0005923392, 
    0.0002440877, 0.0001025401, 1.533864e-05, 5.491815e-06, 5.102534e-06,
  2.343192e-08, 9.298864e-07, 3.42471e-06, 6.888568e-06, 8.162805e-05, 
    0.0002293354, 0.0002908689, 0.0004192111, 0.000764348, 0.0007834257, 
    0.0003439593, 9.559577e-05, 1.525404e-05, 9.058982e-06, 8.274513e-06,
  2.33076e-09, 3.150308e-08, 1.098714e-07, 2.114663e-06, 4.202615e-05, 
    0.0002415244, 0.0003337724, 0.0005384308, 0.0008064988, 0.0008489582, 
    0.0005237455, 0.0001565628, 2.427971e-05, 1.216125e-05, 1.088168e-05,
  3.115119e-09, 2.946884e-09, 2.703552e-09, 2.491788e-07, 2.452453e-05, 
    0.0001796143, 0.0002649738, 0.0004170921, 0.0006841723, 0.0007840727, 
    0.0006426387, 0.0002217474, 4.877331e-05, 1.383368e-05, 1.378814e-05,
  3.636437e-08, 6.200705e-09, 6.6723e-09, 3.43613e-08, 7.621436e-06, 
    0.0001047892, 0.0002077657, 0.0003942716, 0.000646899, 0.0007757781, 
    0.0006518991, 0.0002731872, 7.077885e-05, 2.635757e-05, 1.582856e-05,
  9.791899e-11, 3.491292e-11, 9.0943e-11, 1.003541e-08, 1.811645e-11, 
    2.984032e-09, 1.277749e-08, 3.484923e-07, 1.351118e-06, 7.822297e-06, 
    1.840269e-05, 6.919128e-05, 8.612988e-05, 7.390772e-05, 4.556529e-05,
  6.260754e-10, 2.590712e-10, 1.849587e-11, 3.080166e-09, 3.013746e-08, 
    1.604817e-07, 7.105629e-07, 9.487871e-07, 4.147991e-06, 9.084152e-06, 
    1.696068e-05, 7.303325e-05, 0.0001193881, 8.991601e-05, 7.790276e-05,
  1.431781e-08, 7.258128e-08, 4.211974e-10, 8.139962e-09, 4.463461e-08, 
    1.106973e-07, 2.993237e-07, 7.678067e-07, 2.682743e-06, 6.533522e-06, 
    1.739394e-05, 9.512228e-05, 0.000173644, 0.0001011334, 8.788747e-05,
  1.395718e-06, 4.276399e-07, 2.161193e-09, 3.232414e-11, 1.020698e-07, 
    1.26045e-07, 3.819165e-07, 7.365254e-07, 2.792299e-06, 5.074098e-06, 
    1.821138e-05, 0.0001247881, 0.0002128306, 0.0001007143, 8.010226e-05,
  2.206588e-06, 3.927037e-07, 5.116725e-09, 2.767873e-10, 4.028065e-08, 
    1.631002e-07, 4.00503e-07, 8.865986e-07, 1.475079e-06, 2.910866e-06, 
    4.327592e-05, 0.0001793699, 0.000255034, 0.0001446787, 6.140838e-05,
  1.596751e-05, 2.503051e-06, 4.158941e-08, 2.904011e-08, 8.278658e-08, 
    1.70251e-07, 1.017863e-07, 5.495912e-07, 3.839151e-06, 1.949316e-05, 
    8.123034e-05, 0.0002163403, 0.0002560081, 0.0001861553, 4.432269e-05,
  1.22038e-06, 1.519877e-07, 2.390751e-08, 4.50667e-09, 1.221184e-08, 
    3.831826e-07, 1.12987e-07, 3.825077e-07, 4.990814e-06, 5.069133e-05, 
    0.0001325416, 0.0002136703, 0.0002319766, 0.0001937678, 5.774162e-05,
  1.017503e-05, 1.235288e-06, 4.605564e-08, 3.304997e-08, 4.384906e-08, 
    9.013044e-07, 3.654117e-06, 4.259858e-06, 1.62027e-05, 6.830893e-05, 
    0.0001746522, 0.0002415514, 0.0002100167, 0.0001822035, 0.0001010258,
  1.612603e-05, 3.639186e-06, 1.845128e-06, 1.415926e-06, 9.57931e-06, 
    1.006008e-06, 2.736364e-07, 3.386921e-06, 2.43546e-05, 9.251971e-05, 
    0.0001679651, 0.0002555729, 0.0001975074, 0.0001490899, 0.0001123712,
  1.510417e-05, 7.095347e-06, 4.494789e-06, 3.550654e-06, 9.472096e-06, 
    1.614166e-06, 1.592127e-06, 9.605334e-07, 3.879954e-05, 0.0001105161, 
    0.0001535809, 0.000217704, 0.0001568622, 0.0001239155, 0.0001000997,
  1.196308e-08, 6.49201e-11, 1.271519e-13, 8.33642e-23, 4.365112e-12, 
    6.295498e-22, 3.176284e-10, 6.388811e-08, 1.387911e-08, 1.12556e-07, 
    7.491906e-06, 9.959775e-05, 0.0001468653, 0.0001944198, 0.0001454748,
  9.572318e-08, 1.484384e-09, 1.438467e-11, 1.042872e-23, 2.527569e-11, 
    3.847954e-22, 7.059315e-22, 1.075807e-09, 5.158502e-09, 2.07377e-08, 
    5.584624e-09, 2.556919e-05, 7.836486e-05, 9.499044e-05, 0.0001089481,
  3.062509e-08, 9.57718e-08, 1.748235e-10, 1.712795e-18, 1.38039e-23, 
    1.455125e-22, 5.248915e-22, 3.247058e-10, 9.441117e-10, 9.880111e-09, 
    2.266292e-08, 9.883006e-07, 3.085263e-05, 5.640159e-05, 8.241657e-05,
  9.051713e-08, 1.783558e-07, 4.248174e-09, 1.454068e-11, 2.141784e-24, 
    2.876804e-23, 1.981456e-22, 2.668125e-11, 1.904979e-10, 1.993657e-09, 
    1.157156e-08, 1.339728e-08, 4.554762e-06, 3.549496e-05, 5.257167e-05,
  6.268701e-08, 3.671026e-07, 8.958867e-08, 1.649616e-10, 3.995807e-12, 
    1.472957e-13, 5.206358e-23, 4.869641e-22, 5.189278e-12, 1.810808e-10, 
    4.026385e-09, 1.513012e-08, 7.292565e-08, 9.55996e-06, 2.896627e-05,
  4.354024e-11, 1.249045e-07, 1.777979e-08, 4.864426e-09, 2.957508e-11, 
    1.041738e-10, 2.558599e-12, 4.375496e-12, 4.181324e-11, 3.197037e-13, 
    2.774217e-09, 1.07995e-08, 1.301105e-08, 9.553339e-08, 1.954717e-05,
  8.656635e-11, 8.76537e-09, 1.002582e-08, 2.71017e-08, 2.658916e-09, 
    1.042212e-07, 7.548666e-09, 5.329621e-10, 5.736642e-12, 7.967861e-22, 
    8.082452e-10, 8.505523e-09, 1.920044e-08, 1.815947e-08, 1.210634e-06,
  9.001503e-10, 1.628033e-07, 3.21152e-09, 1.506128e-08, 5.159996e-06, 
    3.684599e-06, 6.878183e-07, 2.32034e-10, 1.375285e-10, 1.102281e-16, 
    9.16988e-15, 2.666764e-09, 1.143552e-08, 1.783595e-08, 5.46499e-08,
  7.734854e-10, 2.915861e-10, 5.010513e-07, 6.812654e-06, 2.678079e-05, 
    6.962595e-06, 2.255026e-08, 1.970783e-09, 2.284016e-11, 1.269258e-17, 
    5.680128e-22, 2.784433e-11, 8.832109e-09, 1.345227e-08, 1.13019e-08,
  1.638409e-07, 1.769348e-07, 6.405293e-07, 7.820498e-06, 3.036779e-05, 
    9.908003e-06, 7.480722e-06, 3.309383e-08, 3.938151e-10, 1.030673e-11, 
    2.248596e-15, 2.403779e-12, 2.08247e-09, 9.67521e-09, 3.496092e-08,
  1.325727e-09, 2.153782e-12, 1.500956e-10, 3.175504e-09, 2.906058e-09, 
    4.317211e-09, 5.547291e-09, 7.847941e-09, 2.597998e-07, 1.242481e-08, 
    5.582446e-07, 2.904155e-05, 6.544063e-05, 0.0003776409, 0.0005267401,
  2.634225e-11, 2.947529e-12, 2.100003e-11, 8.08247e-10, 3.668424e-09, 
    2.474569e-09, 1.171047e-09, 2.893407e-08, 1.61205e-07, 2.214309e-08, 
    6.342775e-09, 1.138961e-08, 2.480292e-06, 7.914189e-05, 0.0004283718,
  3.043228e-10, 1.996275e-09, 1.733673e-11, 8.726023e-12, 3.791489e-12, 
    2.517225e-09, 1.304573e-09, 3.176923e-08, 5.993746e-07, 3.336955e-07, 
    2.479026e-08, 6.705474e-09, 4.393741e-08, 8.886875e-06, 0.0001169977,
  1.07706e-08, 4.493864e-08, 4.058263e-10, 1.83067e-11, 2.476147e-12, 
    2.966953e-10, 1.301579e-09, 8.992916e-10, 3.318667e-08, 1.183108e-07, 
    6.275797e-08, 6.578153e-08, 2.134088e-08, 1.212864e-07, 2.26527e-05,
  9.710554e-09, 1.96075e-08, 6.626215e-10, 1.20283e-10, 4.911091e-11, 
    6.043415e-12, 1.55004e-12, 6.592395e-10, 5.887404e-10, 2.446846e-09, 
    3.002112e-09, 6.316467e-09, 1.293421e-08, 3.85238e-08, 5.644884e-07,
  4.29558e-07, 3.76163e-08, 9.760265e-09, 1.08252e-09, 1.463355e-10, 
    9.627794e-11, 1.020124e-11, 1.011947e-12, 6.244492e-10, 3.312291e-10, 
    7.763497e-10, 1.93493e-09, 2.499976e-09, 2.289547e-08, 3.937844e-08,
  4.173314e-06, 1.065728e-06, 7.434028e-08, 2.778735e-09, 4.593478e-10, 
    1.235572e-10, 4.622483e-11, 4.832837e-13, 3.0918e-13, 7.498162e-10, 
    1.583823e-10, 6.233219e-11, 2.115579e-09, 4.959817e-09, 2.159172e-08,
  1.136151e-05, 7.614803e-06, 2.594633e-06, 6.489699e-09, 2.022254e-09, 
    6.217702e-10, 9.472005e-11, 2.193602e-11, 5.128338e-14, 4.827493e-10, 
    4.327533e-10, 1.579548e-22, 4.572485e-11, 2.895144e-10, 2.938897e-09,
  6.474859e-06, 3.509745e-06, 1.449333e-06, 4.975952e-08, 3.186788e-07, 
    4.384354e-09, 8.894577e-10, 7.496608e-11, 6.828218e-12, 3.276322e-11, 
    7.366797e-11, 3.317896e-10, 1.526636e-11, 6.239793e-11, 1.482094e-09,
  2.069675e-06, 2.109732e-06, 6.716626e-07, 4.603619e-08, 1.174899e-06, 
    3.771531e-09, 5.007875e-10, 1.66319e-10, 1.898918e-11, 1.346192e-10, 
    1.710637e-11, 1.544677e-11, 1.598495e-12, 6.968e-12, 1.631465e-09,
  1.501243e-08, 1.870998e-09, 7.357923e-10, 8.125765e-09, 2.879219e-08, 
    1.399996e-07, 7.94071e-07, 4.04212e-05, 0.0002104777, 0.0004335371, 
    0.0007021811, 0.001045978, 0.0007860472, 0.0002646071, 5.490328e-05,
  1.179636e-06, 9.649966e-08, 1.187664e-09, 2.093249e-08, 6.417237e-09, 
    1.824103e-08, 3.238474e-07, 5.247637e-07, 8.289328e-05, 0.000266516, 
    0.0004385846, 0.0006542978, 0.0008660191, 0.0005075503, 0.0001196915,
  4.097288e-06, 9.571449e-06, 6.281086e-08, 5.814444e-10, 9.775331e-10, 
    3.479588e-09, 4.103888e-06, 6.164052e-06, 7.967919e-06, 0.0001148292, 
    0.0003060928, 0.0003814981, 0.0005332063, 0.0005848057, 0.0002823842,
  1.649364e-05, 2.138765e-05, 1.139063e-06, 3.705864e-09, 3.337125e-09, 
    1.116053e-09, 2.160133e-08, 4.755316e-06, 4.667849e-06, 1.769673e-05, 
    0.0001218606, 0.000296958, 0.0003067905, 0.0004078799, 0.0003696127,
  1.121127e-05, 1.098661e-05, 1.841736e-06, 1.34941e-08, 9.596851e-11, 
    9.920967e-12, 6.710156e-10, 7.345317e-08, 1.075856e-06, 7.419691e-06, 
    3.928016e-05, 0.0001434313, 0.0002563529, 0.0002113527, 0.0003202956,
  1.358984e-05, 1.015769e-05, 5.614765e-08, 3.399291e-08, 3.031146e-09, 
    1.075141e-09, 3.340017e-10, 2.658243e-09, 7.568625e-07, 3.254064e-06, 
    8.277711e-06, 6.255854e-05, 0.0001884959, 0.0001768176, 0.0001204044,
  1.117957e-06, 1.977553e-06, 3.943071e-07, 5.467999e-08, 1.131526e-09, 
    5.219103e-09, 1.70841e-07, 2.706034e-07, 1.147874e-08, 1.860874e-06, 
    3.764801e-06, 3.441788e-06, 7.719895e-05, 0.0001452969, 9.429043e-05,
  3.560028e-07, 9.626306e-07, 1.489075e-06, 4.392461e-07, 1.691559e-08, 
    5.765373e-07, 5.199438e-06, 8.198968e-06, 9.360389e-06, 9.779519e-07, 
    4.155303e-06, 1.520437e-06, 1.509819e-05, 8.980616e-05, 8.600077e-05,
  8.48086e-08, 3.394178e-07, 7.221389e-07, 7.352553e-07, 2.756518e-07, 
    2.031431e-06, 3.34508e-06, 9.201755e-06, 2.024515e-05, 1.400388e-05, 
    6.026041e-06, 6.755909e-06, 1.166741e-06, 3.104781e-05, 7.346404e-05,
  1.748818e-08, 3.147441e-07, 4.979264e-07, 4.643544e-07, 3.701283e-07, 
    8.122412e-07, 4.710486e-06, 5.034879e-06, 1.214904e-05, 1.594143e-05, 
    1.413986e-05, 8.3984e-06, 6.17909e-06, 1.38644e-06, 3.620722e-05,
  1.435918e-09, 2.754849e-09, 4.632431e-10, 1.975949e-09, 1.91981e-08, 
    3.968142e-08, 1.175513e-07, 1.166176e-06, 5.849453e-05, 0.0003255211, 
    0.0004829078, 0.0005150257, 0.0004172259, 0.0002084209, 7.00987e-05,
  1.150514e-10, 3.699819e-11, 2.928547e-10, 1.544213e-09, 1.042107e-08, 
    4.284455e-08, 1.659183e-07, 2.584758e-06, 9.308138e-06, 0.0001581018, 
    0.0004357865, 0.0005982467, 0.0005820283, 0.0004878621, 0.0001410753,
  1.387759e-10, 2.76366e-10, 3.51427e-12, 1.628817e-10, 2.160816e-09, 
    1.430979e-07, 2.777854e-06, 9.501622e-06, 8.040089e-06, 1.946539e-05, 
    0.0002530637, 0.0005486517, 0.0007373451, 0.0006700696, 0.0004469863,
  8.34515e-10, 1.43068e-07, 4.079767e-11, 1.720723e-10, 8.03494e-09, 
    2.384213e-07, 6.202938e-06, 7.084576e-06, 1.541289e-05, 3.013767e-05, 
    6.266632e-05, 0.000427145, 0.0007590407, 0.0008515745, 0.0006376731,
  6.461442e-09, 4.416036e-08, 4.886715e-11, 6.761441e-12, 6.171418e-10, 
    3.344513e-08, 5.611109e-06, 3.873178e-06, 1.755947e-05, 3.773479e-05, 
    3.058734e-05, 0.0001345167, 0.0006864974, 0.0009550976, 0.0008249083,
  2.58233e-08, 1.58252e-07, 1.936799e-12, 8.609066e-14, 3.239671e-09, 
    9.433353e-08, 1.105408e-06, 6.295284e-06, 7.205483e-06, 3.892967e-05, 
    1.886092e-05, 1.319533e-05, 0.0003406976, 0.0009241052, 0.0009729079,
  2.242894e-14, 3.356979e-10, 8.959504e-09, 2.902162e-09, 4.415594e-09, 
    6.05316e-08, 3.342891e-06, 1.765781e-06, 1.920512e-06, 2.903239e-05, 
    3.239878e-05, 1.963998e-05, 1.856052e-05, 0.000663206, 0.001046542,
  6.328094e-17, 1.002573e-09, 3.757567e-08, 1.088984e-08, 9.197203e-11, 
    7.74124e-09, 4.404064e-07, 1.189913e-05, 1.737661e-05, 7.547018e-06, 
    3.867199e-05, 2.952957e-05, 1.582964e-05, 0.0001159055, 0.0008858643,
  2.646871e-23, 1.948949e-09, 1.151082e-07, 2.701067e-08, 8.241077e-10, 
    5.827003e-11, 1.897435e-08, 2.485297e-06, 5.526265e-06, 8.746812e-06, 
    2.079452e-05, 2.60009e-05, 1.026748e-05, 8.527784e-06, 0.0002926412,
  1.681032e-23, 2.735336e-10, 2.624626e-07, 9.016653e-08, 2.567702e-08, 
    5.06824e-09, 1.251683e-08, 4.905048e-07, 3.490024e-06, 7.363774e-06, 
    7.908165e-06, 1.132828e-05, 1.361374e-05, 5.476272e-06, 1.727757e-05,
  2.443611e-07, 8.820515e-08, 3.243488e-08, 3.690268e-08, 2.489741e-07, 
    2.33073e-06, 1.872729e-05, 5.62186e-05, 9.695724e-05, 0.0001102151, 
    5.46465e-05, 4.604842e-05, 0.0002138255, 0.0003110885, 0.0001862754,
  2.382281e-07, 6.085622e-07, 8.916599e-07, 5.650554e-07, 2.298869e-07, 
    5.639725e-07, 2.713942e-06, 1.187411e-05, 3.299715e-05, 5.161988e-05, 
    4.400777e-05, 4.101808e-05, 0.0001166038, 0.0003020948, 0.0002815048,
  4.301413e-07, 9.898104e-07, 1.734011e-06, 2.088188e-06, 1.034466e-06, 
    6.680236e-07, 6.564867e-07, 1.413668e-06, 4.546154e-06, 1.394516e-05, 
    1.959989e-05, 2.285123e-05, 9.420431e-05, 0.0002414411, 0.0002369225,
  7.424919e-08, 8.311025e-07, 1.183705e-07, 5.491075e-07, 2.15841e-07, 
    1.207621e-06, 3.04359e-06, 1.608871e-06, 3.937485e-06, 7.848617e-06, 
    1.673024e-05, 1.943931e-05, 5.26525e-05, 0.0002026139, 0.0002233761,
  2.029745e-08, 1.051199e-07, 5.212764e-08, 2.762837e-07, 1.155594e-06, 
    7.356778e-07, 4.357277e-06, 3.523564e-06, 2.704419e-06, 5.040485e-06, 
    8.804366e-06, 1.272028e-05, 2.571827e-05, 0.0001061128, 0.0001640162,
  6.840277e-10, 3.120614e-09, 6.095626e-09, 2.092594e-08, 3.725952e-07, 
    2.054814e-07, 1.897511e-07, 2.702346e-06, 3.215657e-06, 5.676967e-06, 
    5.072735e-06, 9.086137e-06, 1.367976e-05, 3.545756e-05, 7.998489e-05,
  5.698702e-10, 5.069961e-09, 1.025e-08, 6.471654e-08, 5.040008e-08, 
    2.961277e-07, 6.853838e-08, 3.869922e-07, 7.414772e-07, 1.499117e-06, 
    5.517261e-06, 6.068043e-06, 4.941227e-06, 5.0334e-06, 1.113316e-05,
  1.366906e-09, 3.606197e-09, 1.308435e-08, 5.323875e-07, 1.603954e-07, 
    6.833619e-07, 3.827958e-06, 2.133877e-05, 8.523502e-06, 1.045888e-06, 
    5.706047e-06, 6.696317e-06, 2.97427e-06, 4.510132e-06, 3.283988e-06,
  6.322814e-10, 1.906735e-09, 3.544089e-09, 4.78644e-08, 6.487193e-06, 
    4.782095e-06, 2.643847e-06, 6.994125e-06, 4.204333e-06, 3.748193e-06, 
    3.199111e-06, 6.673337e-06, 4.574074e-06, 5.469482e-06, 5.190592e-06,
  2.660215e-09, 2.019427e-09, 1.112196e-09, 9.324908e-08, 3.772894e-06, 
    2.273317e-06, 9.668332e-06, 1.035931e-05, 7.423038e-06, 8.463448e-06, 
    2.971199e-06, 2.018544e-06, 4.638174e-06, 3.189208e-06, 3.311983e-06,
  3.655431e-05, 5.674995e-05, 6.025464e-05, 3.644657e-05, 4.150216e-05, 
    0.0001090823, 0.0002496122, 0.0003091964, 0.0002147486, 6.336653e-05, 
    1.556581e-06, 2.553991e-07, 2.055448e-06, 3.364329e-06, 6.507519e-06,
  2.309381e-05, 4.65251e-05, 7.119061e-05, 5.134231e-05, 6.860164e-05, 
    0.0001829214, 0.0003473607, 0.0004069422, 0.0002809037, 0.0001144183, 
    1.981485e-05, 3.237908e-06, 5.951426e-06, 9.889018e-06, 1.015027e-05,
  5.414668e-05, 7.741677e-05, 7.267129e-05, 5.051967e-05, 7.619869e-05, 
    0.0002187292, 0.0004085143, 0.0004795931, 0.0003373262, 0.0001390549, 
    3.580412e-05, 8.964523e-06, 1.074821e-05, 1.265294e-05, 1.279419e-05,
  0.0001224649, 0.0001097835, 5.932186e-05, 4.447496e-05, 6.480964e-05, 
    0.0002081288, 0.0004640575, 0.0005759762, 0.0004326541, 0.0001391559, 
    3.261173e-05, 1.881889e-05, 2.787933e-05, 2.989765e-05, 1.712559e-05,
  9.453666e-05, 9.684877e-05, 6.105407e-05, 4.282496e-05, 5.607988e-05, 
    0.0001739073, 0.0004612953, 0.0006709249, 0.0005527751, 0.0002069647, 
    4.813943e-05, 3.537764e-05, 5.516848e-05, 8.206746e-05, 7.06202e-05,
  2.359372e-05, 4.814326e-05, 2.234728e-05, 2.389938e-05, 3.907269e-05, 
    0.0001220469, 0.0003767252, 0.0006663268, 0.0006989518, 0.0003855887, 
    6.650421e-05, 3.840401e-05, 6.762028e-05, 0.0001031421, 0.0001229942,
  8.463091e-08, 2.271301e-06, 1.26525e-05, 1.074449e-05, 1.051278e-05, 
    8.424119e-05, 0.000245401, 0.000497214, 0.00067526, 0.0005489013, 
    0.0001676341, 4.6509e-05, 6.924209e-05, 0.0001118935, 0.0001237034,
  3.1323e-08, 1.279008e-07, 5.036629e-06, 1.118908e-06, 2.078691e-06, 
    1.148772e-05, 0.0001246003, 0.0003613408, 0.0005810912, 0.0005599745, 
    0.0003152788, 8.178656e-05, 5.899072e-05, 9.241072e-05, 0.0001079078,
  1.533087e-08, 2.974369e-08, 2.288707e-06, 1.142727e-06, 9.700969e-06, 
    1.483236e-05, 4.370216e-05, 0.0001264916, 0.0003287116, 0.0004170302, 
    0.0003110424, 0.0001289981, 4.596799e-05, 3.639731e-05, 5.073338e-05,
  5.45621e-09, 1.467549e-07, 3.46942e-07, 1.348227e-06, 7.298023e-06, 
    5.208477e-06, 2.384727e-05, 3.7876e-05, 0.000112661, 0.0002225705, 
    0.0002111821, 0.0001163638, 3.412138e-05, 1.090743e-05, 8.553004e-06,
  0.0001520883, 8.228489e-05, 8.370781e-06, 6.793573e-06, 1.152607e-05, 
    9.857036e-06, 4.606532e-06, 1.071627e-06, 3.58442e-07, 6.371216e-07, 
    6.540546e-08, 3.490508e-09, 1.290341e-06, 1.675049e-06, 2.185869e-06,
  6.464349e-05, 1.55867e-05, 7.493892e-06, 7.073324e-06, 1.222317e-05, 
    8.861555e-06, 6.178231e-06, 4.293377e-06, 1.767696e-06, 8.327748e-07, 
    7.331148e-08, 3.928671e-07, 3.231565e-06, 5.233818e-06, 8.114071e-06,
  5.362187e-05, 2.931772e-05, 1.171653e-05, 9.692669e-06, 1.035646e-05, 
    1.400209e-05, 8.142721e-06, 3.285675e-06, 1.913592e-06, 6.730352e-07, 
    8.87965e-08, 1.876374e-06, 4.34291e-06, 6.688005e-06, 6.785817e-06,
  0.0001115286, 8.647405e-05, 2.850453e-05, 1.985676e-05, 1.096231e-05, 
    1.806087e-05, 1.443313e-05, 6.452603e-06, 3.704647e-06, 8.498619e-07, 
    1.513519e-07, 4.006951e-06, 4.892557e-06, 1.031229e-05, 4.048157e-06,
  0.0001964582, 0.0001208287, 8.169533e-05, 4.535036e-05, 2.470671e-05, 
    3.365858e-05, 4.352332e-05, 3.190274e-05, 8.887831e-06, 1.494706e-06, 
    1.100005e-06, 4.942427e-06, 4.953406e-06, 2.88743e-06, 1.308869e-06,
  0.0002491606, 0.0001562154, 6.903982e-05, 5.586159e-05, 4.408948e-05, 
    4.41613e-05, 0.0001037473, 0.0001519901, 7.553206e-05, 8.199703e-06, 
    2.008676e-06, 3.19661e-06, 4.301805e-06, 7.949528e-07, 1.401041e-07,
  0.0001689011, 8.142029e-05, 4.258327e-05, 4.673763e-05, 4.016321e-05, 
    6.602849e-05, 0.0001540538, 0.0002905068, 0.0002802203, 7.550597e-05, 
    7.799139e-06, 2.471754e-06, 6.294061e-07, 1.780905e-07, 4.344962e-08,
  8.865765e-05, 7.874201e-05, 6.79595e-05, 2.596868e-05, 1.825481e-05, 
    6.643386e-05, 0.0001694813, 0.0004077299, 0.0004518312, 0.0002730957, 
    0.0001207408, 2.190906e-05, 1.742977e-06, 3.457199e-07, 1.530794e-07,
  6.644697e-05, 9.251202e-05, 0.0001090352, 3.178538e-05, 7.372008e-05, 
    0.0001357508, 0.0001840083, 0.0003475202, 0.0004996422, 0.0004790745, 
    0.0003043821, 0.0001679287, 2.200244e-05, 5.331528e-06, 3.135979e-06,
  2.578328e-05, 6.819789e-05, 0.0001055422, 8.717968e-05, 0.0001087035, 
    0.0001183137, 0.0002361996, 0.0003873593, 0.0005575477, 0.0006212585, 
    0.0004784401, 0.0003042609, 0.0001190478, 2.602342e-05, 9.10862e-06,
  0.0001741614, 7.824289e-05, 1.908236e-05, 9.600498e-07, 1.280232e-06, 
    1.864767e-06, 8.387792e-06, 8.337889e-06, 1.260247e-05, 2.570124e-05, 
    1.468126e-05, 2.59424e-08, 6.841032e-06, 2.245543e-06, 1.968233e-07,
  0.000235793, 0.0001547895, 4.793177e-05, 1.149956e-06, 1.038452e-06, 
    1.098729e-06, 5.624965e-06, 8.44565e-06, 1.763842e-05, 4.208033e-05, 
    3.167168e-05, 2.088624e-05, 1.850598e-06, 3.795125e-06, 6.697033e-06,
  0.0002641643, 0.0002368448, 8.885281e-05, 2.935623e-06, 1.590431e-06, 
    1.098696e-06, 3.854823e-06, 6.451628e-06, 1.833422e-05, 4.858304e-05, 
    0.0001352319, 1.831894e-05, 7.951304e-06, 1.258272e-05, 9.944397e-06,
  0.0003364666, 0.0002835941, 0.0001369672, 1.129843e-05, 1.395875e-06, 
    1.735316e-06, 3.137719e-06, 5.193379e-06, 1.937228e-05, 4.969764e-05, 
    0.000120346, 2.118573e-05, 9.748892e-06, 1.185846e-05, 4.903386e-06,
  0.0003956498, 0.0003166989, 0.0001870737, 3.615548e-05, 2.327081e-06, 
    3.887425e-06, 5.235765e-06, 8.570938e-06, 2.053844e-05, 5.451936e-05, 
    0.0002049359, 1.132958e-05, 6.748578e-06, 5.060366e-06, 4.072841e-06,
  0.0004683306, 0.0003768094, 0.0001880461, 5.779105e-05, 7.181032e-06, 
    8.56897e-06, 1.703552e-05, 2.183308e-05, 3.494279e-05, 5.833399e-05, 
    6.049293e-05, 6.644103e-06, 4.987859e-06, 3.452194e-06, 3.082176e-06,
  0.0005365553, 0.0004335395, 0.0002276796, 9.338749e-05, 1.994955e-05, 
    4.423737e-05, 6.566659e-05, 7.751022e-05, 5.819146e-05, 5.345998e-05, 
    2.233689e-05, 8.371106e-07, 1.131943e-06, 3.011412e-06, 1.55739e-06,
  0.0005654584, 0.0005381929, 0.0003080259, 0.0001291149, 3.08895e-05, 
    5.630232e-05, 0.0001244193, 0.0002307418, 0.0001222586, 3.670018e-05, 
    1.317344e-05, 6.917168e-07, 1.223206e-06, 2.174752e-06, 1.129172e-06,
  0.00048522, 0.0006509972, 0.0003846423, 9.498355e-05, 7.487516e-05, 
    6.223562e-05, 7.570363e-05, 4.60469e-05, 1.058493e-05, 2.0703e-05, 
    7.48728e-06, 6.119911e-07, 8.419675e-07, 9.257187e-07, 5.137569e-07,
  0.0003660033, 0.0006716265, 0.0005197002, 6.551683e-05, 4.332836e-05, 
    4.883569e-05, 0.0001642766, 0.0001671114, 0.0001123044, 5.224353e-05, 
    1.352793e-05, 2.262848e-06, 1.578391e-06, 7.229463e-07, 2.868558e-07,
  2.650815e-08, 1.26309e-07, 5.41049e-07, 5.470773e-07, 2.255487e-08, 
    2.028851e-05, 0.0001525876, 0.000221696, 0.0001518654, 7.038292e-05, 
    4.047751e-05, 0.0001982101, 9.536883e-05, 1.205114e-05, 1.821566e-06,
  5.21755e-08, 1.11877e-07, 2.501216e-07, 5.428123e-07, 6.012962e-08, 
    1.673161e-06, 0.0001402737, 0.0002819508, 0.0002199544, 8.316747e-05, 
    7.224161e-05, 0.0001684678, 8.140031e-05, 8.106933e-06, 4.319019e-06,
  2.926394e-07, 5.686278e-07, 9.284577e-08, 2.194725e-07, 4.604691e-08, 
    1.449956e-08, 9.478359e-05, 0.0003100922, 0.0002674807, 0.0001034037, 
    7.511778e-05, 0.0001154918, 1.674695e-05, 1.899373e-06, 6.99228e-07,
  3.14557e-06, 1.226788e-06, 3.152463e-08, 1.870818e-07, 6.298054e-08, 
    1.745016e-07, 6.494777e-05, 0.0002810668, 0.0002967165, 0.0001308145, 
    9.469468e-05, 0.0001485228, 1.709146e-05, 4.035869e-06, 9.916668e-08,
  1.332775e-06, 5.700908e-07, 2.171235e-07, 1.463099e-07, 1.328144e-07, 
    1.970138e-07, 4.200238e-05, 0.0002552726, 0.0002956752, 0.0001621606, 
    0.000126976, 0.0003425309, 1.876324e-05, 4.345441e-07, 2.167029e-07,
  1.74454e-07, 6.97478e-07, 1.577913e-08, 1.205556e-07, 4.23932e-07, 
    5.485616e-07, 9.357144e-06, 0.000220447, 0.0003008004, 0.0002143598, 
    0.0001764558, 0.0002673971, 5.567651e-06, 1.233924e-07, 3.238853e-07,
  6.413342e-09, 3.493107e-09, 1.497884e-09, 1.429206e-07, 6.468205e-07, 
    1.427889e-06, 1.263403e-06, 0.0001501388, 0.0002725582, 0.0002297252, 
    0.0001933508, 9.333991e-05, 1.953297e-06, 5.961664e-07, 9.290002e-07,
  7.741387e-09, 1.252478e-08, 8.709961e-08, 7.430409e-07, 5.746512e-06, 
    4.689422e-06, 1.212332e-06, 0.0001032038, 0.0002414848, 0.0002334981, 
    0.00020403, 7.160664e-05, 2.122049e-06, 2.922749e-07, 5.264639e-07,
  3.718192e-09, 1.132452e-08, 7.598912e-07, 3.019449e-06, 3.096624e-05, 
    5.074047e-06, 2.480854e-07, 3.111864e-05, 0.000174983, 0.0002445697, 
    0.0002312258, 0.0001431276, 4.778586e-06, 4.282651e-07, 3.791782e-07,
  9.062732e-09, 5.802364e-08, 8.848397e-07, 3.814446e-06, 6.72298e-06, 
    2.168951e-06, 7.87742e-07, 2.066392e-05, 0.0001337382, 0.0002364349, 
    0.0002505675, 0.0002258516, 8.402831e-06, 3.182617e-07, 7.537697e-07,
  2.679334e-09, 1.531154e-09, 5.823884e-09, 2.738058e-08, 1.048272e-05, 
    9.560664e-05, 0.0002360551, 0.0004825862, 0.0005107602, 0.000219151, 
    7.039071e-06, 2.300252e-05, 8.968168e-05, 9.609633e-05, 2.424735e-06,
  2.341209e-08, 5.189902e-09, 1.657264e-08, 2.215682e-08, 1.73543e-06, 
    4.51719e-05, 0.0001488502, 0.0004344193, 0.0005323095, 0.0003020222, 
    2.067741e-05, 6.657717e-05, 5.661392e-05, 3.150453e-05, 7.326959e-06,
  3.056324e-08, 8.977401e-08, 3.648659e-08, 5.196712e-08, 2.162175e-08, 
    3.001161e-05, 9.930326e-05, 0.0003191861, 0.0005083451, 0.0003516228, 
    9.655532e-05, 8.116144e-05, 6.172469e-05, 1.314038e-05, 6.541583e-06,
  1.180968e-08, 2.223861e-08, 4.788875e-08, 8.330831e-08, 2.334246e-08, 
    1.10772e-05, 0.0001163145, 0.0002506203, 0.0004778164, 0.0003778803, 
    6.368714e-05, 8.749587e-05, 3.115187e-05, 1.62947e-05, 4.640116e-06,
  9.356052e-09, 1.653288e-08, 1.042718e-07, 2.058255e-08, 6.991755e-08, 
    1.795746e-06, 8.66979e-05, 0.0002356831, 0.0004520173, 0.0004245053, 
    0.0001843553, 9.001559e-05, 3.202037e-05, 1.150531e-05, 1.991907e-06,
  1.081498e-09, 3.376143e-09, 5.716728e-08, 6.382614e-08, 4.512533e-08, 
    1.484208e-07, 6.359879e-05, 0.0002159257, 0.0004418217, 0.0004815023, 
    0.0002649636, 0.0001093561, 7.39101e-06, 7.788071e-06, 4.264566e-07,
  4.228831e-10, 2.168372e-09, 3.197255e-08, 2.278347e-08, 1.00662e-08, 
    4.427502e-08, 2.79284e-05, 0.0001747994, 0.00038762, 0.0005177378, 
    0.0002938368, 0.0001411208, 2.897278e-06, 3.401035e-06, 1.153909e-07,
  2.199887e-10, 3.588096e-09, 2.1426e-08, 2.571638e-08, 2.541523e-08, 
    9.589195e-08, 1.446424e-05, 0.0001907975, 0.0004304343, 0.000561715, 
    0.0003708856, 0.0001689619, 3.097178e-06, 1.696619e-07, 5.017414e-08,
  5.040229e-10, 2.360299e-09, 3.733629e-09, 1.356314e-08, 7.401963e-08, 
    4.467143e-07, 2.563981e-06, 0.0001608551, 0.0004088667, 0.0006002439, 
    0.0004393188, 0.0001974838, 1.333658e-06, 2.52735e-07, 3.447015e-07,
  1.336517e-09, 7.888469e-09, 5.950917e-09, 1.83555e-08, 2.066925e-07, 
    8.093794e-07, 1.329654e-06, 0.0001750005, 0.0004197235, 0.0006440955, 
    0.000555681, 0.0002448544, 4.897147e-06, 4.933258e-07, 6.526357e-07,
  1.410197e-08, 6.190931e-09, 7.661611e-09, 1.114136e-07, 5.402717e-06, 
    3.780287e-05, 0.0002603924, 0.0004522178, 0.0004459436, 0.0001592559, 
    1.754389e-05, 4.842413e-06, 7.370639e-05, 2.307874e-05, 2.190399e-06,
  4.082235e-08, 5.476975e-09, 9.610718e-09, 1.81254e-08, 4.120438e-06, 
    1.513003e-05, 0.0001555866, 0.0004274612, 0.0004720052, 0.0002515263, 
    1.8069e-05, 5.210478e-06, 3.102181e-05, 4.890939e-05, 5.594366e-06,
  1.227666e-08, 2.324464e-08, 1.777216e-09, 3.172133e-09, 9.387845e-07, 
    1.406608e-05, 8.30457e-05, 0.0003176797, 0.0004387145, 0.0002794803, 
    3.411011e-05, 6.318264e-06, 1.710975e-05, 1.028351e-05, 5.668239e-06,
  1.202775e-07, 2.619233e-08, 3.085429e-09, 1.947132e-09, 9.533731e-08, 
    2.729721e-06, 3.785218e-05, 0.0001757199, 0.00033527, 0.0002586997, 
    8.110624e-05, 1.578352e-05, 9.135305e-06, 1.490518e-05, 7.457012e-06,
  1.392472e-08, 6.388391e-09, 1.426104e-09, 6.672088e-10, 1.799913e-07, 
    6.420183e-07, 1.408077e-05, 7.31528e-05, 0.0002118415, 0.0001851363, 
    7.341737e-05, 1.450957e-05, 1.026055e-05, 1.27812e-05, 1.140562e-05,
  8.595491e-09, 8.817981e-08, 9.107258e-10, 3.467335e-10, 3.933629e-08, 
    5.985323e-07, 6.284359e-06, 3.013659e-05, 0.0001176359, 0.0001199278, 
    5.341792e-05, 1.455125e-05, 9.313137e-06, 8.537983e-06, 1.246129e-05,
  3.785968e-09, 3.765178e-09, 4.368855e-10, 1.865624e-10, 2.106798e-09, 
    9.805407e-08, 6.849261e-07, 1.483171e-05, 5.615248e-05, 6.770303e-05, 
    2.929691e-05, 1.496669e-05, 5.111469e-06, 5.376579e-06, 1.442583e-05,
  2.958543e-09, 5.008703e-09, 1.591556e-09, 5.688446e-10, 9.089919e-10, 
    8.11273e-09, 7.362828e-07, 1.350559e-05, 3.236955e-05, 5.305438e-05, 
    2.593913e-05, 1.889694e-05, 1.560286e-06, 5.764153e-06, 1.217998e-05,
  1.890088e-09, 4.999532e-09, 3.603104e-09, 3.403896e-09, 3.917345e-10, 
    6.449581e-09, 2.84294e-08, 1.001905e-07, 1.046507e-05, 4.187433e-05, 
    2.520283e-05, 1.474986e-05, 1.354123e-06, 3.342342e-06, 1.453919e-05,
  6.223536e-10, 3.265295e-09, 3.879929e-09, 1.364625e-07, 1.022512e-09, 
    1.944575e-09, 3.479498e-08, 1.346062e-07, 5.893999e-06, 2.966286e-05, 
    2.877157e-05, 1.22926e-05, 1.59356e-06, 2.654609e-06, 1.432088e-05,
  2.231747e-09, 3.521121e-08, 4.596203e-07, 2.24942e-07, 2.605572e-05, 
    9.871527e-05, 6.927653e-05, 3.483737e-05, 6.068821e-05, 4.760079e-05, 
    2.318519e-06, 1.96287e-05, 5.974527e-05, 1.178819e-05, 2.326803e-09,
  2.892212e-09, 4.93055e-08, 5.485603e-07, 1.46591e-07, 4.284246e-07, 
    1.991241e-05, 2.159844e-05, 4.088313e-05, 0.0001004508, 0.0001064807, 
    1.40716e-05, 7.110439e-05, 6.356472e-05, 1.068182e-06, 1.742887e-08,
  1.451779e-08, 9.075109e-08, 2.387699e-07, 7.256413e-07, 7.094286e-07, 
    4.702543e-06, 1.182734e-05, 5.530698e-05, 0.0001547536, 0.0001735303, 
    4.118641e-05, 4.334976e-05, 4.289479e-05, 4.588439e-06, 9.699092e-08,
  7.258448e-08, 2.738636e-07, 1.097216e-07, 8.724297e-07, 1.179922e-06, 
    3.489654e-06, 1.935958e-05, 8.196005e-05, 0.0002150623, 0.0002579117, 
    0.0001299766, 4.765869e-05, 2.071114e-05, 4.708533e-06, 3.474331e-07,
  2.182735e-08, 1.022127e-07, 1.549598e-07, 9.828042e-07, 5.364976e-07, 
    8.015601e-06, 3.174461e-05, 0.0001159224, 0.0002697106, 0.0003582877, 
    0.0002351255, 4.810511e-05, 1.502631e-05, 4.841048e-06, 1.711254e-06,
  3.742986e-08, 4.389772e-07, 2.313492e-07, 9.293123e-07, 3.563258e-06, 
    1.604368e-05, 5.820524e-05, 0.0001519977, 0.0003424214, 0.0004427656, 
    0.0003122036, 7.050715e-05, 7.485848e-06, 5.118128e-06, 4.97227e-06,
  3.902953e-08, 8.78816e-09, 1.197566e-06, 3.899342e-06, 6.878811e-06, 
    3.651037e-05, 5.079371e-05, 0.0001118294, 0.0003468938, 0.0005079382, 
    0.0003817351, 8.870783e-05, 5.207417e-06, 2.934571e-06, 5.976803e-06,
  2.55952e-08, 4.975743e-08, 2.440983e-06, 5.708654e-06, 8.216351e-06, 
    3.589855e-05, 7.275018e-05, 0.0002174645, 0.0004025476, 0.0005340429, 
    0.0004120409, 9.94619e-05, 6.457929e-06, 7.224612e-06, 8.571535e-06,
  1.993499e-08, 4.548346e-08, 2.947911e-06, 5.10468e-06, 9.121377e-06, 
    2.624347e-05, 3.248791e-05, 0.00014061, 0.0003367609, 0.0005314769, 
    0.0004128547, 0.0001454001, 8.307306e-06, 9.26417e-06, 8.063404e-06,
  1.477017e-08, 2.71812e-08, 2.438579e-06, 5.818148e-06, 7.922014e-06, 
    1.603238e-05, 4.410779e-05, 7.156548e-05, 0.0002805913, 0.0004832486, 
    0.0004090746, 0.0001825814, 1.912635e-05, 1.135932e-05, 1.409646e-05,
  1.87597e-06, 2.706586e-06, 9.223323e-06, 0.0001017567, 0.0003708006, 
    0.0005384845, 0.0004819381, 0.0003329223, 0.0001411269, 4.444973e-05, 
    5.137886e-06, 4.095721e-05, 0.0001605139, 1.968004e-05, 8.932522e-09,
  1.266757e-06, 5.412014e-06, 3.573268e-06, 5.734455e-05, 0.00030458, 
    0.0006557722, 0.000608624, 0.0003719733, 0.0001609383, 4.159001e-05, 
    1.068522e-05, 7.915006e-05, 0.0001816677, 2.49978e-07, 5.675879e-08,
  4.702467e-06, 9.978605e-06, 4.287734e-06, 2.049174e-05, 0.0001994897, 
    0.0006712244, 0.0006918593, 0.0004054323, 0.0001901856, 3.634616e-05, 
    8.040752e-05, 0.0002276445, 0.0001679553, 4.648996e-07, 6.509682e-08,
  3.554186e-06, 1.044901e-05, 1.583432e-06, 1.303659e-05, 0.0001322644, 
    0.0006303775, 0.0007315653, 0.0004193725, 0.0001881543, 4.062292e-05, 
    9.740058e-05, 0.0001977827, 0.0002231773, 1.11446e-05, 1.307515e-07,
  2.031524e-06, 6.421002e-06, 2.587168e-06, 1.479619e-05, 0.0001008755, 
    0.0005884492, 0.0007458376, 0.0004071471, 0.0001604173, 3.196243e-05, 
    0.000155066, 0.0002076707, 0.0001063361, 2.588104e-05, 5.033334e-07,
  5.339624e-06, 4.817055e-06, 2.207844e-06, 1.710084e-05, 0.0001053926, 
    0.0006037283, 0.0007692904, 0.0004386817, 0.000156191, 3.122595e-05, 
    9.82768e-05, 7.572943e-05, 6.960274e-05, 1.611306e-05, 2.018447e-06,
  1.198294e-06, 2.127058e-06, 4.922867e-06, 6.212389e-05, 0.000180567, 
    0.0006791918, 0.0007864712, 0.0003946416, 0.0001195868, 3.112648e-05, 
    1.576784e-05, 6.778939e-06, 1.803975e-06, 2.362548e-06, 3.760439e-06,
  6.009497e-06, 7.323064e-06, 2.3263e-05, 0.0001150783, 0.0002177037, 
    0.0006432915, 0.0007616791, 0.0004629017, 0.0001875123, 3.848686e-05, 
    2.346986e-05, 6.263326e-06, 5.818013e-06, 6.783206e-06, 7.826555e-06,
  1.911352e-05, 1.710066e-05, 4.062313e-05, 6.257881e-05, 0.0002653886, 
    0.0006834922, 0.0007816612, 0.0003076915, 6.711599e-05, 3.306381e-05, 
    2.110809e-05, 6.836457e-06, 7.249822e-06, 9.34557e-06, 8.23983e-06,
  3.611762e-05, 3.669671e-05, 6.973287e-05, 7.965604e-05, 0.000257779, 
    0.0006438264, 0.0008905987, 0.0004079516, 9.547479e-05, 3.013427e-05, 
    2.003549e-05, 9.212103e-06, 9.043233e-06, 7.390965e-06, 7.734864e-06,
  3.164435e-06, 1.862273e-06, 7.560811e-07, 1.034502e-06, 1.864512e-06, 
    1.911272e-06, 1.496761e-06, 1.98117e-06, 2.71772e-05, 0.0001111718, 
    0.0003549617, 0.0007004939, 0.0008451617, 0.0001093826, 4.052791e-05,
  9.089536e-06, 2.212587e-06, 3.473333e-06, 9.396246e-07, 1.236104e-06, 
    1.195283e-06, 1.714201e-06, 6.03812e-06, 1.447289e-05, 0.0001144188, 
    0.0003475481, 0.0007834539, 0.0008898228, 6.390476e-05, 7.131569e-06,
  2.87918e-05, 1.888293e-05, 2.326214e-06, 1.012671e-06, 1.540795e-06, 
    3.000133e-06, 3.033366e-06, 9.641961e-06, 6.749747e-06, 9.564237e-05, 
    0.0003139829, 0.0008178716, 0.0006852873, 9.316752e-05, 7.070748e-06,
  3.939031e-05, 2.266038e-05, 3.947679e-06, 1.59771e-06, 2.644791e-06, 
    4.178592e-06, 3.745593e-06, 1.272945e-05, 9.393937e-06, 6.913704e-05, 
    0.0002710748, 0.0008034359, 0.0007715367, 0.0001259336, 2.234514e-06,
  3.979596e-05, 1.245597e-05, 3.105581e-06, 1.625373e-06, 3.56089e-06, 
    5.976965e-06, 5.182007e-06, 1.644551e-05, 1.348948e-05, 5.839881e-05, 
    0.0002719529, 0.000813292, 0.0008464693, 0.0001845846, 1.025889e-07,
  2.481852e-05, 1.406607e-06, 1.584384e-07, 8.992642e-07, 3.345566e-06, 
    7.389449e-06, 9.2474e-06, 2.304339e-05, 1.62147e-05, 5.469253e-05, 
    0.0002833602, 0.000824129, 0.0008636781, 0.0003025251, 8.675601e-08,
  2.63357e-06, 4.233536e-07, 3.484712e-07, 2.104903e-06, 7.402382e-06, 
    1.19996e-05, 1.054354e-05, 3.063069e-05, 1.358443e-05, 4.500193e-05, 
    0.0003142193, 0.0007398002, 0.0007180519, 9.752146e-06, 1.996302e-07,
  6.68245e-06, 7.420348e-07, 1.081469e-06, 4.490879e-06, 9.131777e-06, 
    1.347553e-05, 2.706525e-05, 3.86052e-05, 1.686348e-05, 4.84187e-05, 
    0.0003542711, 0.0006227202, 0.0005913472, 7.971978e-06, 3.899317e-07,
  1.514876e-05, 1.977322e-06, 4.837257e-06, 5.753704e-06, 2.220035e-05, 
    1.260555e-05, 1.017005e-05, 3.085028e-06, 5.320492e-06, 4.613184e-05, 
    0.0003067386, 0.0005104642, 0.000469692, 4.597398e-06, 1.502352e-06,
  1.835942e-05, 8.400981e-06, 1.222649e-05, 6.290181e-06, 1.718738e-05, 
    2.13395e-05, 4.293805e-05, 1.762492e-05, 1.0113e-05, 4.965337e-05, 
    0.0002431203, 0.0004450129, 0.0003911409, 6.024974e-06, 5.639489e-06,
  1.546832e-11, 2.131757e-11, 4.188e-11, 6.099547e-13, 4.437261e-11, 
    8.42903e-10, 6.494527e-09, 7.303865e-09, 5.218581e-09, 7.859084e-08, 
    2.639164e-07, 3.310067e-07, 1.378847e-06, 1.655522e-06, 5.949359e-06,
  4.671619e-10, 2.160299e-10, 1.085202e-09, 6.672896e-12, 4.987203e-11, 
    4.062645e-10, 1.186416e-09, 8.412455e-11, 6.996394e-09, 2.374874e-08, 
    1.30604e-07, 8.063691e-08, 1.27333e-08, 1.285224e-06, 1.160475e-05,
  6.111816e-09, 8.618126e-10, 1.964848e-10, 5.481494e-12, 3.304805e-11, 
    2.77833e-10, 2.195797e-10, 1.652512e-09, 6.866841e-09, 8.646631e-09, 
    2.400362e-08, 6.50348e-07, 3.220594e-07, 2.921368e-06, 2.057853e-05,
  2.13877e-06, 2.704756e-06, 2.248364e-10, 2.797634e-12, 5.388366e-12, 
    5.978684e-11, 1.30904e-09, 2.811207e-09, 2.498195e-09, 5.384592e-09, 
    1.443094e-08, 6.456248e-07, 1.042651e-06, 1.572686e-05, 2.813146e-05,
  4.157895e-06, 1.823028e-06, 7.039506e-10, 7.248973e-12, 3.631608e-12, 
    1.627648e-10, 1.666104e-09, 2.618529e-09, 4.969306e-09, 6.844245e-09, 
    7.524696e-09, 3.698282e-07, 1.532637e-05, 5.123713e-05, 3.695346e-05,
  1.717853e-05, 1.194513e-06, 7.858786e-10, 6.934243e-12, 2.082622e-12, 
    3.04848e-12, 3.688587e-10, 2.293163e-09, 1.19636e-09, 8.819472e-10, 
    6.745908e-09, 1.037433e-05, 9.855549e-05, 0.0001056878, 4.279974e-05,
  5.385794e-09, 1.107324e-09, 1.195923e-11, 1.386802e-11, 2.131432e-12, 
    5.224964e-12, 8.109049e-11, 7.979903e-10, 1.689465e-10, 3.56347e-09, 
    6.124273e-09, 7.098186e-05, 0.0002349571, 0.00017923, 5.328397e-05,
  2.899464e-07, 1.684234e-08, 5.040186e-09, 4.98472e-09, 6.496696e-10, 
    2.663725e-11, 1.506008e-10, 1.609533e-09, 2.812867e-10, 1.009654e-09, 
    2.261622e-05, 0.0001813954, 0.0003419131, 0.0001802837, 5.559308e-05,
  4.832754e-06, 3.146335e-07, 8.236235e-09, 5.131733e-09, 1.532294e-08, 
    2.375552e-09, 1.625218e-10, 1.717264e-10, 1.868521e-10, 1.793223e-09, 
    0.0001192011, 0.0003279107, 0.0003956307, 0.0001485914, 4.747635e-05,
  4.325353e-06, 5.990677e-07, 2.440594e-08, 9.237886e-09, 9.574656e-09, 
    1.727514e-09, 2.149399e-10, 2.347981e-10, 1.089022e-09, 6.217827e-06, 
    0.0002518062, 0.000433489, 0.0003759629, 0.0001029433, 4.384604e-05,
  2.348521e-09, 2.382661e-08, 5.066694e-08, 6.047154e-08, 2.888915e-07, 
    2.592716e-07, 1.906846e-08, 8.690328e-08, 1.881133e-05, 6.355467e-05, 
    0.0001093663, 0.0001495433, 0.0001745849, 0.0002504186, 1.255407e-05,
  1.712525e-09, 3.608258e-09, 2.61501e-07, 1.918708e-07, 1.122098e-06, 
    1.741364e-07, 4.952664e-08, 1.497977e-08, 1.061925e-06, 3.361052e-05, 
    7.164454e-05, 0.0001009117, 0.0001132805, 0.0001350344, 2.379377e-05,
  5.185011e-08, 2.443989e-07, 1.441973e-07, 2.241558e-07, 3.893562e-07, 
    3.159516e-08, 7.520946e-08, 2.227718e-08, 1.600728e-08, 1.024754e-05, 
    4.703715e-05, 6.200848e-05, 4.988802e-05, 0.0001008039, 9.776486e-05,
  3.696959e-07, 3.696521e-07, 5.062931e-08, 2.023913e-07, 5.896881e-08, 
    2.491139e-08, 6.739112e-08, 2.716575e-08, 4.316938e-07, 3.961837e-08, 
    2.29439e-05, 5.463028e-05, 3.967399e-05, 3.757954e-05, 0.0001328244,
  1.023861e-06, 5.98573e-07, 2.076789e-07, 3.28528e-08, 2.030637e-09, 
    1.035647e-09, 1.515814e-08, 5.105829e-09, 3.097489e-07, 2.628759e-09, 
    2.673214e-06, 3.778578e-05, 3.014239e-05, 1.445017e-05, 0.0001053467,
  1.487337e-05, 5.527541e-07, 3.128044e-09, 4.789094e-10, 1.071231e-10, 
    1.283788e-09, 3.795895e-09, 1.233991e-09, 5.302271e-09, 5.639324e-09, 
    8.950026e-09, 1.455016e-05, 4.250661e-05, 1.006267e-05, 4.097795e-05,
  3.945018e-05, 3.392873e-06, 8.379485e-10, 1.27765e-11, 7.371048e-11, 
    9.919646e-10, 4.25954e-08, 1.093865e-07, 2.036735e-09, 4.207142e-09, 
    5.771564e-09, 1.227424e-06, 2.444141e-05, 1.743948e-05, 5.876125e-06,
  4.688018e-05, 2.921161e-05, 3.66753e-08, 7.27801e-09, 3.123934e-09, 
    8.740904e-11, 1.620137e-07, 2.394237e-07, 1.084289e-09, 1.733924e-09, 
    2.442128e-09, 4.746272e-08, 4.59184e-06, 1.360574e-05, 6.818063e-06,
  2.009603e-05, 2.413884e-05, 1.644778e-06, 3.033636e-08, 1.52239e-08, 
    1.42359e-10, 1.041954e-11, 5.995233e-10, 7.832505e-10, 4.776065e-10, 
    2.915693e-09, 3.116038e-08, 8.175464e-08, 5.640561e-06, 5.050652e-06,
  3.176147e-06, 1.911941e-06, 4.519773e-06, 7.37487e-08, 8.023671e-07, 
    1.209904e-07, 3.053011e-08, 1.685086e-10, 2.261973e-10, 2.274154e-10, 
    1.687411e-09, 6.590928e-09, 1.188337e-08, 8.69548e-07, 2.161726e-06,
  5.237882e-05, 3.979251e-05, 4.832092e-05, 4.593891e-05, 1.474534e-05, 
    5.745647e-05, 0.0002428459, 0.0005481198, 0.0008219758, 0.0008125615, 
    0.000488007, 0.000260512, 0.0002326778, 0.0001709381, 3.592221e-07,
  5.028665e-05, 4.884168e-05, 5.512417e-05, 4.29717e-05, 1.111343e-05, 
    1.911235e-05, 0.0001896905, 0.0005068305, 0.0007893821, 0.0008061898, 
    0.0005257184, 0.0003673553, 0.0003811603, 0.0001744904, 2.902073e-06,
  6.691147e-05, 5.226744e-05, 5.545537e-05, 2.83325e-05, 2.10878e-06, 
    9.562e-06, 0.0001243541, 0.0004457167, 0.000776171, 0.0008266564, 
    0.0005592708, 0.0004216843, 0.0003427017, 0.0002559886, 5.127651e-05,
  8.963329e-05, 4.110225e-05, 3.87793e-05, 7.965071e-06, 5.091391e-07, 
    9.611744e-07, 6.410043e-05, 0.0003440043, 0.0007753696, 0.0007849069, 
    0.0005626482, 0.0005034007, 0.000415814, 0.0003275127, 0.0002126687,
  8.384521e-05, 2.934939e-05, 2.09013e-05, 6.408881e-06, 3.465745e-06, 
    1.886401e-07, 3.433003e-05, 0.0002013918, 0.000689419, 0.0007737905, 
    0.0005969856, 0.0005298188, 0.0005023197, 0.0003462714, 0.0002130286,
  7.582177e-05, 2.313354e-05, 5.28258e-06, 3.393143e-06, 5.514421e-06, 
    1.148951e-06, 2.575327e-05, 0.0001009883, 0.0005006475, 0.0007690861, 
    0.0006499056, 0.0005223142, 0.0004263056, 0.0003029051, 0.0002950777,
  9.97633e-06, 7.866225e-06, 2.161788e-06, 1.358338e-06, 4.365501e-06, 
    9.855653e-06, 2.010514e-05, 6.655862e-05, 0.00030007, 0.0006547787, 
    0.0006117321, 0.0005385504, 0.0004227674, 0.0002287969, 0.0002339746,
  8.659979e-05, 3.178037e-05, 3.213505e-07, 4.506356e-07, 1.175385e-05, 
    1.538072e-05, 2.832458e-05, 4.857324e-05, 0.0001819319, 0.0004942303, 
    0.0006361153, 0.0005498831, 0.0004300053, 0.0002262741, 0.0001318277,
  0.0001352075, 6.086566e-05, 4.374175e-06, 2.234837e-07, 3.479678e-05, 
    2.055395e-05, 7.189143e-06, 1.60697e-05, 3.95237e-05, 0.0003308172, 
    0.0005533951, 0.0006087099, 0.0004818806, 0.0003105923, 0.0001182771,
  0.0001104809, 9.271559e-05, 2.583039e-05, 8.656264e-07, 1.841875e-05, 
    1.183343e-05, 1.198238e-05, 9.464184e-06, 1.061176e-05, 0.0001978805, 
    0.0004504296, 0.0005983079, 0.0005485507, 0.0004108184, 0.000163935,
  8.457447e-09, 7.429657e-07, 1.993714e-06, 5.061005e-06, 1.021171e-05, 
    4.079818e-06, 6.095877e-07, 4.50344e-07, 3.107628e-06, 8.533734e-06, 
    3.472044e-05, 6.049833e-05, 0.0001072176, 0.0002437016, 0.0002257992,
  1.554021e-07, 2.687115e-06, 4.747068e-06, 1.527217e-05, 1.781893e-05, 
    6.04418e-06, 2.004339e-06, 9.565449e-07, 4.600583e-06, 1.791481e-05, 
    5.884453e-05, 9.393509e-05, 8.143613e-05, 0.0001905292, 0.0002246419,
  2.841372e-06, 7.809716e-06, 1.522104e-05, 3.277552e-05, 3.077328e-05, 
    8.365942e-06, 2.110106e-06, 4.04978e-06, 8.890905e-06, 3.617202e-05, 
    0.0001028854, 0.0001337721, 9.442928e-05, 0.0001495185, 0.0002181019,
  4.937256e-06, 1.83163e-05, 4.170609e-05, 5.776717e-05, 2.034264e-05, 
    4.091502e-06, 3.14838e-06, 1.0005e-05, 5.801372e-05, 7.417801e-05, 
    0.0001337978, 0.0001549863, 0.0001066475, 0.000110872, 0.0001795823,
  7.467502e-06, 3.11022e-05, 8.37839e-05, 6.814013e-05, 2.702889e-05, 
    9.293874e-06, 5.047882e-06, 2.801066e-05, 0.0001329335, 0.00017835, 
    0.000201444, 0.0001349991, 0.0001212905, 8.693646e-05, 0.0001436604,
  1.003961e-05, 4.44867e-05, 0.0001143922, 9.633393e-05, 4.884817e-05, 
    1.838042e-05, 1.191846e-05, 5.390463e-05, 0.0002139544, 0.0003282197, 
    0.0001342176, 0.000106371, 0.0001157227, 9.576816e-05, 0.0001210732,
  3.307083e-06, 5.363976e-05, 0.0001195269, 9.244997e-05, 5.451004e-05, 
    2.826289e-05, 1.127389e-05, 6.014013e-05, 0.0002523406, 0.0005142224, 
    0.0002745035, 9.517663e-05, 0.0001008789, 8.691652e-05, 0.0001110508,
  3.744764e-06, 5.353663e-05, 9.02765e-05, 0.0001030396, 6.408425e-05, 
    3.59504e-05, 2.921859e-05, 9.398639e-05, 0.0002889625, 0.0005837294, 
    0.0004317505, 9.712451e-05, 8.600708e-05, 7.74338e-05, 0.0001055419,
  1.234714e-06, 4.685244e-05, 8.059429e-05, 0.0001535583, 0.0001149264, 
    3.556934e-05, 3.293612e-05, 9.530341e-05, 0.0002566397, 0.000595047, 
    0.0005870677, 0.0001250563, 6.194485e-05, 0.00010235, 0.0001024263,
  2.328411e-06, 4.769642e-05, 0.0001130792, 0.000219129, 0.0001654136, 
    5.202601e-05, 2.034763e-05, 0.0001092345, 0.0002353771, 0.0005569701, 
    0.0006933569, 0.0001700383, 4.127874e-05, 8.803955e-05, 9.995307e-05,
  1.167936e-09, 5.466798e-10, 9.657904e-10, 2.183251e-09, 7.621043e-10, 
    6.848796e-10, 1.232726e-10, 8.687221e-10, 5.999249e-09, 1.562981e-06, 
    2.782696e-05, 6.702662e-05, 0.0001172959, 0.0002470278, 0.0003460087,
  8.453329e-10, 7.967552e-10, 1.787115e-09, 1.66916e-09, 2.164528e-09, 
    9.270262e-10, 1.885024e-10, 5.963121e-11, 1.27142e-09, 3.45596e-08, 
    1.699152e-05, 9.27141e-05, 0.0001631866, 0.0002835691, 0.0003118683,
  9.508289e-10, 8.624786e-11, 3.189511e-10, 3.483079e-10, 5.018063e-10, 
    9.050417e-10, 4.713593e-10, 6.553016e-10, 1.131021e-10, 1.041946e-09, 
    1.052318e-06, 6.821234e-05, 0.0001658122, 0.0002739192, 0.0002723424,
  1.058861e-09, 2.891448e-09, 8.025693e-10, 3.111654e-12, 1.208735e-12, 
    3.108921e-10, 5.303278e-10, 6.127299e-10, 3.734933e-10, 1.642659e-10, 
    6.826703e-10, 2.397697e-05, 0.0001325634, 0.0002218185, 0.0002038086,
  8.824763e-10, 1.620261e-09, 1.029659e-09, 9.91181e-22, 1.118517e-10, 
    7.975586e-12, 4.565161e-10, 5.722142e-10, 4.324368e-10, 1.047469e-13, 
    2.038613e-10, 7.307842e-10, 6.551391e-05, 0.00013308, 0.0001104015,
  2.067601e-09, 1.5902e-09, 8.399283e-10, 7.49663e-11, 2.456968e-11, 
    1.958531e-10, 1.756699e-10, 1.428365e-10, 4.074595e-10, 6.067694e-11, 
    2.604168e-11, 7.2188e-10, 2.060807e-06, 5.23278e-05, 3.046065e-05,
  4.238765e-10, 1.257572e-09, 1.328035e-09, 3.172709e-10, 2.391959e-11, 
    3.134086e-15, 9.907908e-11, 5.52075e-11, 1.798266e-10, 7.819164e-11, 
    1.058297e-12, 1.062773e-10, 1.024596e-09, 1.090178e-06, 4.265353e-06,
  4.144394e-07, 7.26984e-09, 1.302634e-09, 4.515234e-10, 2.643594e-11, 
    1.38351e-12, 1.185498e-10, 3.18487e-10, 8.166093e-11, 1.35498e-10, 
    4.80239e-15, 1.040994e-13, 1.189985e-10, 2.737462e-09, 7.824934e-07,
  2.786409e-07, 6.154512e-09, 6.080669e-10, 1.04867e-10, 1.97046e-06, 
    3.39572e-10, 1.905869e-10, 2.556614e-10, 3.596223e-10, 1.495058e-10, 
    1.359411e-10, 2.823129e-16, 1.454448e-11, 7.713466e-09, 3.260505e-07,
  9.612484e-08, 7.018415e-09, 7.792693e-10, 6.625271e-11, 4.366436e-06, 
    4.093312e-07, 5.210237e-07, 1.849199e-10, 5.518738e-10, 3.168941e-10, 
    1.388501e-10, 1.746927e-11, 3.555178e-13, 2.714726e-08, 9.755617e-08,
  8.991361e-06, 8.60279e-06, 5.97308e-06, 1.072623e-06, 3.905232e-07, 
    1.763538e-06, 1.416766e-06, 1.205476e-06, 1.534284e-05, 6.568651e-05, 
    7.369313e-05, 7.449233e-05, 6.048479e-06, 1.263048e-06, 3.307509e-07,
  5.053113e-05, 3.489682e-05, 2.085766e-05, 4.315849e-06, 1.052765e-06, 
    5.747816e-07, 8.530513e-07, 7.917704e-07, 3.860642e-06, 4.516742e-05, 
    9.518127e-05, 0.0002019175, 2.951199e-05, 1.824552e-05, 3.768096e-06,
  8.397042e-05, 6.50599e-05, 3.823164e-05, 1.40041e-05, 1.673443e-06, 
    7.524873e-07, 6.214077e-07, 3.318831e-07, 2.016717e-06, 3.088597e-05, 
    0.0001199148, 0.0002080808, 0.0001352039, 0.0001024916, 5.507612e-05,
  8.743539e-05, 6.991943e-05, 4.381869e-05, 2.117808e-05, 8.259729e-06, 
    2.222402e-06, 2.20067e-06, 2.464168e-07, 1.587376e-06, 1.249814e-05, 
    0.0001257135, 0.0003482501, 0.000302375, 0.000241479, 0.0001524629,
  6.749856e-05, 4.912528e-05, 4.611193e-05, 1.960399e-05, 8.563336e-06, 
    3.226668e-06, 3.479208e-06, 8.361436e-07, 2.23073e-06, 5.611952e-06, 
    0.0001325383, 0.0004126887, 0.0005318146, 0.0004611286, 0.0003412713,
  5.318148e-05, 4.027528e-05, 3.532321e-05, 1.507237e-05, 5.257751e-06, 
    4.215235e-06, 1.655721e-06, 4.368933e-07, 1.426856e-06, 7.333575e-06, 
    0.0001418485, 0.0004406403, 0.0007346055, 0.0006976778, 0.0005217767,
  5.737211e-05, 4.610344e-05, 3.422426e-05, 1.593686e-05, 5.507009e-06, 
    8.12326e-06, 2.727374e-06, 2.085186e-06, 1.546364e-06, 1.447827e-05, 
    0.0001448088, 0.0004645442, 0.0007487203, 0.000817463, 0.0006474215,
  0.0001289322, 6.926938e-05, 4.019147e-05, 1.387664e-05, 5.062128e-06, 
    3.38677e-06, 2.772825e-06, 1.497194e-06, 5.087363e-05, 4.203966e-05, 
    0.0001736008, 0.0004540439, 0.0007134349, 0.0008469131, 0.0006338685,
  0.0001538407, 7.96744e-05, 3.076897e-05, 8.305075e-06, 9.495397e-06, 
    9.813106e-07, 8.555186e-07, 2.645339e-05, 0.0001238134, 7.843972e-05, 
    0.0001869711, 0.0004385813, 0.0006514217, 0.0007889995, 0.0006210055,
  0.0001307533, 6.363137e-05, 1.88264e-05, 2.967843e-06, 3.372e-06, 
    1.595093e-06, 4.269195e-06, 0.0001051614, 0.000192315, 9.457066e-05, 
    0.000151414, 0.0003769684, 0.0005811211, 0.0006701572, 0.0005536096,
  8.029801e-13, 7.641189e-25, 1.665318e-23, 1.199924e-12, 2.636349e-11, 
    8.250253e-10, 2.929078e-08, 2.025464e-06, 6.622433e-05, 0.0002164257, 
    0.0003871885, 0.0004208188, 8.057964e-05, 1.54371e-05, 1.370991e-05,
  1.212611e-11, 2.903205e-12, 7.224255e-14, 7.276151e-12, 2.63921e-11, 
    5.660797e-11, 3.403574e-09, 5.152223e-07, 3.957024e-05, 0.0001746744, 
    0.0003982231, 0.0005303546, 0.0001585857, 2.917879e-05, 1.482456e-05,
  2.189193e-10, 3.984537e-11, 3.345832e-12, 2.675444e-12, 3.696469e-10, 
    5.291473e-11, 6.645688e-10, 2.688673e-07, 2.093791e-05, 0.0001446722, 
    0.0003708391, 0.0004740406, 0.0003208565, 4.591899e-05, 1.51477e-05,
  1.311153e-06, 4.424867e-09, 2.878704e-12, 3.213778e-12, 5.038398e-09, 
    7.39629e-10, 7.081788e-10, 6.463317e-07, 6.151429e-06, 0.0001199032, 
    0.0003086354, 0.0004816141, 0.0004556393, 6.941213e-05, 1.723107e-05,
  9.398202e-08, 2.61401e-09, 1.222189e-09, 1.690724e-09, 1.080467e-07, 
    5.460206e-09, 1.05956e-09, 9.163965e-07, 4.902777e-06, 6.667904e-05, 
    0.0002567871, 0.0004291802, 0.0005195795, 0.0001606099, 2.559232e-05,
  1.748072e-07, 1.091173e-08, 2.244499e-10, 1.249543e-07, 6.154234e-07, 
    2.987736e-08, 9.076027e-08, 4.731873e-07, 1.458563e-06, 3.974516e-05, 
    0.0002238833, 0.000396182, 0.0005774485, 0.0002788716, 3.857734e-05,
  2.64146e-08, 5.503567e-09, 2.579229e-07, 6.358537e-07, 7.535101e-07, 
    9.744475e-07, 3.044527e-06, 1.289296e-05, 5.03971e-06, 1.770344e-05, 
    0.0001747559, 0.0003640775, 0.0006196083, 0.0004025927, 4.593743e-05,
  8.586136e-07, 1.865315e-06, 1.917023e-06, 2.446242e-06, 2.924821e-06, 
    5.772228e-06, 1.206332e-05, 1.357785e-05, 1.116334e-05, 5.012125e-06, 
    0.0001229242, 0.000329527, 0.0005574372, 0.0004867431, 6.380193e-05,
  5.456203e-06, 2.333979e-06, 6.856636e-06, 1.064047e-05, 3.815152e-05, 
    1.27898e-05, 4.1174e-06, 1.51465e-06, 4.558611e-10, 1.20831e-06, 
    8.174501e-05, 0.000289222, 0.0004242218, 0.0005047935, 0.0001187571,
  3.183385e-06, 5.159746e-06, 1.621182e-05, 2.286338e-05, 2.859914e-05, 
    1.504509e-05, 2.097947e-05, 6.693016e-06, 2.826065e-06, 1.591633e-06, 
    5.815492e-05, 0.0002519056, 0.000301312, 0.0004699484, 0.0001976447,
  2.733811e-10, 6.393364e-09, 1.262761e-07, 3.935992e-06, 5.195498e-06, 
    2.08584e-06, 1.062089e-06, 2.105755e-07, 1.389346e-08, 2.146372e-08, 
    2.478021e-08, 3.431817e-06, 3.83249e-05, 5.163089e-05, 2.470583e-05,
  4.466618e-11, 5.927604e-10, 3.32871e-09, 5.491871e-07, 3.725482e-06, 
    2.816528e-06, 6.293108e-07, 6.649807e-08, 1.92699e-08, 1.300977e-09, 
    1.991205e-09, 6.915315e-07, 1.88245e-05, 4.17258e-05, 3.542339e-05,
  1.447011e-11, 4.394002e-11, 1.137448e-09, 3.746782e-09, 1.20247e-06, 
    2.547511e-06, 1.769766e-06, 2.371353e-07, 1.006511e-08, 1.809705e-09, 
    1.46765e-09, 5.764104e-09, 4.107036e-06, 3.172374e-05, 4.060618e-05,
  1.077061e-06, 1.075822e-07, 1.263637e-10, 8.079734e-10, 4.835835e-08, 
    1.412151e-06, 2.019147e-06, 1.027101e-06, 2.108193e-08, 1.677784e-09, 
    5.870155e-10, 6.574588e-10, 4.590576e-07, 1.558874e-05, 3.136214e-05,
  3.611787e-07, 1.421254e-07, 2.48245e-11, 7.969254e-11, 1.58473e-09, 
    2.596113e-07, 1.12743e-06, 1.285744e-06, 1.868275e-07, 2.381004e-09, 
    2.96279e-10, 2.568643e-10, 6.84903e-09, 4.333401e-06, 1.446817e-05,
  7.339876e-08, 9.335134e-10, 5.765177e-10, 3.359813e-11, 9.145811e-11, 
    1.975408e-08, 2.13704e-07, 4.870253e-07, 4.097303e-07, 3.084644e-08, 
    5.216129e-10, 1.211742e-10, 1.977226e-09, 7.622921e-07, 5.480063e-06,
  6.040726e-10, 5.123355e-10, 5.769219e-10, 4.324273e-10, 7.446195e-11, 
    5.715604e-08, 5.498799e-09, 8.978938e-09, 9.561748e-09, 1.191505e-08, 
    1.32498e-09, 2.147033e-10, 4.659143e-10, 2.351314e-08, 2.74267e-06,
  7.246441e-08, 2.570784e-09, 1.477763e-09, 1.24072e-09, 6.529838e-09, 
    3.086278e-07, 4.356828e-07, 3.578565e-09, 1.459031e-09, 1.185247e-09, 
    1.047701e-09, 3.567344e-10, 1.234789e-10, 2.481927e-09, 3.845796e-07,
  2.064775e-08, 1.79307e-09, 8.576546e-08, 6.021256e-08, 8.772221e-06, 
    1.358947e-06, 2.027762e-10, 6.118614e-10, 8.761982e-10, 6.184627e-10, 
    4.600476e-10, 5.425872e-10, 7.303898e-10, 2.969187e-09, 2.382855e-08,
  3.124289e-06, 4.871003e-06, 5.127974e-06, 3.423188e-06, 1.219521e-05, 
    1.158873e-06, 1.096532e-06, 2.451704e-12, 4.857977e-10, 1.104376e-09, 
    7.32893e-10, 4.217248e-10, 5.410604e-08, 1.357243e-09, 5.181926e-09,
  1.798894e-08, 1.893349e-08, 1.798266e-08, 9.782573e-08, 1.236339e-05, 
    3.521301e-05, 4.772808e-05, 6.079544e-05, 6.218667e-05, 3.094335e-05, 
    3.387926e-06, 3.240911e-06, 7.969647e-07, 1.335792e-06, 1.083148e-06,
  5.460158e-08, 2.207017e-07, 4.028019e-08, 1.139134e-08, 7.807647e-07, 
    1.031179e-05, 9.409574e-06, 8.028347e-06, 3.828577e-05, 4.052161e-05, 
    8.045608e-06, 1.15923e-06, 1.287532e-07, 1.966563e-07, 2.781155e-06,
  2.76332e-07, 1.58697e-07, 1.426861e-07, 1.383592e-09, 4.498446e-08, 
    5.391449e-07, 3.087764e-06, 1.328045e-07, 1.156999e-05, 2.821359e-05, 
    2.338314e-05, 5.754463e-07, 4.521398e-07, 3.085173e-08, 2.521131e-06,
  1.37564e-06, 9.636358e-07, 1.500116e-08, 8.368941e-09, 1.284028e-09, 
    3.548957e-07, 8.334092e-07, 3.954883e-08, 6.68438e-08, 9.461868e-06, 
    2.910251e-05, 5.660826e-06, 9.005e-08, 3.711544e-08, 1.21102e-06,
  1.872289e-06, 3.550836e-06, 1.082443e-06, 1.692878e-08, 3.296292e-09, 
    4.316044e-08, 9.532019e-07, 1.117688e-06, 3.114504e-08, 6.358563e-08, 
    1.121805e-05, 1.245395e-05, 4.881234e-07, 2.693167e-08, 2.312555e-07,
  2.280514e-06, 3.483238e-06, 8.30801e-08, 3.231835e-08, 7.816763e-09, 
    2.959307e-09, 2.502793e-07, 1.695831e-06, 1.685196e-06, 1.368426e-08, 
    4.318797e-07, 6.423011e-06, 4.150633e-06, 9.630758e-08, 1.266153e-07,
  1.39248e-09, 1.71568e-08, 4.35098e-08, 9.876272e-08, 4.803312e-08, 
    1.843263e-08, 1.087712e-08, 4.028091e-07, 1.471359e-06, 1.363777e-07, 
    6.112824e-09, 1.55699e-06, 4.751948e-06, 5.951127e-07, 1.83079e-07,
  5.273756e-08, 3.924667e-08, 1.78698e-08, 6.197484e-08, 1.514862e-08, 
    2.220853e-07, 7.91765e-07, 2.1624e-07, 5.803518e-07, 4.294683e-07, 
    5.768885e-09, 3.596597e-07, 2.717108e-06, 1.289217e-06, 4.628383e-08,
  1.340747e-06, 2.773075e-06, 2.824241e-06, 2.525144e-07, 2.465202e-06, 
    5.452091e-08, 1.349632e-08, 2.644796e-09, 1.589815e-07, 4.300078e-07, 
    9.111666e-08, 2.095903e-09, 7.427262e-07, 1.39185e-06, 1.130046e-07,
  2.646963e-06, 5.595623e-06, 4.030006e-06, 3.655169e-06, 9.731575e-06, 
    7.835955e-07, 4.140936e-07, 4.11847e-09, 5.139032e-08, 2.864583e-07, 
    1.377101e-07, 8.212499e-09, 1.175641e-07, 8.920602e-07, 4.972022e-08,
  2.788389e-08, 7.086038e-09, 6.821283e-08, 2.949929e-07, 3.576529e-05, 
    7.617111e-05, 0.0001548973, 0.0002728883, 0.000407231, 0.0006378028, 
    0.0004255622, 0.0001127561, 8.101791e-06, 1.192171e-06, 1.232567e-07,
  1.054112e-06, 1.34779e-07, 4.238562e-08, 2.119377e-07, 4.219378e-06, 
    5.959833e-05, 0.0001166701, 0.00018319, 0.000232423, 0.0003548639, 
    0.0004019447, 0.0002354474, 6.302035e-05, 2.164926e-06, 3.241542e-07,
  1.199084e-05, 1.441256e-05, 6.098236e-06, 2.520419e-07, 8.054154e-08, 
    2.03106e-05, 9.552702e-05, 0.0001484303, 0.0001519087, 0.0001777461, 
    0.000252092, 0.0002226097, 0.000103751, 1.144917e-05, 2.773785e-06,
  1.188499e-05, 1.418038e-05, 5.464765e-06, 6.505564e-08, 3.228449e-08, 
    5.026204e-07, 5.129722e-05, 0.0001316467, 0.0001485456, 0.0001205429, 
    0.0001319159, 0.0001649853, 0.0001092908, 2.824577e-05, 5.051453e-06,
  4.616022e-06, 9.564365e-06, 7.237646e-06, 1.910047e-07, 1.768227e-07, 
    1.086071e-08, 1.019796e-05, 7.769861e-05, 0.0001187406, 9.471796e-05, 
    6.847537e-05, 9.852445e-05, 0.0001075889, 4.474639e-05, 6.166122e-06,
  3.270889e-06, 3.503657e-06, 1.141718e-06, 6.349181e-07, 7.005196e-07, 
    9.607665e-09, 7.80915e-08, 3.906193e-05, 7.806429e-05, 9.361714e-05, 
    5.198784e-05, 4.284178e-05, 8.309303e-05, 7.807204e-05, 1.056368e-05,
  8.865522e-08, 6.231705e-07, 1.468589e-06, 2.248945e-06, 3.202466e-07, 
    9.240964e-08, 4.479125e-09, 4.107491e-06, 5.387281e-05, 8.525045e-05, 
    5.665013e-05, 2.542355e-05, 4.030636e-05, 7.513884e-05, 4.39198e-05,
  9.521054e-08, 2.488734e-07, 1.120583e-06, 2.680823e-06, 2.543581e-07, 
    7.277716e-08, 1.421088e-06, 7.291121e-07, 3.05575e-05, 6.293706e-05, 
    6.773798e-05, 3.150409e-05, 1.518013e-05, 4.965789e-05, 5.12661e-05,
  7.48382e-08, 3.651034e-07, 1.712565e-06, 2.136456e-06, 3.070837e-06, 
    2.025874e-06, 3.527589e-07, 3.179083e-07, 2.364965e-06, 3.320978e-05, 
    4.123448e-05, 2.696408e-05, 1.041392e-05, 1.634669e-05, 3.876872e-05,
  5.751435e-10, 4.086756e-08, 6.688916e-07, 2.320784e-06, 1.433742e-06, 
    3.201532e-06, 1.393468e-06, 8.086366e-07, 3.546988e-06, 8.149869e-06, 
    2.336997e-05, 2.040708e-05, 9.875057e-06, 1.142945e-05, 2.33264e-05,
  1.315986e-08, 3.247387e-08, 4.10296e-08, 4.659292e-08, 6.327282e-08, 
    5.862937e-08, 8.266718e-08, 1.098678e-06, 6.054812e-05, 0.0002246174, 
    0.0002396504, 0.0002223263, 0.0001339599, 2.450301e-06, 2.527872e-07,
  3.310448e-09, 2.939774e-09, 4.369594e-09, 3.415465e-08, 6.591196e-09, 
    1.415149e-08, 2.600475e-08, 8.947762e-08, 5.685148e-06, 0.0001583354, 
    0.0004685021, 0.000561082, 0.0004471408, 9.715863e-05, 4.497071e-06,
  2.48832e-07, 8.184778e-10, 2.632264e-09, 5.378678e-09, 3.53677e-09, 
    3.093255e-09, 6.844336e-09, 2.482475e-07, 3.357586e-06, 3.572592e-05, 
    0.0003940709, 0.001051736, 0.001046374, 0.0005257471, 4.239987e-05,
  5.330187e-10, 4.400841e-10, 4.095111e-10, 8.260649e-10, 1.029077e-09, 
    1.13561e-08, 2.568447e-07, 4.08054e-06, 5.604779e-06, 1.317207e-05, 
    9.188252e-05, 0.0007200027, 0.001522359, 0.001299814, 0.000384911,
  1.058135e-09, 1.058023e-09, 1.643522e-10, 4.550616e-09, 3.305952e-10, 
    2.175539e-08, 2.791433e-07, 3.697685e-06, 1.179592e-05, 1.434765e-05, 
    1.904118e-05, 7.832533e-05, 0.000747797, 0.001201793, 0.000656906,
  6.478093e-10, 1.49195e-09, 1.432333e-11, 4.538042e-10, 8.775634e-10, 
    2.647981e-08, 3.275188e-07, 9.525338e-07, 2.936697e-06, 1.074444e-05, 
    1.468677e-05, 7.033128e-06, 5.386788e-06, 0.0001099294, 0.0002381954,
  2.159024e-10, 4.138902e-10, 3.120263e-10, 4.466827e-10, 1.036648e-09, 
    1.250065e-10, 8.968629e-09, 9.984111e-08, 1.197761e-07, 6.064354e-06, 
    1.132216e-05, 1.053025e-05, 5.11023e-06, 5.623574e-06, 3.120076e-05,
  7.278072e-10, 6.900101e-09, 1.718346e-09, 6.071833e-10, 2.129733e-10, 
    4.777946e-10, 1.681231e-07, 6.140616e-06, 3.528383e-06, 1.399663e-06, 
    9.493277e-06, 1.008252e-05, 4.483451e-06, 2.107277e-06, 5.243992e-06,
  1.626705e-09, 7.619049e-10, 1.437325e-09, 9.028657e-10, 6.203738e-10, 
    1.85656e-08, 1.447291e-09, 2.204426e-07, 3.231298e-07, 1.490088e-06, 
    1.664819e-06, 4.644437e-06, 1.968433e-06, 8.282502e-07, 1.783748e-06,
  2.504537e-09, 2.659475e-10, 1.667102e-08, 1.468674e-08, 7.731306e-08, 
    2.75501e-08, 3.548812e-08, 2.16991e-10, 6.396543e-07, 7.585843e-07, 
    1.059482e-06, 1.542389e-06, 1.59923e-06, 3.802383e-07, 1.295506e-06,
  3.095361e-05, 2.783201e-05, 1.631525e-05, 1.261523e-05, 1.00255e-05, 
    9.002109e-06, 8.4211e-06, 7.649995e-06, 5.470681e-06, 3.532958e-06, 
    2.708944e-06, 3.400874e-05, 0.0001310096, 2.510806e-05, 7.65302e-08,
  1.338762e-05, 1.886036e-05, 2.382763e-05, 1.987788e-05, 1.451878e-05, 
    1.031529e-05, 9.412552e-06, 1.219673e-05, 2.167221e-05, 3.127473e-05, 
    6.159542e-05, 9.338469e-05, 7.501902e-05, 3.75664e-06, 1.995569e-07,
  1.736771e-05, 5.090276e-05, 4.981669e-05, 2.928024e-05, 2.793683e-05, 
    2.387264e-05, 2.404313e-05, 3.081955e-05, 6.461421e-05, 0.0001488699, 
    0.0002278019, 0.0002115102, 9.230985e-05, 5.772844e-06, 6.273514e-07,
  6.53354e-05, 6.926526e-05, 5.117091e-05, 4.389407e-05, 4.333282e-05, 
    4.217516e-05, 4.619033e-05, 4.699397e-05, 6.508585e-05, 0.0001863541, 
    0.0003208347, 0.0003104347, 0.0001634703, 0.0001468649, 4.87215e-05,
  6.853854e-05, 6.114855e-05, 5.128671e-05, 3.274625e-05, 2.596922e-05, 
    3.250023e-05, 4.238345e-05, 6.198083e-05, 7.403139e-05, 0.0001496046, 
    0.0003789652, 0.0005532542, 0.0005275027, 0.0001576311, 7.525048e-07,
  4.744277e-05, 3.704093e-05, 2.224956e-05, 1.632322e-05, 9.879773e-06, 
    1.244749e-05, 2.147695e-05, 4.570705e-05, 8.054038e-05, 0.0001139857, 
    0.0002342003, 0.0005888647, 0.0003273197, 1.212549e-06, 5.226029e-06,
  1.932862e-06, 2.538801e-06, 1.923764e-06, 5.937855e-06, 3.721303e-06, 
    1.007078e-05, 6.308097e-06, 1.172136e-05, 4.862213e-05, 7.823452e-05, 
    1.972082e-05, 0.0001883724, 0.0001287847, 4.159002e-07, 9.596836e-07,
  5.215431e-08, 3.05471e-08, 2.037439e-07, 1.828123e-07, 2.008375e-07, 
    1.529555e-06, 1.000872e-05, 3.91946e-05, 5.426514e-05, 3.619271e-05, 
    8.39154e-06, 2.224395e-06, 5.205576e-07, 2.795279e-07, 5.995166e-07,
  7.088822e-08, 9.034715e-09, 2.782167e-08, 1.337218e-07, 2.226993e-06, 
    4.758395e-06, 3.788941e-06, 3.384851e-06, 4.616213e-06, 9.211675e-06, 
    4.458997e-06, 1.669464e-06, 1.215881e-06, 8.104065e-07, 1.753735e-06,
  2.031932e-07, 1.161027e-08, 4.031181e-08, 4.365662e-07, 1.121037e-06, 
    4.049391e-06, 1.572017e-05, 5.91433e-06, 9.500278e-06, 6.915882e-06, 
    4.465267e-06, 1.469319e-06, 1.116166e-06, 5.514366e-07, 1.817455e-06,
  0.0003341956, 0.0003042115, 0.000176608, 3.95329e-05, 2.561093e-05, 
    4.829344e-05, 8.651305e-05, 0.0001521829, 5.093756e-05, 1.282104e-06, 
    1.934829e-08, 1.030467e-05, 9.704071e-06, 3.641343e-08, 2.676383e-08,
  0.000348338, 0.0003759645, 0.0002704877, 0.0001053541, 6.32327e-05, 
    7.953903e-05, 0.0001163307, 0.0001835669, 8.507378e-05, 4.549728e-07, 
    2.80114e-08, 1.212515e-05, 1.740083e-05, 4.101175e-07, 1.087241e-08,
  0.000363535, 0.0004880313, 0.0003957244, 0.0002012299, 0.0001105883, 
    0.000116309, 0.0001385343, 0.0001982738, 0.0001060448, 5.501511e-07, 
    1.101481e-06, 5.788711e-06, 2.696513e-06, 9.32735e-07, 5.656843e-08,
  0.0003697322, 0.0005890836, 0.000544839, 0.000349301, 0.0001738622, 
    0.000162586, 0.0001527669, 0.0001888059, 0.0001098113, 5.45002e-07, 
    2.152393e-06, 2.998293e-06, 1.283189e-06, 2.050015e-06, 2.032612e-07,
  0.0003713188, 0.000670683, 0.0006973978, 0.0004714626, 0.0002508122, 
    0.0001959539, 0.0001907172, 0.000182956, 0.0001130991, 1.68124e-06, 
    3.642214e-06, 3.83995e-06, 1.51391e-06, 1.607133e-07, 1.526274e-07,
  0.0004707635, 0.0007244647, 0.000768367, 0.0005245481, 0.0003023804, 
    0.0002052559, 0.0002384212, 0.0002171194, 0.0001166074, 3.312377e-06, 
    5.911667e-06, 6.769247e-06, 6.991986e-06, 1.917556e-06, 1.00775e-06,
  0.0005848673, 0.000774068, 0.0007885518, 0.0005520997, 0.0003236958, 
    0.0002781901, 0.0002469204, 0.0002335927, 0.0001166243, 5.04275e-06, 
    4.993719e-06, 8.879137e-06, 6.211279e-06, 2.992022e-06, 1.428011e-06,
  0.0006844501, 0.000896718, 0.0008338032, 0.0006330985, 0.0003508981, 
    0.0002344721, 0.0002652596, 0.0003275154, 0.0001996216, 2.009366e-05, 
    8.549849e-06, 8.541752e-06, 6.58405e-06, 5.081088e-06, 2.530643e-06,
  0.0006970573, 0.0009487399, 0.0008743419, 0.0005894176, 0.0005430861, 
    0.0003431562, 0.0001972384, 0.0001315483, 0.0001330967, 2.837396e-05, 
    1.098306e-05, 9.615545e-06, 6.391425e-06, 4.621336e-06, 5.649553e-06,
  0.0006338623, 0.0009255067, 0.0009504699, 0.0005781421, 0.0004571948, 
    0.0003605382, 0.0003933342, 0.0003214437, 0.0002370277, 5.1568e-05, 
    1.003819e-05, 9.361878e-06, 5.487574e-06, 4.769184e-06, 6.58728e-06,
  3.648939e-06, 5.207614e-06, 2.004701e-06, 1.564398e-06, 7.27173e-06, 
    9.033953e-06, 2.690301e-06, 9.344259e-06, 4.006063e-05, 7.539098e-05, 
    6.217059e-05, 8.153141e-05, 0.0002742616, 3.061714e-05, 1.441994e-08,
  2.484161e-06, 1.957926e-06, 1.305009e-06, 3.048198e-07, 4.363279e-07, 
    4.415091e-07, 1.212735e-06, 1.342175e-06, 1.76708e-05, 4.071188e-05, 
    5.550179e-05, 0.0001553287, 0.0001630061, 3.108142e-08, 8.953347e-09,
  3.072791e-06, 9.571191e-07, 1.397446e-07, 7.175274e-08, 1.776681e-07, 
    1.495684e-06, 2.407849e-06, 2.089236e-06, 1.240764e-05, 2.60267e-05, 
    3.892524e-05, 0.0002013144, 4.154351e-07, 2.49455e-08, 1.098669e-08,
  3.307518e-06, 3.036594e-07, 7.508901e-08, 2.673254e-07, 1.11471e-06, 
    2.265247e-06, 2.200584e-06, 2.639358e-06, 2.037784e-05, 2.886106e-05, 
    5.595619e-05, 0.0001029878, 1.851938e-07, 1.249754e-06, 1.762859e-06,
  6.363163e-07, 6.102222e-08, 5.926004e-07, 2.436194e-06, 2.095591e-06, 
    2.753468e-06, 2.684058e-06, 5.754793e-06, 5.380787e-05, 3.457377e-05, 
    1.796951e-05, 2.512645e-05, 5.562178e-07, 1.566209e-06, 2.625036e-06,
  3.666107e-07, 1.442525e-07, 1.069156e-07, 7.663573e-07, 4.176884e-06, 
    2.435544e-06, 1.299047e-06, 7.878057e-06, 9.377104e-05, 8.427254e-05, 
    2.850584e-05, 4.160781e-05, 4.550501e-08, 2.613199e-07, 2.2446e-06,
  5.117518e-08, 2.508826e-10, 3.603603e-09, 1.965281e-07, 1.643403e-06, 
    3.285837e-06, 2.702032e-07, 7.792315e-07, 8.319454e-05, 0.0001302534, 
    4.769324e-05, 5.087033e-06, 6.905354e-08, 1.263491e-07, 1.655851e-06,
  1.640736e-08, 1.421101e-08, 2.011737e-08, 1.37108e-07, 1.653061e-06, 
    9.660961e-06, 2.382546e-06, 5.300029e-06, 7.396024e-05, 0.0001250375, 
    9.151155e-05, 2.413969e-05, 2.624352e-07, 1.322534e-06, 3.777897e-06,
  1.361773e-07, 1.587803e-07, 3.419094e-08, 2.798879e-07, 5.587082e-06, 
    4.492448e-06, 3.616103e-07, 9.7561e-07, 9.843056e-06, 0.000124631, 
    0.0001202565, 5.541864e-05, 1.577221e-06, 1.989278e-06, 1.855734e-06,
  1.22688e-06, 5.232995e-07, 1.583514e-07, 4.928204e-07, 2.841884e-06, 
    3.810075e-06, 9.736234e-06, 4.695721e-06, 4.081212e-05, 0.0001501419, 
    0.0001443236, 7.877596e-05, 5.832354e-06, 7.368743e-07, 1.498756e-06,
  6.880662e-08, 5.125942e-07, 1.849453e-06, 6.633222e-07, 2.662655e-06, 
    5.523501e-06, 1.886256e-05, 0.0002957818, 0.0002853566, 7.751245e-05, 
    1.347479e-05, 0.00021107, 0.0002006434, 9.117621e-05, 1.692817e-08,
  2.110069e-08, 9.457255e-08, 3.170769e-07, 1.850932e-07, 9.671877e-07, 
    3.812378e-06, 7.137077e-06, 0.0001029585, 0.0003680407, 0.0002402498, 
    0.0002254081, 0.0002074771, 0.0001296628, 2.394363e-05, 4.850409e-08,
  1.689595e-09, 2.768555e-08, 9.989704e-08, 1.183056e-07, 2.548216e-07, 
    1.462156e-06, 5.648666e-06, 1.534156e-05, 0.0003215898, 0.0004435374, 
    0.0003829903, 0.000329312, 0.0001068352, 3.165478e-07, 5.759784e-08,
  4.469773e-10, 1.50164e-09, 2.344396e-08, 8.692027e-08, 6.78266e-08, 
    4.496075e-07, 4.114018e-06, 1.006969e-05, 5.993522e-05, 0.0004906188, 
    0.0004359164, 0.0001377533, 8.772231e-05, 5.17637e-05, 1.538007e-05,
  4.061105e-12, 3.961481e-11, 1.098741e-09, 4.612439e-08, 7.488632e-08, 
    2.72163e-07, 2.027921e-06, 8.770648e-06, 2.011242e-05, 0.0004196949, 
    0.0005201184, 0.0002222647, 4.491599e-05, 6.175638e-06, 2.091004e-06,
  1.119079e-11, 8.837129e-13, 1.374566e-11, 4.144855e-09, 1.01056e-07, 
    9.486401e-08, 2.024226e-07, 3.27982e-06, 1.987644e-05, 0.0001439865, 
    0.0005823128, 0.0004254649, 6.769048e-05, 2.190146e-05, 4.5137e-06,
  1.697799e-16, 2.630202e-21, 6.160302e-21, 3.736953e-14, 6.395189e-08, 
    2.056691e-08, 2.205989e-08, 3.622152e-07, 1.6346e-05, 5.798326e-05, 
    0.0005007769, 0.0005264717, 0.0001240824, 1.207802e-05, 9.561792e-06,
  2.261518e-22, 4.52259e-22, 9.91992e-22, 1.555193e-16, 1.378004e-08, 
    1.223137e-07, 9.294157e-09, 3.864677e-08, 4.970485e-06, 1.831505e-05, 
    0.0001387639, 0.0005705198, 0.0003084966, 3.611402e-05, 8.963876e-06,
  4.460203e-23, 1.673719e-22, 3.627106e-22, 1.629977e-12, 8.529814e-07, 
    3.472162e-08, 4.049399e-09, 3.356829e-09, 2.421578e-08, 6.322872e-06, 
    3.740045e-05, 0.0003206567, 0.0004331115, 0.0001122892, 6.937958e-06,
  2.599546e-15, 1.853629e-23, 5.137784e-23, 2.433471e-12, 1.319924e-06, 
    7.004098e-08, 6.647871e-10, 1.18634e-09, 2.291975e-09, 3.462002e-07, 
    1.730412e-05, 7.616475e-05, 0.0003628157, 0.0002028658, 1.915132e-05,
  3.580643e-08, 3.669886e-07, 6.591888e-05, 8.868174e-05, 3.688661e-05, 
    3.386822e-05, 0.0001625921, 0.0002078227, 0.0001048332, 6.29573e-06, 
    2.323571e-05, 0.0003163985, 0.0002350626, 0.0001213967, 2.255886e-08,
  1.846697e-08, 1.001311e-08, 1.152981e-07, 7.26045e-05, 5.584794e-05, 
    2.00276e-05, 5.110351e-05, 0.0001701202, 0.0001427211, 2.455724e-05, 
    0.0002878554, 0.0005806814, 0.0002837959, 8.504705e-05, 2.574381e-08,
  7.654298e-09, 1.398325e-08, 4.102541e-08, 1.769358e-06, 5.728492e-05, 
    3.206268e-05, 2.007305e-05, 0.0001367114, 0.0001824866, 0.000147745, 
    0.000499394, 0.000446636, 0.000143004, 8.030416e-07, 6.468093e-08,
  1.382147e-09, 5.743116e-09, 9.547918e-09, 6.907461e-08, 5.584449e-06, 
    3.145892e-05, 1.945945e-05, 5.943596e-05, 0.0001617428, 0.0003595983, 
    0.0004723874, 0.000540514, 0.0001265118, 1.526066e-05, 3.945225e-07,
  6.677058e-10, 2.746686e-09, 1.85765e-09, 1.226516e-08, 1.239726e-07, 
    7.85621e-06, 1.649705e-05, 8.719278e-06, 8.144495e-05, 0.0004239874, 
    0.0007354849, 0.0007786416, 0.0002740883, 1.060038e-06, 7.486305e-07,
  5.824246e-10, 1.351958e-09, 1.527529e-08, 4.889171e-09, 9.333284e-08, 
    1.903782e-07, 4.198618e-06, 4.297555e-06, 8.318331e-06, 0.0002177783, 
    0.0007364444, 0.0007870293, 0.0003837607, 5.682141e-05, 8.626221e-06,
  9.908386e-10, 7.687794e-10, 1.502578e-09, 1.737943e-08, 4.563816e-08, 
    6.042252e-08, 5.112047e-07, 2.87833e-06, 7.041858e-06, 3.927457e-05, 
    0.0004911725, 0.0007774047, 0.0005843409, 0.0002109931, 3.630922e-05,
  5.892955e-10, 1.440993e-09, 1.25591e-09, 1.902815e-08, 4.401056e-08, 
    8.22065e-08, 4.056678e-07, 7.49875e-06, 6.393004e-06, 2.916417e-05, 
    0.0001591371, 0.0006219347, 0.000649745, 0.0002513303, 6.572418e-05,
  3.650274e-11, 3.72936e-10, 2.568958e-10, 2.298372e-10, 1.460742e-08, 
    2.006587e-08, 6.326754e-09, 1.55661e-07, 1.57725e-06, 1.293255e-05, 
    5.674453e-05, 0.0004239165, 0.0006252464, 0.0004179128, 6.421607e-05,
  5.71004e-12, 3.287975e-13, 1.888376e-13, 2.227459e-12, 6.258455e-09, 
    1.621607e-08, 9.034553e-09, 1.4035e-08, 1.583353e-06, 9.313453e-06, 
    3.841036e-05, 0.0001831259, 0.0005810864, 0.0005072494, 0.0001896442,
  2.156718e-09, 3.915025e-09, 1.025016e-08, 4.332081e-08, 1.37545e-06, 
    2.344982e-05, 5.909875e-05, 3.538029e-05, 1.069436e-05, 4.070872e-06, 
    3.860702e-06, 9.611459e-05, 0.0004924693, 0.0001187076, 1.318829e-07,
  3.291925e-09, 1.959975e-09, 2.242778e-09, 4.831093e-09, 1.167681e-07, 
    7.027907e-06, 7.018761e-05, 6.778727e-05, 3.802113e-05, 8.623848e-06, 
    3.082308e-05, 0.0001203456, 0.0003675522, 0.0001413861, 3.525073e-07,
  1.171056e-08, 6.283786e-09, 1.321802e-09, 1.354917e-08, 2.365859e-09, 
    7.446719e-07, 4.80013e-05, 0.0001085329, 0.0001087122, 9.764848e-05, 
    0.0001016952, 0.0001562915, 0.0001883094, 6.796744e-05, 5.978177e-07,
  1.036951e-08, 1.963661e-08, 3.459741e-09, 2.111431e-08, 7.059626e-09, 
    9.335624e-08, 3.279434e-06, 7.89718e-05, 0.0001577455, 0.0001986502, 
    0.000307062, 0.0003581588, 0.0001432296, 3.428312e-05, 5.97825e-07,
  1.146532e-08, 1.533568e-08, 1.831024e-08, 7.31593e-10, 2.026941e-08, 
    9.819915e-08, 4.125567e-07, 1.28695e-05, 0.0001187441, 0.0003035211, 
    0.0004808715, 0.0002545813, 0.0002310496, 3.352654e-05, 6.152459e-07,
  4.848912e-09, 1.118793e-08, 1.012434e-08, 1.895289e-09, 3.099842e-09, 
    5.978992e-09, 1.276891e-07, 1.48375e-06, 4.016409e-05, 0.0002166129, 
    0.0004332819, 0.0003485592, 8.39952e-05, 3.338055e-05, 1.210489e-06,
  2.901755e-09, 9.132384e-09, 5.387196e-09, 2.475423e-09, 2.422851e-09, 
    7.307345e-09, 2.961457e-09, 3.586058e-08, 1.393146e-06, 6.048004e-05, 
    0.0003248587, 0.000529161, 0.0003616077, 8.745823e-05, 3.511423e-05,
  3.142836e-09, 5.790012e-09, 4.742585e-09, 2.791086e-09, 9.9901e-10, 
    1.083077e-09, 6.690721e-07, 1.126635e-05, 4.81386e-06, 1.286156e-06, 
    0.0001380362, 0.0004458987, 0.000434097, 0.0001526877, 1.215157e-05,
  2.283443e-09, 3.082507e-09, 4.260394e-09, 3.59818e-09, 2.701022e-09, 
    1.530898e-10, 1.224347e-09, 1.663243e-06, 8.100781e-07, 2.020531e-06, 
    3.193956e-05, 0.0002785224, 0.0003488235, 0.0002009065, 6.909066e-05,
  1.71411e-09, 1.193418e-09, 1.898103e-09, 3.401422e-09, 7.469112e-08, 
    7.307057e-10, 2.622311e-07, 1.742508e-06, 1.874605e-06, 3.482377e-06, 
    9.695234e-06, 0.0001431543, 0.0002330034, 0.0002140466, 0.0001831271,
  5.007285e-10, 8.181102e-10, 5.93046e-09, 7.997485e-09, 1.410221e-07, 
    1.111923e-06, 4.681807e-06, 7.732949e-06, 1.125994e-05, 5.488935e-06, 
    1.786873e-06, 3.039934e-07, 0.0001794084, 0.0001715815, 6.340749e-05,
  9.416978e-10, 3.785917e-09, 3.322974e-09, 2.49296e-10, 9.873801e-10, 
    2.238884e-07, 1.212541e-05, 1.006488e-05, 9.630671e-06, 8.319374e-06, 
    5.113002e-06, 2.357647e-06, 0.0002021047, 0.0001443339, 1.312693e-05,
  1.806294e-08, 8.413244e-07, 1.796114e-06, 2.876686e-10, 8.991467e-11, 
    2.622627e-08, 1.168928e-05, 3.250712e-05, 1.701532e-05, 1.240585e-05, 
    7.708089e-06, 2.731002e-06, 0.0001625703, 0.0001205211, 2.484569e-05,
  5.203676e-07, 5.125057e-06, 1.023932e-06, 3.44156e-10, 2.254163e-10, 
    1.690399e-09, 5.317664e-07, 3.213056e-05, 3.282715e-05, 2.295424e-05, 
    1.334511e-05, 2.336213e-05, 2.055742e-05, 6.612745e-05, 5.738348e-05,
  1.405303e-07, 1.755049e-06, 2.163573e-06, 4.99738e-10, 8.600273e-10, 
    9.093575e-10, 3.228348e-08, 6.404921e-06, 6.164674e-05, 3.286354e-05, 
    5.108617e-05, 5.121567e-05, 4.624892e-05, 4.363547e-05, 3.516912e-05,
  4.943147e-08, 1.202382e-06, 6.419062e-07, 1.341854e-09, 9.696041e-10, 
    4.215609e-09, 2.800452e-08, 1.007147e-06, 6.406813e-05, 0.0001377784, 
    9.38347e-05, 5.013678e-05, 1.154496e-06, 4.039498e-05, 3.180896e-05,
  4.768635e-08, 1.526415e-08, 1.990775e-07, 6.366179e-09, 2.056734e-09, 
    7.981295e-07, 8.107576e-07, 9.318254e-07, 1.545487e-05, 0.0002292543, 
    0.0003135081, 0.0001833571, 4.140463e-05, 2.327933e-05, 2.952298e-05,
  2.330697e-08, 1.280868e-08, 4.379335e-07, 3.711332e-08, 3.859672e-08, 
    2.305886e-06, 1.579399e-05, 3.475411e-05, 1.482525e-05, 0.0001062706, 
    0.0004389893, 0.0005089567, 0.0002089761, 7.255047e-05, 2.844091e-05,
  3.284624e-08, 3.898944e-08, 8.443159e-08, 1.396573e-07, 3.114141e-06, 
    3.763869e-06, 3.829563e-06, 1.172413e-05, 1.042509e-05, 7.101703e-06, 
    0.0001727323, 0.0007413322, 0.0005174826, 0.0001398481, 3.63928e-05,
  2.470353e-08, 2.842346e-08, 4.297483e-08, 1.196756e-07, 4.667783e-06, 
    1.821379e-06, 1.159005e-05, 6.659121e-06, 9.090238e-06, 1.596801e-05, 
    3.76745e-05, 0.0005373252, 0.000752281, 0.0002846084, 6.440345e-05,
  3.423472e-07, 3.867836e-06, 4.563793e-06, 4.709239e-06, 6.2901e-06, 
    7.623743e-06, 3.147212e-06, 5.481992e-07, 1.093527e-06, 1.318562e-06, 
    4.450256e-05, 8.922984e-05, 0.0001687373, 0.0002210373, 0.0001367877,
  2.884839e-08, 7.354921e-07, 2.708334e-06, 2.978637e-06, 4.754789e-06, 
    9.084011e-06, 7.398051e-06, 5.581007e-06, 2.419518e-06, 9.206969e-06, 
    2.157986e-05, 4.299735e-05, 7.285637e-05, 9.223991e-05, 8.963118e-05,
  2.467131e-08, 3.797958e-07, 7.833654e-07, 5.525516e-07, 1.675372e-06, 
    4.979153e-06, 6.979366e-06, 2.729597e-06, 5.765058e-07, 1.547063e-05, 
    2.336116e-05, 1.891916e-05, 4.121776e-05, 6.417591e-05, 5.444077e-05,
  1.775588e-07, 6.134694e-08, 1.371226e-07, 5.727197e-07, 3.260251e-07, 
    1.121085e-06, 2.731866e-06, 3.07077e-06, 2.540075e-06, 1.186525e-05, 
    1.145396e-05, 5.604315e-06, 2.552084e-05, 3.22723e-05, 3.732197e-05,
  2.568139e-07, 6.809846e-08, 1.12988e-06, 3.809789e-07, 9.918426e-08, 
    8.262349e-08, 9.067556e-07, 4.163432e-06, 5.405871e-06, 8.398882e-06, 
    1.352402e-05, 8.188685e-06, 5.659357e-06, 1.022918e-05, 3.673334e-05,
  1.915133e-07, 8.516172e-09, 7.894979e-08, 1.837642e-07, 2.113593e-06, 
    1.207275e-07, 8.590534e-08, 1.106249e-06, 6.454457e-07, 3.855395e-06, 
    1.13304e-05, 1.236262e-05, 4.227404e-06, 2.56796e-06, 1.678341e-05,
  6.980822e-09, 5.497347e-09, 3.343385e-08, 1.483486e-06, 1.036461e-06, 
    9.478975e-07, 5.955272e-07, 1.04569e-06, 2.803904e-07, 1.574074e-06, 
    5.992094e-06, 1.522254e-05, 8.297353e-06, 4.512702e-06, 1.491761e-05,
  9.144144e-09, 5.214536e-09, 9.6582e-09, 8.676465e-07, 5.285139e-07, 
    1.724261e-06, 1.179374e-05, 2.571797e-05, 1.455666e-05, 2.094411e-06, 
    7.962121e-06, 1.214515e-05, 1.061057e-05, 9.636467e-06, 4.916399e-06,
  3.145242e-09, 2.994305e-09, 1.87438e-09, 1.562108e-07, 4.447469e-06, 
    6.073133e-06, 2.365465e-06, 7.06722e-06, 4.064338e-06, 4.182966e-06, 
    6.17682e-06, 9.350078e-06, 9.283453e-06, 9.048601e-06, 7.593648e-06,
  2.652631e-09, 1.059832e-09, 1.786235e-09, 5.211417e-08, 2.693054e-06, 
    1.530392e-06, 9.827508e-06, 8.197905e-06, 2.602069e-06, 3.559242e-06, 
    5.122085e-06, 4.863594e-06, 5.712306e-06, 9.633135e-06, 9.135892e-06,
  1.548521e-05, 3.975169e-05, 0.0007319011, 0.000963346, 0.001008739, 
    0.001008213, 0.0006406887, 0.000240064, 0.0001493706, 0.0001584756, 
    0.0003515292, 0.0008191345, 0.00127173, 0.0008052047, 0.0002434072,
  5.796681e-06, 1.741631e-05, 0.0008895461, 0.001237791, 0.001212559, 
    0.001282405, 0.0008927159, 0.0003043377, 0.0001501521, 0.0001943511, 
    0.0003162097, 0.000675309, 0.001178376, 0.000647128, 0.0001828367,
  2.031282e-05, 1.358118e-05, 0.0002804972, 0.0008393012, 0.0009339248, 
    0.001092762, 0.0009851111, 0.0004891244, 0.0001410718, 0.0001481739, 
    0.0002118607, 0.0004560487, 0.0007577848, 0.0006043865, 0.0002519978,
  7.126492e-06, 2.994248e-05, 1.673198e-05, 0.0002093373, 0.0004842816, 
    0.0007631191, 0.0008920432, 0.0006259494, 0.000198662, 0.0002075113, 
    0.0001669043, 0.0002816476, 0.0004934251, 0.0005722439, 0.000369666,
  1.431977e-06, 1.036474e-05, 8.240936e-06, 5.055959e-05, 0.0001886728, 
    0.0004300356, 0.0006861021, 0.0006284976, 0.0002690204, 0.0002267577, 
    0.0001303878, 0.0001454543, 0.0003374164, 0.0004999845, 0.0005157858,
  5.448693e-06, 4.026619e-06, 1.261239e-06, 3.374958e-06, 7.716818e-05, 
    0.0001682986, 0.0004121411, 0.0004948774, 0.0003195768, 0.000211876, 
    0.0001661191, 0.0001034613, 0.0001246126, 0.0003517538, 0.0004326068,
  1.681683e-08, 2.110139e-08, 4.141695e-08, 2.491547e-07, 4.539401e-06, 
    7.299686e-05, 0.0001698371, 0.0002896198, 0.0003652705, 0.0002654924, 
    0.0002290421, 0.0002241106, 4.423329e-05, 0.0001071773, 0.0002325182,
  3.831784e-08, 1.436945e-08, 2.808234e-08, 1.824929e-07, 2.016591e-07, 
    2.724969e-06, 7.954558e-05, 0.0001946353, 0.0003235867, 0.0003449271, 
    0.0001697107, 0.0001341526, 2.937255e-05, 2.302757e-05, 7.816849e-05,
  2.095538e-08, 1.457393e-08, 1.353463e-08, 1.85092e-08, 2.752337e-06, 
    3.75112e-06, 1.278402e-05, 5.248219e-05, 8.022488e-05, 0.0001664595, 
    0.0001609136, 3.734663e-05, 1.171789e-05, 1.32003e-05, 3.433604e-05,
  2.642895e-08, 1.508634e-08, 1.678153e-08, 1.146615e-08, 1.316299e-06, 
    3.069886e-08, 1.119056e-05, 1.095326e-05, 1.164296e-05, 5.468186e-05, 
    5.569806e-05, 1.377857e-05, 1.157949e-05, 1.31664e-05, 2.646782e-05,
  7.537308e-08, 1.018136e-06, 6.126047e-06, 8.616267e-06, 9.125542e-06, 
    7.807058e-06, 6.263828e-06, 5.792096e-06, 1.135924e-05, 8.844617e-06, 
    3.214526e-06, 3.16367e-05, 0.0002520386, 1.919712e-05, 1.322244e-06,
  1.792464e-09, 1.203471e-06, 1.914898e-05, 4.209666e-05, 4.430646e-05, 
    4.0033e-05, 1.703455e-05, 1.513733e-05, 1.73876e-05, 1.742523e-05, 
    1.342535e-05, 0.0001551445, 0.0003731326, 8.877774e-05, 1.765522e-05,
  2.454907e-06, 2.701355e-06, 4.927218e-06, 8.640124e-05, 0.0001848171, 
    0.000280728, 0.0001791433, 7.231787e-05, 5.676559e-05, 5.869387e-05, 
    8.878417e-05, 0.0001432976, 0.0001548264, 0.0001412996, 4.43091e-05,
  4.000927e-06, 1.36864e-05, 1.122416e-06, 4.088191e-05, 0.00023777, 
    0.0005754241, 0.000534621, 0.0002741076, 0.0001085502, 0.0001167495, 
    0.0001786862, 0.0002631787, 0.0003023329, 0.0002432823, 0.0001106244,
  3.534988e-06, 1.518094e-05, 4.897448e-06, 7.812458e-06, 0.0002393508, 
    0.0006441807, 0.0009161565, 0.0006396519, 0.0002280624, 0.0001575463, 
    0.000283794, 0.0004163438, 0.0004919407, 0.0004903649, 0.0003914781,
  7.783071e-06, 5.880756e-06, 6.351981e-07, 1.816318e-06, 0.0001648405, 
    0.0007630289, 0.001199654, 0.001025049, 0.0006043993, 0.0003443276, 
    0.0004427326, 0.0005829715, 0.000643038, 0.0007313313, 0.0007340939,
  3.190804e-08, 5.749785e-08, 1.213962e-07, 2.723794e-07, 6.343876e-05, 
    0.0008206363, 0.001077027, 0.00136798, 0.00107992, 0.0006308304, 
    0.0005476731, 0.0005556451, 0.0006383632, 0.000810453, 0.0008871215,
  4.201885e-08, 8.405858e-08, 1.52777e-07, 5.339055e-08, 5.242142e-06, 
    0.0006511165, 0.001270869, 0.001668073, 0.001460595, 0.0008354539, 
    0.0005352434, 0.0004472545, 0.0004793148, 0.0006513844, 0.0008097794,
  4.671045e-08, 8.454979e-08, 1.554448e-07, 8.67236e-08, 2.340523e-05, 
    0.0005474665, 0.001252161, 0.001922644, 0.001633733, 0.001005388, 
    0.0005429214, 0.000390649, 0.0004039682, 0.000503476, 0.000655592,
  3.108073e-08, 5.417288e-08, 1.052765e-07, 2.858102e-07, 0.0001019886, 
    0.0006754754, 0.001406481, 0.001964904, 0.001667104, 0.001129504, 
    0.0005905303, 0.0004266085, 0.0004242455, 0.0004345019, 0.0005563018,
  1.837473e-08, 4.669901e-08, 2.220747e-08, 2.187486e-07, 6.231288e-07, 
    4.672315e-07, 6.929688e-08, 1.066391e-07, 1.249157e-06, 1.661299e-06, 
    6.746508e-07, 7.220243e-07, 7.691669e-06, 9.16843e-06, 2.515639e-06,
  2.15066e-08, 2.595494e-08, 5.201971e-09, 1.747879e-09, 2.756905e-08, 
    3.147436e-08, 1.057805e-08, 1.001013e-08, 7.721845e-08, 2.476794e-06, 
    3.407228e-06, 7.315302e-07, 9.1315e-07, 1.149477e-06, 6.048108e-07,
  1.032062e-08, 2.074591e-08, 1.004873e-07, 2.035383e-08, 1.337919e-09, 
    1.195722e-09, 1.197265e-09, 1.156611e-07, 2.410995e-07, 7.020818e-07, 
    3.200953e-06, 2.595404e-06, 8.086826e-07, 1.387125e-07, 3.480717e-07,
  5.952771e-08, 8.406701e-07, 1.052744e-07, 6.292332e-08, 1.95465e-08, 
    7.872051e-10, 7.250168e-10, 1.118239e-07, 9.172284e-08, 1.013374e-06, 
    5.360214e-06, 4.620891e-06, 1.814068e-06, 2.266696e-07, 1.747549e-07,
  5.525736e-08, 9.810321e-07, 8.644097e-07, 7.064358e-08, 1.171358e-07, 
    8.712357e-08, 9.655275e-09, 4.545975e-08, 5.462928e-07, 1.264078e-06, 
    4.322964e-06, 5.542969e-06, 4.80667e-06, 5.59227e-07, 1.907733e-07,
  1.813709e-06, 2.217279e-06, 6.65703e-08, 2.612907e-07, 1.16573e-06, 
    1.336108e-06, 2.547468e-07, 1.805254e-07, 4.573289e-07, 6.012397e-07, 
    3.272309e-06, 5.729513e-06, 1.755342e-06, 1.555786e-06, 3.252771e-07,
  1.898067e-08, 1.679659e-07, 3.633676e-07, 4.190866e-06, 5.020649e-06, 
    5.638503e-06, 9.571299e-07, 1.246472e-07, 3.598479e-07, 5.609646e-07, 
    3.483651e-06, 5.896664e-06, 3.064146e-06, 1.086631e-07, 5.629324e-07,
  6.086732e-09, 2.282508e-08, 7.200164e-07, 3.740064e-06, 7.634933e-07, 
    3.212005e-06, 1.411605e-05, 1.876907e-05, 1.049973e-05, 3.02508e-07, 
    1.586136e-06, 7.039837e-06, 3.025631e-06, 4.536856e-08, 2.029641e-06,
  2.30887e-09, 3.231363e-08, 6.232348e-07, 7.282784e-07, 7.339847e-06, 
    6.381574e-06, 1.133705e-06, 1.951215e-06, 7.247926e-07, 7.893869e-07, 
    4.064188e-06, 4.136593e-06, 2.26782e-06, 1.242803e-07, 5.964584e-06,
  1.430825e-09, 1.181981e-08, 3.125409e-07, 1.159581e-06, 2.610368e-05, 
    4.791436e-05, 6.731833e-05, 2.772879e-05, 2.570735e-05, 1.375919e-05, 
    3.462561e-06, 8.198103e-07, 2.41678e-07, 7.216327e-07, 1.648643e-05,
  1.330166e-06, 4.31866e-06, 3.147234e-06, 4.248357e-06, 2.520317e-05, 
    5.359278e-05, 8.076953e-05, 0.0001321568, 0.0001828865, 0.0001048876, 
    2.476564e-05, 1.692362e-06, 9.197014e-05, 1.264711e-05, 1.281569e-07,
  1.822935e-05, 3.083531e-05, 2.604425e-05, 9.513549e-06, 2.331861e-05, 
    5.844524e-05, 9.916892e-05, 0.0001316254, 0.0002139481, 0.0001296041, 
    2.483129e-05, 4.570355e-05, 5.391433e-05, 9.318913e-07, 4.856683e-07,
  3.983724e-05, 6.382776e-05, 5.322203e-05, 2.785601e-05, 2.326241e-05, 
    7.787585e-05, 0.0001286052, 0.0001356972, 0.0002176668, 0.0001295317, 
    1.883625e-05, 7.872382e-05, 6.038411e-06, 7.015639e-07, 5.389013e-07,
  3.828797e-05, 6.985389e-05, 6.19596e-05, 3.985286e-05, 2.542443e-05, 
    8.691721e-05, 0.0001241484, 0.0001163526, 0.0001828941, 0.0001088407, 
    6.278501e-06, 4.179681e-05, 2.321074e-06, 9.911067e-06, 6.124135e-07,
  1.361242e-05, 3.82107e-05, 6.756846e-05, 5.969448e-05, 5.037841e-05, 
    9.126126e-05, 9.768244e-05, 8.127758e-05, 0.0001387244, 7.914882e-05, 
    4.618242e-06, 1.736773e-06, 4.158493e-06, 2.201237e-06, 5.559577e-07,
  1.070859e-05, 2.359992e-05, 5.22946e-05, 7.733809e-05, 8.296816e-05, 
    0.0001030207, 9.42857e-05, 7.50599e-05, 9.806137e-05, 5.052487e-05, 
    7.566678e-06, 2.034877e-06, 4.591298e-06, 3.050886e-06, 5.418229e-07,
  7.155159e-07, 5.971074e-06, 4.986687e-05, 7.743593e-05, 9.386914e-05, 
    0.0001283388, 9.50027e-05, 0.0001293897, 6.946475e-05, 2.779923e-05, 
    1.508274e-06, 2.633864e-06, 3.796234e-06, 3.408185e-06, 1.359937e-06,
  2.534558e-06, 1.014323e-05, 4.886031e-05, 8.031212e-05, 8.752679e-05, 
    8.431929e-05, 0.0001066161, 0.0001201136, 0.0001254262, 1.193503e-05, 
    1.001778e-06, 1.238194e-06, 3.865723e-06, 3.545659e-06, 1.664638e-06,
  3.624365e-06, 1.05709e-05, 3.62136e-05, 5.604983e-05, 0.0001143022, 
    7.273275e-05, 5.374875e-05, 1.272823e-05, 7.515796e-07, 4.47665e-06, 
    6.561692e-07, 1.353035e-06, 3.294824e-06, 4.593768e-06, 2.175781e-06,
  8.93846e-06, 1.695265e-05, 3.287203e-05, 5.060642e-05, 7.817899e-05, 
    7.294965e-05, 0.0001139409, 4.604911e-05, 6.013251e-06, 3.524784e-06, 
    1.069469e-06, 2.086828e-06, 2.598948e-06, 3.829097e-06, 8.511099e-07,
  3.083802e-11, 6.991818e-11, 1.485156e-10, 1.389881e-09, 4.488867e-07, 
    1.103398e-05, 1.69645e-05, 2.8014e-05, 5.850242e-05, 2.953127e-05, 
    2.264029e-05, 6.207653e-05, 0.000321591, 0.0006299235, 0.000280297,
  9.988682e-10, 3.762484e-11, 1.305937e-10, 1.840677e-08, 1.583075e-06, 
    1.699763e-05, 2.443478e-05, 4.563713e-05, 8.710326e-05, 6.52859e-05, 
    4.229702e-05, 0.0001389934, 0.0002373767, 0.0004784852, 0.0003348251,
  1.476889e-08, 1.411157e-11, 6.947039e-10, 5.305473e-08, 2.541144e-06, 
    1.745167e-05, 3.298518e-05, 7.349026e-05, 0.0001012685, 8.459232e-05, 
    6.820285e-05, 8.281441e-05, 0.0001468095, 0.0003468754, 0.0002360534,
  4.035224e-07, 4.770819e-07, 5.529052e-07, 1.776973e-08, 2.051142e-06, 
    2.287338e-05, 5.59026e-05, 0.0001046447, 0.0001152237, 9.294657e-05, 
    7.264768e-05, 5.628703e-05, 0.0001056822, 0.0002751142, 0.0001804104,
  2.599229e-06, 5.530686e-06, 2.986698e-06, 2.736108e-08, 3.448387e-06, 
    4.107027e-05, 8.91499e-05, 0.0001341799, 0.0001338353, 0.0001095043, 
    7.849615e-05, 5.71551e-05, 0.0001064203, 0.0002269245, 0.0001744738,
  9.99632e-06, 7.678742e-06, 1.346637e-06, 1.36667e-07, 7.203213e-06, 
    7.157791e-05, 0.0001307328, 0.0001594054, 0.000161069, 0.0001349111, 
    8.306518e-05, 5.790558e-05, 0.0001308451, 0.0002094484, 0.0001761344,
  2.185595e-08, 2.668433e-07, 3.289882e-07, 3.178768e-07, 1.199332e-05, 
    0.0001000058, 0.0001640269, 0.0001622987, 0.0001646825, 0.0001535385, 
    7.573528e-05, 5.539577e-05, 0.0001532336, 0.000239173, 0.0001720234,
  1.586726e-07, 2.117888e-07, 7.604838e-08, 3.799945e-07, 1.692062e-05, 
    0.0001322771, 0.0001869592, 0.0001586849, 0.0001762585, 0.0001640597, 
    9.099484e-05, 5.561349e-05, 0.0001593449, 0.0002698178, 0.0001589896,
  2.674237e-07, 4.096595e-07, 2.642382e-07, 2.761912e-07, 2.826595e-05, 
    0.0001512367, 0.0001732184, 0.0001417145, 0.0002222699, 0.0002092015, 
    0.0001169966, 6.90458e-05, 0.0001530309, 0.0002798281, 0.0001289372,
  3.042448e-07, 6.698097e-07, 3.335977e-07, 1.505084e-07, 4.955457e-05, 
    0.0001879168, 0.000212907, 0.0001624134, 0.0002735327, 0.0002133614, 
    0.0001121347, 7.774306e-05, 0.0001433161, 0.0002549427, 7.890662e-05,
  8.449912e-11, 5.636046e-14, 1.725182e-19, 1.094319e-17, 6.033123e-13, 
    3.414703e-10, 1.527428e-07, 1.184238e-06, 2.972345e-06, 5.593443e-06, 
    1.664329e-05, 6.984034e-05, 0.0002423917, 0.0004639893, 0.0003935152,
  1.722322e-09, 1.725322e-09, 1.570386e-10, 8.892121e-20, 2.169489e-13, 
    9.103259e-12, 8.049027e-08, 1.247063e-06, 2.040329e-06, 3.537844e-06, 
    1.611456e-05, 4.964616e-05, 0.0001868267, 0.0006269357, 0.0005708889,
  7.177382e-08, 4.898902e-10, 4.098439e-11, 7.646548e-22, 1.593152e-18, 
    9.037175e-13, 2.60219e-08, 1.268103e-06, 1.837094e-06, 4.002267e-06, 
    1.874108e-05, 6.789865e-05, 0.000216434, 0.0006264425, 0.0006451632,
  3.897777e-06, 1.572847e-09, 2.47861e-11, 2.970138e-13, 7.738553e-18, 
    9.958624e-11, 1.74855e-08, 1.3738e-06, 1.651032e-06, 4.523508e-06, 
    2.953765e-05, 8.853427e-05, 0.000251884, 0.0005745873, 0.0006583141,
  2.489274e-06, 2.543574e-07, 7.06564e-10, 1.299712e-14, 2.098468e-15, 
    5.92123e-11, 1.581082e-08, 8.085744e-07, 2.769356e-06, 4.677947e-06, 
    2.831446e-05, 0.0001028331, 0.0002308654, 0.0005104208, 0.000700474,
  6.695554e-06, 6.593756e-07, 6.540244e-12, 2.392035e-12, 1.9452e-14, 
    4.829142e-10, 2.529187e-08, 2.465566e-06, 3.130756e-06, 4.789766e-06, 
    2.965391e-05, 9.384592e-05, 0.0002187366, 0.0004967579, 0.0007486917,
  2.797161e-07, 2.737186e-09, 2.503453e-09, 9.104823e-10, 1.004272e-08, 
    1.011413e-06, 1.486693e-05, 2.266608e-05, 2.148939e-06, 3.038358e-06, 
    2.294978e-05, 8.571288e-05, 0.0002033224, 0.0004921212, 0.0007371282,
  8.304529e-08, 2.442076e-08, 2.329244e-08, 1.139778e-08, 1.695871e-08, 
    4.181084e-06, 2.259797e-05, 1.128961e-05, 9.603973e-06, 2.39222e-06, 
    2.315228e-05, 9.236348e-05, 0.0002145594, 0.0004557543, 0.0007307368,
  5.106094e-08, 3.621305e-08, 1.598189e-08, 2.975731e-08, 5.745641e-06, 
    7.56364e-06, 3.079761e-07, 4.619973e-07, 1.627758e-06, 2.269141e-06, 
    3.158289e-05, 0.0001109505, 0.0002116651, 0.0004408297, 0.0007114759,
  2.416983e-08, 8.922281e-09, 9.220095e-09, 3.151173e-08, 5.24934e-06, 
    9.479526e-06, 1.493657e-05, 5.959207e-07, 2.366635e-06, 1.559142e-06, 
    2.922159e-05, 0.0001025632, 0.0001811482, 0.0004411984, 0.000673846,
  4.44109e-11, 1.431734e-10, 5.995355e-09, 6.278424e-09, 3.833808e-09, 
    2.646346e-10, 2.334862e-09, 8.621805e-08, 1.799561e-06, 5.272225e-06, 
    4.547309e-06, 8.510209e-06, 0.0001836624, 0.0005553715, 0.0007218131,
  7.818125e-10, 6.066577e-10, 8.136117e-11, 8.014501e-09, 3.969431e-09, 
    1.868145e-10, 6.726014e-10, 5.076257e-08, 1.380287e-06, 1.148268e-05, 
    1.852102e-05, 6.233485e-05, 0.0001829727, 0.0006665651, 0.0007500139,
  3.383343e-07, 2.244532e-09, 2.106614e-09, 1.998951e-08, 3.028003e-09, 
    5.7136e-11, 4.79841e-11, 2.904084e-09, 4.126186e-07, 2.32509e-05, 
    5.818989e-05, 9.846417e-05, 0.0001333173, 0.0005910656, 0.000702015,
  7.380604e-06, 1.591763e-06, 8.451189e-10, 5.278955e-09, 8.092083e-10, 
    9.849472e-10, 1.746031e-10, 6.092997e-10, 8.960505e-08, 1.05804e-05, 
    7.213395e-05, 0.0001373246, 0.0001629315, 0.0004109485, 0.0005224936,
  8.729457e-06, 4.087044e-06, 2.942603e-09, 2.877448e-08, 3.885514e-08, 
    1.326864e-07, 1.537325e-08, 8.685756e-09, 7.433741e-09, 1.912987e-06, 
    3.264551e-05, 0.0001045424, 0.0001656135, 0.0002698415, 0.0003463053,
  1.254095e-05, 8.20608e-06, 4.911756e-09, 2.156057e-07, 2.531723e-06, 
    1.518051e-06, 9.761891e-07, 2.187645e-07, 3.756819e-07, 1.022926e-06, 
    7.469625e-06, 4.475337e-05, 0.0001274862, 0.0001756292, 0.0002376692,
  1.05289e-07, 3.556335e-08, 2.425972e-08, 1.900445e-07, 1.652601e-06, 
    5.693824e-06, 5.524164e-06, 1.73983e-06, 1.812284e-06, 3.214583e-07, 
    2.286842e-06, 1.081773e-05, 7.596514e-05, 0.000141273, 0.0001896662,
  1.274255e-07, 7.478796e-08, 6.102954e-08, 1.124146e-07, 2.477745e-07, 
    2.458029e-06, 2.218212e-05, 1.870138e-05, 3.699245e-06, 3.462492e-07, 
    1.764517e-06, 2.75344e-06, 2.538956e-05, 0.0001121607, 0.0001688765,
  8.77606e-08, 1.616456e-08, 4.419486e-08, 1.765501e-07, 3.386184e-06, 
    1.622024e-06, 1.436004e-06, 1.112329e-06, 3.140555e-07, 6.945054e-07, 
    2.496772e-06, 1.176863e-06, 6.214906e-06, 7.087798e-05, 0.0001367496,
  6.075339e-08, 8.807142e-09, 3.942879e-08, 1.118065e-07, 6.631794e-06, 
    4.616915e-07, 3.698222e-06, 5.981673e-07, 7.372283e-07, 1.336919e-06, 
    3.229175e-07, 1.557173e-06, 5.156136e-06, 5.679559e-05, 0.0001376965,
  2.569472e-07, 1.17667e-06, 9.189966e-08, 5.09926e-07, 8.953083e-06, 
    6.788704e-06, 3.121424e-05, 8.621901e-05, 6.095695e-05, 2.267161e-05, 
    1.099946e-05, 0.000116797, 0.0002698149, 0.0002085239, 0.0001201224,
  6.700908e-08, 7.678163e-07, 1.626381e-06, 2.55405e-07, 1.679683e-06, 
    5.658836e-06, 1.939609e-05, 5.64592e-05, 5.997514e-05, 3.700805e-05, 
    7.120309e-05, 0.0001194973, 0.0003490949, 0.0002823237, 0.0001555231,
  3.41034e-07, 1.606878e-06, 1.554106e-06, 1.437321e-06, 3.813015e-06, 
    1.283684e-05, 2.274205e-05, 3.167041e-05, 8.888826e-05, 8.949299e-05, 
    0.0001104141, 0.0003218687, 0.0003212806, 0.0003701988, 0.0001745144,
  5.128517e-07, 1.575422e-06, 2.788629e-06, 3.901078e-06, 1.465577e-06, 
    1.005263e-05, 3.27843e-05, 0.000164761, 0.0003222605, 0.0003996796, 
    0.0004294944, 0.0007304483, 0.0005065134, 0.0004134516, 0.0002347527,
  5.07185e-08, 8.61207e-07, 4.464264e-06, 5.427209e-06, 2.832795e-06, 
    1.905473e-05, 0.0002812905, 0.0005061267, 0.0004743518, 0.0004986041, 
    0.0007722625, 0.001048808, 0.0005152806, 0.0003709359, 0.0002884831,
  2.840916e-06, 3.800303e-06, 4.16091e-06, 7.138872e-07, 1.652882e-06, 
    0.0001668252, 0.0004975356, 0.0006287108, 0.0005579917, 0.0005457897, 
    0.0008750012, 0.0007723634, 0.0004967852, 0.0002808086, 0.0001914622,
  4.786782e-06, 5.315945e-06, 5.828776e-06, 2.111351e-06, 2.361074e-06, 
    0.0002973053, 0.0005309857, 0.0008077379, 0.0007456542, 0.0006747271, 
    0.0008734482, 0.001062747, 0.0005308227, 0.0002145663, 9.480747e-05,
  1.990746e-06, 2.719254e-06, 2.937431e-06, 1.778089e-06, 8.509765e-06, 
    0.0004378834, 0.0008043825, 0.001046066, 0.0009569051, 0.000683655, 
    0.0007852967, 0.000798782, 0.0004902948, 0.0002131184, 6.88721e-05,
  2.51222e-06, 2.173721e-07, 3.344092e-07, 5.859193e-07, 8.121895e-05, 
    0.0006168312, 0.001129586, 0.001178664, 0.0008259692, 0.0005902519, 
    0.0006519856, 0.0006144784, 0.0003774557, 0.0001864764, 6.649503e-05,
  3.094763e-06, 2.456585e-07, 4.899968e-09, 3.380166e-08, 0.0001386094, 
    0.000574452, 0.001145361, 0.001051651, 0.0005767173, 0.0003511823, 
    0.0003930591, 0.0003674951, 0.0002334878, 0.0001230132, 4.912104e-05,
  7.801367e-06, 9.361751e-06, 2.359806e-06, 9.802346e-06, 6.621321e-05, 
    0.0005703786, 0.0009062419, 0.0006528007, 0.0002691628, 0.0001354177, 
    7.89445e-05, 4.577734e-05, 3.528901e-05, 1.123303e-05, 7.613648e-06,
  4.562851e-06, 1.905652e-06, 3.121901e-06, 4.101463e-06, 4.312965e-05, 
    0.0005071189, 0.001006064, 0.0008354727, 0.0004018848, 0.0001262812, 
    8.074537e-05, 0.0001666185, 4.874509e-05, 1.956928e-05, 1.140778e-05,
  5.4554e-06, 1.238097e-06, 1.723364e-07, 2.497823e-06, 3.762781e-05, 
    0.0003649367, 0.0009750566, 0.0009340002, 0.0004793144, 0.0001374657, 
    0.0005136519, 0.0004032498, 3.332661e-05, 1.680966e-05, 7.696336e-06,
  3.575729e-06, 1.792003e-06, 4.406943e-08, 1.69579e-06, 3.619202e-05, 
    0.0002838562, 0.0008976102, 0.001028302, 0.0006212401, 0.0006055292, 
    0.0007120425, 0.0001969227, 2.167248e-05, 1.22607e-05, 3.516436e-06,
  8.002432e-07, 1.620555e-07, 5.081904e-07, 6.909693e-07, 9.879088e-06, 
    0.0001566928, 0.0007817142, 0.001097723, 0.0007731025, 0.000434233, 
    0.0005796247, 0.0002903042, 2.049203e-05, 1.190162e-05, 4.667292e-06,
  9.763378e-09, 6.122102e-08, 2.443948e-07, 2.082971e-07, 7.485171e-06, 
    3.920445e-05, 0.0006748866, 0.001118466, 0.0008632591, 0.0003877582, 
    0.000446373, 0.0004161411, 5.90562e-05, 1.040023e-05, 3.464314e-06,
  1.632375e-06, 1.244814e-06, 1.058528e-07, 2.466738e-08, 1.108532e-05, 
    3.153097e-05, 0.0005043797, 0.0009745823, 0.0008241732, 0.0003806224, 
    0.0005425251, 0.0005125841, 0.0001272594, 4.128874e-06, 4.305747e-07,
  3.86122e-07, 5.56993e-08, 4.09936e-08, 2.694631e-08, 8.555471e-06, 
    3.695335e-05, 0.0003507832, 0.0008343736, 0.0007805971, 0.0004558442, 
    0.0007114431, 0.0006295019, 0.0001971363, 2.698923e-06, 5.664565e-08,
  2.9394e-06, 4.965195e-06, 5.669673e-06, 5.286566e-06, 7.190672e-05, 
    0.0001499581, 0.0001836745, 0.0005976611, 0.0006053107, 0.0007361129, 
    0.0009127298, 0.0006927015, 0.0001785262, 8.138163e-06, 1.571678e-06,
  1.983007e-06, 2.95287e-06, 4.736985e-06, 8.825432e-06, 0.0002632253, 
    0.0004047564, 0.0004764829, 0.0005049902, 0.00066919, 0.0008826663, 
    0.000991072, 0.0006889356, 0.0001203999, 3.450878e-05, 9.418968e-06,
  3.588092e-08, 3.869531e-07, 9.86454e-09, 3.868445e-08, 1.017655e-06, 
    2.61646e-07, 1.080404e-05, 0.0001835791, 0.0003737773, 0.0003852857, 
    0.0002880599, 0.0002934709, 0.0001166866, 9.834989e-07, 6.872445e-08,
  1.120936e-08, 6.177984e-07, 1.036783e-07, 9.513601e-09, 3.702105e-09, 
    1.633792e-09, 9.066265e-08, 5.510679e-05, 0.0002530669, 0.0003701785, 
    0.0004742357, 0.0004899036, 7.316657e-05, 9.224989e-07, 4.748924e-08,
  1.350964e-08, 2.282069e-08, 2.786259e-08, 2.876255e-09, 2.03423e-09, 
    4.27727e-09, 1.188989e-08, 2.066064e-05, 0.0001106018, 0.0003078987, 
    0.0006400814, 0.0006645446, 4.894087e-06, 1.63734e-06, 1.291421e-07,
  3.023794e-07, 3.133278e-08, 9.245569e-08, 1.079436e-08, 6.840975e-09, 
    2.368726e-09, 6.168995e-09, 1.408381e-05, 6.241467e-05, 0.0001821503, 
    0.0006949032, 0.0007079833, 1.557855e-05, 8.201276e-06, 1.601951e-06,
  5.81784e-07, 5.738451e-08, 5.722801e-08, 6.162287e-09, 7.794331e-09, 
    3.602556e-09, 6.480361e-08, 7.657375e-06, 4.170609e-05, 0.0001361151, 
    0.0006347246, 0.000478601, 2.911552e-05, 1.812632e-05, 7.618915e-06,
  7.491134e-07, 3.470822e-07, 1.018149e-08, 3.506366e-09, 7.331189e-10, 
    4.360141e-09, 7.649319e-07, 2.599838e-05, 6.185419e-05, 0.0001205506, 
    0.000353324, 0.0005528586, 6.921952e-05, 2.663928e-05, 1.129741e-05,
  4.667349e-07, 2.91922e-08, 4.162214e-09, 1.021116e-09, 6.981088e-10, 
    4.419336e-09, 2.057025e-06, 0.0001139674, 0.0001958317, 0.0001891587, 
    0.0002001347, 0.0005442848, 0.0001319396, 3.000985e-05, 1.048863e-05,
  1.888932e-06, 1.168219e-07, 2.402555e-08, 9.955591e-08, 7.262449e-09, 
    1.079556e-08, 7.046951e-06, 0.0003488597, 0.0005084376, 0.0004200143, 
    0.0002692321, 0.0007928311, 0.0002513894, 3.823239e-05, 6.58108e-06,
  2.230103e-06, 2.101104e-06, 3.684027e-06, 1.488684e-06, 6.894156e-07, 
    8.600101e-08, 9.614135e-06, 0.0003779954, 0.0007409601, 0.0007049734, 
    0.0003966241, 0.0005764521, 0.0003272869, 5.469656e-05, 3.827826e-06,
  1.081416e-05, 4.748793e-06, 3.865623e-06, 4.11788e-06, 4.301452e-06, 
    9.079677e-08, 4.52665e-06, 0.0002746522, 0.0008109937, 0.0008429969, 
    0.0005059351, 0.0006000101, 0.0003155982, 9.011108e-05, 5.304998e-06,
  1.860961e-06, 6.157171e-07, 7.492508e-07, 1.971407e-07, 7.940954e-07, 
    7.239623e-06, 0.0003901315, 0.000681916, 0.0006707409, 0.0005162296, 
    0.0003987511, 0.0002584592, 0.0001311396, 8.721136e-05, 4.769588e-05,
  3.744666e-07, 3.447932e-09, 2.975231e-08, 3.045459e-07, 2.183791e-07, 
    1.065086e-06, 8.342387e-05, 0.0006003706, 0.0007519263, 0.0006922896, 
    0.0006921751, 0.0005268924, 0.0002260659, 0.0001105012, 6.816353e-05,
  1.642498e-07, 3.708589e-08, 1.136783e-07, 8.106101e-08, 8.998509e-08, 
    1.774384e-07, 4.739148e-05, 0.0003778076, 0.0007693826, 0.0008688831, 
    0.0009743535, 0.0008466018, 0.0003592815, 0.0001316989, 7.796613e-05,
  3.303659e-06, 4.408678e-06, 5.478751e-07, 4.148905e-08, 2.704014e-08, 
    1.278693e-06, 6.759585e-05, 0.0002481304, 0.0007444557, 0.0009679768, 
    0.001166293, 0.0009524496, 0.0004040213, 0.000155749, 7.300865e-05,
  6.844588e-06, 1.037067e-05, 3.212931e-06, 1.591752e-07, 2.584717e-08, 
    4.088834e-06, 0.0001489806, 0.0003125913, 0.0006996836, 0.0009373972, 
    0.001191829, 0.0009110051, 0.0003944271, 0.0001711078, 8.242043e-05,
  2.321172e-05, 1.997764e-05, 1.882801e-06, 2.822709e-07, 2.919098e-08, 
    7.182015e-06, 0.0002594275, 0.00047473, 0.000680368, 0.0009255043, 
    0.001099608, 0.0008198068, 0.0003823022, 0.000186122, 9.096123e-05,
  7.966424e-06, 8.164442e-06, 3.770781e-06, 5.757724e-07, 1.315679e-08, 
    3.91773e-05, 0.0002957748, 0.0005620308, 0.000708374, 0.0008844336, 
    0.001004099, 0.0007356416, 0.0003962825, 0.0001856231, 8.317026e-05,
  8.403423e-06, 8.760572e-06, 5.710753e-06, 6.968127e-07, 2.021726e-07, 
    4.405646e-05, 0.000262272, 0.0006086021, 0.0008001444, 0.00090405, 
    0.001002523, 0.0007821873, 0.0004092458, 0.0001747153, 5.784687e-05,
  8.487028e-06, 1.030016e-05, 7.805334e-06, 1.607724e-06, 1.995984e-07, 
    3.437444e-06, 0.0001615812, 0.0004938444, 0.0006679885, 0.0008375474, 
    0.0009576931, 0.0007321861, 0.0004381494, 0.0001303895, 4.916806e-05,
  9.52561e-06, 1.150278e-05, 9.399503e-06, 5.15824e-06, 6.742815e-07, 
    4.195406e-07, 4.941147e-05, 0.0002953916, 0.0005078238, 0.0006135538, 
    0.0007393558, 0.0005721514, 0.0004413216, 0.0001294599, 4.763426e-05,
  3.84211e-06, 3.525644e-06, 9.799277e-06, 8.559986e-07, 1.151216e-06, 
    1.195154e-07, 4.902258e-09, 7.773617e-08, 3.31113e-07, 1.735304e-06, 
    2.183708e-06, 5.88571e-06, 4.671287e-06, 5.321891e-05, 0.0001365521,
  9.694644e-06, 1.660766e-05, 4.899562e-06, 1.402705e-06, 3.491621e-07, 
    3.811594e-07, 2.159643e-08, 3.065063e-07, 1.20454e-06, 2.142933e-06, 
    3.357411e-06, 5.505085e-06, 4.746888e-06, 1.955784e-06, 9.9971e-05,
  6.341448e-05, 4.321326e-05, 4.425633e-06, 7.719406e-07, 7.217246e-07, 
    7.560727e-08, 2.776503e-07, 5.280028e-08, 3.118758e-07, 1.236248e-06, 
    6.237647e-06, 6.768017e-06, 3.859206e-06, 2.789285e-06, 0.0001190096,
  1.309077e-05, 1.577442e-05, 1.308535e-07, 5.908181e-08, 4.981727e-07, 
    7.630184e-07, 7.218751e-08, 2.353212e-07, 1.408437e-06, 2.110605e-06, 
    7.39022e-06, 8.268566e-06, 4.056375e-06, 2.507974e-05, 0.0001022913,
  4.139335e-06, 4.17351e-06, 2.786546e-06, 6.221478e-07, 1.013522e-06, 
    1.168434e-06, 6.442056e-07, 1.526477e-06, 7.803273e-07, 2.611562e-06, 
    5.714626e-06, 9.330493e-06, 3.759242e-06, 5.72117e-07, 3.966147e-05,
  3.048042e-05, 2.127935e-05, 2.480134e-06, 2.97779e-06, 2.937714e-06, 
    2.801632e-07, 2.589889e-06, 2.506888e-06, 1.19212e-06, 9.957881e-07, 
    6.070572e-06, 9.170722e-06, 3.802702e-06, 1.073655e-06, 5.477453e-06,
  1.365578e-05, 1.258234e-05, 5.566151e-06, 6.974196e-06, 2.351972e-06, 
    5.240538e-06, 1.812941e-05, 1.833472e-05, 8.465195e-06, 3.125152e-06, 
    5.093126e-06, 1.22085e-05, 1.016402e-05, 2.144777e-06, 4.360614e-06,
  7.687952e-06, 8.707048e-06, 7.134492e-06, 9.445862e-06, 4.790315e-08, 
    2.722967e-05, 0.0001120666, 0.000172865, 0.0001139243, 3.315302e-05, 
    3.290575e-05, 4.151118e-05, 1.294125e-05, 2.850144e-06, 4.988029e-06,
  6.082781e-06, 7.025867e-06, 7.238819e-06, 1.072864e-05, 5.271306e-06, 
    3.278996e-05, 0.0001891834, 0.0003917822, 0.0003636659, 0.00021029, 
    0.0001594452, 0.0001047792, 2.231341e-05, 3.233927e-06, 6.4637e-06,
  3.342157e-06, 3.879823e-06, 7.438204e-06, 1.183951e-05, 5.710109e-06, 
    4.815651e-05, 0.0002459602, 0.0005730285, 0.0006300052, 0.0004768919, 
    0.0003543016, 0.0002252929, 4.44316e-05, 4.119657e-06, 9.301689e-06,
  1.4405e-06, 4.47131e-07, 8.654495e-07, 3.321648e-07, 6.660164e-07, 
    6.967277e-08, 2.042136e-05, 6.794366e-05, 0.0001215998, 0.0001272977, 
    0.0002834344, 0.0005718635, 0.0006118233, 0.0001543128, 7.79022e-05,
  7.399988e-06, 1.325787e-07, 5.27245e-07, 1.772257e-07, 7.689763e-07, 
    8.635673e-08, 2.672489e-06, 3.588211e-05, 0.0001104442, 0.0001460006, 
    0.0002866753, 0.0005646267, 0.0004674367, 0.0001261783, 3.39871e-05,
  1.742878e-05, 8.139783e-06, 2.716068e-08, 6.711483e-08, 4.731575e-07, 
    2.519097e-07, 3.010426e-07, 1.763431e-05, 0.0001026632, 0.0001371752, 
    0.0002161164, 0.0004405959, 0.0004625155, 0.0001489009, 0.0001028057,
  1.234711e-05, 7.365632e-06, 7.50089e-07, 3.940926e-09, 2.892889e-09, 
    3.890587e-08, 3.806204e-07, 2.688043e-06, 6.579606e-05, 0.0001216845, 
    0.0001065812, 0.0003046301, 0.0003835009, 0.000154619, 0.0001657951,
  2.288718e-06, 5.183032e-06, 5.556746e-06, 6.259261e-08, 8.879434e-08, 
    4.97762e-09, 9.637122e-08, 2.667904e-07, 3.580185e-05, 9.42662e-05, 
    7.285793e-05, 0.0001275437, 0.0002956461, 0.0002230747, 0.0001039753,
  5.447572e-06, 7.696681e-06, 1.59374e-06, 5.341503e-08, 3.691532e-07, 
    3.062322e-09, 4.072073e-09, 2.332763e-06, 8.588467e-06, 8.305321e-05, 
    6.02934e-05, 6.087571e-05, 0.0002287781, 0.000204313, 0.0001227996,
  1.322801e-06, 1.656765e-06, 1.008859e-07, 2.959099e-07, 8.895093e-08, 
    3.426393e-08, 1.435563e-06, 5.070575e-06, 5.207955e-06, 5.876265e-05, 
    5.042917e-05, 2.683226e-05, 0.0001800233, 0.0001965465, 6.035929e-05,
  2.076156e-07, 3.222852e-07, 9.438952e-08, 7.607636e-07, 3.821809e-09, 
    5.243402e-07, 3.010303e-06, 4.421332e-06, 1.051007e-05, 2.148303e-05, 
    1.458103e-05, 1.184823e-05, 0.000126216, 0.0001671929, 3.675557e-05,
  7.381623e-09, 2.378079e-07, 1.278603e-07, 1.416814e-07, 1.267179e-06, 
    9.983303e-07, 1.435843e-06, 2.369728e-06, 4.357417e-06, 1.330054e-05, 
    1.051543e-05, 5.632329e-06, 7.539292e-05, 0.0001553074, 8.193058e-05,
  3.698844e-09, 1.211119e-08, 2.814558e-07, 5.345499e-07, 1.980556e-06, 
    3.506345e-07, 2.004916e-06, 2.399131e-06, 4.172895e-06, 8.084947e-06, 
    5.984434e-06, 5.020102e-06, 2.279931e-05, 0.0001287046, 8.828455e-05,
  2.709127e-09, 6.65242e-08, 3.218916e-06, 5.682686e-07, 2.9549e-07, 
    0.0001405384, 0.0004216085, 0.000567065, 0.0005125941, 0.0002042845, 
    8.31967e-05, 0.0002191249, 0.0002499911, 7.674241e-05, 2.727254e-06,
  8.752873e-10, 8.139112e-09, 5.767574e-08, 2.895083e-06, 4.903962e-06, 
    4.907382e-05, 0.0004127725, 0.0005482738, 0.0004818949, 0.0002292853, 
    0.0001723326, 0.0003936177, 0.0004388226, 6.017583e-05, 1.109953e-05,
  3.583016e-10, 1.151012e-08, 9.738485e-08, 1.107133e-06, 6.895106e-06, 
    2.362008e-05, 0.0002789519, 0.0004904102, 0.0004692202, 0.0002426196, 
    0.0002312479, 0.000448311, 0.0007004698, 4.150546e-05, 1.636751e-05,
  1.565638e-10, 1.075097e-08, 6.59862e-08, 8.738331e-08, 3.968707e-06, 
    1.454123e-05, 0.0001402381, 0.0003831584, 0.0003942759, 0.0003033964, 
    0.0003180365, 0.0004908683, 0.0003601998, 9.880619e-05, 3.568719e-07,
  4.066545e-10, 1.514319e-08, 1.013656e-07, 1.929213e-07, 2.97099e-07, 
    1.127978e-05, 0.0001006649, 0.0002801247, 0.0003688191, 0.0003454594, 
    0.0004147058, 0.0005439525, 0.0005276008, 9.784893e-05, 5.852619e-07,
  3.675057e-10, 4.224738e-08, 4.085561e-08, 1.721393e-07, 1.742881e-07, 
    1.55494e-05, 0.0001002882, 0.0002321614, 0.0003488945, 0.0004014226, 
    0.0005636104, 0.0006459073, 0.0004196381, 4.32534e-05, 4.642445e-05,
  3.021138e-09, 1.098667e-08, 4.177442e-08, 5.078064e-08, 5.54917e-07, 
    4.580371e-05, 8.785279e-05, 0.0001433761, 0.0002886547, 0.0004988768, 
    0.0006834865, 0.0008193626, 0.0005486332, 7.519445e-05, 4.160319e-07,
  1.542892e-10, 8.206311e-09, 1.87151e-08, 1.739692e-08, 1.082839e-07, 
    2.596718e-05, 0.0001024433, 0.0003026795, 0.0004501191, 0.0006341549, 
    0.0008409085, 0.0007935349, 0.000687302, 0.0001519394, 5.581746e-07,
  1.887875e-11, 8.795211e-10, 8.522629e-09, 4.393286e-07, 8.270029e-06, 
    2.594988e-05, 6.426396e-05, 0.0003146003, 0.0005397702, 0.0007433151, 
    0.0007561857, 0.0005660205, 0.0005578176, 0.0001551242, 7.639202e-07,
  1.120444e-12, 2.431869e-10, 5.906378e-09, 1.031211e-08, 1.768187e-06, 
    6.897024e-06, 9.311763e-05, 0.0003459326, 0.000642177, 0.000821719, 
    0.0006493821, 0.0003328264, 0.0003320822, 0.0001407783, 2.01096e-06,
  3.170864e-09, 7.85446e-09, 7.922883e-09, 5.95179e-08, 4.500031e-07, 
    8.806926e-06, 9.81636e-05, 0.0002308818, 0.0003602551, 0.0003133604, 
    0.0001757172, 0.0002309255, 0.0001752569, 4.253913e-05, 2.850518e-05,
  4.800233e-09, 3.268056e-06, 2.216528e-08, 1.403178e-06, 6.008377e-07, 
    2.910372e-06, 0.0001485105, 0.0003548963, 0.0004916649, 0.000404846, 
    0.0002636318, 0.0002089117, 0.0002806845, 2.567559e-05, 1.774041e-05,
  9.147777e-06, 1.627175e-05, 2.083956e-06, 1.688035e-06, 6.376914e-07, 
    1.379843e-06, 9.418547e-05, 0.0004466088, 0.0005995722, 0.000527462, 
    0.0003721847, 0.0002229519, 0.000244094, 4.996627e-05, 1.615893e-05,
  2.988216e-06, 1.705786e-05, 4.349915e-06, 3.221153e-08, 1.324984e-06, 
    1.124901e-06, 5.410108e-05, 0.0005054686, 0.000730027, 0.0005900169, 
    0.000308898, 0.0001588174, 5.404827e-05, 3.503876e-05, 5.929204e-06,
  7.158973e-07, 1.395023e-05, 1.627254e-05, 6.49711e-08, 9.695713e-08, 
    1.418311e-06, 6.913838e-05, 0.0004809685, 0.0008323191, 0.0006686923, 
    0.000324317, 0.0001540098, 0.0002668788, 5.303449e-05, 4.630454e-06,
  2.116592e-06, 6.607412e-06, 2.262268e-06, 6.365467e-07, 4.903892e-08, 
    5.115691e-06, 0.000118789, 0.000530549, 0.0009065844, 0.0007010501, 
    0.0002365789, 0.0002776474, 0.0001388893, 9.531048e-06, 7.026044e-06,
  2.060181e-08, 3.875642e-08, 1.567983e-07, 1.346138e-08, 1.792118e-06, 
    1.415303e-05, 0.0001136552, 0.0005375891, 0.0009245005, 0.0006877441, 
    0.0002412865, 0.0001228916, 0.0001223305, 6.722164e-06, 1.712988e-06,
  2.435278e-09, 1.556642e-08, 3.766078e-08, 2.981241e-08, 3.85007e-06, 
    3.119908e-05, 0.0001681029, 0.0005601537, 0.0008486896, 0.0006030036, 
    0.0001876864, 0.0002431591, 0.000167799, 4.041101e-06, 7.014774e-07,
  1.006573e-09, 5.801996e-09, 9.811679e-09, 5.327568e-08, 2.875707e-05, 
    6.152835e-05, 0.0001318116, 0.0004688935, 0.0006220378, 0.000493972, 
    0.0003602577, 0.0002245867, 9.067732e-05, 1.928859e-06, 9.473501e-07,
  7.825386e-10, 4.574805e-09, 4.730702e-07, 1.402235e-06, 8.52354e-05, 
    0.0001346235, 0.0002492123, 0.0004904463, 0.0007149332, 0.000444099, 
    0.000395225, 0.0002158541, 7.64484e-06, 4.558138e-06, 9.780998e-07,
  3.571094e-07, 6.700304e-07, 2.685432e-06, 5.961329e-06, 5.465361e-06, 
    4.691954e-06, 6.061615e-06, 7.13147e-06, 5.329869e-06, 5.842029e-06, 
    1.518469e-05, 7.079569e-05, 0.0001181821, 5.794067e-05, 2.730543e-05,
  9.438757e-08, 2.484826e-07, 3.036132e-07, 2.245016e-06, 4.313674e-06, 
    4.460234e-06, 6.044522e-06, 4.900021e-06, 9.138299e-07, 1.825878e-05, 
    3.30583e-05, 6.047495e-05, 0.000111153, 6.249342e-05, 7.369822e-05,
  1.277993e-07, 1.649233e-06, 6.556444e-08, 3.490003e-07, 1.661485e-06, 
    2.198074e-06, 4.756446e-06, 5.357681e-06, 1.360521e-06, 6.42142e-05, 
    0.0001125388, 8.539532e-05, 0.0001293989, 0.0001664752, 0.0001373814,
  3.341135e-08, 2.060025e-06, 1.011963e-07, 2.285355e-07, 4.979688e-09, 
    3.051171e-07, 2.852369e-06, 2.469153e-05, 4.224671e-05, 9.0211e-05, 
    0.0001187979, 0.0001127305, 0.0001282803, 0.0001120417, 4.39109e-05,
  9.561562e-08, 2.618184e-06, 2.343859e-06, 7.338163e-09, 5.344629e-09, 
    2.464017e-08, 3.1678e-06, 2.059778e-05, 8.407065e-05, 0.0001559175, 
    0.0001384095, 0.0001346583, 0.0001530078, 6.530514e-05, 3.460671e-05,
  2.380441e-06, 4.849217e-06, 1.924358e-07, 2.399571e-08, 4.259367e-08, 
    2.073336e-07, 5.966249e-06, 3.452385e-05, 0.0001375995, 0.0002370212, 
    0.0001624384, 0.0001210297, 8.380417e-05, 6.171389e-05, 2.894594e-05,
  1.927339e-08, 3.441845e-08, 1.389913e-08, 6.309302e-08, 9.446267e-07, 
    1.948696e-05, 3.692684e-05, 6.489461e-05, 0.0001256228, 0.0001237065, 
    0.0001183096, 9.69556e-05, 8.539706e-05, 4.266746e-05, 1.840798e-05,
  4.689074e-09, 3.787929e-08, 4.368762e-09, 2.295431e-08, 2.616124e-06, 
    2.018204e-05, 6.675719e-05, 0.0001560984, 0.0002027989, 0.0001128532, 
    0.0001116005, 0.0001717792, 0.0001653547, 3.367188e-05, 8.574013e-06,
  5.292704e-09, 6.97014e-09, 1.839245e-08, 1.251959e-07, 1.101087e-05, 
    3.202995e-05, 9.356839e-05, 9.405211e-05, 0.0001412226, 0.0001588566, 
    0.0001493374, 0.0001589946, 0.0002591082, 6.18675e-05, 4.081043e-06,
  4.056295e-08, 6.288258e-08, 8.70157e-07, 6.360982e-08, 1.262147e-05, 
    3.775469e-05, 0.0001918089, 0.000216635, 0.0002806311, 0.0002767493, 
    0.0002415279, 0.0002691524, 9.743108e-05, 1.177639e-05, 1.787964e-06,
  0.0003891907, 0.0003903742, 0.0003108858, 0.0001962179, 0.0001775297, 
    0.0002192583, 0.0002451586, 0.0002169196, 0.000128755, 6.454039e-05, 
    3.17954e-05, 5.304008e-05, 0.0001063308, 1.739054e-05, 2.664748e-07,
  0.0003542315, 0.0003508814, 0.0003185036, 0.0002320991, 0.0001841745, 
    0.0001978113, 0.000204927, 0.0001942822, 0.0001486842, 8.143501e-05, 
    4.578758e-05, 0.0001343022, 9.988554e-05, 1.722515e-06, 3.41716e-05,
  0.0003323296, 0.0003532185, 0.0003080121, 0.0002823242, 0.0002102157, 
    0.000178054, 0.0001721333, 0.0001697278, 0.0001655301, 0.0001306088, 
    0.000112418, 0.0001130611, 8.669548e-05, 7.144807e-05, 2.917926e-05,
  0.0003449661, 0.000335737, 0.0002501455, 0.0002525074, 0.0002008696, 
    0.0001825299, 0.0001676055, 0.0001681531, 0.0001576483, 0.0001676302, 
    0.0001581513, 8.8669e-05, 6.816487e-05, 3.959533e-05, 1.155421e-05,
  0.0002876105, 0.0002725002, 0.0002576846, 0.0002100924, 0.0002024154, 
    0.0002154747, 0.0002020636, 0.0001671342, 0.0002084586, 0.0001709557, 
    0.000117816, 0.000109283, 8.976016e-05, 3.667617e-05, 1.710023e-05,
  0.0002516763, 0.0002174457, 0.0001913531, 0.0002167197, 0.0002145962, 
    0.0003245046, 0.0002632442, 0.000197174, 0.000154109, 0.0002197299, 
    0.0001400572, 0.000194052, 2.071327e-05, 2.238907e-05, 2.637673e-05,
  0.0001609151, 0.0001625886, 0.0001971532, 0.0002253927, 0.0001723108, 
    0.000357631, 0.0003746464, 0.0003150576, 0.0001812679, 0.0001262465, 
    0.0001550829, 8.94236e-05, 4.716512e-05, 2.132885e-05, 1.475017e-05,
  0.0001759913, 0.0002104247, 0.0002103013, 0.0002111292, 0.0001307301, 
    0.0001564364, 0.0002495983, 0.0002963227, 0.000318387, 0.0001113364, 
    3.888088e-05, 5.52198e-05, 4.305392e-05, 3.507396e-05, 1.315147e-05,
  0.0001735523, 0.0002251377, 0.0002198277, 0.0001200886, 0.0002273113, 
    0.0001444122, 0.0001138384, 3.521171e-05, 9.15718e-05, 0.0001411995, 
    8.081019e-05, 5.684812e-05, 5.797297e-05, 4.948799e-05, 7.150311e-06,
  0.0001810728, 0.0002222716, 0.0002221057, 0.0001095993, 0.0001284909, 
    8.294126e-05, 0.0002000046, 0.0001044316, 0.0002187223, 0.0002025683, 
    0.0001089107, 8.731281e-05, 0.0001049821, 1.692928e-05, 1.612495e-06,
  1.912482e-06, 1.040869e-06, 6.200187e-07, 3.916351e-06, 5.090026e-06, 
    0.0001987148, 0.0002877579, 0.0006454687, 0.0003755193, 1.766636e-05, 
    6.245534e-06, 1.133381e-05, 9.243799e-06, 1.807971e-05, 1.275459e-05,
  3.96553e-06, 1.472621e-06, 3.339126e-07, 1.363952e-06, 1.574603e-06, 
    0.0001495925, 0.0003348537, 0.0007463333, 0.0004480735, 3.870622e-05, 
    1.193405e-05, 5.45824e-05, 3.470037e-05, 1.465181e-05, 1.023433e-05,
  1.205121e-05, 5.238052e-06, 1.665119e-07, 1.065799e-06, 1.580018e-06, 
    3.107618e-05, 0.0002820263, 0.000374578, 0.0004198246, 0.0001464571, 
    3.18302e-05, 5.831599e-05, 3.173287e-05, 2.814341e-05, 1.614355e-05,
  1.115149e-05, 4.631757e-06, 9.265723e-07, 1.370878e-06, 3.107732e-06, 
    6.443892e-06, 8.963347e-05, 0.0002442132, 0.0004430448, 0.0002017923, 
    0.0001034061, 5.987681e-05, 1.007506e-05, 1.258384e-05, 1.645727e-05,
  8.316827e-06, 2.615622e-06, 9.871939e-07, 3.060959e-07, 4.655374e-06, 
    4.68184e-06, 5.623773e-05, 0.0002026908, 0.0005164426, 0.0001966884, 
    8.578326e-05, 0.0001110043, 2.595108e-05, 1.963733e-05, 2.563436e-08,
  9.474868e-06, 4.557087e-06, 7.368548e-09, 2.274657e-07, 4.861942e-06, 
    8.629424e-06, 6.945586e-05, 0.0002104559, 0.0004187449, 0.0002382386, 
    9.523304e-05, 0.0001250848, 3.382656e-05, 4.843757e-06, 1.135083e-05,
  9.3214e-09, 2.491069e-09, 2.561009e-08, 6.104872e-07, 2.537551e-06, 
    2.554807e-05, 8.768103e-05, 0.0002027396, 0.0002949356, 0.0003057929, 
    0.000104774, 8.823836e-05, 3.552038e-05, 1.560693e-06, 4.709111e-07,
  6.874184e-07, 6.309445e-07, 5.017358e-07, 1.702169e-06, 4.485522e-06, 
    2.356983e-05, 8.049762e-05, 0.0001791578, 0.0001999174, 0.0002339047, 
    9.39961e-05, 0.0001042242, 7.978723e-05, 1.07115e-05, 3.304096e-07,
  8.738769e-06, 9.309164e-06, 5.888787e-06, 1.510355e-06, 4.51368e-05, 
    3.270332e-05, 5.110852e-05, 6.077417e-05, 7.536708e-05, 0.0001932093, 
    0.0002264348, 0.000145952, 8.088555e-05, 2.544766e-05, 6.547818e-07,
  2.556456e-05, 2.367538e-05, 1.481884e-05, 3.178949e-06, 3.318312e-05, 
    5.133961e-05, 0.0001258716, 0.0001328928, 0.0001156894, 0.0001296427, 
    0.0002543663, 0.0001486295, 4.414483e-05, 7.551605e-06, 3.598331e-07,
  1.6316e-08, 5.946337e-08, 1.736694e-06, 6.344313e-05, 0.0003163622, 
    0.0008513401, 0.0007800093, 0.0002275892, 5.336513e-05, 2.883846e-05, 
    8.85603e-07, 8.413277e-06, 1.042964e-07, 1.480178e-06, 2.432397e-06,
  1.341568e-08, 2.553965e-08, 2.837471e-07, 2.968109e-05, 0.0004234336, 
    0.001118431, 0.001224419, 0.0004428879, 3.620307e-05, 4.617394e-05, 
    1.42758e-05, 3.787503e-06, 4.286044e-06, 3.77304e-06, 3.828814e-06,
  6.168735e-08, 1.924711e-08, 5.01902e-08, 3.91907e-06, 0.0004762699, 
    0.001168084, 0.001697055, 0.0007517722, 3.361189e-05, 4.494391e-05, 
    3.249839e-05, 6.045721e-06, 8.089432e-06, 6.660134e-06, 6.87572e-06,
  3.244539e-06, 3.505168e-07, 6.753243e-08, 1.593807e-06, 0.0003141747, 
    0.0009674912, 0.001591785, 0.001032736, 0.0001373278, 0.0001051323, 
    5.318229e-05, 1.02869e-05, 7.941923e-06, 1.499026e-06, 1.269606e-05,
  4.110486e-06, 1.856769e-06, 3.803893e-07, 8.303562e-07, 6.194203e-05, 
    0.0006749824, 0.001112439, 0.001247422, 0.0004502731, 8.926892e-05, 
    5.030525e-05, 1.745272e-05, 9.503403e-06, 8.631403e-06, 6.658508e-06,
  1.206356e-06, 7.316666e-06, 2.335757e-08, 9.615937e-08, 1.382145e-05, 
    0.0002697275, 0.0008267691, 0.001111452, 0.0007569469, 0.0001458978, 
    7.442641e-05, 1.466195e-05, 5.770961e-06, 8.500925e-07, 1.069129e-05,
  5.777578e-09, 6.401375e-08, 5.883684e-08, 9.96209e-08, 1.747724e-06, 
    7.626083e-05, 0.0004369614, 0.0006905378, 0.0008291878, 0.0003204472, 
    5.170049e-05, 3.220476e-05, 1.883409e-05, 7.925633e-06, 1.256984e-05,
  2.868229e-09, 1.438221e-08, 1.494227e-07, 1.616024e-07, 1.930011e-08, 
    8.092761e-06, 0.0001451847, 0.0004364744, 0.0007421249, 0.000453683, 
    0.000103605, 5.217265e-05, 1.716394e-05, 1.260217e-05, 1.91682e-06,
  4.737485e-10, 3.005176e-09, 1.267739e-07, 2.443691e-07, 1.512177e-05, 
    3.646234e-06, 1.732867e-05, 0.0002770453, 0.0005194229, 0.0005667983, 
    0.0001642789, 6.132507e-05, 3.58394e-05, 2.989802e-05, 5.144925e-06,
  1.658382e-07, 6.666449e-09, 1.862613e-08, 3.63489e-07, 2.663453e-05, 
    6.95157e-06, 4.058939e-06, 0.0001147821, 0.0004674913, 0.0005816778, 
    0.0002841655, 4.802471e-05, 1.785376e-05, 1.799735e-05, 3.330398e-08,
  2.239049e-08, 9.65425e-09, 8.572803e-07, 2.563129e-05, 0.0001376935, 
    0.0003155969, 0.0004085506, 0.0001722773, 4.91272e-06, 2.897755e-06, 
    5.418904e-05, 0.0003105897, 0.0003652205, 5.678535e-06, 3.519902e-06,
  3.54439e-08, 9.519207e-07, 1.285982e-07, 5.964505e-06, 0.0001389899, 
    0.0002375899, 0.0003987899, 0.0002517859, 2.618283e-05, 9.436207e-06, 
    8.776849e-05, 0.0004664131, 0.0003156508, 1.260723e-05, 4.149811e-06,
  2.012267e-05, 5.965635e-06, 3.858662e-07, 1.792752e-06, 0.0001404623, 
    0.0001711308, 0.0003155056, 0.0002726961, 6.433798e-05, 1.781267e-05, 
    0.0001448289, 0.0003568385, 0.0001742069, 4.864413e-05, 1.140372e-05,
  1.130403e-05, 1.400861e-05, 2.58882e-08, 1.817165e-06, 0.0001350276, 
    0.0002588489, 0.0002600848, 0.0002589883, 0.0001380602, 7.8028e-05, 
    0.0001643689, 0.0003751238, 0.0002445363, 1.121681e-05, 1.120512e-05,
  3.279122e-06, 1.215437e-05, 2.434328e-06, 5.093791e-07, 5.492852e-05, 
    0.0004600695, 0.0005009493, 0.0003348833, 0.0001813062, 0.0001620801, 
    0.0001341749, 0.0002204381, 0.0001618056, 1.148118e-05, 2.399344e-06,
  7.061504e-06, 9.824682e-06, 1.939296e-06, 5.791531e-07, 6.672097e-06, 
    0.0005922573, 0.0009045849, 0.0006188664, 0.0003380498, 0.000210243, 
    0.0002061712, 0.0001134374, 3.397748e-05, 1.497851e-06, 2.699599e-06,
  6.291988e-06, 3.855085e-06, 1.314849e-06, 7.488258e-07, 8.019788e-06, 
    0.0005667755, 0.001155343, 0.001164909, 0.0006856929, 0.0002074544, 
    5.841773e-05, 0.0001477281, 5.408288e-05, 6.451254e-07, 5.000003e-07,
  5.125117e-06, 2.777122e-06, 1.381456e-06, 1.071056e-06, 5.45133e-07, 
    0.0001732347, 0.001157174, 0.001434979, 0.001060532, 0.0004590214, 
    0.0001256034, 0.0001334446, 4.692471e-05, 1.000335e-05, 1.509734e-08,
  5.785953e-06, 3.906659e-06, 1.717612e-06, 1.181804e-06, 3.899111e-06, 
    6.139487e-05, 0.0008651171, 0.001497318, 0.001038002, 0.0006329985, 
    0.0003223496, 0.0001215748, 4.800221e-05, 2.088189e-05, 2.980902e-08,
  5.174466e-06, 4.067748e-06, 3.483337e-06, 2.246534e-06, 1.62091e-05, 
    2.384791e-05, 0.0006185924, 0.001459313, 0.001413353, 0.000950942, 
    0.0004780167, 0.0001812534, 5.389298e-05, 4.812898e-06, 5.675111e-06,
  7.223008e-09, 1.922246e-09, 6.720886e-09, 2.740888e-08, 1.399052e-06, 
    7.826934e-07, 1.132003e-08, 9.936224e-08, 2.400833e-07, 5.167504e-07, 
    2.209579e-06, 9.002857e-05, 0.0002026291, 0.0001972062, 0.0001201852,
  1.255001e-09, 1.997281e-06, 1.836102e-07, 4.076024e-06, 3.939542e-06, 
    1.505979e-06, 1.249431e-07, 4.183703e-07, 7.999461e-07, 1.047341e-06, 
    7.01654e-07, 5.790932e-05, 0.0001656089, 0.0001802791, 0.0001282497,
  2.471896e-06, 5.443243e-06, 1.129989e-06, 2.144087e-06, 6.747264e-06, 
    5.742742e-06, 2.703649e-06, 2.076057e-06, 1.970353e-06, 2.073853e-06, 
    1.767662e-06, 2.671833e-05, 0.0001572268, 0.0001699546, 0.0001828315,
  4.128395e-06, 7.509395e-06, 9.155975e-07, 1.35624e-06, 2.337639e-06, 
    1.535645e-06, 1.51785e-06, 2.037168e-06, 2.057979e-06, 3.528475e-06, 
    2.447082e-06, 7.505487e-06, 0.0001315633, 0.0001196828, 0.0001060107,
  2.446517e-06, 5.95329e-06, 2.905617e-06, 2.753192e-07, 1.248942e-06, 
    1.045446e-06, 4.478477e-07, 1.789523e-06, 8.562955e-07, 2.276699e-06, 
    3.20261e-06, 1.394662e-06, 8.511783e-05, 8.936894e-05, 0.0001183577,
  2.241276e-05, 1.868875e-05, 2.400149e-06, 6.108247e-06, 8.806861e-06, 
    3.104513e-06, 1.512702e-06, 5.209481e-07, 5.361496e-07, 4.465755e-07, 
    3.120276e-06, 1.699548e-06, 3.472251e-05, 4.953747e-05, 0.0001137451,
  2.654839e-05, 2.990594e-05, 2.049496e-05, 1.552057e-05, 1.539698e-05, 
    6.698401e-06, 4.019654e-07, 8.779122e-08, 6.945717e-08, 3.292274e-07, 
    1.206178e-06, 3.111489e-06, 2.342638e-05, 3.110155e-05, 4.961768e-05,
  2.274401e-05, 2.903258e-05, 2.397704e-05, 2.492019e-05, 5.274363e-06, 
    7.728473e-06, 5.765277e-06, 9.554551e-06, 7.716736e-07, 2.313548e-07, 
    4.79521e-07, 3.986357e-06, 2.31282e-05, 2.867087e-05, 4.696716e-05,
  2.122116e-05, 2.646775e-05, 2.935471e-05, 2.353457e-05, 4.235941e-05, 
    1.932397e-06, 5.876636e-08, 1.073592e-07, 5.601032e-07, 1.999918e-06, 
    3.253915e-06, 8.193697e-06, 1.097872e-05, 2.233144e-05, 3.066891e-05,
  1.757708e-05, 2.129808e-05, 2.464706e-05, 1.903347e-05, 3.375021e-05, 
    5.851709e-06, 2.495396e-06, 3.981315e-08, 1.440042e-07, 2.342728e-06, 
    5.60964e-06, 1.219758e-05, 1.021549e-05, 1.448667e-05, 2.22429e-05,
  6.790033e-10, 8.042869e-09, 8.056317e-07, 6.503645e-07, 6.47799e-06, 
    4.06981e-06, 7.777188e-07, 2.244294e-06, 2.804035e-06, 5.797835e-06, 
    3.690092e-06, 9.711277e-05, 0.0006698889, 0.0005910269, 0.0002547153,
  1.246151e-08, 9.06529e-08, 1.395128e-06, 2.198241e-06, 4.145548e-06, 
    1.466963e-06, 2.347431e-06, 2.004837e-06, 4.136487e-06, 8.590815e-06, 
    7.764842e-06, 4.73056e-05, 0.0006834513, 0.0005686387, 0.0001319015,
  1.786269e-06, 3.532825e-06, 1.563048e-06, 8.143254e-07, 1.269722e-07, 
    1.601365e-06, 1.805149e-06, 4.454443e-06, 2.918159e-06, 7.249389e-06, 
    1.196624e-05, 1.140197e-05, 0.0005931061, 0.0005400151, 0.0001374354,
  1.570737e-05, 1.340515e-05, 1.812918e-06, 2.312639e-06, 7.124061e-07, 
    2.807118e-07, 9.451079e-07, 3.78966e-06, 4.832145e-06, 4.949094e-06, 
    9.979663e-06, 3.004873e-06, 0.0004764929, 0.0005158241, 0.0001008958,
  4.775433e-06, 9.553847e-06, 9.305851e-06, 1.693721e-06, 6.658813e-07, 
    5.848996e-07, 1.046039e-06, 1.534469e-06, 4.232597e-06, 5.35679e-06, 
    4.001499e-06, 1.334674e-06, 0.0003666795, 0.0004614901, 9.026313e-05,
  1.229016e-05, 1.455751e-05, 3.811072e-06, 1.629235e-06, 2.878445e-06, 
    2.099247e-06, 6.574876e-07, 2.846866e-06, 6.397152e-06, 4.814643e-06, 
    5.448189e-06, 1.887357e-06, 0.0002562609, 0.0004249624, 9.255835e-05,
  4.628854e-06, 7.868009e-06, 7.199658e-06, 6.335088e-06, 4.244935e-06, 
    7.791284e-06, 1.27178e-07, 1.322962e-07, 2.65475e-09, 6.521905e-08, 
    3.274283e-07, 3.740669e-06, 0.0001502089, 0.0003439276, 8.397534e-05,
  6.726467e-06, 9.150366e-06, 9.010699e-06, 1.204904e-05, 3.151681e-06, 
    1.403678e-05, 9.875415e-06, 1.265063e-05, 9.319445e-07, 3.384566e-09, 
    2.446077e-08, 3.012771e-08, 4.684143e-05, 0.0002298872, 7.22706e-05,
  9.06235e-06, 1.293508e-05, 9.432237e-06, 2.042893e-05, 2.823107e-05, 
    5.765256e-06, 1.225217e-06, 1.039959e-06, 1.239319e-06, 1.115875e-06, 
    1.671613e-06, 3.027682e-06, 1.044544e-05, 0.0001412165, 6.725732e-05,
  1.291622e-05, 1.16932e-05, 1.213634e-05, 1.853941e-05, 2.847359e-05, 
    1.296747e-05, 8.747625e-06, 2.163494e-06, 2.115938e-06, 2.219729e-06, 
    4.25696e-06, 6.265634e-06, 3.829014e-06, 7.980994e-05, 6.111316e-05 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.2466774, 0.6143242, 0.0668168, 0.2301621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.4924844, 0.2132108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.600569, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1560082, 0,
  1, 1, 0.7132517, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02739768, 0,
  0.6230268, 0.6280472, 0.3043983, 0.08344039, 0, 0.3148882, 0.01188002, 0, 
    0, 0, 0, 0.08803581, 0, 0, 0,
  0, 0, 0, 0, 0.01144353, 0.8597386, 0.8205094, 0.5086318, 0.1258651, 
    0.08909279, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.291879, 0.6933324, 1, 0.9996726, 0.6666086, 0.08008575, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0.611689, 0.7180831, 0.4623523, 0.2838529, 0.02767258, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0.002817577, 0.8915156, 0.5654301, 0.7485356, 0.3018697, 0, 0, 0, 
    0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0.04916316, 0.5638732, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3486554,
  2.316188, 6.745579, 0.5592819, 0.3199724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  147.4583, 171.3604, 6.513342, 0.3383408, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03840884, 0.4204801, 0,
  316.1323, 305.6766, 15.46485, 0.007546596, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1807817, 1.695307, 0,
  309.9182, 276.4409, 123.1236, 0.0108671, 0, 1.460928, 0.05467265, 0, 0, 0, 
    0.009753421, 0.03281464, 0.7768181, 0.4781904, 0,
  365.1592, 241.1036, 8.988194, 1.559117, 0.4356286, 6.775464, 0.2077458, 
    1.032432, 0.002793631, 0.1432027, 0.862155, 4.338077, 0.2366837, 0, 0,
  0, 0, 0, 0, 0.1289662, 151.094, 22.45284, 14.93281, 5.254983, 2.574013, 
    0.002986824, 0.1528066, 0.0002596498, 0, 0,
  0, 0, 0, 0, 13.93511, 217.993, 380.8379, 455.4515, 234.498, 2.407733, 0, 0, 
    0, 0, 0,
  0, 0.0003258124, 0, 0, 414.0298, 282.8423, 143.9435, 10.21257, 0.1187258, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 1.536109, 363.0271, 340.0019, 397.2344, 11.61882, 0, 0, 0, 0, 0, 
    0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
