netcdf \00010101.atmos_daily.tile1.pr {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pr(time, grid_yt, grid_xt) ;
		pr:_FillValue = 1.e+20f ;
		pr:missing_value = 1.e+20f ;
		pr:units = "kg m-2 s-1" ;
		pr:long_name = "Precipitation" ;
		pr:cell_methods = "time: mean" ;
		pr:cell_measures = "area: area" ;
		pr:time_avg_info = "average_T1,average_T2,average_DT" ;
		pr:standard_name = "precipitation_flux" ;
		pr:interp_method = "conserve_order1" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:53:52 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile1.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile1.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0.1986115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9611561, 0.1583273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7949425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7552791, 0.2484612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.9872221, 0.4156101, 0.04560489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.8345782, 0.2958934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.7792858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9990003, 0.3505592, 0.06537855, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.8140894, 0.2409153, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.9453563, 0.02902743, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pr =
  4.713877e-13, 7.623415e-23, 1.094407e-16, 5.411814e-12, 4.371689e-10, 
    4.574633e-08, 8.971883e-08, 5.92099e-07, 7.415822e-07, 8.13993e-07, 
    1.521001e-06, 3.25465e-06, 4.845844e-06, 9.333253e-06, 1.533958e-05,
  1.307887e-11, 2.614716e-12, 4.076838e-09, 1.749993e-09, 6.943567e-10, 
    9.121751e-08, 1.02796e-07, 5.407937e-07, 1.260665e-06, 2.253785e-06, 
    2.570465e-06, 2.20713e-06, 2.518911e-06, 4.927645e-06, 7.92354e-06,
  4.432859e-08, 8.004712e-08, 1.323674e-07, 7.168814e-07, 1.946835e-07, 
    9.554856e-08, 1.00618e-08, 2.925152e-07, 9.07921e-07, 2.149117e-06, 
    3.983875e-06, 4.24042e-06, 3.577846e-06, 4.591651e-06, 5.575831e-06,
  4.380032e-08, 1.446408e-07, 1.040673e-07, 5.737196e-07, 9.73707e-08, 
    5.109993e-08, 6.407722e-08, 1.189671e-07, 4.564454e-07, 9.621059e-07, 
    5.289973e-06, 5.856591e-06, 6.162211e-06, 7.608057e-06, 9.071532e-06,
  1.241064e-09, 7.999288e-08, 9.823052e-08, 3.230392e-07, 3.230251e-07, 
    7.671547e-08, 3.343474e-09, 1.065378e-07, 2.367578e-07, 4.816728e-07, 
    2.265674e-06, 5.460699e-06, 6.235727e-06, 7.727407e-06, 9.210525e-06,
  1.657459e-08, 1.900403e-07, 4.35982e-07, 1.354921e-06, 3.947626e-07, 
    2.073009e-09, 5.655901e-08, 1.109221e-07, 8.968339e-08, 7.198781e-08, 
    2.353743e-07, 9.998564e-07, 2.354925e-06, 4.022495e-06, 3.955327e-06,
  1.682562e-07, 8.702764e-07, 1.510579e-06, 1.515561e-06, 2.066967e-06, 
    3.865159e-08, 2.015108e-09, 7.837757e-08, 1.230101e-08, 1.667335e-08, 
    5.03192e-08, 8.387853e-09, 7.097881e-08, 1.767566e-06, 1.52184e-06,
  3.98545e-08, 1.898403e-07, 1.168277e-06, 5.189688e-07, 1.607883e-06, 
    1.335701e-07, 1.275158e-10, 2.940066e-10, 6.371817e-09, 1.522944e-08, 
    5.204957e-09, 1.905618e-08, 1.561021e-07, 1.319636e-06, 1.919886e-06,
  1.807929e-08, 1.299799e-07, 3.405e-07, 1.905012e-07, 6.470196e-08, 
    5.464742e-07, 4.637246e-08, 4.871953e-08, 1.773214e-09, 1.720455e-08, 
    3.775314e-09, 5.04769e-09, 2.737376e-07, 7.825954e-07, 1.008179e-06,
  2.979097e-08, 6.609277e-07, 2.631709e-06, 1.4838e-06, 1.841989e-07, 
    1.202036e-06, 3.439532e-06, 3.541429e-07, 6.532102e-09, 1.824395e-10, 
    8.173432e-10, 8.511517e-09, 1.439338e-07, 2.016906e-07, 4.059634e-07,
  3.570241e-10, 1.236705e-10, 2.10963e-11, 1.127075e-08, 3.506159e-09, 
    1.265325e-09, 6.905553e-10, 9.069178e-08, 1.289595e-07, 6.288454e-08, 
    5.904377e-08, 1.964804e-08, 1.315653e-08, 5.144306e-08, 2.389312e-07,
  1.146023e-09, 4.570676e-10, 5.751075e-12, 4.657599e-09, 4.279986e-09, 
    1.098509e-09, 1.127733e-09, 3.134024e-09, 2.108004e-08, 3.388571e-08, 
    1.101111e-07, 1.456028e-07, 3.165758e-07, 3.821766e-09, 2.833876e-09,
  1.625789e-11, 5.68487e-12, 2.19784e-11, 2.772807e-09, 7.583093e-09, 
    1.63208e-09, 9.107021e-10, 1.151476e-09, 5.590674e-09, 4.170046e-08, 
    2.743508e-07, 3.130205e-07, 1.978662e-07, 2.706646e-07, 2.719436e-07,
  5.871971e-16, 5.41227e-11, 6.055648e-11, 1.328153e-10, 7.420104e-09, 
    1.756159e-09, 6.623585e-10, 1.206608e-10, 3.059063e-09, 5.977702e-09, 
    3.470887e-08, 3.606064e-07, 6.287792e-07, 5.869474e-07, 5.349424e-07,
  7.984912e-16, 2.807502e-22, 7.874488e-12, 1.868994e-10, 9.391697e-09, 
    1.25603e-09, 6.740541e-10, 1.115987e-10, 6.433406e-12, 1.039018e-09, 
    1.647429e-07, 1.37765e-07, 3.506403e-07, 7.574462e-07, 1.087979e-06,
  5.472269e-13, 1.17755e-13, 8.972099e-10, 1.398424e-08, 7.383153e-09, 
    7.793102e-09, 6.339365e-10, 3.090747e-10, 3.886903e-09, 2.754778e-09, 
    1.368256e-07, 5.076107e-08, 8.574499e-08, 5.828646e-07, 8.817524e-07,
  5.974804e-11, 4.446316e-11, 1.278278e-11, 2.85276e-09, 3.450835e-09, 
    4.2977e-09, 9.202986e-10, 1.678644e-08, 1.891791e-09, 5.890082e-09, 
    1.170619e-07, 3.413478e-07, 1.154285e-07, 1.721844e-07, 3.445025e-07,
  1.075132e-08, 1.238393e-10, 9.971823e-13, 2.614042e-10, 1.412689e-09, 
    3.29384e-08, 1.026952e-08, 1.116053e-07, 8.86098e-08, 1.800053e-07, 
    5.232827e-07, 1.120892e-06, 6.071893e-07, 1.104081e-06, 1.691692e-06,
  1.162949e-09, 3.339387e-08, 9.663285e-10, 1.326929e-10, 2.052626e-11, 
    6.819459e-08, 3.31869e-07, 8.445144e-08, 4.901772e-07, 9.945421e-07, 
    2.292411e-06, 1.838409e-06, 8.561883e-07, 5.055317e-07, 5.504102e-07,
  4.064694e-09, 6.002017e-09, 6.234302e-09, 2.734803e-09, 5.331263e-09, 
    1.786961e-07, 1.619225e-06, 7.09295e-07, 9.283149e-07, 9.218822e-07, 
    1.434678e-06, 1.456668e-06, 1.439723e-06, 9.335477e-07, 8.868772e-07,
  2.539641e-05, 4.757459e-05, 6.702002e-05, 0.0001126005, 0.0001287644, 
    7.914239e-05, 2.558e-05, 2.853044e-05, 5.23497e-05, 8.052649e-05, 
    0.0001016242, 0.0001104305, 0.0001375222, 0.0001348319, 0.00013537,
  3.044356e-05, 3.992164e-05, 5.189187e-05, 7.275015e-05, 9.076096e-05, 
    8.426573e-05, 6.084289e-05, 5.001943e-05, 7.366722e-05, 7.470533e-05, 
    8.895733e-05, 0.0001003459, 0.0001117212, 9.217492e-05, 5.441309e-05,
  0.0001441953, 7.542242e-05, 5.955345e-05, 6.221768e-05, 5.027576e-05, 
    4.61781e-05, 4.668726e-05, 5.828207e-05, 6.419196e-05, 7.744091e-05, 
    9.561895e-05, 9.118026e-05, 6.395178e-05, 2.675633e-05, 2.359483e-06,
  0.0003992957, 0.0003214781, 0.0002422536, 0.0001724118, 8.874897e-05, 
    5.468394e-05, 6.247683e-05, 7.697882e-05, 6.612849e-05, 6.854517e-05, 
    4.864093e-05, 1.763831e-05, 1.970478e-06, 1.456354e-06, 5.244804e-06,
  0.0004184796, 0.0004355258, 0.000411861, 0.0003289353, 0.0002072125, 
    0.0001137792, 9.578376e-05, 7.729134e-05, 4.721465e-05, 1.270113e-05, 
    8.935332e-06, 4.253785e-06, 2.627248e-06, 2.497327e-06, 4.877933e-06,
  0.0002874765, 0.0003734751, 0.0004308898, 0.0003975663, 0.0002835789, 
    0.0001982046, 0.000149481, 0.0001586161, 0.0001253816, 6.343928e-05, 
    4.599896e-05, 1.711311e-05, 6.654757e-06, 3.228206e-06, 5.357712e-06,
  0.0001963908, 0.0002613277, 0.0003636777, 0.0003960597, 0.0003576006, 
    0.0002489375, 0.0002100835, 0.0002139134, 0.0001898182, 0.0001297365, 
    6.581436e-05, 8.905912e-06, 3.230794e-06, 2.739039e-06, 3.212613e-06,
  0.0001046082, 0.0001540267, 0.0001677099, 0.0002807907, 0.0003090369, 
    0.0002817333, 0.0002170489, 0.0001973097, 0.0001799561, 0.0001547716, 
    7.212733e-05, 1.144959e-05, 3.168641e-06, 1.782153e-06, 2.891762e-06,
  4.907107e-05, 7.5509e-05, 7.667409e-05, 7.941778e-05, 0.0001505076, 
    0.0002072558, 0.0002043358, 0.0001662076, 0.0001476071, 9.178101e-05, 
    2.490889e-05, 2.215546e-06, 2.523952e-06, 1.370738e-06, 2.856033e-06,
  4.900648e-06, 3.105502e-05, 6.428511e-05, 8.303252e-05, 0.0001204833, 
    9.594042e-05, 9.543775e-05, 6.759742e-05, 3.232116e-05, 3.643562e-06, 
    8.343094e-07, 1.107333e-06, 2.042937e-06, 1.247999e-06, 1.915924e-06,
  5.047698e-15, 6.380513e-26, 6.208879e-26, 2.918254e-26, 5.843112e-27, 
    8.286024e-28, 5.57467e-28, 3.908885e-17, 1.669465e-15, 2.072365e-10, 
    1.141425e-07, 4.064316e-07, 6.671243e-07, 1.442064e-06, 1.840529e-05,
  3.656328e-26, 3.426695e-26, 2.928347e-26, 2.234321e-26, 9.945387e-27, 
    5.106206e-27, 1.077141e-27, 5.37527e-27, 1.005319e-10, 2.938954e-10, 
    4.652897e-09, 4.613477e-08, 6.143924e-07, 2.231264e-05, 6.071635e-05,
  2.215293e-11, 5.987436e-11, 1.387742e-26, 1.638007e-26, 7.933489e-13, 
    4.413985e-18, 1.164589e-16, 6.344507e-13, 1.119045e-08, 1.738634e-08, 
    2.86074e-06, 2.492582e-05, 6.264885e-05, 9.661885e-05, 0.0001261205,
  1.245951e-07, 1.555979e-10, 1.509649e-11, 2.542474e-11, 3.180536e-12, 
    5.749187e-13, 6.438884e-10, 4.00815e-08, 6.465598e-07, 2.324157e-05, 
    6.785004e-05, 0.0001181368, 0.0001550261, 0.0001579467, 0.000156942,
  2.753739e-06, 1.279047e-06, 6.525629e-08, 1.473413e-07, 1.123998e-07, 
    1.716191e-07, 5.920414e-07, 4.535055e-06, 2.499482e-05, 5.889068e-05, 
    8.205975e-05, 0.0001039999, 0.0001141231, 0.0001346624, 0.0001450661,
  5.619353e-06, 4.861884e-06, 8.227292e-06, 3.525182e-06, 1.974844e-06, 
    8.69375e-07, 1.402711e-05, 1.283477e-05, 2.602149e-05, 8.305239e-05, 
    8.047823e-05, 5.706262e-05, 8.906943e-05, 0.0001207763, 0.0001403614,
  3.044211e-05, 4.055863e-05, 4.575999e-05, 2.180644e-05, 5.132713e-06, 
    3.517275e-06, 8.155036e-06, 8.726262e-06, 4.199798e-05, 3.664225e-05, 
    5.199926e-05, 4.600019e-05, 6.341009e-05, 9.337591e-05, 0.0001207924,
  3.21345e-05, 0.0001118133, 0.0001665859, 0.0001842468, 7.625924e-05, 
    1.884228e-05, 6.091191e-06, 9.93092e-06, 2.185254e-05, 2.073451e-05, 
    9.332911e-05, 8.502694e-05, 7.653567e-05, 7.824299e-05, 9.214861e-05,
  8.881975e-05, 7.009487e-05, 0.0001770817, 0.0002646617, 0.000269789, 
    0.0001408252, 3.116121e-05, 1.260195e-05, 1.744475e-05, 6.69058e-05, 
    0.0001297478, 0.00016912, 0.0001065704, 9.65887e-05, 9.291572e-05,
  0.000102338, 6.398546e-05, 6.250992e-05, 0.0002195563, 0.0003024039, 
    0.0002963752, 0.0002002861, 8.663801e-05, 9.269218e-05, 0.0001340208, 
    0.0001882771, 0.0002182947, 0.0001548552, 9.203207e-05, 7.009213e-05,
  0.000107137, 0.000151098, 0.0001702924, 0.0001581288, 0.0001603369, 
    0.0001461988, 8.495757e-05, 1.158041e-05, 7.569019e-06, 5.519092e-06, 
    1.669142e-06, 1.074165e-07, 2.529464e-08, 2.264507e-09, 4.736162e-09,
  0.0004441065, 0.0001213593, 0.0001510662, 0.000143461, 9.785439e-05, 
    4.407528e-05, 7.072485e-06, 5.534495e-06, 7.248146e-06, 6.846001e-06, 
    1.764414e-06, 4.156354e-07, 8.073365e-08, 3.372913e-08, 6.381357e-08,
  0.0002623056, 0.0004282682, 0.0001900373, 0.000124289, 2.695389e-05, 
    8.383653e-07, 2.996225e-06, 5.914294e-06, 8.394106e-06, 9.486316e-06, 
    3.006921e-06, 1.049082e-06, 4.195156e-07, 1.845025e-07, 5.908971e-07,
  0.0004155431, 0.0002642279, 0.0001170994, 1.04333e-05, 6.440324e-07, 
    5.672823e-07, 4.275495e-07, 2.737218e-06, 6.713739e-06, 8.861014e-06, 
    6.266042e-06, 2.102372e-06, 2.096421e-07, 8.032805e-08, 8.686092e-07,
  0.00018387, 0.0001555353, 1.438497e-07, 9.337053e-07, 8.051682e-07, 
    6.820684e-07, 1.036357e-06, 2.412639e-06, 4.871078e-06, 6.225143e-06, 
    6.561423e-06, 2.421054e-06, 8.891901e-07, 2.704343e-07, 4.934058e-07,
  0.0001041873, 9.072241e-05, 7.948367e-05, 2.615521e-06, 2.454836e-06, 
    1.709172e-06, 1.770291e-06, 2.436009e-06, 3.290734e-06, 5.052899e-06, 
    7.09042e-06, 2.847624e-06, 1.218253e-06, 7.916906e-07, 4.422563e-07,
  9.673143e-05, 9.003704e-05, 7.602293e-05, 6.703628e-05, 1.953482e-06, 
    4.370108e-07, 1.635883e-06, 3.608887e-06, 4.484979e-06, 2.629428e-05, 
    1.481152e-05, 7.753426e-06, 4.63924e-06, 1.739769e-06, 1.015992e-06,
  8.122877e-05, 7.736123e-05, 7.05552e-05, 6.468158e-05, 1.532001e-06, 
    9.979452e-07, 2.238092e-06, 2.339087e-06, 3.916921e-06, 1.723354e-05, 
    2.923249e-05, 3.027776e-05, 9.174702e-06, 6.766596e-06, 4.781999e-06,
  6.454889e-05, 6.379729e-05, 5.358728e-05, 6.335963e-05, 4.864575e-05, 
    1.474643e-06, 2.307318e-06, 3.686614e-06, 5.325368e-06, 4.495645e-05, 
    4.447719e-05, 2.194086e-05, 1.674229e-05, 9.463281e-06, 5.382232e-06,
  4.784251e-05, 6.523104e-05, 6.98478e-05, 6.79665e-05, 6.170182e-05, 
    5.86171e-05, 3.529599e-06, 3.521845e-06, 8.199197e-06, 4.785513e-05, 
    4.83457e-05, 1.786767e-05, 1.017299e-05, 2.504368e-06, 2.844729e-06,
  2.352029e-07, 6.074454e-08, 2.620991e-07, 1.650327e-07, 9.651503e-07, 
    3.67711e-05, 0.0001248283, 0.0002442737, 0.0002799977, 0.0003163933, 
    0.0003645752, 0.0003923468, 0.0003928253, 0.0003624913, 0.0003189644,
  2.256775e-08, 2.610394e-07, 9.151107e-07, 1.220806e-05, 8.199314e-05, 
    0.0002005419, 0.000292006, 0.0003227297, 0.0003369618, 0.0003950212, 
    0.0003893997, 0.0003627372, 0.0002847405, 0.000236858, 0.0002033174,
  7.567883e-07, 9.263693e-06, 6.888723e-05, 0.0001962125, 0.0003183788, 
    0.0003605067, 0.0003784887, 0.0003625451, 0.0003817462, 0.0003662993, 
    0.000313344, 0.0002313837, 0.0002061469, 0.0001897867, 0.000183259,
  4.36981e-05, 0.0001065937, 0.0002166434, 0.0003398526, 0.000353123, 
    0.0003537899, 0.000340941, 0.0003187266, 0.0002953661, 0.0002579766, 
    0.0002297745, 0.0002323448, 0.0002280449, 0.0002316562, 0.0002133332,
  0.0001367538, 0.0002265753, 0.000305076, 0.0003438386, 0.000337591, 
    0.0003026749, 0.0002564576, 0.0002310165, 0.0002326634, 0.0002640735, 
    0.0003286581, 0.0003217189, 0.0002523181, 0.0002150378, 0.00019629,
  0.000220615, 0.0002913846, 0.0003139367, 0.0003051344, 0.000305965, 
    0.0002601387, 0.0002274205, 0.0002771846, 0.0003797432, 0.0004657631, 
    0.0003814271, 0.0002746688, 0.0002232938, 0.000192599, 0.0001499691,
  0.0003577624, 0.0004477784, 0.0004583481, 0.0004783759, 0.0004486654, 
    0.0003963548, 0.0004118278, 0.0004636051, 0.000471047, 0.0003647799, 
    0.0002448562, 0.000196219, 0.0001694191, 0.0001289914, 9.344549e-05,
  0.0004456415, 0.000558276, 0.0006130761, 0.0006538086, 0.0006033861, 
    0.000523834, 0.0004450972, 0.0003543167, 0.0002776854, 0.0002200422, 
    0.0001726428, 0.0001348472, 9.68317e-05, 7.440833e-05, 5.510167e-05,
  0.0003828816, 0.0004541211, 0.0004878961, 0.0005305281, 0.0005265977, 
    0.0004307505, 0.0003089133, 0.0002045851, 0.0001543212, 0.0001207061, 
    9.59e-05, 7.777182e-05, 6.079117e-05, 4.837849e-05, 4.236585e-05,
  0.0003070195, 0.000312847, 0.0002794545, 0.0002405528, 0.0002301759, 
    0.0002414236, 0.0001873033, 0.0001183134, 6.576611e-05, 5.665755e-05, 
    5.124239e-05, 4.762179e-05, 5.039976e-05, 4.2653e-05, 2.026129e-05,
  7.838408e-24, 7.368411e-24, 1.603196e-23, 4.409803e-11, 4.788847e-11, 
    5.335584e-08, 2.765348e-07, 5.514875e-07, 1.127793e-06, 2.29024e-06, 
    2.493209e-06, 2.829639e-06, 6.401796e-06, 6.447221e-06, 4.684512e-06,
  4.449365e-11, 1.212799e-10, 8.172756e-23, 2.73564e-07, 1.071941e-06, 
    4.535555e-09, 8.063486e-08, 1.502607e-07, 3.339292e-07, 7.160232e-07, 
    1.318447e-06, 2.130653e-06, 2.228368e-06, 2.128471e-06, 1.530467e-06,
  4.15815e-08, 4.012496e-09, 6.411904e-11, 1.684565e-07, 7.074998e-06, 
    7.775639e-06, 5.932438e-06, 7.716058e-07, 1.172745e-06, 8.762597e-07, 
    5.298015e-07, 1.246255e-07, 2.529794e-07, 3.172264e-07, 3.840393e-07,
  2.680849e-09, 1.111022e-09, 2.744013e-10, 8.902038e-07, 6.573372e-06, 
    1.139814e-05, 1.556559e-06, 9.142821e-07, 2.418951e-07, 1.433951e-08, 
    7.372007e-09, 4.422443e-09, 4.442388e-08, 2.749301e-07, 1.542891e-06,
  3.0406e-10, 1.211685e-08, 1.431895e-08, 1.827664e-06, 2.694889e-06, 
    1.780139e-06, 4.599949e-07, 1.008647e-07, 5.543004e-08, 2.891769e-08, 
    7.760359e-08, 3.361844e-07, 9.756224e-07, 2.90389e-06, 1.064289e-05,
  7.838797e-11, 1.457951e-08, 1.458438e-06, 1.006054e-06, 1.76834e-06, 
    3.158089e-06, 3.856588e-07, 3.04114e-07, 3.415926e-07, 6.472051e-07, 
    1.203462e-06, 3.215894e-06, 8.237986e-06, 2.134241e-05, 1.819383e-05,
  1.333303e-08, 1.071569e-06, 9.881337e-06, 1.641118e-05, 3.301794e-06, 
    1.381701e-06, 1.567153e-06, 1.292264e-06, 2.698446e-06, 6.331579e-06, 
    1.208439e-05, 1.354266e-05, 9.524391e-06, 1.144542e-05, 1.480334e-05,
  8.633205e-07, 2.130484e-06, 8.036071e-06, 2.138401e-05, 9.039245e-06, 
    7.187576e-06, 7.28233e-06, 8.748051e-06, 1.289314e-05, 1.695998e-05, 
    1.375255e-05, 1.649372e-05, 2.432042e-05, 3.083699e-05, 5.535042e-05,
  1.316394e-06, 3.344114e-06, 2.701285e-06, 3.635504e-06, 5.875099e-06, 
    6.721311e-06, 2.087804e-05, 3.544426e-05, 3.618694e-05, 5.484844e-05, 
    8.864796e-05, 9.934585e-05, 0.0001099368, 0.0001201386, 0.0001753715,
  1.723449e-06, 9.145423e-06, 1.615103e-05, 2.405871e-05, 3.132399e-05, 
    6.072912e-05, 7.392982e-05, 9.018803e-05, 0.0001277901, 0.0001438099, 
    0.0001339047, 0.0001278286, 0.0001470496, 0.000203029, 0.0002571794,
  3.720651e-11, 6.660686e-11, 3.471295e-11, 1.465501e-09, 1.698107e-09, 
    1.729889e-09, 7.260981e-10, 4.438489e-10, 1.162654e-10, 7.1057e-11, 
    6.684913e-11, 1.154398e-10, 2.855021e-08, 1.056989e-07, 1.281511e-07,
  2.520261e-07, 6.838655e-10, 7.395631e-08, 2.131308e-08, 9.590909e-08, 
    2.171828e-07, 9.366111e-08, 7.232626e-08, 1.043341e-07, 4.146522e-09, 
    1.953032e-08, 5.68858e-10, 3.376063e-08, 2.520369e-07, 5.074938e-07,
  3.487186e-07, 6.255815e-07, 1.943273e-07, 3.084938e-07, 3.006223e-07, 
    2.348418e-07, 3.375096e-07, 2.271349e-07, 1.133608e-08, 1.26617e-07, 
    7.04394e-08, 1.628013e-08, 1.763532e-07, 7.136149e-07, 9.553183e-07,
  4.82696e-07, 1.579009e-07, 5.295345e-07, 4.20192e-07, 6.700031e-07, 
    4.76585e-07, 5.516855e-07, 3.964936e-07, 7.171117e-07, 3.62439e-07, 
    3.539156e-07, 3.364512e-07, 3.985085e-07, 5.739722e-07, 5.152064e-07,
  3.683453e-06, 2.215725e-06, 8.467136e-07, 5.185337e-07, 1.223062e-06, 
    1.794157e-06, 2.619053e-06, 2.21477e-06, 2.219949e-06, 1.956163e-06, 
    2.35072e-06, 2.114233e-06, 1.475123e-06, 1.120455e-06, 8.706511e-07,
  9.627109e-06, 5.702768e-06, 5.041968e-06, 2.203766e-06, 1.782597e-06, 
    3.192364e-06, 3.839215e-06, 3.188829e-06, 3.247464e-06, 2.631763e-06, 
    3.293678e-06, 3.137842e-06, 2.18463e-06, 1.568194e-06, 1.406187e-06,
  3.559241e-05, 1.070016e-05, 1.543543e-05, 5.612019e-06, 4.146036e-06, 
    5.232936e-06, 6.40823e-06, 5.479602e-06, 2.711133e-06, 1.857241e-06, 
    2.707148e-06, 3.430765e-07, 2.921395e-07, 1.029439e-08, 2.109702e-08,
  0.0002095094, 7.838065e-05, 3.967243e-05, 4.257387e-05, 1.222295e-05, 
    6.118602e-06, 7.324473e-06, 9.418341e-06, 6.219657e-06, 3.838799e-06, 
    1.389291e-06, 1.959579e-06, 7.747735e-07, 7.100203e-07, 8.215447e-07,
  0.000505517, 0.0002971707, 0.0001356304, 0.0001443533, 0.0001632941, 
    7.84625e-05, 1.654813e-05, 1.083899e-05, 6.613483e-06, 4.89936e-06, 
    5.226352e-06, 9.924463e-06, 1.605955e-05, 1.383582e-05, 9.91559e-06,
  0.0004767881, 0.0003584054, 0.0002225343, 0.0002065023, 0.0002267942, 
    0.0002318939, 0.0001858258, 6.324035e-05, 1.656545e-05, 1.305572e-05, 
    1.996856e-05, 4.229124e-05, 0.0001039652, 0.0001250508, 0.0001053922,
  1.35002e-07, 1.513516e-08, 1.301168e-07, 5.935403e-07, 1.836741e-07, 
    4.528093e-07, 1.272709e-06, 3.069317e-06, 1.899964e-06, 4.170883e-07, 
    4.002443e-07, 3.977897e-07, 2.337747e-06, 2.576227e-06, 3.073192e-06,
  5.496714e-06, 2.72247e-07, 5.26422e-07, 2.349547e-06, 1.733375e-06, 
    4.436211e-07, 2.923438e-06, 3.375705e-06, 9.777176e-07, 3.195163e-07, 
    4.503487e-07, 4.933869e-07, 7.877388e-07, 5.42715e-07, 8.454979e-07,
  1.410514e-05, 9.259647e-06, 1.015241e-06, 6.151598e-06, 5.411571e-06, 
    8.113866e-06, 4.717319e-06, 2.691059e-06, 5.283441e-07, 9.545078e-07, 
    2.199183e-06, 1.052689e-06, 6.022244e-07, 4.318032e-07, 2.648116e-07,
  5.470841e-05, 1.989773e-05, 4.493342e-06, 5.277876e-06, 1.806304e-05, 
    1.182883e-05, 7.47778e-06, 2.070012e-06, 1.134354e-06, 1.913477e-06, 
    2.820925e-06, 2.136552e-06, 8.246948e-07, 4.080348e-07, 2.624154e-07,
  0.0003474164, 0.0002998635, 0.0001715639, 4.690924e-05, 3.170729e-05, 
    4.31041e-05, 3.741547e-05, 1.487128e-05, 4.383044e-06, 2.309325e-06, 
    2.286263e-06, 3.126799e-06, 1.246885e-06, 5.297691e-07, 2.561733e-07,
  0.000421176, 0.0004131921, 0.0003415029, 0.0002745093, 0.0002326936, 
    0.0002088464, 0.0002227202, 0.0001247576, 4.415523e-05, 1.850333e-05, 
    1.220154e-05, 3.547264e-06, 1.783012e-06, 7.143809e-07, 3.257272e-07,
  0.0003734882, 0.0002970023, 0.0002307347, 0.0001866361, 0.0002334837, 
    0.0003813283, 0.0004370821, 0.0003042483, 0.0001430773, 7.04953e-05, 
    5.063905e-05, 2.480853e-05, 5.587786e-06, 5.135721e-07, 1.14428e-06,
  0.0001983083, 0.0002239852, 0.0001035704, 0.0001772117, 0.0002970264, 
    0.0004382181, 0.0004473219, 0.0003207214, 0.0001878743, 0.0001087884, 
    0.0001086532, 8.090435e-05, 2.72332e-05, 5.661658e-06, 5.044788e-06,
  0.000162785, 0.0002680081, 0.0001531168, 0.0001726087, 0.0003422668, 
    0.0003903188, 0.0002773138, 0.0001666308, 0.0001414848, 0.0001168521, 
    5.082862e-05, 5.087271e-05, 3.078956e-05, 1.340258e-05, 6.8694e-06,
  0.0001171359, 0.0002559461, 0.0001584575, 0.0001717176, 0.0002005625, 
    0.0001360706, 6.986167e-05, 6.768807e-05, 4.892269e-05, 4.530527e-05, 
    6.680936e-05, 2.854048e-05, 8.417999e-06, 1.916256e-05, 1.315104e-05,
  4.724467e-09, 3.22687e-09, 2.510181e-09, 2.454878e-08, 4.08251e-06, 
    4.093414e-06, 2.166869e-06, 2.314317e-06, 3.758498e-06, 5.010266e-06, 
    4.650617e-06, 1.910048e-06, 3.232093e-06, 3.659649e-06, 3.312686e-06,
  1.37257e-06, 6.899335e-09, 1.53813e-09, 5.004925e-07, 2.092775e-06, 
    1.732263e-06, 2.233781e-06, 1.817646e-06, 5.041136e-06, 3.89553e-06, 
    8.695804e-07, 1.421519e-06, 1.955286e-06, 3.66097e-06, 4.680964e-06,
  4.980564e-07, 4.923898e-08, 9.536262e-09, 4.794899e-07, 1.601569e-06, 
    4.585143e-06, 4.943117e-06, 8.863553e-06, 1.219163e-05, 1.216228e-05, 
    3.102047e-06, 1.433832e-06, 3.770452e-06, 5.639464e-06, 5.968198e-06,
  4.41519e-06, 2.780871e-06, 2.206468e-07, 1.400936e-06, 4.199634e-06, 
    1.151181e-05, 3.86861e-05, 7.845011e-05, 0.0001075151, 8.818856e-05, 
    4.55245e-05, 1.969475e-05, 1.395319e-05, 2.495141e-05, 1.456064e-05,
  2.4473e-05, 5.342842e-06, 5.749956e-07, 5.455212e-06, 1.55358e-05, 
    5.145146e-05, 0.0001220244, 0.0002311531, 0.0003369656, 0.0003936856, 
    0.0003567916, 0.0002150775, 0.0001149978, 7.139729e-05, 4.800515e-05,
  3.820235e-05, 5.283975e-05, 5.369675e-05, 3.497109e-06, 3.701111e-05, 
    9.344593e-05, 0.0001884256, 0.0003350606, 0.0004957109, 0.0006678503, 
    0.0007607368, 0.00076878, 0.0006362845, 0.0004216575, 0.0002575505,
  2.911532e-05, 5.172926e-05, 5.660718e-05, 6.848327e-05, 3.300365e-07, 
    2.222584e-05, 6.098818e-05, 0.0001435981, 0.0003141912, 0.0005342683, 
    0.0007294655, 0.0008997651, 0.001003827, 0.001009447, 0.0008567642,
  2.077218e-05, 3.192753e-05, 4.485483e-05, 5.888776e-05, 3.535137e-06, 
    2.688907e-08, 1.305729e-06, 1.040962e-05, 3.649146e-05, 0.000118791, 
    0.0002684172, 0.0005060149, 0.0007091085, 0.0007881144, 0.0008206079,
  5.351193e-05, 5.203987e-05, 5.672591e-05, 8.733154e-05, 5.631494e-05, 
    1.174878e-05, 1.049654e-06, 4.0503e-06, 1.287427e-05, 2.274682e-05, 
    2.489199e-05, 7.916659e-05, 0.0002881685, 0.0003948406, 0.0003665549,
  7.580047e-05, 0.0001190849, 0.0001721263, 0.0001998681, 0.0001756729, 
    0.0001249669, 6.006299e-06, 1.450995e-05, 1.553394e-05, 1.587973e-05, 
    1.274819e-05, 1.771263e-05, 7.604181e-05, 0.0001547023, 8.416592e-05,
  7.9091e-12, 3.235947e-12, 1.457314e-24, 1.709623e-10, 4.687164e-08, 
    2.539861e-08, 1.345853e-09, 3.355746e-09, 2.295988e-06, 2.924387e-06, 
    3.852448e-06, 2.831993e-06, 1.647589e-06, 3.05237e-06, 4.13943e-06,
  2.362824e-10, 2.121602e-23, 4.311468e-24, 9.035026e-10, 2.52436e-09, 
    3.90968e-09, 3.536395e-09, 1.188744e-09, 8.344884e-08, 2.73492e-06, 
    5.276547e-06, 2.575369e-06, 6.33942e-07, 1.431583e-06, 5.558965e-06,
  2.068594e-08, 2.16511e-08, 1.07412e-23, 9.03885e-17, 1.947307e-11, 
    5.37953e-10, 1.346594e-09, 1.202642e-10, 2.464708e-08, 9.088662e-07, 
    3.885672e-06, 3.397451e-06, 2.412997e-06, 3.543709e-06, 6.88423e-06,
  3.872825e-10, 6.831773e-11, 2.01083e-15, 7.28454e-24, 1.857884e-13, 
    1.306719e-10, 4.821791e-10, 7.711807e-10, 5.283025e-07, 3.373803e-06, 
    4.293067e-06, 5.724324e-06, 5.130848e-06, 3.7484e-06, 5.070364e-06,
  2.491882e-15, 4.611326e-13, 2.599416e-09, 1.280418e-16, 4.005235e-12, 
    7.19776e-12, 1.266892e-11, 5.940644e-09, 1.76636e-07, 4.364222e-06, 
    6.914196e-06, 7.60029e-06, 6.644796e-06, 6.045446e-06, 9.034284e-06,
  3.692495e-10, 4.905245e-12, 6.560589e-12, 3.599162e-12, 2.535607e-11, 
    1.992551e-11, 1.502018e-11, 3.30149e-08, 5.325052e-08, 4.214947e-06, 
    6.152352e-06, 7.411485e-06, 7.850162e-06, 7.751263e-06, 1.084161e-05,
  7.756078e-07, 4.50163e-07, 7.452051e-09, 1.50833e-08, 1.574556e-10, 
    8.031385e-11, 2.407147e-11, 8.280592e-12, 3.558153e-08, 1.131642e-06, 
    2.544782e-06, 4.076046e-06, 5.347008e-06, 8.725156e-06, 2.03324e-05,
  1.256787e-06, 1.973335e-06, 9.393463e-07, 1.076929e-06, 2.781115e-08, 
    5.292372e-10, 7.621454e-11, 1.490652e-11, 2.975801e-10, 6.504829e-07, 
    6.152273e-07, 2.175247e-06, 4.276855e-06, 1.039696e-05, 2.787376e-05,
  1.353309e-05, 1.014336e-05, 5.841107e-06, 4.955301e-06, 3.645055e-06, 
    7.41644e-10, 2.280766e-10, 1.047831e-10, 1.967282e-10, 1.692332e-08, 
    7.879462e-08, 3.430216e-06, 5.319643e-06, 9.407107e-06, 2.388143e-05,
  3.439502e-05, 5.806888e-05, 4.95914e-05, 3.874224e-05, 3.129241e-05, 
    1.508974e-05, 1.431078e-09, 4.139793e-10, 7.989083e-10, 5.82082e-10, 
    1.168563e-08, 2.251537e-07, 7.213191e-07, 2.408517e-06, 8.614568e-06,
  5.144889e-10, 2.972777e-11, 8.700467e-12, 1.905569e-11, 6.341737e-11, 
    3.519468e-11, 1.989364e-08, 2.211342e-07, 5.490749e-07, 5.239609e-07, 
    2.941466e-06, 6.904638e-06, 9.997107e-06, 9.700464e-06, 1.350703e-05,
  3.845789e-10, 5.060099e-11, 1.073408e-10, 6.025842e-13, 1.364338e-16, 
    9.922443e-12, 7.76057e-11, 8.185626e-08, 4.564745e-08, 1.158873e-07, 
    5.16715e-06, 4.978019e-06, 5.026543e-06, 4.414918e-06, 4.119609e-06,
  8.222926e-07, 6.865396e-08, 8.546288e-15, 2.849619e-22, 4.205925e-16, 
    2.68455e-13, 1.01285e-12, 1.405946e-09, 1.983474e-09, 3.377317e-08, 
    5.432236e-06, 6.900892e-06, 5.096227e-06, 3.78912e-06, 3.181931e-06,
  4.721204e-06, 1.544106e-06, 1.420847e-17, 4.002489e-17, 2.520805e-15, 
    3.31581e-13, 1.359822e-11, 4.964138e-09, 5.431898e-09, 5.234022e-08, 
    7.518704e-06, 7.998995e-06, 5.011455e-06, 5.071233e-06, 6.717943e-06,
  1.554583e-05, 8.844864e-06, 1.221558e-14, 1.016149e-14, 2.150534e-13, 
    4.470981e-13, 6.210752e-11, 4.468437e-09, 5.171771e-09, 7.415772e-08, 
    3.702567e-06, 4.009561e-06, 3.843529e-06, 7.877886e-06, 6.057835e-06,
  3.066687e-05, 2.579424e-05, 1.43273e-05, 9.634346e-13, 8.76949e-13, 
    8.896805e-13, 2.417596e-11, 1.962489e-09, 3.060453e-09, 8.646465e-08, 
    8.766381e-07, 2.051287e-06, 4.404686e-06, 6.713868e-06, 6.647037e-06,
  5.587292e-05, 5.051596e-05, 3.881691e-05, 7.304187e-06, 2.26613e-12, 
    2.211136e-12, 7.367252e-12, 5.678578e-10, 2.144003e-09, 1.312739e-07, 
    1.452424e-06, 1.021397e-06, 5.041322e-06, 4.148705e-06, 4.526576e-06,
  7.01508e-05, 5.591442e-05, 5.630426e-05, 2.304326e-05, 8.186981e-11, 
    1.183183e-11, 4.106816e-12, 1.682763e-11, 3.970301e-09, 2.550321e-07, 
    3.402624e-06, 2.19921e-06, 6.152436e-06, 3.868816e-06, 3.278059e-06,
  8.89573e-05, 7.857529e-05, 6.690306e-05, 2.90191e-05, 1.561888e-06, 
    4.92157e-10, 9.566944e-12, 2.888284e-12, 3.53838e-10, 1.511057e-07, 
    1.182565e-06, 3.206133e-06, 2.244869e-06, 3.828293e-06, 2.541792e-06,
  0.0001163551, 0.0001274489, 8.449322e-05, 4.222649e-05, 2.216578e-06, 
    7.761508e-07, 3.042152e-11, 3.836478e-12, 1.072159e-11, 1.940462e-11, 
    4.255382e-11, 1.316777e-10, 1.682436e-10, 5.931053e-09, 1.412003e-06,
  2.291428e-09, 1.877253e-09, 2.189353e-08, 2.5346e-07, 8.301897e-07, 
    6.182211e-07, 1.095069e-06, 2.046655e-06, 4.28156e-06, 4.384195e-06, 
    6.40466e-06, 5.8842e-06, 7.023023e-06, 8.55412e-06, 9.442353e-06,
  5.807622e-05, 2.041723e-10, 7.560008e-10, 2.743035e-10, 2.847524e-09, 
    3.306021e-08, 1.123418e-07, 8.927526e-07, 2.580824e-06, 3.894218e-06, 
    4.746592e-06, 6.896685e-06, 6.473938e-06, 8.900733e-06, 9.96519e-06,
  6.278623e-05, 5.904981e-05, 1.029996e-09, 4.899398e-10, 3.01162e-10, 
    6.533111e-09, 2.780086e-08, 2.062202e-07, 6.421457e-07, 2.132864e-06, 
    5.583291e-06, 5.557272e-06, 6.772299e-06, 7.233162e-06, 8.391656e-06,
  0.0001060564, 6.624874e-05, 2.226002e-08, 2.930674e-10, 1.57264e-10, 
    4.581271e-10, 8.495553e-09, 4.798304e-08, 1.851698e-07, 4.976559e-07, 
    4.244778e-06, 5.313921e-06, 5.209215e-06, 4.340252e-06, 6.070378e-06,
  0.0001365404, 9.967291e-05, 1.11853e-07, 2.676633e-10, 3.175147e-11, 
    2.84175e-11, 2.298501e-09, 3.275774e-08, 7.680534e-08, 2.493497e-07, 
    3.65908e-06, 3.398897e-06, 4.826167e-06, 5.58552e-06, 5.050259e-06,
  0.0002102202, 0.0001649139, 7.955062e-05, 4.757611e-10, 1.675216e-11, 
    8.912184e-11, 3.859007e-10, 5.861341e-09, 2.577261e-08, 4.141847e-08, 
    2.878801e-07, 7.282422e-07, 2.038307e-06, 3.816006e-06, 3.338262e-06,
  0.0001560361, 0.0001983576, 0.00010559, 3.376822e-05, 4.206295e-11, 
    1.074593e-11, 4.006074e-11, 1.376183e-10, 6.950265e-10, 1.766161e-08, 
    5.642764e-08, 8.257756e-08, 3.414196e-07, 5.885759e-07, 2.254037e-06,
  0.0001926979, 0.0001782946, 9.576872e-05, 3.526846e-05, 7.165337e-10, 
    9.375636e-11, 5.58007e-13, 1.292425e-11, 1.18137e-10, 7.982278e-10, 
    3.805177e-10, 4.106668e-09, 3.924747e-08, 8.22765e-08, 3.067621e-07,
  0.0001268803, 0.0001318919, 6.559144e-05, 3.326358e-05, 3.316945e-05, 
    1.231468e-09, 2.170812e-11, 1.658397e-10, 1.806013e-10, 1.61944e-09, 
    6.116985e-10, 3.244196e-11, 2.939767e-09, 2.695054e-08, 3.502236e-09,
  0.0001602146, 0.0001155101, 8.794235e-05, 5.370715e-05, 5.875807e-05, 
    2.68217e-05, 5.126063e-11, 8.342972e-09, 8.139458e-10, 1.569372e-09, 
    3.999e-11, 1.065544e-11, 2.110176e-10, 1.041971e-09, 4.15915e-09,
  8.470118e-06, 1.036739e-09, 8.03199e-10, 9.450535e-09, 2.702199e-08, 
    1.605036e-07, 2.446763e-07, 5.7666e-07, 1.16299e-06, 1.235245e-06, 
    9.387246e-07, 1.224732e-06, 4.943685e-06, 1.986191e-05, 3.715018e-05,
  0.000127142, 2.703316e-09, 9.710188e-09, 1.01834e-07, 1.293333e-07, 
    9.145194e-08, 5.282433e-07, 6.075286e-07, 5.886894e-07, 6.158131e-07, 
    3.780791e-07, 1.730504e-07, 6.757516e-07, 3.688879e-06, 8.012039e-06,
  0.0001637536, 0.0001788752, 6.853186e-08, 3.999725e-07, 1.30367e-07, 
    1.268102e-07, 2.960129e-07, 7.311996e-08, 3.578817e-08, 9.237159e-09, 
    2.666741e-08, 4.154496e-08, 6.782935e-08, 2.066778e-06, 6.735638e-06,
  0.0002141189, 0.0002121248, 1.322532e-05, 4.829345e-07, 1.019967e-07, 
    7.81671e-08, 8.823431e-08, 1.239166e-08, 3.861973e-09, 8.878721e-09, 
    1.985322e-08, 1.409672e-08, 2.653686e-08, 1.350949e-07, 5.14597e-06,
  0.000236176, 0.0002314477, 1.265299e-05, 9.594327e-07, 8.097051e-08, 
    1.368389e-08, 3.576545e-08, 1.164633e-09, 4.54769e-09, 3.048344e-09, 
    1.288356e-08, 4.488923e-09, 1.233063e-08, 1.458898e-07, 3.124384e-06,
  0.0001898527, 0.0002076694, 0.0001557399, 5.729991e-06, 1.838812e-06, 
    1.903229e-07, 1.185165e-09, 2.172269e-10, 1.050448e-09, 2.049606e-09, 
    1.469734e-09, 1.144734e-09, 1.775282e-09, 1.815288e-08, 2.174605e-07,
  0.0001930184, 0.0001595848, 0.00018341, 0.0001722128, 4.421003e-06, 
    7.377257e-08, 4.120303e-10, 1.270525e-10, 2.999154e-10, 7.489286e-10, 
    3.898011e-10, 2.391965e-10, 9.003512e-10, 2.683155e-09, 2.54766e-08,
  0.0001512908, 0.0001600121, 0.0001627449, 0.0001619772, 7.794681e-07, 
    2.4889e-09, 3.331733e-10, 4.930014e-10, 2.044363e-10, 9.851612e-11, 
    2.335778e-10, 3.963886e-10, 6.090947e-10, 1.430545e-09, 2.253397e-09,
  0.0001817971, 0.0001223307, 8.81181e-05, 9.595455e-05, 0.000103323, 
    8.945636e-09, 3.044203e-10, 1.035467e-10, 3.506335e-12, 1.235733e-10, 
    3.887506e-10, 3.251168e-10, 2.418196e-10, 3.218953e-10, 1.237093e-09,
  0.0001536245, 0.0001277169, 6.974931e-05, 4.789005e-05, 4.34813e-05, 
    1.730917e-05, 4.934685e-10, 3.948784e-09, 1.35001e-07, 5.618808e-10, 
    8.045244e-10, 6.252603e-11, 6.760265e-11, 1.396359e-10, 7.895303e-08,
  2.532981e-07, 6.764144e-06, 7.740924e-06, 7.90316e-07, 3.130617e-08, 
    6.947585e-08, 1.453223e-07, 1.491969e-06, 1.000417e-05, 1.045275e-05, 
    8.461155e-06, 5.432591e-06, 1.36387e-05, 3.04106e-05, 6.585913e-05,
  0.0001822891, 2.406521e-06, 4.004944e-06, 9.324743e-07, 9.581939e-09, 
    4.949085e-08, 1.987126e-07, 3.717836e-07, 1.218072e-06, 1.02189e-06, 
    6.138363e-07, 3.770241e-07, 1.979441e-07, 1.59694e-07, 3.356666e-07,
  0.0002027784, 0.0001604808, 1.624396e-06, 6.212617e-07, 7.379664e-09, 
    2.93869e-07, 1.924855e-07, 2.904703e-07, 5.247209e-07, 1.183757e-07, 
    5.812976e-08, 3.693233e-08, 2.510689e-08, 3.141223e-08, 4.482753e-08,
  0.0001707315, 0.0001562374, 1.788674e-06, 7.27402e-09, 1.321135e-09, 
    7.391625e-08, 8.16424e-09, 3.616046e-09, 2.144753e-09, 2.299384e-08, 
    4.038948e-08, 7.278445e-09, 1.336144e-08, 2.173047e-08, 5.739695e-08,
  0.0001630742, 0.0001043786, 5.651669e-07, 9.228754e-08, 1.189349e-08, 
    2.169043e-09, 3.641437e-09, 8.626123e-10, 3.123456e-09, 1.444604e-08, 
    6.691191e-09, 3.94327e-09, 6.916227e-09, 1.395791e-08, 4.418482e-08,
  0.0001273014, 0.0001013201, 7.014766e-05, 4.3323e-07, 2.544916e-09, 
    2.610965e-10, 6.454027e-10, 3.316778e-09, 7.083214e-09, 9.643196e-09, 
    4.484331e-09, 1.031831e-09, 6.446336e-09, 5.318372e-09, 9.551214e-09,
  0.0001253303, 7.816432e-05, 7.485e-05, 5.161014e-05, 2.625666e-09, 
    3.080005e-10, 6.711517e-10, 6.186174e-09, 1.765323e-09, 9.106554e-09, 
    1.00855e-08, 1.986852e-09, 7.846766e-08, 6.686094e-09, 6.348279e-09,
  4.733825e-05, 4.267292e-05, 5.262492e-05, 4.439113e-05, 5.369252e-09, 
    5.219304e-10, 4.91505e-10, 6.762483e-10, 1.589176e-09, 2.457828e-08, 
    5.580474e-09, 3.969501e-09, 6.10818e-08, 1.971704e-07, 1.657124e-07,
  5.753585e-05, 3.94719e-05, 2.650816e-05, 2.701146e-05, 9.612497e-06, 
    8.60679e-10, 5.560178e-10, 2.617778e-09, 2.225677e-08, 4.922728e-09, 
    1.524629e-07, 1.116017e-08, 9.843003e-08, 7.036321e-08, 2.610319e-07,
  4.764929e-05, 2.629642e-05, 2.048553e-05, 1.104678e-05, 3.200105e-06, 
    2.068967e-06, 8.621232e-11, 5.071433e-07, 3.827208e-07, 7.101922e-07, 
    2.877492e-07, 8.363314e-07, 2.272459e-07, 5.868911e-07, 7.238951e-07,
  0.0002575203, 0.0002800088, 0.0002753707, 0.0002611368, 0.000267443, 
    0.0002985077, 0.0003177874, 0.0003461701, 0.0003763729, 0.0003866534, 
    0.0003735033, 0.0003751063, 0.0003368236, 0.0003255822, 0.0003123429,
  0.0003584523, 0.0003060699, 0.0003299085, 0.0003385088, 0.000332959, 
    0.0003421204, 0.0003588204, 0.0003829889, 0.0003909718, 0.0003665547, 
    0.0003501131, 0.0003432623, 0.000306145, 0.0002918046, 0.0002655679,
  0.0004666423, 0.0004983561, 0.0003797026, 0.0002956436, 0.000268578, 
    0.0002512221, 0.0002411858, 0.0002449857, 0.0002415821, 0.0002382878, 
    0.0002277674, 0.0002158194, 0.0002101332, 0.0001867737, 0.0001615863,
  0.0004255408, 0.0004576148, 0.0003008722, 0.0002321997, 0.0002308307, 
    0.0002001173, 0.0001815091, 0.0001629654, 0.0001453304, 0.00014159, 
    0.0001211023, 0.0001092656, 9.152611e-05, 6.402862e-05, 4.285121e-05,
  0.0001992204, 0.0001899753, 9.278533e-05, 0.0001025512, 0.0001522937, 
    3.650409e-05, 9.442968e-06, 1.906477e-06, 2.327521e-06, 6.215927e-06, 
    1.796806e-05, 3.226844e-05, 4.020349e-05, 4.315874e-05, 3.512756e-05,
  0.0001175631, 9.862326e-05, 0.0001131649, 7.809888e-06, 3.590763e-06, 
    4.679432e-07, 5.263417e-08, 2.22588e-08, 3.892963e-08, 2.961616e-07, 
    1.754169e-06, 5.212647e-06, 6.11243e-06, 5.001903e-06, 4.376132e-06,
  6.994088e-05, 6.37259e-05, 6.269137e-05, 4.743938e-05, 1.874183e-06, 
    5.986506e-09, 9.978318e-09, 6.128897e-08, 2.107672e-07, 1.605793e-07, 
    1.416278e-07, 3.927948e-08, 9.929168e-09, 2.934415e-09, 8.09821e-10,
  4.174604e-05, 3.077848e-05, 2.802723e-05, 2.507009e-05, 1.414914e-08, 
    9.426806e-10, 2.575536e-09, 2.093585e-09, 1.497872e-10, 5.116717e-11, 
    1.098441e-10, 8.011092e-10, 2.702594e-08, 3.446451e-08, 4.734655e-08,
  3.606077e-05, 1.113142e-05, 1.226131e-05, 1.574012e-05, 1.209889e-05, 
    6.300466e-10, 1.093004e-09, 5.542383e-10, 1.382975e-09, 1.208206e-09, 
    1.073501e-08, 1.264264e-08, 7.028552e-08, 7.280699e-08, 7.03652e-08,
  9.471932e-06, 6.860224e-06, 1.600438e-06, 7.174597e-07, 9.357352e-08, 
    7.281157e-07, 2.085118e-14, 4.194291e-09, 2.150577e-07, 2.761037e-08, 
    2.212767e-07, 8.382008e-08, 7.759197e-07, 5.393858e-07, 6.960054e-07,
  5.751305e-05, 6.178729e-05, 6.35838e-05, 6.121012e-05, 8.197041e-05, 
    8.991732e-05, 0.0001263136, 0.0001490335, 0.0001584242, 0.0001905463, 
    0.0001970498, 0.0002096197, 0.0002118304, 0.0002043058, 0.0001588851,
  0.0002878474, 0.0002401678, 0.000247812, 0.0002658576, 0.0002879172, 
    0.0003366338, 0.000352007, 0.0004225214, 0.0004814008, 0.0005135107, 
    0.0004786408, 0.0004222832, 0.0003442799, 0.0002738135, 0.000218215,
  0.0005796311, 0.0005479824, 0.0004667965, 0.0004632047, 0.0004983979, 
    0.000560724, 0.0006742786, 0.0008066603, 0.0009161211, 0.0008929675, 
    0.0007805283, 0.0005768763, 0.0003983102, 0.0002764038, 0.0001701681,
  0.0006520892, 0.0006258656, 0.0005478357, 0.000536401, 0.0005975605, 
    0.0007172831, 0.0007555676, 0.0007916139, 0.000790241, 0.0006417272, 
    0.0005283628, 0.0004595108, 0.000386608, 0.0002925019, 0.0002168914,
  0.0003385153, 0.0003832745, 0.0003710114, 0.0002893046, 0.0004151192, 
    0.0002497536, 0.0001372459, 9.420625e-05, 6.546237e-05, 4.86719e-05, 
    5.238449e-05, 5.553251e-05, 5.080149e-05, 6.867567e-05, 9.777504e-05,
  6.350363e-05, 8.04564e-05, 0.0001226625, 4.683439e-05, 1.499456e-05, 
    1.008433e-05, 8.120648e-06, 1.028533e-05, 8.942306e-06, 4.513755e-06, 
    4.088223e-06, 8.289681e-06, 4.499931e-06, 3.089113e-06, 3.366915e-06,
  4.295673e-05, 4.880039e-05, 5.622867e-05, 4.152584e-05, 1.070232e-05, 
    2.30487e-06, 1.541077e-06, 7.761701e-07, 3.815309e-07, 3.28125e-07, 
    2.666406e-07, 2.487933e-07, 1.431153e-07, 9.362915e-08, 5.303434e-08,
  7.125671e-05, 5.66104e-05, 3.959113e-05, 3.022058e-05, 3.748661e-07, 
    2.408759e-08, 5.01862e-09, 6.914485e-10, 1.295735e-10, 2.211485e-10, 
    1.66102e-08, 8.41961e-08, 7.034184e-08, 7.567555e-08, 5.339311e-08,
  4.745556e-05, 2.234636e-05, 1.710108e-05, 3.034695e-05, 2.92018e-05, 
    2.199304e-09, 7.850231e-10, 1.81778e-09, 1.484018e-10, 2.374889e-10, 
    1.759059e-08, 1.518635e-08, 5.867241e-07, 3.595548e-08, 3.541318e-07,
  2.160343e-05, 1.370329e-05, 7.511465e-06, 8.438912e-06, 1.140682e-05, 
    8.64702e-06, 1.219861e-09, 1.112937e-09, 2.518068e-10, 1.927624e-09, 
    2.905775e-07, 1.42674e-06, 1.366566e-06, 1.505552e-06, 2.098175e-06,
  1.205373e-06, 2.720445e-06, 3.215903e-06, 4.000746e-06, 2.914093e-06, 
    2.894991e-06, 4.217993e-06, 3.105844e-06, 2.696477e-06, 1.029241e-06, 
    1.173276e-06, 8.871327e-07, 7.520241e-07, 2.013527e-06, 2.300018e-05,
  1.189281e-05, 6.400108e-06, 5.48159e-06, 7.941392e-06, 5.296942e-06, 
    4.686478e-06, 4.075953e-06, 2.02267e-06, 1.559254e-06, 2.34577e-06, 
    8.322366e-06, 2.246034e-05, 5.199671e-05, 0.0001131924, 0.000199152,
  3.12269e-06, 7.386603e-06, 7.694329e-06, 1.205538e-05, 1.159187e-05, 
    6.209252e-06, 5.382959e-06, 5.907131e-06, 8.204602e-06, 2.049731e-05, 
    5.487503e-05, 0.0001235556, 0.0002242246, 0.000349273, 0.0004634982,
  0.000243642, 6.159522e-05, 6.63829e-06, 9.993436e-06, 1.612974e-05, 
    1.563837e-05, 1.411143e-05, 1.797197e-05, 6.479827e-05, 0.0001611917, 
    0.0002793502, 0.0003761618, 0.000455933, 0.0005032148, 0.0005022123,
  0.0007956981, 0.0007115733, 0.0004007484, 0.0001449509, 0.0001003998, 
    0.0001335118, 0.0002073348, 0.0003248056, 0.0004560424, 0.0005343097, 
    0.0005242578, 0.0004305223, 0.0002993758, 0.0001912423, 0.0001409299,
  0.0005938286, 0.0004226485, 0.0003036487, 0.00018194, 0.0001420853, 
    0.0001882774, 0.0002822664, 0.0003866225, 0.0003789216, 0.000217846, 
    0.0001535315, 6.297464e-05, 4.438059e-05, 3.984641e-05, 3.23778e-05,
  3.79258e-05, 2.641153e-05, 6.64032e-05, 5.351649e-05, 2.436617e-05, 
    2.248279e-05, 6.931859e-05, 0.0001058137, 4.792101e-05, 5.218866e-05, 
    4.062286e-05, 1.420467e-05, 2.19667e-06, 3.03004e-06, 5.835802e-06,
  0.0001326572, 0.0001289205, 2.400911e-05, 5.239738e-05, 1.815025e-05, 
    3.323869e-06, 8.545385e-06, 8.811665e-05, 1.404103e-05, 2.93861e-06, 
    5.161115e-06, 3.546109e-06, 1.020871e-06, 1.461889e-06, 1.764571e-06,
  8.760281e-05, 7.562468e-05, 0.0001348676, 0.0001300349, 0.0001628687, 
    1.511752e-06, 3.302171e-08, 2.999517e-06, 1.355461e-05, 3.13177e-06, 
    1.026701e-05, 1.511954e-05, 1.203079e-05, 5.358364e-06, 4.077074e-06,
  6.777627e-05, 7.698279e-06, 8.657981e-06, 9.225401e-05, 0.0001053444, 
    0.0001050005, 4.473016e-09, 3.572173e-10, 1.422251e-06, 5.37989e-06, 
    1.234522e-05, 1.962095e-05, 1.67659e-05, 1.401514e-05, 1.126014e-05,
  1.037931e-07, 1.439346e-06, 2.23199e-06, 6.287531e-06, 6.343079e-06, 
    7.798703e-06, 9.408923e-06, 5.808978e-06, 1.325823e-06, 2.498304e-06, 
    3.947691e-05, 0.0001672761, 0.0003693962, 0.0005577152, 0.000687853,
  0.0001564144, 0.0001518686, 3.354521e-05, 5.031635e-06, 5.796397e-06, 
    7.736495e-06, 1.045673e-05, 1.021775e-05, 9.926211e-06, 5.230114e-05, 
    0.0001894349, 0.000383072, 0.0005414763, 0.0006201686, 0.0006160145,
  0.0002754753, 0.0004295566, 0.0004646991, 0.0003128139, 0.0001060462, 
    2.60362e-05, 1.49545e-05, 1.502223e-05, 5.116397e-05, 0.0001214467, 
    0.0002681952, 0.0003887601, 0.0004025641, 0.0003517723, 0.0002754269,
  0.0002390945, 0.0004017952, 0.0004595182, 0.0005205274, 0.0004443524, 
    0.0003604878, 0.0003251785, 0.0003121143, 0.0003270605, 0.0003950791, 
    0.0003956154, 0.0003489782, 0.0002413116, 0.0001464724, 0.0001158513,
  0.0001366983, 0.0001641354, 0.0001907214, 0.0001931807, 0.0003186636, 
    0.0005997932, 0.0004712798, 0.0005006175, 0.000524151, 0.0004813926, 
    0.0003730125, 0.0002375407, 0.0001493805, 9.96653e-05, 7.715774e-05,
  8.274923e-05, 4.188976e-05, 5.584176e-05, 3.933288e-05, 3.603802e-05, 
    0.0002538451, 0.0003607912, 0.0002814549, 0.0002487616, 0.0002081699, 
    0.0001583727, 0.0001138511, 7.452602e-05, 6.149176e-05, 4.287078e-05,
  0.0001109893, 5.85338e-05, 3.644635e-05, 7.080146e-05, 9.025595e-06, 
    3.267278e-05, 0.0001746577, 9.314877e-05, 5.249155e-05, 7.252182e-05, 
    6.843506e-05, 7.826358e-05, 7.830853e-05, 7.315844e-05, 5.434802e-05,
  0.0001001954, 5.92713e-05, 6.8876e-05, 7.313395e-05, 9.934141e-06, 
    1.018494e-05, 2.935398e-05, 6.33137e-05, 2.908001e-05, 3.628636e-05, 
    5.753873e-05, 4.434424e-05, 5.351068e-05, 5.330385e-05, 4.126669e-05,
  0.0001308143, 7.188263e-05, 0.0001163253, 0.0001158957, 0.0001439599, 
    2.621921e-05, 3.55781e-05, 4.050803e-05, 3.716077e-05, 1.154865e-05, 
    2.200377e-05, 3.99145e-05, 3.099345e-05, 8.120517e-06, 2.11423e-05,
  0.0001461952, 0.0001204983, 0.0001292336, 0.0001236752, 0.0001567297, 
    0.0001032897, 1.609777e-05, 1.296664e-05, 1.372293e-05, 3.046842e-05, 
    2.742607e-05, 4.04809e-05, 1.85753e-05, 2.296572e-05, 3.403993e-06,
  2.376259e-23, 5.30548e-12, 1.328914e-10, 7.393255e-11, 5.407719e-12, 
    1.082174e-10, 1.81811e-09, 7.034382e-08, 5.341487e-07, 5.471174e-07, 
    3.963356e-06, 6.432324e-06, 6.471663e-06, 7.785918e-06, 3.059111e-05,
  8.724715e-24, 2.92814e-23, 2.540423e-12, 3.414858e-11, 1.718409e-10, 
    7.559582e-08, 1.594316e-07, 4.565407e-07, 8.428441e-07, 9.73061e-07, 
    2.79177e-06, 3.602477e-06, 2.668979e-06, 2.976812e-06, 2.35803e-05,
  8.448974e-14, 5.221606e-10, 1.231593e-08, 2.239825e-09, 8.275186e-11, 
    1.746132e-09, 4.322461e-09, 2.161962e-09, 5.462683e-07, 1.394743e-06, 
    3.635118e-06, 9.067431e-06, 2.341146e-05, 4.205266e-05, 4.130954e-05,
  1.126849e-10, 1.469702e-10, 1.657679e-09, 9.983276e-14, 3.291234e-11, 
    2.385949e-10, 1.030647e-10, 8.073804e-09, 1.793862e-06, 7.136317e-06, 
    4.184079e-05, 7.591036e-05, 9.772523e-05, 0.0001021155, 0.0001103603,
  1.037927e-08, 5.591196e-08, 4.281034e-10, 6.031775e-12, 1.011145e-09, 
    1.061048e-08, 3.389434e-09, 5.081652e-07, 1.990313e-05, 6.485836e-05, 
    0.0001138788, 0.0001310775, 0.0001066771, 9.805746e-05, 0.0001500517,
  1.378401e-06, 1.39602e-06, 3.44831e-07, 1.57358e-07, 1.967351e-07, 
    5.980246e-07, 1.675137e-06, 1.169651e-05, 5.478081e-05, 0.0001101772, 
    0.0001532943, 0.0001824424, 0.00018466, 0.0001527818, 0.0001999017,
  5.655038e-06, 3.231111e-06, 3.367287e-06, 3.828567e-06, 3.090501e-06, 
    3.50942e-06, 1.602405e-05, 4.642659e-05, 4.631572e-05, 6.917783e-05, 
    9.812252e-05, 0.0001400686, 0.0001946956, 0.0002555289, 0.000325276,
  1.774398e-05, 5.667791e-06, 4.880886e-06, 8.377129e-06, 5.367697e-06, 
    8.409028e-06, 2.426929e-05, 1.902414e-05, 1.575154e-05, 5.334641e-06, 
    1.409738e-05, 9.589072e-06, 4.983587e-05, 0.0001600601, 0.0002757203,
  5.401836e-06, 1.440978e-05, 1.154038e-05, 1.236123e-05, 8.875885e-06, 
    1.492692e-05, 2.128612e-05, 1.247397e-05, 3.432258e-05, 7.380832e-06, 
    9.360881e-06, 1.112212e-05, 1.263049e-05, 1.798752e-05, 0.0001335092,
  1.835157e-05, 1.168149e-05, 9.398107e-06, 9.290393e-06, 9.790698e-06, 
    2.665603e-05, 3.7864e-06, 2.067705e-07, 1.746616e-05, 3.474075e-05, 
    7.859852e-06, 4.104232e-05, 8.249142e-05, 3.505967e-05, 3.501422e-05,
  6.05976e-10, 9.614779e-11, 6.339824e-13, 6.370495e-11, 4.420517e-10, 
    1.60361e-09, 2.583345e-09, 5.017787e-09, 4.196421e-09, 6.505678e-09, 
    1.043369e-08, 8.495753e-09, 1.304338e-08, 1.954367e-08, 1.926448e-07,
  4.630149e-09, 4.81379e-09, 1.682308e-09, 4.007163e-10, 2.985419e-09, 
    2.406229e-09, 1.324827e-09, 1.310173e-09, 2.075623e-09, 2.373593e-09, 
    1.22664e-08, 1.388974e-08, 1.466485e-07, 2.781786e-07, 3.229469e-07,
  3.261377e-09, 6.61119e-10, 2.072055e-09, 5.290336e-10, 1.364922e-09, 
    1.115078e-09, 2.992321e-09, 5.924285e-09, 7.830893e-09, 2.224026e-09, 
    3.022273e-09, 8.72983e-08, 2.184115e-08, 3.102975e-07, 4.811055e-08,
  2.842552e-09, 1.161495e-08, 4.681521e-08, 2.166324e-09, 1.540208e-09, 
    2.141571e-10, 5.0384e-10, 1.774098e-09, 1.336731e-09, 5.250758e-09, 
    2.340363e-09, 2.181617e-08, 2.843496e-07, 2.12795e-07, 8.996755e-08,
  2.391954e-09, 7.31642e-09, 1.262716e-08, 2.239363e-09, 7.563603e-10, 
    1.655696e-09, 6.983033e-10, 1.03044e-08, 1.774309e-08, 1.024847e-08, 
    1.238813e-09, 1.609975e-08, 5.918822e-07, 1.728342e-07, 9.611246e-09,
  4.331336e-09, 1.31933e-08, 3.807775e-08, 9.594655e-08, 2.457056e-07, 
    2.743624e-08, 2.127135e-08, 3.128723e-09, 1.048436e-08, 2.54242e-08, 
    1.857052e-09, 9.724956e-08, 6.30815e-08, 1.022758e-08, 5.897502e-09,
  1.904697e-09, 4.900635e-09, 1.310602e-08, 3.394198e-10, 9.943277e-10, 
    3.764997e-10, 6.036345e-10, 1.394926e-09, 3.769354e-09, 2.925964e-09, 
    1.285763e-09, 1.300073e-08, 3.174831e-09, 4.891224e-10, 7.688672e-10,
  9.285811e-08, 3.690954e-08, 1.057261e-08, 2.711057e-08, 3.919064e-10, 
    4.837262e-10, 2.162476e-10, 2.777217e-09, 2.958987e-09, 5.29883e-10, 
    5.041064e-10, 7.806525e-10, 1.126636e-08, 1.021427e-09, 1.359163e-09,
  6.355678e-07, 1.143692e-06, 1.533139e-07, 1.390698e-09, 1.100005e-07, 
    1.16068e-08, 2.801416e-08, 1.303703e-08, 2.528638e-09, 6.908182e-10, 
    5.460593e-10, 1.004095e-09, 2.620622e-09, 2.417232e-10, 3.481442e-10,
  1.501749e-06, 1.019711e-06, 3.549628e-06, 3.538808e-06, 2.814002e-07, 
    1.023795e-06, 1.582045e-06, 2.004244e-07, 4.823196e-07, 4.158226e-08, 
    4.071038e-08, 1.550564e-08, 6.986854e-10, 1.550408e-09, 2.456766e-09,
  6.313078e-09, 4.666022e-06, 4.442686e-06, 1.038153e-05, 3.734816e-06, 
    1.564068e-06, 1.663503e-06, 3.365285e-07, 6.806744e-08, 2.631009e-08, 
    2.679931e-09, 6.759142e-09, 1.441443e-08, 4.603038e-08, 1.073998e-07,
  2.408908e-06, 2.450167e-06, 1.756097e-06, 2.783961e-06, 4.249104e-06, 
    3.735946e-06, 2.843487e-06, 8.398201e-07, 2.554624e-07, 2.492697e-09, 
    1.159159e-09, 2.481633e-09, 2.925207e-09, 3.604269e-09, 4.251482e-09,
  1.097006e-05, 9.221073e-06, 3.577299e-07, 3.048824e-06, 2.002476e-06, 
    3.015194e-06, 2.75102e-06, 2.71334e-06, 2.589872e-06, 4.169395e-07, 
    1.054038e-08, 5.003913e-09, 1.384276e-09, 2.082835e-09, 2.561903e-09,
  3.18158e-05, 1.842286e-05, 1.852041e-06, 1.118973e-06, 2.35901e-06, 
    2.105954e-06, 1.670762e-06, 6.146649e-06, 2.769753e-06, 2.142922e-06, 
    1.695321e-06, 4.65639e-07, 9.575668e-08, 4.501188e-08, 1.298075e-07,
  5.615448e-05, 3.65652e-05, 2.346066e-06, 3.578717e-07, 5.410938e-07, 
    2.482024e-06, 3.530587e-06, 2.507247e-06, 4.438556e-06, 3.606785e-06, 
    3.280391e-06, 2.444968e-06, 1.760121e-06, 1.893122e-06, 1.526152e-06,
  3.921117e-05, 2.742514e-05, 2.236398e-05, 5.052422e-07, 1.342183e-07, 
    1.585472e-06, 8.69878e-07, 2.257563e-06, 2.739037e-06, 3.334124e-06, 
    3.851422e-06, 5.396153e-06, 1.392434e-06, 1.141815e-06, 9.695151e-07,
  2.624292e-05, 1.678601e-05, 1.459292e-05, 9.964097e-06, 3.359998e-07, 
    1.362245e-07, 1.215521e-06, 1.09592e-06, 2.038812e-06, 2.123013e-06, 
    2.024767e-06, 1.862795e-06, 3.368394e-06, 2.185202e-06, 9.328118e-07,
  1.600395e-05, 8.783785e-06, 4.685087e-06, 5.606191e-06, 1.393691e-07, 
    1.228403e-06, 5.493294e-07, 5.109173e-07, 6.233761e-07, 7.74769e-07, 
    2.545764e-06, 1.136208e-06, 5.944948e-06, 2.278173e-06, 1.744174e-06,
  1.843026e-05, 8.859628e-06, 2.476055e-06, 4.555105e-06, 6.507132e-06, 
    8.174193e-07, 1.828656e-06, 5.894482e-07, 8.845668e-07, 1.129476e-06, 
    1.63148e-06, 4.139589e-06, 4.38799e-06, 3.491441e-06, 1.563542e-06,
  2.539364e-05, 1.389105e-05, 1.490151e-05, 5.116029e-06, 3.264063e-06, 
    9.419317e-06, 3.667701e-06, 2.659808e-06, 3.158399e-06, 2.074934e-06, 
    2.074288e-06, 2.644344e-06, 4.379712e-06, 3.049001e-06, 3.667581e-06,
  8.706799e-05, 0.0001599341, 0.0002879784, 0.0003626202, 0.0003583888, 
    0.0003386678, 0.0003503926, 0.000370136, 0.0003579827, 0.0003200044, 
    0.0002630558, 0.0002042766, 0.0001588042, 0.0001261278, 0.0001010793,
  0.000168082, 0.0002687486, 0.0002899049, 0.0002549889, 0.000202989, 
    0.0002060835, 0.0002442101, 0.0002955701, 0.0003421478, 0.0003546995, 
    0.0003648319, 0.0003451316, 0.0003225942, 0.0002796075, 0.0002878923,
  0.0003042695, 0.0002724508, 8.037056e-05, 0.0002047662, 9.076553e-05, 
    8.906342e-05, 0.0001171565, 0.0001619772, 0.0002106718, 0.0002500527, 
    0.0002897943, 0.0003217537, 0.000326599, 0.0003388203, 0.0003448551,
  0.000308242, 0.0002149488, 1.468515e-05, 1.111285e-05, 4.748847e-05, 
    1.245957e-05, 2.092735e-05, 3.450651e-05, 6.647054e-05, 9.677801e-05, 
    0.0001331596, 0.0001773499, 0.0002132056, 0.0002350924, 0.0002775843,
  8.149919e-05, 6.315862e-05, 2.666153e-05, 1.826099e-05, 1.147154e-05, 
    1.153697e-05, 5.148531e-06, 6.443207e-06, 1.012753e-05, 1.035297e-05, 
    2.034468e-05, 2.622445e-05, 4.323512e-05, 5.768304e-05, 5.308093e-05,
  0.0001074912, 0.0001448252, 0.0001160396, 2.323888e-05, 3.069927e-06, 
    7.92168e-07, 1.254469e-06, 2.633216e-06, 2.779687e-06, 1.504174e-06, 
    3.843713e-06, 6.28524e-06, 1.032303e-05, 2.039544e-05, 2.570559e-05,
  0.0003916358, 0.0003115872, 0.0002337916, 0.0001392702, 0.0001147795, 
    1.5505e-05, 1.769873e-05, 1.853583e-05, 7.572418e-06, 1.34409e-07, 
    2.424038e-07, 4.617939e-07, 3.1809e-06, 3.812919e-06, 5.584613e-06,
  0.0008369737, 0.0006290954, 0.0003459247, 0.0001787866, 3.473432e-05, 
    1.83113e-05, 4.21361e-05, 4.566557e-05, 2.093326e-05, 5.169088e-08, 
    4.774872e-07, 4.518512e-08, 1.269716e-07, 1.460365e-07, 1.089759e-07,
  0.0008257233, 0.0005574157, 0.0004493313, 0.0002024341, 0.0001572082, 
    6.503913e-06, 2.651917e-05, 3.129177e-05, 4.412409e-06, 7.152007e-07, 
    2.851585e-06, 1.309442e-06, 2.389488e-06, 1.966197e-08, 1.733436e-06,
  0.0005013969, 0.0004457944, 0.0002450837, 0.0001694191, 0.0001683349, 
    0.0001398916, 1.450412e-05, 6.298336e-06, 1.101638e-06, 1.750745e-06, 
    2.458653e-06, 2.483675e-06, 4.442351e-06, 3.903952e-06, 5.293355e-06,
  5.501245e-06, 6.826853e-06, 3.057393e-05, 6.168084e-05, 9.112214e-05, 
    9.271812e-05, 8.258878e-05, 0.000101097, 0.0001262294, 0.0001262778, 
    0.000127874, 0.000124797, 0.0001120534, 0.0001173336, 0.0001277562,
  2.928808e-05, 5.785599e-05, 6.245271e-05, 8.62634e-05, 0.0001022179, 
    0.000112801, 0.0001238595, 0.000160244, 0.0002193425, 0.0002888882, 
    0.000352449, 0.0003996778, 0.0004494272, 0.0004817046, 0.0005076498,
  4.518787e-05, 4.2179e-05, 4.020424e-05, 3.798843e-05, 3.98238e-05, 
    5.223196e-05, 0.0001021805, 0.0001656281, 0.0002467699, 0.0003473733, 
    0.000446198, 0.000502357, 0.0005723716, 0.0006436689, 0.000687382,
  5.834957e-05, 6.472859e-05, 4.855757e-05, 4.629179e-05, 4.858294e-05, 
    6.359457e-05, 9.457667e-05, 0.000142187, 0.0002673423, 0.0004961449, 
    0.0006568761, 0.0007401683, 0.0007671427, 0.0007895298, 0.0007599007,
  3.46913e-05, 5.634703e-05, 4.30561e-05, 3.796077e-05, 3.344366e-05, 
    4.735599e-05, 0.0001113354, 0.0005100411, 0.001025779, 0.001286465, 
    0.001187437, 0.001049092, 0.0009558033, 0.0007509268, 0.0005934422,
  2.212719e-05, 6.008477e-05, 9.815619e-05, 9.198426e-05, 0.0001305182, 
    0.0003477332, 0.0007668673, 0.001449814, 0.00188811, 0.001914644, 
    0.001885137, 0.001799837, 0.001481684, 0.0008116908, 0.0003539191,
  3.534035e-05, 0.0001712488, 0.0003613853, 0.0005027166, 0.0006596245, 
    0.0008891753, 0.001267369, 0.001549175, 0.001897775, 0.0018424, 
    0.001833142, 0.001715449, 0.001379175, 0.0008604168, 0.0003899664,
  9.888468e-05, 0.000442197, 0.0007193884, 0.0009140249, 0.001298334, 
    0.000959203, 0.001257202, 0.0009855705, 0.0008693071, 0.000813526, 
    0.0009164395, 0.0009403506, 0.0008233518, 0.0006055172, 0.0003928381,
  0.0001392939, 0.0004771053, 0.0006798301, 0.0007731016, 0.0007660635, 
    0.0005116157, 0.000545577, 0.0004464607, 0.0002994848, 0.000344574, 
    0.0003753127, 0.0003627062, 0.0002958535, 0.0002684199, 0.0002270737,
  8.818252e-05, 0.0002701942, 0.0004234802, 0.0004437678, 0.0003976669, 
    0.0003609062, 0.0003516267, 0.0003583776, 0.0002021292, 0.0001719927, 
    0.0001075277, 7.331427e-05, 4.162824e-05, 2.604262e-05, 4.134222e-05,
  6.114019e-06, 4.802073e-06, 8.985783e-06, 4.830866e-06, 2.558502e-06, 
    1.625354e-06, 2.029739e-06, 6.381509e-06, 6.32471e-06, 5.198591e-06, 
    2.462963e-06, 9.193381e-07, 4.953935e-07, 1.16456e-07, 1.352913e-08,
  1.475426e-05, 1.044967e-05, 9.24039e-06, 6.958704e-06, 3.39906e-06, 
    4.076251e-06, 6.144493e-06, 9.32552e-06, 2.599076e-06, 1.159653e-06, 
    2.914848e-07, 8.774941e-08, 4.447909e-08, 1.68142e-07, 3.553788e-08,
  7.031392e-06, 1.47238e-05, 1.084783e-05, 8.520749e-06, 5.614535e-06, 
    6.097909e-06, 7.135581e-06, 4.095882e-06, 1.442023e-06, 1.834161e-07, 
    9.721997e-08, 9.617947e-08, 3.154407e-07, 2.197064e-07, 2.276311e-06,
  7.998626e-06, 9.198221e-06, 1.026857e-05, 1.206127e-05, 9.526923e-06, 
    9.754745e-06, 7.733745e-06, 2.622284e-06, 1.951889e-07, 2.165141e-07, 
    2.855186e-07, 2.449097e-08, 8.624547e-08, 1.380642e-07, 4.508485e-07,
  8.890261e-06, 9.986928e-06, 1.210562e-05, 1.166491e-05, 1.151205e-05, 
    9.710693e-06, 5.990872e-06, 1.27076e-06, 8.133006e-08, 4.882399e-08, 
    8.445592e-08, 5.379287e-05, 0.0003758563, 0.0003573252, 0.0001189304,
  5.6064e-06, 1.078653e-05, 1.799467e-05, 1.508378e-05, 1.224657e-05, 
    1.020523e-05, 4.048379e-06, 7.613274e-07, 1.420089e-06, 1.022156e-06, 
    5.994221e-05, 0.0006059263, 0.001414326, 0.001720604, 0.001928144,
  4.514827e-06, 1.02247e-05, 1.099824e-05, 1.40346e-05, 1.488916e-05, 
    1.092351e-05, 4.119679e-06, 5.824551e-06, 4.64717e-06, 5.211841e-06, 
    8.103823e-05, 0.0004307978, 0.001093707, 0.001594316, 0.001866416,
  7.732301e-07, 6.823468e-06, 7.758049e-06, 1.264448e-05, 1.475618e-05, 
    1.171326e-05, 1.298727e-05, 1.539627e-05, 1.094447e-05, 7.453245e-06, 
    5.552098e-05, 0.0001016447, 0.0002276936, 0.0004526463, 0.0007344051,
  6.170469e-07, 7.779125e-07, 4.81645e-06, 5.10585e-06, 1.147969e-05, 
    1.475117e-05, 1.587415e-05, 1.832016e-05, 1.634864e-05, 9.071392e-06, 
    3.749415e-05, 5.86158e-05, 8.033455e-05, 0.0001552097, 0.0003373917,
  8.848361e-09, 7.446837e-08, 2.39772e-06, 1.073293e-05, 1.317071e-05, 
    2.04014e-05, 2.148142e-05, 2.584823e-05, 2.271355e-05, 1.791878e-05, 
    1.954402e-05, 4.358769e-05, 6.420478e-05, 9.236294e-05, 0.0001631246,
  1.941464e-09, 1.585914e-08, 2.795023e-09, 2.600019e-10, 3.32588e-12, 
    4.035284e-11, 3.177972e-12, 6.643578e-12, 4.456602e-09, 2.617083e-07, 
    3.754975e-07, 2.568886e-07, 6.696832e-07, 9.855817e-07, 1.13453e-06,
  3.182628e-07, 9.341792e-07, 6.973256e-07, 3.765048e-09, 2.771763e-10, 
    6.026876e-11, 3.00816e-10, 1.770784e-10, 9.553085e-09, 1.10577e-07, 
    2.610571e-07, 3.676461e-08, 4.25762e-08, 1.367087e-07, 7.198405e-07,
  1.991926e-07, 1.165805e-06, 3.06991e-06, 1.338216e-08, 1.492847e-09, 
    4.079668e-11, 2.794023e-10, 1.962017e-10, 9.542868e-10, 3.289868e-09, 
    4.177407e-08, 9.33787e-08, 4.690157e-08, 1.254961e-08, 5.745632e-08,
  3.446758e-07, 9.373726e-08, 5.918851e-07, 4.110344e-06, 1.318909e-08, 
    1.120305e-09, 2.163368e-10, 8.044545e-10, 4.347357e-09, 3.04443e-09, 
    3.144573e-08, 1.050346e-07, 9.388895e-08, 9.631327e-09, 1.608838e-10,
  6.913778e-07, 1.055558e-06, 1.657532e-06, 2.054466e-06, 1.086145e-06, 
    7.902496e-08, 1.823196e-07, 1.400015e-07, 1.209016e-09, 5.4777e-09, 
    1.16881e-07, 5.326314e-08, 2.333295e-07, 8.184494e-08, 1.382533e-09,
  7.097756e-07, 8.374624e-07, 3.191304e-06, 4.269919e-06, 2.708827e-06, 
    1.481988e-06, 1.607108e-07, 6.378793e-08, 7.490159e-09, 8.629054e-08, 
    1.087581e-08, 3.346977e-07, 2.407609e-07, 3.671797e-08, 4.945974e-09,
  2.681412e-07, 1.433926e-06, 6.368999e-06, 1.08905e-05, 5.811957e-06, 
    4.573875e-06, 1.584027e-06, 4.355055e-07, 9.177122e-07, 4.850256e-08, 
    7.649584e-07, 6.445521e-07, 4.069251e-07, 4.95751e-08, 1.06888e-08,
  1.010667e-07, 6.285647e-07, 4.143993e-06, 1.137504e-05, 1.143469e-05, 
    9.211785e-06, 1.858425e-06, 1.153065e-06, 2.241409e-06, 4.905785e-07, 
    2.018574e-06, 1.2506e-06, 6.004554e-07, 2.642633e-07, 1.546542e-07,
  1.945919e-08, 3.265667e-07, 8.507397e-07, 3.213224e-06, 9.48514e-06, 
    7.847432e-06, 7.368873e-06, 9.25772e-06, 3.009119e-06, 2.009971e-06, 
    9.318964e-07, 1.461327e-06, 1.2863e-06, 4.094348e-07, 7.616889e-07,
  2.248951e-07, 4.457104e-07, 1.321307e-06, 3.240345e-06, 5.336292e-06, 
    1.082451e-05, 6.949223e-06, 1.039824e-05, 1.194673e-05, 4.00623e-06, 
    1.019465e-06, 5.217806e-07, 2.978319e-07, 3.329046e-08, 1.127641e-06,
  6.106536e-08, 2.532748e-08, 9.852279e-09, 6.194541e-08, 1.083489e-08, 
    8.805971e-10, 2.20611e-09, 1.019049e-08, 4.42822e-07, 3.824658e-06, 
    1.666503e-06, 1.462842e-06, 1.060504e-06, 1.016658e-06, 3.241979e-07,
  2.841484e-07, 7.409304e-08, 1.782407e-07, 2.978042e-07, 2.713905e-08, 
    8.057575e-09, 1.436924e-09, 1.467027e-09, 3.275749e-09, 9.194025e-07, 
    1.578544e-06, 1.798723e-06, 2.255158e-06, 1.849168e-06, 7.308112e-07,
  6.379565e-07, 1.188603e-06, 2.193107e-06, 1.546916e-06, 4.434461e-07, 
    1.201309e-07, 5.115363e-08, 6.689002e-09, 6.518916e-10, 4.544769e-08, 
    5.938749e-07, 1.185607e-06, 1.71214e-06, 7.391122e-07, 1.787893e-06,
  1.453157e-06, 1.321857e-06, 3.479002e-06, 2.564211e-06, 1.208594e-06, 
    8.194608e-07, 3.950716e-07, 1.332812e-07, 5.405155e-09, 3.837971e-08, 
    2.125445e-08, 9.670434e-08, 6.502067e-07, 8.46922e-07, 2.083274e-06,
  1.062612e-06, 1.774501e-06, 3.26667e-06, 3.158375e-06, 3.139298e-06, 
    2.224526e-06, 1.846359e-06, 8.966106e-07, 6.992088e-08, 5.54037e-08, 
    1.145193e-07, 1.382655e-08, 8.091649e-08, 3.191724e-07, 6.143237e-07,
  6.906379e-07, 1.495062e-06, 3.281941e-06, 3.950453e-06, 2.110491e-06, 
    3.940006e-06, 3.721709e-06, 2.86313e-06, 1.864576e-06, 4.244106e-07, 
    4.03888e-07, 2.264952e-07, 1.557599e-07, 2.150994e-08, 1.553394e-07,
  5.210898e-07, 1.275324e-06, 4.739035e-06, 6.226626e-06, 3.177869e-06, 
    3.512352e-06, 6.919149e-06, 5.221098e-06, 4.727081e-06, 4.598386e-06, 
    2.452007e-06, 1.63373e-06, 5.384418e-07, 1.17631e-07, 2.186303e-08,
  3.762764e-07, 6.670689e-07, 2.19926e-06, 5.941373e-06, 3.49451e-06, 
    6.11317e-06, 2.90463e-06, 4.724682e-06, 5.216106e-06, 5.92602e-06, 
    5.775519e-06, 5.880356e-06, 3.08655e-06, 2.138483e-06, 8.112969e-08,
  4.280683e-07, 9.624307e-08, 5.300179e-07, 3.843796e-06, 5.484575e-06, 
    5.12256e-06, 4.893887e-06, 5.116557e-06, 5.913559e-06, 5.71791e-06, 
    6.690542e-06, 8.676887e-06, 9.286676e-06, 2.663796e-06, 1.701201e-06,
  4.780949e-07, 4.475897e-08, 1.607882e-06, 2.424043e-06, 2.4061e-06, 
    4.734902e-06, 6.204995e-06, 8.42274e-06, 2.948237e-05, 2.929337e-05, 
    4.930676e-06, 1.167753e-05, 7.048009e-06, 1.244448e-06, 3.766043e-06,
  1.267921e-09, 6.192973e-07, 3.682479e-06, 3.529314e-06, 1.541028e-06, 
    3.886284e-06, 2.113329e-06, 1.245148e-06, 3.385385e-06, 1.678331e-06, 
    2.175133e-06, 2.074644e-06, 1.608941e-06, 2.33599e-06, 1.768506e-06,
  4.268544e-07, 1.420169e-07, 2.770128e-06, 7.409657e-06, 5.121579e-06, 
    9.570661e-06, 2.403411e-06, 1.317018e-06, 1.81559e-06, 2.708688e-06, 
    2.70782e-06, 1.969247e-06, 2.581955e-06, 3.07325e-06, 2.842905e-06,
  7.678381e-07, 2.225019e-06, 1.045262e-06, 9.323448e-06, 8.479162e-06, 
    1.005707e-05, 3.168278e-06, 7.736774e-07, 2.24149e-06, 4.727491e-06, 
    3.448082e-06, 4.371267e-06, 3.680833e-06, 4.592372e-06, 4.968014e-06,
  2.259756e-06, 2.674912e-06, 4.10645e-06, 4.620638e-06, 2.156118e-05, 
    7.21196e-06, 4.539164e-06, 1.560474e-06, 2.286187e-06, 5.100028e-06, 
    4.075493e-06, 2.076777e-06, 3.246474e-06, 3.955142e-06, 5.236048e-06,
  2.498569e-06, 3.572307e-06, 6.94654e-06, 5.079093e-06, 6.693508e-06, 
    1.094788e-05, 5.496446e-06, 8.086597e-07, 1.328178e-06, 3.251436e-06, 
    2.962653e-06, 2.747232e-06, 4.649436e-06, 4.922799e-06, 3.261764e-06,
  2.442938e-06, 3.736839e-06, 8.9926e-06, 5.664471e-06, 1.714643e-06, 
    7.719003e-06, 5.078027e-06, 2.64366e-06, 1.874632e-06, 1.244266e-06, 
    2.805001e-06, 5.031866e-06, 3.570691e-06, 4.351953e-06, 2.420211e-06,
  3.941667e-06, 3.116783e-06, 1.155134e-05, 1.465689e-05, 3.057489e-06, 
    4.398272e-06, 7.344681e-06, 9.305909e-06, 5.905373e-06, 2.352526e-06, 
    2.915635e-06, 6.476461e-06, 4.655799e-06, 3.481443e-06, 4.393354e-06,
  3.169132e-06, 2.407518e-06, 1.317522e-05, 2.1718e-05, 2.26669e-06, 
    1.667358e-06, 6.50266e-06, 1.348844e-05, 1.00491e-05, 1.266777e-05, 
    6.156148e-06, 6.391517e-06, 6.747503e-06, 5.790643e-06, 5.825182e-06,
  2.947173e-06, 2.860164e-06, 8.195335e-06, 1.579552e-05, 1.041638e-05, 
    2.095069e-06, 7.260729e-06, 1.263533e-05, 2.11529e-05, 1.311246e-05, 
    2.364178e-05, 1.208914e-05, 7.278667e-06, 8.283564e-06, 1.013665e-05,
  2.514511e-06, 4.315191e-06, 9.044587e-06, 1.632892e-05, 5.226172e-06, 
    8.361848e-06, 1.759784e-05, 3.074738e-05, 1.73319e-05, 2.650577e-05, 
    3.561323e-05, 2.111434e-05, 1.723406e-05, 1.873169e-05, 1.66314e-05,
  5.596316e-06, 5.623634e-08, 1.552296e-06, 8.502246e-06, 1.6227e-05, 
    1.392794e-05, 6.11723e-06, 2.467685e-06, 1.465107e-06, 1.262479e-06, 
    1.083102e-06, 7.774941e-07, 1.37756e-06, 2.43062e-06, 6.157799e-06,
  2.291564e-05, 1.922079e-08, 3.119611e-07, 7.549623e-07, 1.149788e-07, 
    1.255876e-08, 3.146282e-08, 2.919506e-07, 2.033292e-07, 3.737529e-07, 
    4.023742e-07, 7.920418e-07, 8.286761e-07, 2.564079e-06, 8.090742e-06,
  1.73306e-05, 6.287104e-06, 5.560625e-09, 4.383662e-07, 9.880131e-09, 
    4.705766e-09, 1.607279e-08, 3.784979e-08, 5.498484e-08, 7.615685e-08, 
    1.58181e-07, 4.59107e-07, 4.443112e-07, 2.713025e-06, 7.531904e-06,
  6.157466e-06, 1.981527e-06, 7.25231e-09, 2.376725e-09, 7.344095e-07, 
    8.428074e-09, 5.893404e-09, 2.648463e-07, 9.32643e-08, 9.538425e-08, 
    2.190045e-08, 7.584449e-08, 2.884935e-07, 1.629821e-06, 4.012969e-06,
  9.242238e-06, 8.071842e-06, 4.528624e-10, 6.975268e-08, 1.058578e-06, 
    1.481663e-06, 7.353395e-09, 1.055293e-08, 2.349257e-07, 4.008743e-07, 
    4.125546e-07, 2.509104e-07, 1.761345e-07, 1.548487e-06, 2.524374e-06,
  9.510457e-06, 1.005308e-05, 8.918594e-06, 1.103267e-08, 4.445271e-07, 
    9.36371e-07, 2.738935e-07, 1.492886e-08, 3.330568e-07, 8.258048e-07, 
    8.342722e-07, 5.551311e-07, 1.811159e-07, 1.017587e-06, 1.410906e-06,
  8.84912e-06, 1.04351e-05, 1.739649e-05, 1.876986e-05, 2.196845e-07, 
    6.711753e-07, 1.101323e-06, 2.363618e-07, 5.271625e-07, 6.304024e-07, 
    1.302832e-06, 1.496573e-06, 2.432958e-06, 5.284612e-06, 5.371799e-06,
  5.211112e-06, 1.282495e-05, 1.852717e-05, 3.25716e-05, 2.468832e-09, 
    7.982429e-07, 9.621399e-07, 1.268157e-06, 1.392796e-06, 5.646507e-07, 
    2.002955e-06, 2.09349e-06, 4.00316e-06, 3.477332e-06, 4.168307e-06,
  7.4963e-06, 6.375537e-06, 1.762175e-05, 4.01387e-05, 3.378935e-05, 
    1.953709e-07, 2.362241e-06, 1.553131e-06, 1.2744e-06, 1.540567e-06, 
    2.124061e-06, 2.242626e-06, 1.970574e-06, 2.917361e-06, 7.992188e-06,
  6.148711e-06, 8.17099e-06, 1.174273e-05, 2.774158e-05, 4.530275e-05, 
    3.308114e-05, 2.695078e-06, 3.000915e-06, 1.330009e-06, 2.6445e-06, 
    3.763354e-06, 5.40679e-06, 4.906246e-06, 1.044771e-05, 1.736105e-05,
  3.443892e-07, 4.817037e-06, 1.557231e-05, 3.261036e-05, 5.965672e-05, 
    0.0001031751, 0.0001475072, 0.0002251557, 0.0002770464, 0.0003131161, 
    0.0003244205, 0.0002644334, 0.0001983033, 0.0001553452, 0.0001391564,
  1.117693e-07, 4.34378e-07, 1.640191e-05, 6.436582e-05, 0.0001269619, 
    0.0001927182, 0.0002618997, 0.0002929436, 0.0002722298, 0.0002611479, 
    0.000216541, 0.0001829559, 0.0001592924, 0.0001361283, 0.0001086097,
  1.673333e-06, 2.593595e-06, 7.875874e-06, 4.673968e-05, 0.0001249716, 
    0.0001850696, 0.000224912, 0.0002386542, 0.000222265, 0.0001928137, 
    0.0001666432, 0.00015967, 0.0001401352, 0.0001150047, 9.17704e-05,
  4.343396e-06, 6.940724e-06, 8.963578e-06, 2.563752e-05, 7.55974e-05, 
    9.715659e-05, 0.0001094128, 0.0001211374, 0.0001264805, 0.0001108706, 
    0.0001049554, 0.0001003738, 9.623148e-05, 7.823432e-05, 5.683833e-05,
  6.694975e-06, 1.051937e-05, 1.016562e-05, 1.19637e-05, 1.819637e-05, 
    4.921907e-05, 4.623914e-05, 5.521131e-05, 6.007512e-05, 7.164105e-05, 
    8.404596e-05, 7.230008e-05, 7.858254e-05, 5.792803e-05, 3.889933e-05,
  2.963139e-06, 7.79334e-06, 1.327914e-05, 6.986094e-06, 4.85071e-06, 
    1.048878e-05, 2.349017e-05, 3.220979e-05, 3.646027e-05, 5.197715e-05, 
    6.573694e-05, 5.980986e-05, 6.176298e-05, 4.036687e-05, 4.180261e-05,
  3.298379e-05, 8.128586e-06, 1.080348e-05, 2.888662e-05, 3.69839e-06, 
    6.755803e-06, 2.45193e-05, 2.527583e-05, 5.480725e-05, 3.56215e-05, 
    4.47916e-05, 4.442913e-05, 6.546265e-05, 4.667327e-05, 3.70631e-05,
  2.566057e-05, 2.962861e-05, 4.245035e-05, 1.650379e-05, 8.022193e-06, 
    1.913962e-06, 3.539113e-06, 6.676986e-06, 1.306609e-05, 1.870574e-05, 
    3.974194e-05, 2.53338e-05, 4.291508e-05, 3.925918e-05, 3.730153e-05,
  2.335875e-05, 2.932732e-05, 3.74527e-05, 2.540217e-05, 2.951817e-05, 
    6.880033e-06, 3.668574e-06, 1.183537e-06, 1.751586e-06, 2.599219e-05, 
    2.711516e-05, 2.682343e-05, 3.992363e-05, 4.896844e-05, 4.454591e-05,
  7.187969e-06, 2.263677e-05, 3.545901e-05, 3.003607e-05, 3.777722e-05, 
    4.624748e-05, 6.514026e-06, 2.36066e-06, 1.659513e-06, 1.794429e-05, 
    2.46237e-05, 6.082847e-05, 6.53056e-05, 5.371673e-05, 3.932715e-05,
  1.072184e-14, 4.000246e-09, 1.774638e-07, 2.455055e-07, 5.288589e-09, 
    5.342899e-07, 8.417499e-07, 1.615463e-06, 1.430616e-06, 2.165204e-06, 
    2.229511e-06, 2.610036e-06, 3.086038e-06, 3.561471e-06, 4.945161e-06,
  3.436727e-12, 3.453621e-09, 6.543563e-08, 2.294705e-06, 3.489328e-07, 
    5.622726e-07, 2.829156e-07, 3.284101e-07, 6.302505e-07, 6.806376e-07, 
    1.593755e-06, 3.118574e-06, 2.979339e-06, 3.802701e-06, 4.038087e-06,
  1.386742e-11, 8.449602e-09, 6.412933e-08, 4.233937e-07, 1.180382e-07, 
    2.158282e-07, 2.235794e-07, 1.243385e-07, 1.675289e-07, 4.791368e-07, 
    6.474019e-07, 7.583392e-07, 1.630935e-06, 2.642958e-06, 3.043861e-06,
  5.44808e-11, 5.492976e-08, 3.57428e-07, 4.425789e-08, 6.814662e-09, 
    4.659005e-08, 1.604435e-07, 2.748329e-07, 2.518784e-07, 1.301298e-07, 
    2.316245e-07, 3.128426e-07, 1.130857e-06, 1.396066e-06, 1.186086e-06,
  1.42327e-09, 1.169979e-07, 2.575404e-08, 3.686215e-07, 6.484997e-07, 
    7.103915e-07, 6.748654e-09, 3.189672e-08, 1.686132e-07, 4.330673e-07, 
    5.482014e-08, 2.897994e-07, 6.577643e-07, 5.361657e-07, 9.290076e-07,
  9.610909e-07, 4.587354e-07, 1.377365e-07, 1.942791e-07, 1.072044e-07, 
    3.998826e-07, 1.4037e-07, 2.938633e-07, 6.92983e-07, 8.232681e-07, 
    1.941358e-06, 5.358583e-07, 1.101696e-06, 8.085569e-07, 4.706874e-07,
  8.37483e-07, 1.1538e-06, 2.913923e-06, 2.349013e-06, 6.261758e-07, 
    1.938436e-06, 1.655978e-06, 2.573034e-07, 9.130517e-08, 4.667662e-07, 
    7.954126e-07, 2.211895e-06, 1.859999e-06, 9.260747e-07, 7.705312e-07,
  3.379185e-07, 1.194456e-06, 7.028598e-06, 1.102221e-05, 1.873548e-06, 
    1.578865e-06, 1.34569e-06, 1.117747e-06, 3.160138e-07, 1.09888e-06, 
    1.342813e-06, 2.168591e-06, 2.77206e-06, 2.03596e-06, 1.89916e-06,
  9.822929e-07, 2.439698e-06, 1.833391e-06, 2.918908e-06, 8.642778e-06, 
    5.247083e-06, 1.119663e-06, 5.11745e-07, 7.313577e-07, 7.862107e-07, 
    1.751642e-06, 1.997564e-06, 1.650613e-06, 5.816496e-06, 2.578457e-05,
  6.236027e-07, 3.509727e-06, 1.074161e-05, 1.148628e-05, 5.748806e-06, 
    9.687463e-06, 2.25811e-06, 3.266231e-06, 3.533315e-06, 3.115143e-06, 
    3.70222e-06, 3.963096e-06, 6.733928e-06, 1.62339e-05, 4.06935e-05,
  1.589173e-07, 1.115381e-06, 5.034068e-06, 1.222113e-05, 8.058772e-06, 
    6.537827e-06, 4.214839e-06, 3.451263e-06, 3.041079e-06, 2.500392e-06, 
    7.704745e-07, 4.252479e-07, 1.190757e-08, 2.892001e-09, 1.62386e-09,
  7.419576e-06, 1.172686e-06, 6.18071e-06, 1.257946e-05, 9.117311e-06, 
    6.628371e-06, 5.758063e-06, 5.851478e-06, 5.482704e-06, 3.061218e-06, 
    8.065747e-07, 6.815836e-07, 7.834837e-08, 3.698927e-09, 4.209993e-10,
  9.553644e-06, 9.994103e-06, 2.043933e-06, 6.585278e-06, 9.636263e-06, 
    5.614584e-06, 3.606429e-06, 1.283001e-06, 2.261993e-06, 2.839015e-06, 
    2.003483e-06, 1.684267e-06, 7.081845e-08, 1.687073e-09, 1.017831e-09,
  1.351473e-05, 6.183448e-06, 3.670271e-06, 3.659694e-06, 4.415074e-06, 
    2.064347e-06, 9.668159e-07, 6.637582e-07, 4.444184e-07, 1.913108e-06, 
    2.287781e-06, 8.201272e-07, 5.124086e-07, 3.516162e-08, 5.70445e-09,
  3.718626e-05, 6.293031e-05, 1.502661e-06, 3.358334e-06, 2.245727e-06, 
    3.098548e-06, 1.760399e-06, 9.588814e-07, 7.64291e-07, 7.781791e-07, 
    1.093766e-06, 2.05304e-06, 2.566267e-06, 3.535901e-07, 1.805505e-07,
  4.700899e-05, 6.901372e-05, 5.542691e-05, 4.201566e-06, 1.549452e-06, 
    1.250344e-06, 1.43298e-06, 2.088457e-06, 1.265592e-06, 1.502162e-06, 
    2.310475e-06, 3.275888e-06, 2.575614e-06, 1.489488e-06, 6.251447e-07,
  5.18063e-05, 8.192467e-05, 7.484694e-05, 3.327571e-05, 3.302673e-06, 
    2.790944e-06, 3.635256e-06, 4.406659e-06, 3.228129e-06, 1.107862e-06, 
    1.856219e-06, 3.418465e-06, 3.653633e-06, 3.080598e-06, 9.938864e-07,
  6.219219e-05, 8.631217e-05, 7.475688e-05, 4.383942e-05, 1.795326e-06, 
    6.025244e-06, 5.411731e-06, 4.28944e-06, 5.537154e-06, 4.276236e-06, 
    2.189438e-06, 1.838686e-06, 5.830197e-06, 7.284063e-06, 7.188339e-06,
  6.050175e-05, 0.0001417966, 0.0001341182, 0.0001025213, 5.956084e-05, 
    5.193415e-06, 2.688431e-06, 2.209594e-06, 2.102024e-06, 3.150396e-06, 
    2.867432e-06, 4.562658e-06, 5.124582e-06, 5.934509e-06, 1.119934e-05,
  0.0001095497, 0.000204886, 0.0001380449, 0.0001860468, 0.0001050814, 
    2.305481e-05, 7.291366e-06, 3.662078e-06, 1.062552e-06, 2.393597e-06, 
    3.609525e-06, 3.167895e-06, 3.139714e-06, 5.454913e-06, 1.229188e-05,
  7.006117e-06, 5.318039e-06, 3.403001e-05, 0.0001349576, 7.300775e-05, 
    0.0001202518, 0.0001863468, 0.0002944951, 0.0003769476, 0.0004058782, 
    0.0003505463, 0.0002505442, 0.0001454283, 0.0001050042, 8.313239e-05,
  1.815397e-05, 9.149726e-06, 8.934559e-06, 0.0001570543, 3.090245e-05, 
    6.216377e-05, 8.78952e-05, 0.0001306678, 0.0002276922, 0.000314249, 
    0.0003688191, 0.0003481688, 0.0002458167, 0.0001690585, 0.0001142496,
  1.913312e-05, 4.015139e-05, 1.096229e-05, 2.563432e-05, 9.935522e-05, 
    3.593284e-05, 5.58902e-05, 5.685387e-05, 5.036973e-05, 5.845284e-05, 
    0.0001170603, 0.0001844674, 0.0001603818, 0.0001148205, 7.017583e-05,
  1.90999e-05, 2.398486e-05, 1.217806e-05, 1.239005e-05, 4.026546e-05, 
    3.757037e-05, 5.258058e-05, 4.35644e-05, 3.510665e-05, 1.462544e-05, 
    1.164014e-05, 1.882297e-05, 2.251716e-05, 3.360309e-05, 4.987261e-05,
  2.73766e-05, 5.839532e-05, 2.730956e-05, 1.360277e-05, 2.397723e-05, 
    5.573489e-05, 4.254665e-05, 3.816202e-05, 3.477025e-05, 2.514085e-05, 
    1.560274e-05, 1.073761e-05, 1.088859e-05, 2.326826e-05, 2.702983e-05,
  7.264419e-05, 0.0001006657, 0.0001129657, 1.375434e-06, 6.527973e-06, 
    1.764452e-05, 1.651183e-05, 2.914934e-05, 2.570278e-05, 1.232793e-05, 
    5.843571e-06, 7.803564e-06, 1.366367e-05, 2.004995e-05, 2.193956e-05,
  0.0001183259, 0.0001780975, 0.0002318772, 0.0001970626, 1.357604e-05, 
    1.348423e-05, 6.269397e-06, 3.398639e-06, 9.109988e-07, 3.563053e-06, 
    4.071379e-06, 1.062887e-05, 1.050912e-05, 1.435837e-05, 2.961982e-05,
  0.0002314064, 0.0003789589, 0.0005198476, 0.0004274711, 1.160897e-05, 
    7.997533e-06, 1.01831e-06, 2.016934e-07, 6.106961e-07, 1.471495e-06, 
    4.673247e-06, 6.323319e-06, 9.747583e-06, 1.130339e-05, 3.797453e-05,
  0.0003114355, 0.0004284355, 0.0004808664, 0.0003276594, 0.000161572, 
    2.996133e-06, 1.483235e-06, 1.796874e-07, 2.736487e-07, 9.751759e-07, 
    5.319552e-06, 5.870736e-06, 6.775375e-06, 8.582459e-06, 2.792049e-05,
  0.0003619132, 0.0003423049, 0.0003411974, 0.000223873, 0.0001848039, 
    0.0001681423, 7.70567e-07, 9.721686e-07, 3.021396e-07, 1.579225e-06, 
    3.722788e-06, 2.886014e-06, 4.039589e-06, 8.372638e-06, 2.859732e-05,
  2.513358e-06, 3.530518e-06, 2.389868e-06, 2.048121e-06, 1.510268e-06, 
    2.43153e-06, 3.33783e-06, 2.585049e-06, 6.45253e-06, 4.660712e-06, 
    3.603532e-06, 6.00339e-06, 1.148764e-05, 1.459177e-05, 1.367052e-05,
  7.571016e-06, 2.411611e-06, 3.193851e-06, 1.841691e-06, 6.67338e-07, 
    2.900422e-07, 9.84105e-07, 3.041182e-06, 4.534443e-06, 3.356522e-06, 
    6.860293e-06, 3.831597e-05, 7.137108e-05, 8.661105e-05, 0.0001459077,
  7.165479e-06, 6.792642e-06, 1.00346e-05, 4.007667e-06, 2.492385e-06, 
    1.023502e-06, 2.785613e-06, 5.379303e-06, 1.07178e-05, 2.132503e-05, 
    4.779776e-05, 0.0001029429, 0.0001818314, 0.0002691108, 0.0003194575,
  4.13826e-05, 7.806993e-05, 0.0001004306, 5.599896e-05, 1.092577e-05, 
    3.800352e-06, 7.87431e-06, 1.476143e-05, 2.04164e-05, 3.592926e-05, 
    3.213006e-05, 4.193596e-05, 0.0001696093, 0.0003033816, 0.0002557669,
  0.0003643893, 0.0004660275, 0.0003841523, 0.0002182568, 5.867469e-05, 
    7.296973e-06, 1.28585e-05, 8.447464e-05, 0.0002899959, 0.0005292244, 
    0.0007370125, 0.0009260366, 0.001089253, 0.001144247, 0.0009558888,
  0.0008995585, 0.0009228542, 0.0007883689, 0.0005283033, 0.000282732, 
    0.0001503181, 0.0001776736, 0.0003566916, 0.0005764879, 0.0007523234, 
    0.0008233148, 0.0008537115, 0.0009064269, 0.0009075738, 0.0009490813,
  0.0009177942, 0.0008191693, 0.0006239332, 0.0004455002, 0.0002193189, 
    9.704437e-05, 0.0001017641, 0.0001278777, 0.0001223445, 8.663631e-05, 
    5.899282e-05, 6.863097e-05, 9.228213e-05, 0.0002013456, 0.00033581,
  0.0006596156, 0.0006093156, 0.000312295, 0.0002798088, 9.856755e-05, 
    1.096937e-05, 1.904106e-05, 1.696172e-05, 7.879627e-06, 3.038797e-06, 
    6.314561e-06, 8.812523e-06, 9.680535e-06, 8.872665e-06, 1.194103e-05,
  0.000581739, 0.0003088805, 0.0002673046, 0.0003446855, 0.0002516524, 
    1.943897e-05, 2.57889e-05, 2.463615e-05, 8.738794e-06, 8.189312e-07, 
    8.540127e-07, 1.598188e-06, 1.035123e-06, 1.740399e-06, 2.69354e-06,
  0.0002705198, 0.0001976895, 0.0001903194, 0.0001633744, 0.0001627152, 
    0.0001837434, 2.805754e-05, 2.71289e-05, 8.407262e-06, 1.400277e-06, 
    2.374148e-07, 9.738635e-08, 1.980886e-07, 3.146074e-07, 5.25034e-06,
  3.392071e-07, 4.616826e-08, 2.956647e-08, 2.159847e-07, 7.412391e-07, 
    6.74059e-07, 5.840302e-07, 3.221437e-07, 1.410957e-06, 1.203024e-06, 
    2.360169e-06, 6.271918e-07, 8.701714e-07, 1.138192e-06, 1.722738e-06,
  1.789264e-06, 5.350282e-07, 3.983607e-06, 4.426639e-06, 2.286409e-06, 
    5.509009e-06, 7.838947e-06, 2.710909e-05, 2.634644e-05, 3.199448e-05, 
    4.1897e-05, 4.086982e-05, 5.780247e-05, 5.063802e-05, 7.270605e-05,
  6.250767e-07, 1.108167e-06, 6.842156e-06, 2.377771e-05, 5.648481e-05, 
    9.063278e-05, 0.0001214101, 0.0001520003, 0.0001962587, 0.0002206594, 
    0.0002441492, 0.0002371504, 0.0002323831, 0.0002182055, 0.0001953209,
  1.885689e-06, 7.992159e-06, 1.946487e-05, 9.572016e-05, 0.0001675798, 
    0.0001998354, 0.0002589234, 0.0002950168, 0.00032971, 0.0003547832, 
    0.0003589626, 0.0003503417, 0.0003187162, 0.0003258098, 0.0003347661,
  1.053828e-05, 3.009303e-05, 8.633023e-05, 0.0002152301, 0.0003572968, 
    0.0005009947, 0.0005676276, 0.0006380178, 0.0007092619, 0.0007827724, 
    0.0007933237, 0.0007623813, 0.0007374636, 0.0007750383, 0.000863366,
  1.595771e-05, 4.029596e-05, 0.00018433, 0.0003693899, 0.0005652652, 
    0.000668156, 0.000700577, 0.0007114925, 0.0007438639, 0.0007666954, 
    0.0007838199, 0.0007636498, 0.0007470916, 0.0007997868, 0.0008829256,
  1.46045e-05, 3.151052e-05, 0.0001326979, 0.0002822154, 0.0003823719, 
    0.0004054081, 0.0003480983, 0.0003165267, 0.000295736, 0.0002611627, 
    0.0002544532, 0.000266584, 0.0003038814, 0.000353907, 0.0003473182,
  1.523481e-05, 2.854749e-05, 3.937065e-05, 0.0001081558, 6.291449e-05, 
    3.853356e-05, 4.608477e-05, 5.928466e-05, 6.204663e-05, 5.830741e-05, 
    5.98993e-05, 7.289898e-05, 0.0001475192, 0.0001954245, 0.0001680384,
  2.958677e-05, 4.716442e-05, 4.036634e-05, 4.413874e-05, 3.910834e-05, 
    1.707968e-05, 1.507512e-05, 3.395027e-05, 5.544069e-05, 5.253452e-05, 
    6.206133e-05, 0.0001705441, 0.0002589283, 0.0002401012, 0.0001401739,
  6.901066e-05, 9.415617e-05, 8.826197e-05, 0.0001250184, 8.311658e-05, 
    4.310455e-05, 1.622342e-05, 2.759493e-05, 3.552144e-05, 6.820871e-05, 
    0.0001980452, 0.0002852457, 0.0003065777, 0.0001751328, 5.432052e-05,
  9.885639e-26, 8.855201e-26, 6.793632e-26, 5.124128e-11, 8.501155e-09, 
    7.02228e-08, 2.404526e-07, 2.206708e-06, 1.3586e-06, 2.446568e-06, 
    2.424137e-06, 2.518635e-06, 2.257856e-06, 2.599544e-06, 3.869456e-06,
  8.777834e-26, 5.007406e-26, 2.125133e-18, 2.056722e-18, 3.844528e-11, 
    6.829306e-11, 9.232184e-09, 3.303698e-09, 8.256198e-08, 7.32766e-07, 
    2.996991e-07, 1.046461e-06, 1.501557e-06, 2.691102e-06, 4.252966e-06,
  4.029808e-26, 3.498955e-26, 3.973063e-15, 2.496967e-20, 1.624224e-26, 
    1.628522e-11, 8.607855e-11, 3.500655e-11, 8.472014e-09, 1.944812e-09, 
    1.224529e-09, 1.325246e-08, 7.713182e-09, 4.782561e-07, 1.174274e-06,
  6.663661e-11, 2.35717e-16, 1.920287e-14, 4.146492e-13, 9.467795e-13, 
    1.754855e-13, 2.742816e-14, 1.093777e-12, 6.814957e-11, 1.394628e-10, 
    6.835676e-11, 7.030361e-10, 6.169623e-10, 4.123017e-10, 7.343295e-10,
  1.591622e-10, 1.265398e-10, 2.028398e-13, 9.633472e-13, 1.495615e-12, 
    2.046732e-11, 1.575488e-11, 3.970015e-10, 2.116581e-08, 2.70203e-11, 
    4.310185e-10, 3.302664e-09, 8.329206e-08, 2.616671e-08, 1.411997e-07,
  7.036662e-12, 1.780159e-11, 5.747535e-08, 5.361525e-10, 8.017894e-12, 
    3.242249e-12, 1.722515e-09, 1.528176e-08, 5.861089e-08, 1.620054e-08, 
    2.93098e-07, 9.408141e-07, 2.169003e-07, 5.069664e-07, 1.315378e-06,
  1.368139e-12, 4.580003e-11, 5.259155e-08, 6.569218e-08, 2.400793e-09, 
    3.233942e-07, 4.676152e-07, 1.616812e-07, 3.217911e-07, 9.908831e-08, 
    1.250183e-06, 3.420388e-06, 4.310417e-06, 3.00067e-06, 1.844258e-06,
  7.08165e-09, 1.282944e-07, 1.194642e-07, 5.384937e-07, 1.135321e-06, 
    5.413519e-07, 5.81896e-07, 7.657763e-07, 1.147305e-06, 1.391983e-06, 
    1.433624e-06, 7.481925e-06, 9.949925e-06, 6.73074e-06, 7.591525e-06,
  1.325263e-07, 3.245169e-07, 9.512268e-07, 1.953678e-06, 3.536956e-06, 
    2.544271e-06, 3.387724e-06, 3.399681e-06, 4.113628e-06, 5.486484e-06, 
    5.926096e-06, 6.408029e-06, 1.11659e-05, 1.303808e-05, 8.818044e-06,
  3.414182e-08, 2.972934e-07, 2.747835e-06, 9.936773e-06, 7.820597e-06, 
    8.35804e-06, 4.709043e-06, 5.541644e-06, 6.859653e-06, 8.499971e-06, 
    9.604166e-06, 8.813859e-06, 6.335212e-06, 2.556802e-06, 2.961621e-06,
  1.108673e-25, 2.81432e-11, 4.730808e-11, 2.040717e-11, 1.077261e-11, 
    6.943034e-12, 2.113419e-11, 1.388629e-10, 3.845769e-07, 8.851098e-07, 
    1.419735e-06, 1.21352e-06, 7.422609e-07, 6.165975e-07, 3.263197e-07,
  1.410508e-26, 1.261486e-12, 1.821371e-12, 2.57515e-12, 2.180752e-11, 
    7.686891e-11, 4.103694e-11, 3.663876e-10, 4.274148e-08, 3.379168e-07, 
    3.152877e-07, 1.856732e-07, 1.395228e-06, 1.088009e-06, 1.527874e-06,
  1.192029e-26, 2.903674e-26, 3.803831e-26, 5.120163e-26, 1.101364e-25, 
    3.437112e-25, 1.094269e-12, 9.19089e-12, 6.297127e-11, 1.795896e-11, 
    4.41981e-11, 1.081826e-09, 1.174191e-08, 4.645001e-07, 5.589074e-07,
  8.852464e-27, 9.847912e-27, 6.533117e-27, 1.778275e-27, 4.753814e-27, 
    1.179037e-26, 3.802347e-26, 1.8197e-25, 2.452866e-11, 2.943192e-11, 
    1.41591e-11, 1.320823e-11, 5.863588e-12, 1.939182e-10, 5.17026e-10,
  3.022937e-27, 2.774513e-27, 1.621248e-19, 4.469577e-20, 2.653387e-34, 
    1.826643e-33, 3.411951e-28, 1.682715e-27, 1.292831e-27, 1.275439e-12, 
    1.734444e-12, 1.716398e-19, 1.413265e-27, 1.675043e-17, 5.278416e-15,
  4.598873e-14, 1.204494e-12, 1.52496e-08, 9.619578e-13, 0, 1.135967e-30, 
    2.782682e-29, 1.737154e-33, 2.889751e-33, 0, 2.263563e-29, 0, 0, 0, 
    1.710305e-15,
  1.654348e-11, 2.239931e-08, 5.029548e-08, 1.734546e-08, 2.068537e-12, 
    7.731447e-12, 2.794685e-11, 1.341118e-15, 2.813053e-28, 1.523702e-28, 0, 
    0, 0, 8.551659e-23, 3.414661e-14,
  9.917348e-08, 1.740364e-09, 6.803905e-08, 1.39652e-07, 6.343063e-08, 
    1.004782e-08, 1.418117e-09, 1.243929e-10, 3.881724e-11, 1.881832e-10, 
    1.203676e-12, 2.230904e-12, 1.651055e-13, 1.071267e-12, 4.147608e-11,
  3.996002e-06, 4.571412e-09, 1.665604e-13, 3.547289e-08, 2.358598e-07, 
    3.193546e-08, 4.84195e-09, 9.535182e-08, 5.935189e-08, 2.527232e-07, 
    5.02174e-08, 8.019494e-08, 1.736404e-08, 8.098319e-10, 8.067433e-10,
  7.000384e-06, 4.139594e-06, 2.078699e-09, 2.196252e-10, 5.467211e-08, 
    1.306842e-07, 7.949264e-08, 7.827904e-08, 8.142174e-08, 8.910799e-08, 
    1.989127e-07, 2.890372e-07, 9.212947e-08, 2.679824e-07, 5.240482e-08,
  5.689761e-05, 5.823934e-05, 4.627465e-05, 3.25433e-05, 2.118044e-05, 
    2.639026e-05, 1.931103e-05, 2.267266e-05, 2.872258e-05, 8.324389e-06, 
    5.639698e-06, 1.844067e-06, 2.597528e-06, 8.54872e-06, 1.547042e-06,
  1.784892e-05, 2.325638e-05, 2.525237e-05, 2.165624e-05, 1.46975e-05, 
    1.034907e-05, 4.902583e-06, 3.698544e-06, 3.14786e-06, 1.692691e-06, 
    1.054398e-06, 1.539915e-06, 3.741189e-06, 5.63978e-06, 7.890312e-06,
  2.263621e-06, 5.135446e-06, 3.399563e-06, 5.492032e-06, 5.605052e-06, 
    5.57711e-06, 5.911899e-06, 6.922657e-06, 7.544591e-06, 4.929156e-06, 
    6.215424e-06, 7.905769e-06, 7.834478e-06, 8.365326e-06, 4.961211e-06,
  6.904196e-06, 7.199104e-06, 5.477979e-06, 5.558906e-06, 6.052963e-06, 
    7.144198e-06, 7.703599e-06, 9.226414e-06, 8.651919e-06, 1.19995e-05, 
    8.863844e-06, 7.198231e-06, 3.883079e-06, 1.534305e-06, 5.576806e-08,
  8.443243e-06, 9.307591e-06, 4.83022e-06, 2.705335e-06, 3.049514e-06, 
    5.129399e-06, 7.945198e-06, 7.028747e-06, 7.574259e-06, 6.837184e-06, 
    4.241857e-06, 2.232239e-06, 7.067071e-07, 2.892062e-07, 8.362541e-07,
  3.630023e-06, 7.345066e-06, 1.973366e-06, 1.187155e-06, 2.00193e-06, 
    3.488811e-06, 3.841059e-06, 3.905621e-06, 5.808815e-06, 3.609619e-06, 
    1.657903e-06, 8.908671e-07, 2.037249e-06, 8.217818e-06, 3.094428e-05,
  4.301361e-07, 9.313099e-07, 4.108293e-07, 1.052246e-06, 1.702897e-06, 
    2.109746e-06, 4.146339e-06, 5.469181e-06, 5.830279e-06, 2.880856e-06, 
    4.012025e-06, 3.130552e-06, 1.212653e-05, 3.227976e-05, 4.114299e-05,
  3.314573e-06, 2.65098e-06, 1.49076e-06, 1.802507e-06, 2.289139e-06, 
    1.082446e-06, 2.723783e-06, 4.070409e-06, 6.520384e-06, 3.754379e-06, 
    4.643997e-06, 7.517529e-06, 3.066925e-05, 2.562435e-05, 1.747777e-05,
  8.249822e-06, 7.261909e-06, 7.48927e-06, 1.002523e-05, 7.668672e-06, 
    2.002491e-06, 2.008715e-06, 3.134498e-06, 6.619027e-06, 5.577016e-06, 
    5.846122e-06, 1.950495e-05, 3.411631e-05, 1.509732e-05, 1.604137e-05,
  1.547647e-05, 8.900358e-06, 2.330747e-05, 1.838984e-05, 2.514793e-05, 
    3.105972e-05, 1.517954e-08, 1.932156e-06, 6.41315e-06, 1.183336e-05, 
    2.578859e-05, 4.319299e-05, 4.101714e-05, 5.407539e-05, 5.45421e-05,
  5.20458e-10, 2.302512e-10, 1.651802e-06, 5.384939e-06, 4.427946e-06, 
    7.60353e-06, 7.059115e-06, 6.449525e-06, 5.951667e-06, 6.379556e-06, 
    6.566427e-06, 5.686896e-06, 4.353194e-06, 5.39025e-06, 1.098948e-05,
  7.917048e-09, 9.445764e-08, 1.527433e-06, 3.954868e-06, 5.36639e-06, 
    6.558766e-06, 6.790145e-06, 6.566372e-06, 5.703909e-06, 5.022298e-06, 
    4.58612e-06, 4.605776e-06, 5.524644e-06, 7.020161e-06, 8.278029e-06,
  2.850208e-09, 2.100571e-08, 1.674207e-06, 2.76662e-06, 3.893039e-06, 
    6.591666e-06, 4.916431e-06, 6.453294e-06, 6.658923e-06, 5.148054e-06, 
    3.998829e-06, 3.604343e-06, 3.080236e-06, 3.90783e-06, 1.035702e-05,
  5.182571e-08, 3.220305e-08, 7.367541e-07, 3.453337e-06, 4.714248e-06, 
    1.883126e-06, 2.477007e-06, 4.866985e-06, 6.198865e-06, 7.250444e-06, 
    6.136992e-06, 6.075079e-06, 6.863208e-06, 1.127181e-05, 1.120628e-05,
  4.720398e-06, 2.651836e-06, 3.225458e-06, 7.270466e-06, 9.429283e-06, 
    9.601985e-06, 6.372145e-06, 9.297494e-06, 1.853287e-05, 3.648926e-05, 
    2.499708e-05, 1.703147e-05, 1.839111e-05, 1.345509e-05, 1.062267e-05,
  1.042742e-05, 7.71358e-06, 3.756001e-06, 7.18868e-06, 1.08928e-05, 
    1.591087e-05, 2.059062e-05, 1.233201e-05, 1.78375e-05, 1.924897e-05, 
    3.528423e-05, 3.414665e-05, 2.090613e-05, 2.143258e-05, 2.019584e-05,
  5.552727e-06, 1.019507e-05, 1.331941e-05, 8.326007e-06, 4.422792e-06, 
    6.041483e-06, 8.38981e-06, 7.47595e-06, 9.658741e-06, 1.712197e-05, 
    2.3516e-05, 2.586722e-05, 1.726416e-05, 2.284182e-05, 3.621548e-05,
  7.649766e-06, 7.437877e-06, 7.2133e-06, 1.504648e-05, 8.582358e-06, 
    2.738058e-06, 4.279082e-06, 7.803936e-06, 1.118583e-05, 1.143936e-05, 
    1.153776e-05, 1.134506e-05, 2.024267e-05, 2.161689e-05, 3.105173e-05,
  1.207221e-05, 8.983397e-06, 7.07098e-06, 7.00308e-06, 1.525092e-05, 
    9.221998e-06, 5.460582e-06, 5.922244e-06, 9.500724e-06, 8.520315e-06, 
    6.064626e-06, 7.628842e-06, 1.723552e-05, 2.95572e-05, 2.527989e-05,
  7.551715e-06, 1.033285e-05, 6.691169e-06, 6.384974e-06, 8.585685e-06, 
    1.690526e-05, 5.392051e-06, 9.874988e-06, 1.472215e-05, 1.008434e-05, 
    8.109992e-06, 6.781434e-06, 9.783253e-06, 1.168292e-05, 3.010615e-05,
  5.590107e-12, 3.862901e-10, 2.231402e-07, 2.443631e-06, 2.897672e-06, 
    3.017247e-06, 3.834492e-06, 2.658064e-06, 2.450857e-06, 3.255182e-06, 
    5.215807e-06, 4.449069e-06, 4.206732e-06, 5.044914e-06, 5.381247e-06,
  6.439665e-09, 6.121144e-09, 5.665566e-08, 1.536387e-06, 2.405814e-06, 
    3.591991e-06, 4.440136e-06, 3.311482e-06, 3.440686e-06, 4.516896e-06, 
    5.160701e-06, 5.791975e-06, 4.074429e-06, 4.48449e-06, 6.696428e-06,
  1.148624e-08, 7.014447e-08, 1.006119e-06, 2.876353e-06, 2.981437e-06, 
    3.327632e-06, 4.601638e-06, 3.77585e-06, 2.865822e-06, 3.582733e-06, 
    4.425156e-06, 4.951471e-06, 4.055548e-06, 4.192912e-06, 6.297414e-06,
  1.831982e-08, 1.001728e-07, 1.409041e-08, 9.311336e-07, 2.021801e-06, 
    3.039062e-06, 3.259612e-06, 3.176013e-06, 2.742041e-06, 2.54914e-06, 
    3.390398e-06, 3.641049e-06, 3.585147e-06, 4.40374e-06, 6.45253e-06,
  1.56706e-11, 7.827055e-08, 3.20736e-07, 7.450203e-07, 1.724672e-06, 
    4.183467e-06, 4.368727e-06, 3.675156e-06, 2.757913e-06, 3.390812e-06, 
    3.738646e-06, 3.509795e-06, 3.832796e-06, 6.16721e-06, 8.583166e-06,
  5.185561e-10, 4.16821e-08, 4.738695e-07, 1.442581e-06, 1.741799e-06, 
    5.256708e-06, 6.000835e-06, 4.717854e-06, 3.894554e-06, 2.960951e-06, 
    3.26222e-06, 3.70565e-06, 3.11017e-06, 5.791172e-06, 9.234998e-06,
  4.415499e-09, 4.882054e-08, 6.466993e-07, 7.46216e-07, 1.716185e-06, 
    3.253087e-06, 5.314765e-06, 4.999903e-06, 5.02926e-06, 3.964656e-06, 
    3.952437e-06, 5.187151e-06, 8.435777e-06, 8.241496e-06, 1.02748e-05,
  1.567025e-08, 3.972363e-07, 3.999698e-07, 4.12857e-06, 5.592981e-07, 
    1.090023e-06, 3.238739e-06, 4.024364e-06, 5.79159e-06, 6.947443e-06, 
    8.158087e-06, 1.269881e-05, 1.710766e-05, 1.43306e-05, 1.289601e-05,
  1.038493e-05, 3.742981e-06, 3.135105e-06, 1.172883e-06, 5.00299e-06, 
    1.008678e-06, 2.198715e-06, 3.715854e-06, 5.742507e-06, 8.945352e-06, 
    1.381844e-05, 1.740438e-05, 1.883767e-05, 1.506433e-05, 1.095788e-05,
  8.803817e-06, 1.142164e-05, 7.68376e-06, 5.286673e-06, 4.635073e-06, 
    4.961228e-06, 7.333431e-07, 2.326003e-06, 5.63764e-06, 1.02752e-05, 
    1.402118e-05, 1.669642e-05, 2.342801e-05, 1.645198e-05, 7.877081e-06,
  6.249765e-11, 7.294028e-14, 5.822393e-11, 6.058074e-12, 1.554147e-11, 
    3.56269e-11, 1.013796e-10, 1.305621e-08, 3.609166e-08, 1.169539e-07, 
    1.992643e-07, 5.103435e-07, 3.639606e-07, 7.891072e-07, 7.792839e-07,
  4.733595e-13, 1.05507e-17, 4.508979e-19, 2.985344e-12, 1.310815e-13, 
    7.510981e-11, 1.264664e-09, 1.306844e-07, 6.669779e-08, 6.391406e-08, 
    1.284059e-07, 1.832001e-07, 1.978555e-07, 1.688821e-07, 2.612535e-07,
  4.589874e-11, 3.696563e-08, 1.364725e-12, 5.118908e-10, 4.310313e-10, 
    7.968197e-08, 3.628788e-07, 4.534129e-07, 2.110056e-07, 5.603941e-08, 
    1.346452e-07, 1.783644e-07, 4.979128e-08, 1.44688e-07, 2.322001e-07,
  1.088716e-07, 7.350559e-08, 1.245752e-08, 9.876026e-10, 7.892294e-08, 
    2.758373e-07, 3.813927e-07, 3.296431e-07, 2.200214e-07, 3.533654e-07, 
    4.615188e-07, 5.1327e-07, 9.277368e-08, 7.323563e-07, 8.580469e-07,
  3.476648e-07, 8.22869e-07, 7.79594e-07, 6.2372e-07, 1.020118e-06, 
    4.35107e-07, 2.713135e-07, 1.74231e-07, 2.60217e-07, 6.241648e-07, 
    1.145858e-06, 9.086687e-07, 1.120029e-06, 1.107882e-06, 1.65055e-06,
  5.528369e-07, 8.015303e-07, 1.53856e-06, 1.793157e-06, 1.297942e-06, 
    1.081889e-06, 3.274602e-07, 2.043301e-07, 2.86504e-07, 7.013997e-07, 
    1.543012e-06, 1.192188e-06, 1.207167e-06, 1.669738e-06, 2.361087e-06,
  2.103881e-06, 1.287222e-06, 4.007443e-06, 4.100507e-06, 3.602789e-06, 
    1.927137e-06, 7.80348e-07, 4.193714e-07, 7.911705e-07, 1.308244e-06, 
    1.376902e-06, 1.518172e-06, 1.718448e-06, 2.404657e-06, 3.748615e-06,
  3.696142e-06, 3.693144e-06, 4.452111e-06, 7.529453e-06, 4.429717e-06, 
    3.746754e-06, 2.53511e-06, 1.336638e-06, 1.48841e-06, 1.673156e-06, 
    1.801044e-06, 2.244911e-06, 2.47704e-06, 3.325127e-06, 4.352989e-06,
  1.157476e-05, 5.330643e-06, 5.146431e-06, 5.167485e-06, 8.474435e-06, 
    7.439137e-06, 5.561683e-06, 3.575942e-06, 2.915972e-06, 2.392802e-06, 
    2.464689e-06, 3.226432e-06, 4.31933e-06, 5.603214e-06, 5.525232e-06,
  2.765574e-05, 1.313261e-05, 7.066865e-06, 7.506909e-06, 6.432434e-06, 
    1.036977e-05, 9.441014e-06, 4.168086e-06, 4.684341e-06, 4.511476e-06, 
    5.003777e-06, 6.215958e-06, 7.202219e-06, 9.31968e-06, 7.93107e-06,
  6.61791e-15, 5.803523e-13, 1.142328e-11, 4.391869e-09, 2.991549e-11, 
    1.44608e-11, 1.489383e-11, 4.514061e-09, 4.499846e-07, 8.427945e-07, 
    3.026361e-06, 3.305443e-06, 3.197167e-06, 6.593747e-06, 2.036765e-05,
  1.122599e-18, 7.927645e-10, 1.367001e-08, 4.534307e-08, 1.054038e-08, 
    3.027362e-09, 2.852668e-12, 4.223651e-13, 8.933791e-08, 1.40534e-07, 
    6.799645e-08, 3.492706e-07, 5.346308e-07, 2.290594e-06, 5.506022e-06,
  3.040489e-12, 1.297178e-08, 2.512599e-07, 2.744593e-07, 6.767551e-08, 
    5.962129e-08, 1.204387e-09, 2.740989e-09, 2.386941e-10, 2.544247e-08, 
    3.898448e-08, 3.733804e-08, 1.63354e-07, 9.683945e-07, 1.746343e-06,
  4.631156e-08, 1.117967e-08, 6.37994e-08, 6.484311e-07, 1.802813e-07, 
    4.888041e-07, 9.238065e-08, 1.352482e-07, 5.395382e-08, 1.25166e-07, 
    3.330403e-08, 2.137802e-08, 9.639337e-11, 1.311145e-09, 1.867283e-08,
  5.027035e-07, 1.475219e-07, 1.192192e-08, 9.031624e-08, 3.243725e-07, 
    1.297087e-06, 6.90303e-07, 8.808352e-07, 5.644245e-07, 3.422139e-07, 
    1.924493e-07, 2.869741e-08, 2.125123e-09, 2.793943e-09, 1.558417e-09,
  2.682828e-06, 1.976627e-06, 1.47026e-06, 3.433924e-07, 6.643738e-07, 
    1.256154e-07, 4.295059e-07, 1.957386e-07, 5.06141e-08, 1.904749e-07, 
    6.739979e-07, 2.703889e-07, 2.99767e-08, 5.680369e-08, 6.111504e-08,
  7.465955e-06, 3.795271e-06, 4.942913e-06, 4.623444e-06, 2.448934e-06, 
    2.15251e-06, 5.279048e-07, 3.210948e-07, 4.015774e-07, 1.507369e-06, 
    1.02774e-06, 1.834263e-06, 1.72231e-06, 6.383493e-07, 9.011271e-08,
  1.203289e-05, 7.033521e-06, 5.089189e-06, 7.07012e-06, 4.256333e-06, 
    4.493834e-06, 2.697931e-06, 1.998741e-06, 3.456161e-06, 3.221818e-07, 
    3.14658e-06, 3.345318e-06, 3.742369e-06, 2.283285e-06, 3.160219e-06,
  1.15732e-05, 7.257061e-06, 3.636195e-06, 4.163172e-06, 6.073772e-06, 
    6.802962e-06, 9.381982e-06, 5.860693e-06, 4.084795e-06, 2.366749e-06, 
    2.680418e-06, 3.51306e-06, 4.391353e-06, 3.659174e-06, 3.258962e-06,
  1.309552e-05, 4.483651e-06, 4.420178e-06, 3.178765e-06, 1.845318e-06, 
    7.065681e-06, 1.199722e-05, 1.015865e-05, 9.813363e-06, 7.091073e-06, 
    5.91398e-06, 5.322079e-06, 5.029087e-06, 6.813641e-06, 7.55651e-06,
  6.371522e-08, 7.120987e-07, 1.596614e-06, 2.925363e-07, 6.121792e-08, 
    1.188471e-09, 1.250182e-11, 1.082256e-10, 6.760467e-07, 1.578359e-06, 
    1.090265e-06, 9.707478e-07, 4.495991e-07, 1.197253e-07, 1.194347e-07,
  3.909039e-07, 1.024688e-07, 1.088411e-06, 9.431306e-07, 2.089761e-07, 
    2.844804e-08, 2.10298e-09, 2.208221e-10, 1.241865e-08, 4.148474e-07, 
    1.244456e-06, 1.874219e-06, 1.751301e-06, 1.79719e-06, 1.940662e-06,
  2.068904e-06, 4.017288e-06, 2.627368e-06, 2.277019e-06, 3.521455e-06, 
    1.357778e-06, 5.683187e-08, 2.560917e-08, 3.802242e-08, 1.207971e-07, 
    2.375355e-08, 4.839301e-07, 1.726162e-06, 3.061271e-06, 4.120311e-06,
  3.793425e-06, 4.158042e-06, 3.511532e-06, 3.543036e-06, 2.145954e-06, 
    1.796398e-06, 1.736302e-06, 4.452016e-07, 4.287146e-08, 2.959303e-08, 
    1.893894e-08, 6.684308e-10, 1.056302e-08, 5.605852e-07, 1.677629e-06,
  2.570619e-06, 4.352531e-06, 5.114827e-06, 4.195179e-06, 3.214227e-06, 
    4.207518e-06, 2.743412e-06, 1.437014e-06, 5.599825e-07, 3.510665e-08, 
    6.293952e-08, 1.370242e-09, 6.424746e-10, 5.149875e-09, 7.047137e-09,
  1.581874e-06, 3.784472e-06, 6.143941e-06, 3.891749e-06, 6.534008e-06, 
    5.544291e-06, 2.309617e-06, 1.366124e-06, 1.77303e-06, 1.136425e-06, 
    2.137929e-07, 2.235079e-08, 2.761953e-09, 1.261358e-09, 1.675222e-09,
  8.88738e-07, 2.738682e-06, 9.073198e-06, 9.226087e-06, 8.296854e-06, 
    5.204723e-06, 5.763125e-06, 2.124985e-06, 3.007893e-06, 1.750425e-06, 
    1.90588e-06, 7.331481e-07, 2.474101e-07, 3.532771e-08, 1.626078e-08,
  2.555261e-07, 1.813406e-06, 4.227071e-06, 1.091064e-05, 6.27818e-06, 
    7.296246e-06, 9.119208e-06, 7.126515e-06, 7.053807e-06, 4.223811e-06, 
    4.251818e-06, 4.433011e-06, 3.159649e-06, 3.059145e-06, 3.016312e-06,
  4.123825e-07, 7.63035e-07, 1.551544e-06, 5.149539e-06, 1.141572e-05, 
    9.544172e-06, 9.836472e-06, 9.972478e-06, 7.939309e-06, 8.109975e-06, 
    7.120773e-06, 4.41255e-06, 3.881381e-06, 3.065695e-06, 3.37409e-06,
  1.238467e-07, 2.179922e-07, 6.192865e-07, 3.912153e-06, 5.14362e-06, 
    1.229548e-05, 1.15733e-05, 9.023471e-06, 1.028103e-05, 1.000444e-05, 
    1.051596e-05, 8.506479e-06, 8.462835e-06, 6.293133e-06, 5.626927e-06,
  3.78488e-09, 4.433477e-07, 2.170279e-07, 1.038855e-06, 2.710159e-07, 
    4.076032e-07, 1.293355e-07, 6.167879e-07, 1.692347e-06, 2.938019e-06, 
    2.353969e-06, 3.283282e-06, 2.377828e-07, 1.510529e-07, 5.681182e-08,
  3.009783e-06, 5.04916e-07, 1.344763e-06, 1.226342e-06, 3.527734e-07, 
    4.562802e-07, 3.706695e-07, 1.735138e-07, 2.651408e-07, 1.045045e-06, 
    2.623009e-06, 2.027763e-06, 3.864067e-06, 2.282153e-06, 5.160262e-07,
  5.59539e-06, 8.049467e-06, 2.653636e-06, 2.939726e-06, 5.952348e-07, 
    1.743911e-07, 6.729196e-07, 3.586102e-07, 1.429053e-07, 9.937477e-08, 
    1.47058e-06, 2.080402e-06, 2.748164e-06, 2.277841e-06, 1.395142e-06,
  6.571554e-06, 6.609177e-06, 6.174422e-06, 5.977593e-06, 2.681292e-06, 
    1.089357e-07, 3.273231e-07, 7.587607e-07, 6.013269e-07, 3.317577e-07, 
    3.861871e-07, 1.050495e-06, 1.411546e-06, 4.157286e-06, 3.059829e-06,
  4.728836e-06, 6.384372e-06, 7.158938e-06, 5.135316e-06, 5.174156e-06, 
    1.363017e-06, 5.037862e-08, 4.068141e-07, 1.082619e-06, 5.412624e-07, 
    2.309229e-07, 1.315857e-06, 1.255828e-06, 1.661655e-06, 2.892142e-06,
  2.22412e-06, 4.239057e-06, 8.326124e-06, 6.702711e-06, 4.787123e-06, 
    3.782088e-06, 2.448632e-06, 4.261935e-07, 1.087777e-06, 7.490123e-07, 
    4.417216e-07, 5.450611e-07, 7.444605e-07, 2.281597e-06, 2.925825e-06,
  2.750113e-06, 3.290149e-06, 8.616546e-06, 1.437095e-05, 9.438275e-06, 
    5.948921e-06, 5.681229e-06, 1.747754e-06, 2.088461e-06, 7.899937e-07, 
    7.822488e-07, 5.997554e-07, 5.952849e-07, 5.994361e-07, 5.107785e-07,
  4.061179e-06, 1.993285e-06, 3.918113e-06, 1.384795e-05, 8.724636e-06, 
    7.383686e-06, 8.375753e-06, 5.552279e-06, 4.237073e-06, 4.330855e-06, 
    1.553438e-06, 1.871588e-06, 1.671726e-06, 1.08153e-06, 4.997902e-07,
  5.788158e-06, 2.334981e-06, 1.366031e-06, 9.444841e-06, 1.346309e-05, 
    1.037202e-05, 1.083357e-05, 9.268068e-06, 8.392175e-06, 4.757759e-06, 
    5.356909e-06, 4.444887e-06, 1.728615e-06, 7.547144e-07, 7.370394e-07,
  5.905078e-06, 2.722147e-06, 1.228701e-06, 4.092104e-06, 6.680184e-06, 
    1.312216e-05, 1.117071e-05, 1.042481e-05, 9.918234e-06, 8.017535e-06, 
    7.507651e-06, 5.037562e-06, 3.335837e-06, 3.775892e-06, 1.211009e-06,
  7.887989e-09, 4.52725e-09, 2.729784e-07, 1.918911e-06, 9.652925e-07, 
    6.370348e-07, 2.490996e-06, 3.274039e-06, 3.935693e-06, 2.431583e-06, 
    1.825632e-06, 3.834635e-06, 3.729503e-06, 2.24826e-06, 1.206908e-06,
  1.199135e-06, 1.938576e-07, 1.299242e-06, 1.237729e-06, 1.564267e-06, 
    1.534796e-06, 1.444796e-06, 7.669982e-07, 4.375952e-07, 1.258787e-06, 
    1.574205e-06, 4.536742e-06, 2.74907e-06, 2.206304e-06, 1.555304e-07,
  3.080095e-06, 2.326159e-06, 2.024774e-06, 8.59325e-07, 5.170704e-07, 
    1.389248e-06, 1.441953e-06, 3.768746e-07, 6.317263e-07, 1.339139e-06, 
    3.387134e-06, 3.725339e-06, 2.890309e-06, 3.123002e-06, 1.294726e-06,
  5.847848e-06, 3.217096e-06, 1.486138e-06, 1.174059e-06, 2.189938e-06, 
    1.048992e-06, 1.997334e-06, 2.603041e-06, 7.640901e-07, 2.605738e-06, 
    4.375361e-06, 5.007588e-06, 4.098676e-06, 6.041362e-06, 5.339442e-06,
  8.508688e-06, 4.381246e-06, 1.66186e-06, 2.436016e-06, 2.030075e-06, 
    2.627891e-06, 2.889298e-06, 3.492921e-06, 1.445293e-06, 2.098763e-06, 
    2.841831e-06, 1.656917e-06, 2.381057e-06, 3.943725e-06, 2.401472e-06,
  8.278112e-06, 7.453933e-06, 4.15422e-06, 1.023397e-06, 2.081454e-06, 
    2.242807e-06, 4.278897e-06, 4.341149e-06, 2.865098e-06, 2.036893e-06, 
    2.230646e-06, 3.189312e-06, 3.645843e-06, 4.563787e-06, 6.463446e-06,
  1.024646e-05, 1.005687e-05, 7.557968e-06, 4.188937e-06, 2.819383e-06, 
    3.885152e-06, 2.965934e-06, 3.989677e-06, 3.587064e-06, 1.737766e-06, 
    2.767294e-06, 2.718774e-06, 4.769836e-06, 4.814825e-06, 7.126906e-06,
  7.637289e-06, 1.248074e-05, 1.223084e-05, 4.277872e-06, 1.380807e-06, 
    2.518274e-06, 3.954304e-06, 2.746243e-06, 3.413259e-06, 2.224344e-06, 
    2.819273e-06, 5.179559e-06, 3.631915e-06, 7.359103e-06, 1.323057e-05,
  8.779989e-06, 1.142505e-05, 7.886722e-06, 5.121695e-06, 3.014255e-06, 
    1.689869e-06, 4.209546e-06, 6.625672e-06, 1.027062e-05, 6.582978e-06, 
    5.982196e-06, 1.008703e-05, 2.023249e-05, 3.178102e-05, 2.661191e-05,
  8.818663e-06, 1.227576e-05, 1.119076e-05, 8.675398e-06, 2.546158e-06, 
    4.113715e-06, 3.841724e-06, 7.254329e-06, 9.885664e-06, 1.838833e-05, 
    2.187876e-05, 2.548463e-05, 3.213961e-05, 2.997596e-05, 3.786153e-05,
  7.788177e-08, 4.992571e-07, 4.438609e-07, 2.536914e-06, 4.510342e-06, 
    3.913131e-06, 2.25051e-06, 4.830612e-06, 5.414311e-06, 5.331557e-06, 
    4.066031e-06, 3.852384e-06, 3.226196e-06, 2.52355e-06, 1.618563e-06,
  5.384241e-07, 1.230821e-06, 1.473027e-06, 3.035211e-06, 3.182008e-06, 
    3.687425e-06, 2.827312e-06, 8.702747e-06, 8.717164e-06, 8.360752e-06, 
    9.165704e-06, 7.329124e-06, 4.724642e-06, 5.295255e-06, 5.387864e-06,
  6.976841e-07, 1.198089e-06, 1.62693e-06, 3.042298e-06, 2.227563e-06, 
    4.623423e-06, 4.797409e-06, 9.687811e-06, 9.552845e-06, 7.755727e-06, 
    7.082866e-06, 7.764061e-06, 8.547566e-06, 6.987613e-06, 7.19581e-06,
  1.380646e-06, 2.353579e-06, 1.845126e-06, 3.804732e-06, 4.298055e-06, 
    6.075902e-06, 6.76217e-06, 7.36946e-06, 1.03622e-05, 1.167193e-05, 
    9.543341e-06, 4.165459e-06, 3.018951e-06, 1.705441e-06, 2.489192e-06,
  1.205682e-06, 2.441744e-06, 4.313747e-06, 5.222223e-06, 4.475861e-06, 
    6.961382e-06, 8.070128e-06, 7.355719e-06, 9.501683e-06, 8.464841e-06, 
    1.237958e-05, 5.226056e-06, 4.017582e-06, 2.934582e-06, 4.308447e-06,
  1.071068e-06, 4.321059e-06, 7.583976e-06, 6.450505e-06, 6.234888e-06, 
    6.231366e-06, 7.902329e-06, 8.064962e-06, 1.113032e-05, 9.010629e-06, 
    1.280126e-05, 8.614508e-06, 5.730409e-06, 7.393071e-06, 4.4078e-06,
  1.099783e-07, 2.582919e-06, 8.106466e-06, 2.061141e-05, 8.681366e-06, 
    6.400578e-06, 1.221923e-05, 1.070153e-05, 1.202953e-05, 2.066732e-05, 
    1.580328e-05, 1.046692e-05, 1.256657e-05, 1.186521e-05, 8.771574e-06,
  2.227623e-08, 9.404573e-07, 4.896041e-06, 1.47366e-05, 1.065996e-05, 
    1.097255e-05, 1.343521e-05, 1.004046e-05, 1.181968e-05, 9.36759e-06, 
    2.020976e-05, 2.729188e-05, 2.188847e-05, 3.613681e-05, 2.246561e-05,
  3.653337e-07, 1.147377e-07, 7.332627e-07, 7.741663e-06, 2.054785e-05, 
    1.839417e-05, 1.259775e-05, 1.306651e-05, 1.469105e-05, 1.129059e-05, 
    9.844352e-06, 9.046401e-06, 1.470901e-05, 1.984898e-05, 3.489599e-05,
  3.259788e-07, 6.494467e-08, 8.081251e-08, 2.263122e-06, 1.052778e-05, 
    1.761287e-05, 1.500383e-05, 1.473786e-05, 1.388892e-05, 1.263922e-05, 
    1.043204e-05, 1.232755e-05, 1.17259e-05, 9.596242e-06, 1.333026e-05,
  9.385281e-09, 6.174373e-07, 4.874867e-06, 4.470513e-06, 3.803055e-06, 
    3.002304e-06, 3.939269e-06, 4.713536e-06, 3.467143e-06, 3.227737e-06, 
    1.354239e-06, 3.201169e-07, 1.29921e-06, 4.686533e-06, 6.069131e-06,
  1.106215e-05, 5.964204e-08, 2.302637e-06, 4.991197e-06, 3.417207e-06, 
    2.308009e-06, 1.310045e-06, 2.555876e-06, 2.479584e-06, 2.126053e-06, 
    8.403532e-07, 6.6221e-07, 2.657774e-07, 3.044632e-06, 3.403871e-06,
  1.07041e-05, 1.235441e-05, 4.804833e-06, 4.318801e-06, 3.376478e-06, 
    1.100362e-06, 9.886887e-07, 6.328805e-07, 1.556674e-06, 1.800978e-06, 
    1.476152e-06, 8.353504e-07, 7.093412e-07, 2.137635e-06, 2.858155e-06,
  1.202216e-05, 1.146664e-05, 6.589556e-06, 4.022036e-06, 3.757666e-06, 
    1.723111e-06, 2.151202e-06, 3.588023e-07, 9.930798e-07, 1.829852e-06, 
    8.725453e-07, 1.258354e-06, 1.505341e-06, 3.024853e-06, 3.662367e-06,
  8.016488e-06, 1.134762e-05, 6.582654e-06, 6.597073e-06, 4.184069e-06, 
    2.1383e-06, 1.132734e-06, 5.262999e-07, 5.366019e-07, 1.042381e-06, 
    1.731776e-06, 1.179018e-06, 1.62379e-06, 2.831852e-06, 3.851932e-06,
  3.599832e-06, 1.10903e-05, 1.188972e-05, 7.398536e-06, 4.28514e-06, 
    1.805331e-06, 5.391004e-07, 7.824074e-07, 1.036079e-06, 1.90276e-06, 
    9.723071e-07, 1.406148e-06, 1.575504e-06, 1.86874e-06, 3.793683e-06,
  1.879038e-06, 9.445357e-06, 2.588124e-05, 2.896627e-05, 8.645043e-06, 
    3.852157e-06, 2.211526e-06, 1.965856e-07, 9.859647e-07, 1.257648e-06, 
    2.769013e-06, 2.549266e-06, 3.587925e-06, 4.871376e-06, 3.484654e-06,
  2.396814e-06, 5.680887e-06, 1.747642e-05, 3.526628e-05, 1.532831e-05, 
    8.783203e-06, 6.631803e-06, 2.35816e-06, 4.071255e-06, 3.475402e-06, 
    4.259219e-06, 4.574553e-06, 6.598789e-06, 5.324362e-06, 8.299315e-06,
  8.325184e-07, 3.407734e-06, 1.084443e-05, 3.13651e-05, 3.657368e-05, 
    2.292968e-05, 7.924758e-06, 7.863637e-06, 1.228901e-05, 1.238855e-05, 
    9.988808e-06, 9.121485e-06, 9.761278e-06, 1.717254e-05, 2.454593e-05,
  7.096981e-08, 8.774332e-07, 5.237111e-06, 2.989438e-05, 3.039061e-05, 
    4.499791e-05, 3.090285e-05, 1.711963e-05, 1.522737e-05, 1.667508e-05, 
    2.152066e-05, 3.018938e-05, 2.414685e-05, 1.753045e-05, 2.082516e-05,
  1.556698e-09, 2.463176e-07, 1.734899e-06, 3.69695e-06, 3.142288e-06, 
    3.04273e-06, 2.531263e-06, 2.092334e-06, 2.49675e-06, 1.118364e-06, 
    7.970265e-07, 7.155118e-07, 1.163627e-06, 3.684438e-07, 1.005495e-06,
  4.46685e-06, 6.975707e-07, 1.940592e-06, 2.898734e-06, 3.258529e-06, 
    2.330015e-06, 1.891109e-06, 9.744516e-07, 9.138805e-07, 1.062216e-06, 
    9.812364e-07, 1.158215e-06, 4.144328e-07, 2.193311e-06, 1.13942e-06,
  8.280143e-06, 6.269884e-06, 2.058054e-06, 1.713656e-06, 2.402092e-06, 
    1.037958e-06, 1.400144e-06, 1.631135e-06, 1.994063e-06, 8.055893e-07, 
    1.938784e-06, 2.098228e-06, 2.617525e-06, 4.259704e-06, 4.378722e-06,
  1.433167e-05, 1.593313e-06, 8.218205e-07, 2.386542e-06, 2.931711e-06, 
    3.948875e-07, 2.319047e-07, 2.752938e-07, 7.863909e-07, 3.717648e-06, 
    3.029026e-06, 4.549421e-06, 7.006733e-06, 7.144608e-06, 7.375755e-06,
  7.631445e-06, 2.524072e-06, 7.698914e-07, 1.868541e-06, 4.807727e-07, 
    6.267928e-07, 1.312832e-07, 1.549267e-06, 2.826705e-06, 4.731633e-06, 
    8.824128e-06, 1.211589e-05, 1.000885e-05, 8.545864e-06, 8.429738e-06,
  5.875558e-06, 3.461259e-06, 3.383181e-06, 1.65554e-06, 1.72405e-06, 
    1.014951e-06, 3.165008e-06, 3.723349e-06, 8.942443e-06, 1.19035e-05, 
    1.213455e-05, 1.069723e-05, 5.545079e-06, 6.475695e-06, 5.216044e-06,
  7.205052e-06, 7.244215e-06, 1.033471e-05, 3.808995e-06, 9.162292e-06, 
    4.75465e-06, 6.784093e-06, 7.490851e-06, 6.239409e-06, 1.261943e-05, 
    1.383895e-05, 1.053816e-05, 6.946079e-06, 6.377869e-06, 4.918436e-06,
  8.092699e-06, 1.113253e-05, 1.263585e-05, 1.754978e-05, 1.075982e-05, 
    1.144896e-05, 1.62636e-05, 1.26899e-05, 1.806375e-05, 1.298836e-05, 
    1.33403e-05, 1.030903e-05, 9.072385e-06, 7.453375e-06, 4.853663e-06,
  9.14356e-06, 1.759621e-05, 2.032408e-05, 2.185692e-05, 3.749243e-05, 
    3.156986e-05, 2.275832e-05, 2.085601e-05, 2.173323e-05, 1.621513e-05, 
    1.801212e-05, 1.616598e-05, 1.842139e-05, 1.813133e-05, 1.26015e-05,
  5.057061e-06, 1.685995e-05, 1.507661e-05, 2.758404e-05, 3.827631e-05, 
    6.236354e-05, 3.754684e-05, 3.184054e-05, 2.817885e-05, 2.490051e-05, 
    2.491383e-05, 3.876738e-05, 3.412326e-05, 2.234401e-05, 1.354912e-05,
  1.041312e-07, 1.740219e-06, 5.065962e-06, 1.023829e-05, 1.061943e-05, 
    1.292521e-05, 1.169792e-05, 1.262432e-05, 1.385516e-05, 1.978969e-05, 
    2.060183e-05, 2.257142e-05, 2.029591e-05, 1.861237e-05, 1.883961e-05,
  6.74877e-07, 2.173895e-06, 5.387923e-06, 4.903676e-06, 5.670686e-06, 
    1.015021e-05, 1.258449e-05, 1.129091e-05, 1.548349e-05, 1.336843e-05, 
    1.71409e-05, 1.627423e-05, 2.027284e-05, 1.709088e-05, 1.666266e-05,
  4.599517e-07, 3.923762e-06, 4.413412e-06, 4.027671e-06, 2.589516e-06, 
    3.552242e-06, 4.978584e-06, 7.272637e-06, 1.074262e-05, 1.33151e-05, 
    1.256621e-05, 1.416406e-05, 1.477174e-05, 1.207942e-05, 1.217271e-05,
  5.464947e-07, 1.236434e-06, 4.305679e-06, 4.320734e-06, 1.33907e-06, 
    1.670092e-06, 2.49394e-06, 1.791937e-06, 3.79062e-06, 9.08643e-06, 
    8.425641e-06, 7.800373e-06, 7.432369e-06, 7.370548e-06, 8.746117e-06,
  2.135743e-06, 2.364776e-06, 1.805811e-06, 2.62395e-06, 2.813432e-06, 
    2.399713e-06, 1.76649e-06, 1.623162e-06, 3.604889e-06, 4.099498e-06, 
    4.085925e-06, 3.950083e-06, 4.277135e-06, 4.871131e-06, 5.524545e-06,
  2.426819e-06, 1.065513e-05, 1.675266e-05, 6.208108e-06, 3.221772e-06, 
    7.243363e-06, 4.25997e-06, 3.100529e-06, 2.833035e-06, 3.430629e-06, 
    4.832894e-06, 2.255383e-06, 3.513645e-06, 3.397113e-06, 3.188245e-06,
  2.615861e-06, 1.132929e-05, 2.614866e-05, 3.403359e-05, 1.846024e-05, 
    1.242504e-05, 9.763387e-06, 5.45226e-06, 4.230591e-06, 4.125401e-06, 
    4.608423e-06, 5.126984e-06, 4.95084e-06, 3.969612e-06, 3.580149e-06,
  2.296219e-06, 1.215294e-05, 2.220171e-05, 4.085658e-05, 3.364199e-05, 
    2.217702e-05, 1.521222e-05, 9.597301e-06, 7.110667e-06, 6.863083e-06, 
    6.079566e-06, 9.767682e-06, 6.587726e-06, 6.192269e-06, 5.979456e-06,
  5.477602e-06, 9.860117e-06, 1.243752e-05, 2.372496e-05, 4.385617e-05, 
    3.771515e-05, 2.142966e-05, 1.079096e-05, 8.918247e-06, 6.248285e-06, 
    6.899733e-06, 7.613607e-06, 7.523085e-06, 5.579372e-06, 5.131082e-06,
  8.296163e-06, 9.794387e-06, 1.58664e-05, 2.059327e-05, 3.243646e-05, 
    5.265023e-05, 2.496803e-05, 1.870441e-05, 1.339016e-05, 1.253289e-05, 
    1.365748e-05, 1.169361e-05, 1.044254e-05, 9.442846e-06, 1.985187e-05,
  4.918494e-07, 3.332314e-06, 8.407646e-06, 1.114193e-05, 7.748437e-06, 
    5.659473e-06, 5.707909e-06, 3.219698e-06, 4.553746e-06, 4.194339e-06, 
    4.272112e-06, 3.992781e-06, 4.306959e-06, 4.73528e-06, 4.047987e-06,
  2.621982e-06, 2.331931e-06, 8.592049e-06, 1.030616e-05, 8.345995e-06, 
    8.005863e-06, 8.448454e-06, 8.205575e-06, 7.493805e-06, 7.310472e-06, 
    4.422322e-06, 4.573225e-06, 4.788968e-06, 5.685995e-06, 6.952028e-06,
  2.724805e-06, 3.934367e-06, 7.923828e-06, 9.839846e-06, 9.387823e-06, 
    6.766696e-06, 9.000999e-06, 8.109322e-06, 8.115962e-06, 7.630109e-06, 
    4.617084e-06, 5.487344e-06, 6.944687e-06, 7.915201e-06, 1.134877e-05,
  3.245501e-06, 2.759979e-06, 7.299904e-06, 9.702644e-06, 7.178589e-06, 
    8.422213e-06, 9.864561e-06, 7.825925e-06, 9.533729e-06, 8.799996e-06, 
    8.557427e-06, 9.778197e-06, 1.053882e-05, 1.179667e-05, 1.615852e-05,
  1.999767e-06, 2.188553e-06, 3.308847e-06, 7.873673e-06, 7.545153e-06, 
    9.772917e-06, 8.544889e-06, 1.08002e-05, 8.488149e-06, 8.209759e-06, 
    1.253974e-05, 1.419133e-05, 1.35784e-05, 1.424596e-05, 1.833777e-05,
  8.546463e-07, 9.320599e-07, 2.973511e-06, 5.704232e-06, 6.926859e-06, 
    6.322311e-06, 6.116656e-06, 7.533732e-06, 7.609798e-06, 8.446407e-06, 
    9.199151e-06, 1.064545e-05, 1.097213e-05, 1.357109e-05, 1.433945e-05,
  1.172055e-06, 9.462723e-07, 1.783417e-06, 5.657624e-06, 4.342549e-06, 
    8.147762e-06, 9.660851e-06, 7.113654e-06, 1.004467e-05, 9.176795e-06, 
    8.571714e-06, 9.386117e-06, 9.992046e-06, 1.172869e-05, 1.132428e-05,
  1.829457e-06, 8.459547e-07, 1.776255e-06, 3.903542e-06, 4.216746e-06, 
    3.805564e-06, 4.748289e-06, 4.680712e-06, 7.749749e-06, 8.808624e-06, 
    8.735293e-06, 9.516647e-06, 9.508652e-06, 9.917099e-06, 1.130514e-05,
  1.285344e-05, 9.282548e-06, 1.212315e-06, 4.762062e-06, 5.127167e-06, 
    6.671924e-06, 6.027529e-06, 5.443654e-06, 7.483944e-06, 7.853392e-06, 
    7.131686e-06, 7.958197e-06, 1.038037e-05, 9.934909e-06, 1.728273e-05,
  2.600369e-05, 2.044194e-05, 4.991334e-07, 2.282073e-06, 7.438915e-06, 
    1.229949e-05, 7.583313e-06, 7.308803e-06, 7.455195e-06, 9.362323e-06, 
    8.824585e-06, 8.744327e-06, 1.735711e-05, 1.48901e-05, 1.968549e-05,
  1.895358e-10, 1.830784e-06, 1.940997e-06, 3.082561e-06, 3.188816e-06, 
    2.839472e-06, 2.265318e-06, 2.118127e-06, 2.599944e-06, 2.138245e-06, 
    2.151867e-06, 2.946699e-06, 6.201342e-06, 6.978818e-06, 6.220842e-06,
  9.943564e-07, 4.02764e-07, 3.216028e-06, 3.364197e-06, 2.36498e-06, 
    3.178543e-06, 3.100323e-06, 2.345294e-06, 2.497391e-06, 2.222084e-06, 
    2.40929e-06, 3.463682e-06, 5.570117e-06, 5.801743e-06, 8.387967e-06,
  9.999789e-07, 2.072476e-06, 4.694858e-06, 4.164534e-06, 3.629858e-06, 
    2.662149e-06, 3.184066e-06, 3.081066e-06, 3.06477e-06, 3.415761e-06, 
    3.514954e-06, 4.862145e-06, 6.094636e-06, 6.874953e-06, 6.469075e-06,
  1.727524e-06, 3.22296e-06, 3.101435e-06, 5.358111e-06, 3.29856e-06, 
    3.227119e-06, 3.633342e-06, 3.524517e-06, 3.979445e-06, 4.125006e-06, 
    3.470623e-06, 3.611722e-06, 5.614269e-06, 4.293316e-06, 5.760803e-06,
  4.04175e-06, 5.637228e-06, 1.896233e-06, 4.739092e-06, 2.757558e-06, 
    3.913608e-06, 4.02939e-06, 3.860047e-06, 3.906729e-06, 4.07723e-06, 
    5.186238e-06, 5.756531e-06, 6.897093e-06, 6.630523e-06, 4.284635e-06,
  1.428738e-06, 2.457255e-06, 4.469845e-06, 1.82635e-06, 3.21544e-06, 
    3.108122e-06, 3.597044e-06, 2.764635e-06, 3.897516e-06, 4.554627e-06, 
    5.469684e-06, 7.262911e-06, 9.386376e-06, 8.358342e-06, 6.501343e-06,
  6.838175e-06, 2.528796e-06, 4.550914e-06, 6.86156e-06, 5.210053e-06, 
    3.622501e-06, 3.376566e-06, 2.220162e-06, 4.494342e-06, 5.447747e-06, 
    7.944083e-06, 9.629602e-06, 8.93215e-06, 1.018475e-05, 9.132584e-06,
  1.145097e-05, 4.397234e-06, 1.166349e-06, 6.879843e-06, 3.526397e-06, 
    7.46945e-06, 3.564597e-06, 2.354958e-06, 4.730392e-06, 5.300462e-06, 
    7.331015e-06, 8.387371e-06, 1.012637e-05, 1.085788e-05, 9.616345e-06,
  1.847518e-05, 1.348809e-05, 1.075605e-06, 1.55843e-06, 5.304691e-06, 
    6.524989e-06, 1.051542e-05, 7.636961e-06, 5.751709e-06, 5.079624e-06, 
    7.188981e-06, 1.123727e-05, 1.380735e-05, 8.960265e-06, 9.156851e-06,
  3.370369e-05, 3.35714e-05, 9.790164e-06, 3.047033e-07, 1.378887e-07, 
    5.896278e-06, 1.446158e-05, 1.484505e-05, 1.234142e-05, 8.084857e-06, 
    9.538195e-06, 9.360467e-06, 1.085286e-05, 7.649509e-06, 9.317785e-06,
  2.832863e-08, 3.181827e-06, 2.489499e-06, 2.725017e-06, 4.252553e-06, 
    5.699091e-06, 7.057436e-06, 7.227695e-06, 1.697697e-05, 8.000139e-06, 
    1.434707e-05, 1.326276e-05, 6.680619e-06, 3.959593e-06, 1.844308e-06,
  7.705241e-07, 3.467794e-07, 1.685744e-06, 2.367345e-06, 3.346167e-06, 
    5.441638e-06, 6.192688e-06, 6.681501e-06, 6.001416e-06, 8.275228e-06, 
    1.117407e-05, 9.379675e-06, 4.150629e-06, 2.691643e-06, 1.633903e-06,
  1.095285e-06, 6.897291e-07, 2.408603e-06, 2.965135e-06, 3.046719e-06, 
    3.164966e-06, 3.682011e-06, 6.821695e-06, 1.12012e-05, 1.238975e-05, 
    1.342233e-05, 7.875382e-06, 5.035504e-06, 3.877069e-06, 2.345319e-06,
  3.522447e-06, 5.649677e-07, 1.441328e-06, 2.082086e-06, 2.955424e-06, 
    3.377279e-06, 4.847718e-06, 6.10721e-06, 1.427419e-05, 1.569444e-05, 
    1.54495e-05, 9.31232e-06, 6.449352e-06, 3.288432e-06, 1.377566e-06,
  2.328186e-06, 1.821132e-06, 2.812785e-07, 2.528652e-06, 2.517424e-06, 
    4.481543e-06, 5.74193e-06, 5.162331e-06, 7.288491e-06, 2.033587e-05, 
    1.445417e-05, 1.0686e-05, 7.788815e-06, 3.68498e-06, 2.756016e-06,
  4.49864e-06, 3.783869e-06, 6.874879e-07, 1.604844e-08, 1.695534e-06, 
    3.761331e-06, 6.606e-06, 4.436324e-06, 7.863211e-06, 1.184009e-05, 
    1.156327e-05, 1.124348e-05, 7.414486e-06, 5.436341e-06, 2.380398e-06,
  8.876775e-06, 3.597851e-06, 1.89602e-06, 1.291686e-06, 3.407023e-06, 
    3.033332e-06, 6.702104e-06, 2.11081e-06, 4.793081e-06, 7.909397e-06, 
    7.620778e-06, 1.049007e-05, 7.746102e-06, 7.123627e-06, 4.499218e-06,
  1.468521e-05, 4.04326e-06, 7.258479e-07, 1.017495e-06, 2.10905e-08, 
    2.234175e-06, 4.921757e-06, 4.14637e-06, 1.121721e-05, 7.016075e-06, 
    6.860048e-06, 9.004024e-06, 7.611353e-06, 7.751194e-06, 4.91049e-06,
  3.061147e-05, 7.52503e-06, 6.565348e-07, 1.079798e-07, 6.155581e-07, 
    7.126949e-07, 4.468414e-06, 6.37102e-06, 1.100133e-05, 5.807224e-06, 
    6.525092e-06, 3.902692e-06, 2.031149e-06, 4.085537e-06, 5.295358e-06,
  4.676263e-05, 1.171034e-05, 9.490492e-07, 3.417696e-09, 5.500302e-08, 
    8.085985e-07, 3.604721e-06, 4.844005e-06, 7.068813e-06, 1.324449e-05, 
    7.916219e-06, 5.835673e-06, 5.870486e-06, 1.604662e-06, 5.997942e-06,
  5.95437e-10, 1.847885e-07, 2.234217e-06, 5.04048e-06, 1.231264e-05, 
    1.089773e-05, 7.295552e-06, 1.189805e-05, 1.473903e-05, 4.877705e-06, 
    4.281924e-06, 3.879387e-06, 1.101111e-06, 4.586869e-07, 2.085307e-07,
  1.311428e-07, 2.71545e-07, 1.912255e-06, 5.234475e-06, 4.68362e-06, 
    7.187394e-06, 1.40177e-05, 1.429353e-05, 2.526615e-05, 1.229353e-05, 
    3.097877e-06, 4.344438e-06, 8.982977e-07, 1.188344e-07, 6.634226e-08,
  9.781493e-09, 8.699187e-07, 1.915906e-06, 3.674519e-06, 3.537822e-06, 
    2.000469e-06, 3.540665e-06, 1.374558e-05, 2.214098e-05, 1.563537e-05, 
    1.076292e-06, 2.251172e-06, 2.589944e-07, 5.371214e-08, 2.024398e-07,
  1.507444e-09, 8.931557e-07, 1.30729e-06, 2.922756e-06, 6.128889e-06, 
    2.559657e-06, 5.839608e-06, 6.500614e-06, 7.642315e-06, 4.288065e-06, 
    5.291561e-06, 1.238698e-06, 1.683624e-07, 4.528756e-09, 5.877162e-07,
  9.535674e-10, 3.474404e-07, 8.593382e-07, 2.591057e-06, 3.637223e-06, 
    5.920991e-06, 6.887018e-06, 6.599953e-06, 1.098283e-06, 8.561337e-06, 
    7.714435e-06, 3.404895e-06, 1.538771e-06, 7.368291e-07, 9.24508e-07,
  1.030327e-09, 2.356185e-07, 1.283455e-06, 1.058018e-06, 1.38472e-06, 
    4.338623e-06, 7.434501e-06, 2.313506e-06, 4.896728e-06, 1.292419e-05, 
    1.184387e-05, 7.007558e-06, 2.32802e-06, 1.771653e-06, 8.022348e-07,
  6.756272e-10, 1.860899e-07, 1.825892e-06, 8.226044e-07, 1.445492e-06, 
    4.762333e-06, 4.217957e-06, 1.27718e-06, 3.948394e-06, 6.177002e-06, 
    5.725251e-06, 5.973417e-06, 3.394977e-06, 5.758796e-07, 7.396707e-07,
  8.240487e-09, 5.85935e-08, 6.06841e-08, 5.314402e-07, 2.504356e-07, 
    2.59758e-06, 4.146028e-06, 4.029989e-07, 6.354788e-06, 2.260292e-06, 
    7.615e-06, 3.442258e-06, 2.851323e-06, 1.747555e-06, 1.684364e-06,
  5.312014e-07, 1.32297e-07, 4.700405e-10, 7.268575e-11, 4.226164e-10, 
    1.586926e-07, 3.265643e-06, 4.261929e-06, 9.015669e-06, 4.910881e-06, 
    6.018073e-06, 1.688775e-06, 4.983277e-06, 2.119255e-06, 6.11219e-07,
  8.372531e-07, 1.324815e-07, 1.397986e-08, 6.060973e-11, 2.436795e-10, 
    1.02943e-09, 8.715679e-07, 3.599228e-06, 7.117126e-06, 7.451612e-06, 
    1.098951e-05, 1.018467e-05, 3.547203e-06, 3.469865e-06, 1.5982e-06,
  1.67222e-07, 1.889487e-06, 1.137985e-05, 9.847175e-06, 2.395422e-05, 
    4.651234e-05, 0.0001052643, 7.467251e-05, 0.0001209255, 3.003971e-05, 
    1.02959e-05, 5.710939e-06, 4.993575e-06, 7.337469e-06, 5.834107e-06,
  8.26627e-06, 1.23452e-06, 2.100344e-05, 2.353591e-05, 2.217071e-05, 
    7.257387e-05, 8.286244e-05, 0.0001136791, 9.145999e-05, 6.531444e-05, 
    2.562791e-06, 1.409577e-06, 4.985451e-07, 5.560329e-07, 5.500911e-08,
  1.52697e-05, 1.378033e-05, 2.123829e-05, 1.114037e-05, 7.098424e-05, 
    4.039126e-05, 8.180651e-05, 9.687086e-05, 7.310636e-05, 1.657472e-05, 
    1.100286e-06, 7.757942e-07, 1.602809e-07, 2.463602e-09, 8.663774e-09,
  1.530297e-05, 1.847162e-05, 3.38532e-06, 1.686128e-05, 2.495492e-05, 
    2.419466e-06, 1.605107e-05, 2.782932e-05, 4.928344e-05, 3.033063e-05, 
    6.784561e-06, 5.25813e-07, 2.407147e-07, 2.578271e-07, 1.401816e-07,
  6.864673e-06, 1.640746e-05, 9.573741e-07, 1.214999e-05, 1.38218e-05, 
    1.321855e-05, 1.139799e-05, 3.737981e-05, 4.011258e-05, 3.859685e-05, 
    1.019057e-05, 1.517231e-06, 5.595376e-08, 7.185099e-07, 9.518184e-07,
  5.362717e-06, 1.26215e-05, 2.137222e-05, 8.421906e-07, 1.277834e-05, 
    2.942619e-05, 4.543335e-05, 2.108026e-05, 1.482847e-05, 4.28973e-05, 
    1.036531e-05, 1.342612e-06, 8.454124e-07, 1.833637e-06, 1.66829e-06,
  5.123499e-09, 1.182517e-06, 7.619078e-06, 1.784948e-05, 4.694096e-06, 
    3.091835e-05, 5.450514e-05, 3.225652e-05, 3.116406e-05, 1.986608e-05, 
    1.157481e-05, 1.282067e-06, 6.885309e-07, 1.285664e-06, 2.386092e-06,
  1.093044e-08, 3.054829e-07, 1.971837e-06, 1.196316e-05, 1.293191e-06, 
    2.273966e-05, 4.137691e-05, 1.25642e-05, 3.751847e-05, 3.064289e-05, 
    7.281008e-06, 1.097119e-06, 8.705085e-07, 1.279399e-06, 2.824912e-06,
  2.513824e-08, 1.890469e-07, 1.061732e-08, 1.1624e-05, 3.806848e-05, 
    3.565498e-06, 2.174219e-05, 4.167094e-05, 5.95709e-05, 1.902044e-05, 
    4.732882e-06, 1.142562e-06, 1.582795e-06, 1.299942e-06, 2.698668e-06,
  4.940064e-08, 4.043074e-08, 3.463734e-07, 2.71028e-06, 1.581762e-05, 
    1.413643e-05, 1.22613e-05, 1.774265e-05, 5.608593e-05, 2.611097e-05, 
    8.767956e-06, 4.87164e-06, 3.503739e-06, 1.85326e-06, 2.315264e-06,
  1.979123e-09, 1.404271e-08, 3.809731e-05, 1.099875e-05, 1.237171e-05, 
    6.942655e-06, 2.959812e-05, 1.24306e-05, 1.293551e-06, 1.287142e-06, 
    3.875076e-07, 4.630527e-07, 1.321262e-07, 3.146463e-07, 5.590126e-07,
  7.366615e-05, 3.42512e-06, 4.564682e-05, 8.282554e-05, 4.377512e-06, 
    3.368342e-06, 2.878545e-06, 9.642442e-07, 1.013344e-06, 9.386201e-07, 
    8.838211e-07, 7.388458e-07, 2.830786e-07, 3.755711e-07, 2.381225e-07,
  9.626026e-05, 7.201199e-05, 4.260748e-05, 9.050293e-05, 3.430656e-05, 
    2.032692e-06, 1.823112e-06, 9.56393e-07, 1.102216e-06, 2.004839e-06, 
    2.532399e-06, 1.5538e-06, 1.068154e-06, 7.736534e-07, 8.144673e-07,
  9.308186e-05, 8.133156e-05, 3.25607e-05, 8.080461e-05, 0.0001059377, 
    1.60732e-05, 2.475383e-06, 1.315688e-06, 1.141856e-06, 2.448809e-06, 
    2.584407e-06, 3.397873e-06, 2.623062e-06, 1.805438e-06, 2.131276e-06,
  7.75828e-05, 7.680753e-05, 7.636551e-06, 8.372161e-05, 9.020448e-05, 
    2.026192e-05, 3.921572e-06, 2.394073e-06, 9.639313e-07, 2.406971e-06, 
    4.030072e-06, 4.922016e-06, 5.485338e-06, 2.949399e-06, 2.876167e-06,
  7.252019e-05, 4.353957e-05, 6.928499e-05, 6.736105e-09, 3.63894e-05, 
    7.293422e-05, 3.836723e-05, 3.29406e-06, 1.509202e-06, 2.971761e-06, 
    4.48067e-06, 7.980909e-06, 6.607862e-06, 4.256681e-06, 3.540712e-06,
  5.321098e-05, 3.753314e-05, 7.544426e-05, 7.950909e-05, 8.465371e-05, 
    7.78689e-05, 0.0001123159, 3.594789e-05, 2.12848e-06, 2.328387e-06, 
    4.214559e-06, 7.992461e-06, 9.509143e-06, 7.796726e-06, 4.440464e-06,
  4.814879e-05, 1.940549e-05, 3.306388e-05, 8.455156e-05, 1.3842e-08, 
    2.197877e-05, 8.52517e-05, 5.817567e-05, 1.936311e-05, 3.132339e-06, 
    4.509634e-06, 7.823091e-06, 1.300665e-05, 1.766561e-05, 2.417671e-05,
  5.193529e-05, 1.905474e-05, 7.705366e-06, 4.990626e-05, 5.549083e-05, 
    2.220432e-06, 5.497621e-05, 6.998557e-05, 8.135201e-05, 2.65754e-05, 
    3.346041e-06, 5.712089e-06, 1.026865e-05, 2.349614e-05, 3.301875e-05,
  2.399481e-05, 1.557904e-05, 5.564506e-06, 1.239838e-05, 5.327507e-05, 
    4.573863e-05, 2.801107e-05, 7.092657e-05, 8.416972e-05, 6.368417e-05, 
    8.604288e-06, 5.587498e-06, 1.000024e-05, 1.718201e-05, 2.278226e-05,
  8.130214e-09, 3.866904e-06, 1.166419e-05, 2.752205e-06, 3.280707e-06, 
    3.199312e-06, 5.20308e-06, 9.243881e-06, 1.731823e-05, 9.985243e-06, 
    8.733627e-06, 5.81809e-06, 6.839698e-06, 1.941587e-05, 4.105833e-05,
  5.765595e-05, 2.209972e-07, 2.730461e-05, 2.052166e-05, 2.446789e-06, 
    2.552451e-06, 3.565342e-06, 1.042717e-05, 2.463203e-05, 1.230425e-05, 
    1.58517e-05, 4.206331e-06, 7.756641e-06, 1.886673e-05, 5.714132e-05,
  3.39666e-05, 4.945626e-05, 3.309394e-05, 2.132589e-05, 1.069728e-05, 
    1.38578e-06, 3.349246e-06, 6.804978e-06, 2.242206e-05, 1.620226e-05, 
    1.650816e-05, 2.017974e-05, 4.97562e-05, 8.764462e-06, 5.328352e-05,
  7.367356e-05, 4.571564e-05, 8.273081e-06, 4.755452e-05, 5.965956e-06, 
    1.173678e-05, 2.745305e-06, 5.874886e-06, 1.268592e-05, 2.569037e-05, 
    2.71849e-05, 3.936852e-05, 2.401978e-05, 2.449999e-05, 2.534855e-05,
  7.182986e-05, 6.473018e-05, 1.68076e-06, 6.425286e-05, 2.206344e-05, 
    1.164797e-05, 2.176492e-06, 2.958878e-06, 7.004031e-06, 1.389655e-05, 
    2.228547e-05, 3.331575e-05, 5.162107e-05, 4.83135e-05, 5.49702e-05,
  8.901754e-05, 3.820272e-05, 6.025895e-05, 1.102834e-05, 5.629611e-05, 
    7.264572e-06, 7.655668e-06, 1.124651e-05, 4.908982e-06, 8.154499e-06, 
    2.467537e-05, 1.643688e-05, 5.69879e-05, 5.415701e-05, 0.0001069935,
  7.42801e-05, 5.269689e-05, 8.667379e-05, 7.899875e-05, 3.455019e-05, 
    2.911345e-05, 2.620667e-05, 7.312803e-06, 1.080908e-05, 1.142779e-05, 
    1.797536e-05, 3.075331e-05, 4.293655e-05, 9.647293e-05, 0.0001562531,
  6.604827e-05, 4.463343e-05, 5.106797e-05, 6.262586e-05, 4.962173e-07, 
    2.555458e-05, 3.176918e-05, 1.421919e-05, 3.490872e-05, 3.191184e-05, 
    3.610236e-05, 2.967289e-05, 4.672928e-05, 0.0001180241, 9.364571e-05,
  6.824766e-05, 4.415039e-05, 1.151519e-05, 1.644731e-05, 2.65719e-05, 
    9.69549e-08, 2.185353e-05, 5.004155e-05, 5.788067e-05, 4.636743e-05, 
    3.741904e-05, 3.982698e-05, 4.573289e-05, 3.568573e-05, 7.952043e-05,
  7.600513e-05, 4.109272e-05, 2.855164e-06, 1.68489e-06, 1.153894e-06, 
    1.644315e-05, 6.957781e-06, 6.315864e-05, 5.447263e-05, 7.676184e-05, 
    5.428162e-05, 4.429267e-05, 5.67214e-05, 9.762118e-05, 0.0001304219,
  4.889501e-10, 9.987512e-09, 3.305375e-06, 3.564955e-06, 1.952442e-06, 
    3.085674e-06, 7.432056e-06, 1.588774e-05, 2.420087e-05, 3.997995e-05, 
    3.156451e-05, 1.989481e-05, 6.953082e-06, 1.029863e-05, 2.369605e-05,
  8.707e-06, 1.345236e-08, 6.017283e-07, 4.426363e-06, 7.829091e-06, 
    4.231169e-06, 1.08396e-05, 2.71618e-05, 3.396907e-05, 4.950432e-05, 
    3.386835e-05, 1.938424e-05, 2.640452e-05, 3.368308e-06, 2.087226e-05,
  9.330309e-06, 9.341852e-06, 4.195292e-07, 5.248315e-06, 1.578082e-05, 
    1.18456e-05, 1.075361e-05, 2.96966e-05, 9.858234e-05, 6.898852e-05, 
    3.140057e-05, 2.956312e-05, 5.407371e-06, 2.00395e-06, 2.885191e-06,
  4.891887e-06, 5.508236e-06, 7.814553e-08, 2.583206e-06, 9.05851e-06, 
    8.761006e-06, 1.156384e-05, 2.12374e-05, 0.0001285405, 0.000100369, 
    4.979689e-05, 3.973599e-05, 5.431176e-05, 2.106137e-05, 3.14387e-05,
  7.886983e-06, 2.437771e-06, 3.594639e-07, 6.279834e-06, 1.035221e-05, 
    1.943064e-05, 1.405872e-05, 3.819945e-05, 9.445013e-05, 0.0001599291, 
    0.0001032818, 5.846026e-05, 4.575318e-05, 6.990782e-05, 7.391476e-05,
  7.281566e-06, 2.8436e-06, 3.286041e-06, 8.343171e-07, 6.235885e-06, 
    1.531988e-05, 2.75107e-05, 4.657996e-05, 9.080743e-05, 0.0001886534, 
    0.0002171462, 0.0001132852, 8.729771e-05, 7.360873e-05, 6.65889e-05,
  1.620258e-05, 9.984828e-06, 3.62451e-06, 7.031447e-06, 3.29263e-06, 
    1.14021e-05, 2.083513e-05, 4.763761e-05, 8.361732e-05, 0.0002437093, 
    0.0003375378, 0.0002751483, 0.0001007201, 6.629878e-05, 3.555342e-05,
  4.348192e-05, 9.730722e-06, 3.850288e-06, 4.157396e-06, 1.247508e-08, 
    5.155021e-06, 1.312407e-05, 2.131983e-05, 6.75655e-05, 0.0002225562, 
    0.000348054, 0.0002318602, 0.0002488231, 0.0001422412, 1.727596e-05,
  5.614118e-05, 1.521261e-05, 2.986944e-06, 3.975193e-06, 2.415614e-06, 
    1.80234e-06, 1.354413e-05, 1.974718e-05, 4.929668e-05, 5.785942e-05, 
    0.0001035565, 0.0002187858, 0.0003493357, 0.0001776974, 7.866934e-05,
  3.001595e-05, 2.067764e-05, 6.387359e-06, 1.243734e-06, 1.492223e-06, 
    4.690186e-06, 1.090818e-05, 4.181856e-05, 4.230031e-05, 5.527874e-05, 
    3.024006e-05, 6.890472e-05, 0.0002801089, 0.0003077148, 8.671647e-05,
  4.570615e-06, 2.738203e-05, 2.270588e-05, 3.758345e-05, 4.858476e-05, 
    6.903463e-05, 0.0001077515, 8.845834e-05, 5.386854e-05, 4.299998e-05, 
    6.310566e-05, 9.010886e-05, 4.019682e-06, 3.333378e-06, 2.546621e-06,
  2.75278e-05, 1.398207e-05, 4.96954e-05, 6.383929e-05, 8.753939e-05, 
    6.680957e-05, 8.815047e-05, 8.220408e-05, 8.860244e-05, 9.119883e-05, 
    9.67577e-05, 5.096251e-05, 5.74549e-06, 2.830602e-06, 3.036792e-06,
  1.746036e-05, 2.187391e-05, 2.456075e-05, 5.165364e-05, 0.0001060002, 
    4.419932e-05, 6.313336e-05, 5.187561e-05, 6.938818e-05, 7.385591e-05, 
    9.147687e-05, 0.0001947019, 7.938161e-05, 5.489272e-06, 3.091702e-06,
  4.489212e-05, 2.007964e-05, 1.175571e-05, 5.547613e-05, 5.383514e-05, 
    4.509569e-05, 5.097539e-05, 5.048978e-05, 4.441569e-05, 5.000178e-05, 
    7.325375e-05, 0.0002089321, 0.0001195155, 1.3275e-05, 1.072491e-05,
  7.61398e-05, 3.832538e-05, 2.002256e-06, 3.064581e-05, 6.958659e-05, 
    7.244463e-05, 3.411022e-05, 2.896562e-05, 1.678759e-05, 1.278976e-05, 
    5.87843e-05, 0.0001365234, 6.275241e-05, 4.511428e-05, 3.004917e-05,
  8.644883e-05, 7.976455e-05, 1.270531e-05, 1.212582e-06, 1.849619e-05, 
    6.017558e-05, 4.73889e-05, 4.085505e-05, 1.660799e-05, 1.75224e-05, 
    2.747895e-05, 4.90295e-05, 5.761939e-05, 2.25519e-05, 2.434344e-05,
  0.0001010417, 6.488251e-05, 4.024302e-05, 2.635294e-05, 7.356542e-06, 
    2.630817e-05, 3.977929e-05, 4.573225e-05, 5.734675e-05, 5.028199e-05, 
    3.339742e-05, 4.24238e-05, 2.728595e-05, 6.070435e-05, 1.895023e-05,
  6.549012e-05, 7.612361e-05, 4.306557e-05, 2.508511e-05, 7.904415e-09, 
    6.971396e-06, 2.616764e-05, 5.440562e-05, 7.846141e-05, 6.701372e-05, 
    6.202739e-05, 4.210168e-05, 7.216037e-05, 8.160791e-06, 1.118505e-05,
  4.539367e-05, 8.583516e-05, 2.508675e-05, 8.419067e-06, 6.625214e-06, 
    6.06985e-09, 1.118283e-05, 4.805067e-05, 0.0001101531, 7.735246e-05, 
    8.860177e-05, 5.433048e-05, 1.410191e-05, 7.250706e-06, 3.255395e-05,
  2.575491e-05, 2.737913e-05, 9.491541e-06, 5.32685e-06, 1.716503e-06, 
    1.811582e-07, 3.327225e-07, 1.514785e-05, 6.177564e-05, 9.455017e-05, 
    0.0001035345, 5.532466e-05, 5.84778e-05, 2.494289e-05, 2.340042e-05,
  1.246935e-07, 3.222164e-05, 8.065372e-05, 0.0001346145, 0.0002280224, 
    0.0001536978, 5.277427e-05, 6.129132e-05, 8.1618e-05, 7.842873e-05, 
    7.182311e-05, 7.753444e-05, 5.405485e-05, 9.830124e-06, 7.321622e-06,
  0.0001033973, 3.943473e-08, 7.901622e-05, 0.0001449819, 0.0001848886, 
    0.0001338023, 0.000100829, 7.513611e-05, 5.373406e-05, 3.887393e-05, 
    2.865685e-05, 3.949513e-05, 2.002341e-05, 8.649661e-06, 1.039131e-05,
  0.0001216697, 0.0001062593, 6.538534e-05, 0.0001302908, 0.0001706886, 
    6.767488e-05, 8.569511e-05, 9.678893e-05, 4.101103e-05, 1.488803e-05, 
    2.603182e-05, 1.220498e-05, 1.847276e-05, 1.392637e-05, 1.131215e-05,
  0.0001132944, 0.0001059817, 9.990256e-07, 6.763348e-05, 9.359449e-05, 
    0.0001303118, 8.849093e-05, 7.378608e-05, 2.903501e-05, 1.844852e-05, 
    6.524036e-06, 1.544995e-05, 1.649857e-05, 2.960572e-05, 1.136962e-05,
  0.000138545, 0.0001215625, 1.476751e-05, 3.178193e-05, 8.454028e-05, 
    3.389508e-05, 7.525543e-05, 9.78729e-05, 3.724065e-05, 2.70807e-05, 
    3.046431e-05, 6.53287e-06, 1.941987e-05, 2.768759e-05, 3.722001e-05,
  0.0001174712, 0.0001173262, 9.928359e-05, 1.430092e-06, 2.767216e-05, 
    2.819316e-05, 8.304228e-05, 5.935297e-05, 1.36415e-05, 3.092032e-05, 
    2.772943e-05, 2.12058e-05, 4.070344e-05, 4.446146e-05, 7.771442e-05,
  0.000116721, 0.0001073516, 4.55437e-05, 5.432255e-05, 2.862607e-06, 
    1.20682e-05, 6.207615e-05, 7.082809e-06, 2.856436e-05, 4.032883e-05, 
    2.705329e-05, 1.450114e-05, 2.810915e-05, 3.724419e-05, 4.942884e-05,
  7.027666e-05, 0.0001085909, 7.551219e-05, 3.653009e-05, 4.003033e-08, 
    4.041722e-06, 1.678043e-05, 4.587163e-07, 1.928283e-05, 9.35646e-06, 
    1.560468e-05, 1.540708e-05, 8.385819e-06, 4.013725e-05, 3.731492e-05,
  5.779476e-05, 9.432593e-05, 7.465101e-05, 4.983592e-05, 2.725229e-05, 
    1.323967e-07, 1.790576e-05, 4.387913e-06, 1.04815e-05, 8.546613e-06, 
    2.036667e-05, 2.064327e-05, 1.590161e-05, 3.687124e-05, 5.443723e-05,
  1.835862e-05, 4.246801e-05, 1.941053e-05, 7.507212e-06, 2.648752e-05, 
    2.331965e-05, 9.735425e-07, 6.494315e-06, 6.402502e-06, 6.045897e-06, 
    1.52668e-05, 1.897816e-05, 2.224089e-05, 1.529504e-05, 4.391715e-05,
  2.821733e-05, 1.203799e-05, 9.964903e-05, 0.0001768089, 0.0001735896, 
    9.685129e-05, 5.35931e-05, 5.946059e-08, 5.964016e-07, 4.590489e-06, 
    6.556977e-06, 2.074205e-06, 4.401183e-07, 2.213673e-06, 7.193043e-06,
  0.000263957, 1.225248e-06, 4.822965e-05, 0.0001163165, 9.913772e-05, 
    4.208825e-05, 3.136172e-05, 2.041388e-07, 1.85129e-06, 4.530662e-06, 
    1.861244e-06, 2.93924e-06, 1.978563e-07, 1.900305e-06, 5.468866e-06,
  0.0002109344, 0.0002366328, 2.825984e-06, 5.895046e-05, 7.736974e-05, 
    9.610463e-06, 2.37499e-05, 1.165691e-05, 8.193741e-07, 1.628772e-06, 
    5.50769e-06, 5.222882e-06, 2.143945e-05, 6.972241e-06, 3.512332e-06,
  0.0001543339, 0.0001513379, 1.85038e-06, 1.223564e-06, 2.372253e-05, 
    3.577134e-05, 2.260575e-05, 7.16771e-06, 2.364613e-06, 1.533525e-06, 
    6.973926e-06, 1.225182e-05, 7.418149e-06, 8.852563e-06, 3.567999e-06,
  0.0001314876, 0.0001532638, 6.74538e-07, 2.31294e-08, 2.097345e-06, 
    8.187158e-06, 1.54752e-05, 8.73949e-06, 1.101395e-05, 1.692762e-05, 
    1.387957e-05, 1.372724e-05, 2.122385e-05, 2.467352e-05, 1.486151e-05,
  9.473543e-05, 0.0001528993, 0.0001793462, 6.91317e-08, 1.056266e-06, 
    4.766771e-06, 5.203658e-06, 3.256296e-06, 9.207088e-06, 1.419924e-05, 
    1.398778e-05, 2.478687e-05, 1.91711e-05, 2.006007e-05, 1.336452e-05,
  0.0001211304, 0.0001840641, 0.0001784264, 9.208019e-05, 4.429652e-07, 
    8.314668e-07, 6.591617e-07, 1.574653e-08, 2.489191e-05, 1.818175e-05, 
    1.322116e-05, 2.653599e-05, 2.641654e-05, 2.063249e-05, 2.578173e-05,
  0.0001695359, 0.0001806144, 0.0001900014, 9.517305e-05, 4.447051e-08, 
    4.751707e-09, 5.372009e-07, 1.207049e-09, 1.942951e-05, 1.325699e-05, 
    1.550545e-05, 2.759065e-05, 3.616892e-05, 3.286964e-05, 4.379458e-05,
  0.0001740193, 0.0001841174, 0.0001783117, 0.0001141221, 3.25095e-05, 
    2.790059e-08, 9.718599e-07, 4.737176e-06, 4.057513e-06, 6.737736e-06, 
    1.993284e-05, 2.632306e-05, 3.404064e-05, 5.315314e-05, 4.796442e-05,
  0.0002306536, 0.0001640913, 0.0001469711, 0.0001439558, 0.0001180356, 
    2.773935e-05, 5.413043e-10, 5.486225e-06, 5.124173e-06, 6.181045e-06, 
    1.122807e-05, 2.504072e-05, 2.771204e-05, 2.855312e-05, 5.144639e-05,
  1.019045e-05, 8.358862e-06, 8.318018e-06, 4.859153e-05, 3.950434e-05, 
    0.000120488, 0.0001954096, 0.0002863586, 0.0003669331, 0.0004394091, 
    0.0004377163, 0.0003958378, 0.0003046147, 0.0002034386, 0.0001251397,
  7.870254e-05, 4.45104e-06, 1.457353e-05, 2.790504e-05, 5.669777e-05, 
    5.53287e-05, 8.592236e-05, 9.107461e-05, 8.768185e-05, 8.699413e-05, 
    7.726101e-05, 5.859919e-05, 3.405348e-05, 1.71693e-05, 1.845565e-05,
  6.981686e-05, 0.0001005994, 2.184038e-05, 3.157164e-05, 6.986972e-05, 
    4.748247e-05, 1.54279e-05, 6.257777e-07, 2.844249e-07, 9.927247e-07, 
    6.683113e-07, 4.495779e-06, 7.886083e-06, 6.741855e-06, 5.917992e-06,
  0.0001074701, 0.0001348485, 5.603984e-05, 1.996683e-05, 2.036692e-05, 
    2.408448e-05, 7.316687e-06, 7.3474e-07, 7.787808e-07, 2.160354e-06, 
    5.595495e-07, 1.827608e-06, 2.357995e-06, 3.100391e-06, 1.477803e-06,
  9.914227e-05, 0.0001315617, 3.754917e-05, 1.271362e-06, 4.901748e-06, 
    1.879916e-05, 1.017314e-05, 1.176977e-05, 4.470655e-06, 5.78278e-06, 
    6.162561e-06, 1.702452e-06, 9.838011e-06, 4.557941e-07, 1.338427e-06,
  7.038545e-05, 0.0001214346, 0.0001410611, 3.417149e-06, 3.938304e-05, 
    8.772193e-05, 6.439938e-05, 3.256309e-05, 1.865051e-05, 1.564999e-05, 
    1.51522e-05, 1.621337e-06, 3.559658e-06, 1.65277e-06, 1.75356e-07,
  5.8507e-05, 0.0001412991, 0.0001791999, 0.0001274461, 0.00010078, 
    0.0001387899, 0.0001070841, 5.299637e-05, 2.145149e-05, 1.096461e-05, 
    5.613755e-06, 5.403823e-06, 2.447923e-06, 1.300977e-05, 1.518305e-06,
  5.95166e-05, 0.0001667147, 0.000282062, 0.0002563118, 5.181009e-05, 
    4.401865e-05, 2.90463e-05, 1.504105e-05, 1.776194e-06, 3.554131e-07, 
    2.758123e-06, 5.805964e-06, 5.478768e-06, 1.141912e-05, 6.944211e-06,
  7.681713e-05, 0.0001688295, 0.0003645043, 0.0003748771, 0.0001334491, 
    1.013999e-06, 1.934862e-07, 1.933805e-08, 1.459791e-07, 4.783258e-07, 
    6.214958e-06, 1.704166e-06, 7.875052e-06, 3.642486e-06, 1.079855e-05,
  0.0001610184, 0.0001534925, 0.0002165625, 0.0002375899, 0.0002303711, 
    0.0001267079, 1.107616e-07, 2.150528e-09, 2.818949e-07, 2.96606e-06, 
    2.569061e-06, 8.617984e-06, 1.331014e-05, 1.719153e-05, 1.634597e-05,
  4.589764e-06, 6.043737e-06, 5.150702e-06, 5.838574e-06, 5.341302e-06, 
    8.614372e-06, 1.68445e-05, 3.178319e-05, 8.664999e-05, 0.0001660889, 
    0.0003235604, 0.000488563, 0.0007065006, 0.0009352234, 0.001026727,
  1.006981e-05, 4.434491e-06, 6.582547e-06, 9.659784e-06, 3.308981e-05, 
    5.430188e-05, 9.826676e-05, 0.000165092, 0.0002563909, 0.0003634517, 
    0.0004602095, 0.0004941385, 0.0005266404, 0.0005553741, 0.0004541197,
  1.182408e-05, 1.828028e-05, 3.007724e-05, 3.791918e-05, 3.530037e-05, 
    4.698992e-05, 6.672785e-05, 7.534851e-05, 0.0001744575, 0.0003147409, 
    0.0004885303, 0.0006432094, 0.0006967422, 0.0005713627, 0.0002240721,
  3.178366e-05, 4.118591e-05, 4.920796e-05, 4.072552e-05, 7.023569e-05, 
    7.668383e-05, 7.530856e-05, 5.30344e-05, 8.705465e-05, 0.0002243189, 
    0.0004279893, 0.0007118776, 0.000884256, 0.0008667912, 0.0004166921,
  5.586033e-05, 5.968226e-05, 8.4696e-05, 2.948012e-05, 6.757722e-05, 
    0.000155231, 0.0001910131, 6.119189e-05, 2.571747e-05, 6.934609e-05, 
    0.0002277807, 0.0004713945, 0.0006981796, 0.0007169275, 0.0005789294,
  5.526535e-05, 0.0001020893, 6.053193e-05, 1.069059e-05, 2.303048e-05, 
    1.645971e-05, 3.353458e-05, 1.91566e-06, 1.446594e-06, 1.409994e-05, 
    5.76995e-05, 0.0001636377, 0.0002686834, 0.0003296252, 0.0002945549,
  5.196992e-05, 7.954834e-05, 8.79962e-05, 5.269774e-05, 3.636781e-07, 
    9.024979e-07, 1.50475e-06, 9.251296e-07, 1.196851e-06, 1.241981e-05, 
    1.263243e-05, 2.795666e-05, 2.803276e-05, 2.888821e-05, 2.08272e-05,
  8.517588e-05, 0.0001227269, 0.0001186425, 0.0001323048, 3.237085e-07, 
    1.550638e-06, 3.280368e-06, 4.319648e-06, 5.450165e-06, 2.756211e-06, 
    7.213491e-06, 4.761952e-06, 1.07315e-05, 5.391433e-06, 1.230439e-05,
  0.0001815624, 0.0002614852, 0.0002824248, 0.0001917976, 0.000115023, 
    1.447514e-06, 2.75775e-06, 1.727666e-06, 5.171341e-07, 1.131522e-06, 
    5.942575e-06, 2.096804e-06, 5.628985e-06, 4.4981e-06, 4.573596e-06,
  0.0002285449, 0.0003197501, 0.0003260378, 0.0002751515, 0.0001120428, 
    0.0001108844, 6.144865e-08, 3.830659e-08, 4.104425e-07, 9.66682e-07, 
    1.539785e-07, 1.742923e-05, 2.036798e-05, 2.284276e-05, 8.036094e-06,
  1.941246e-06, 1.883025e-05, 1.254114e-05, 1.355151e-05, 4.142915e-06, 
    2.832196e-06, 2.54345e-06, 3.489538e-06, 5.033542e-06, 7.039783e-06, 
    9.516988e-06, 1.488273e-05, 8.674774e-05, 0.0005952108, 0.0009640421,
  3.323356e-05, 1.740395e-05, 1.867512e-05, 1.062484e-05, 1.238104e-05, 
    4.650623e-06, 3.959625e-06, 4.373592e-06, 4.911872e-06, 5.125157e-06, 
    8.495858e-06, 1.243911e-05, 6.921669e-05, 0.0003046439, 0.0005125834,
  4.189657e-05, 3.910235e-05, 2.619267e-05, 3.765547e-05, 2.470773e-05, 
    2.453128e-05, 2.146274e-05, 1.324284e-05, 8.515579e-06, 1.321732e-05, 
    3.636719e-05, 1.545748e-05, 5.916862e-05, 0.0001184175, 0.0001075323,
  3.085573e-05, 2.744675e-05, 2.760716e-05, 3.685704e-05, 4.716308e-05, 
    6.810528e-05, 7.627875e-05, 5.964889e-05, 6.09606e-05, 4.781271e-05, 
    2.996054e-05, 2.353985e-05, 5.183295e-05, 3.907004e-05, 3.64233e-05,
  3.869185e-05, 3.588185e-05, 2.342911e-05, 8.321364e-06, 1.913413e-05, 
    3.191417e-05, 5.37324e-05, 5.317271e-05, 3.258677e-05, 4.759003e-05, 
    5.797064e-05, 5.374659e-05, 5.963771e-05, 9.277486e-05, 9.629171e-05,
  3.411778e-05, 2.749005e-05, 2.792495e-05, 6.277441e-06, 5.430979e-06, 
    4.974452e-06, 1.886627e-05, 1.263548e-05, 1.506455e-07, 4.004343e-05, 
    5.11839e-05, 4.869306e-05, 7.506121e-05, 0.0001218198, 0.0001530695,
  8.209391e-05, 5.155439e-05, 4.6073e-05, 1.783659e-05, 1.951952e-06, 
    3.895305e-07, 2.589031e-06, 2.153313e-06, 8.541558e-06, 1.496965e-05, 
    3.230438e-05, 7.289287e-05, 9.684172e-05, 0.0001355367, 0.0001155653,
  0.0001357949, 9.874668e-05, 0.0001061501, 6.825706e-05, 8.034908e-07, 
    5.770489e-09, 3.613901e-06, 9.911228e-09, 8.329496e-06, 1.135272e-05, 
    1.980389e-05, 5.366016e-05, 7.257889e-05, 6.923333e-05, 4.065068e-05,
  0.0001790792, 0.0002012736, 0.0001141485, 0.0001292184, 7.487123e-05, 
    9.683087e-08, 2.899034e-06, 2.448704e-08, 1.557292e-05, 1.400393e-05, 
    1.266392e-05, 3.242787e-05, 4.988041e-05, 3.499059e-05, 4.370729e-05,
  0.0001626752, 0.0001618871, 0.0002691837, 0.0001728943, 0.0001057775, 
    6.105095e-05, 3.783133e-07, 2.078463e-05, 1.552876e-05, 1.285774e-05, 
    1.708633e-05, 3.339415e-05, 3.370747e-05, 4.096425e-05, 2.291003e-05,
  5.807102e-08, 3.004356e-06, 6.668535e-06, 7.648691e-06, 3.945925e-05, 
    5.311245e-05, 4.500956e-05, 1.369094e-05, 5.035707e-06, 6.397674e-06, 
    1.43535e-05, 7.325091e-06, 7.377864e-06, 9.006695e-06, 1.380527e-05,
  1.635076e-05, 3.6623e-06, 7.090122e-06, 3.258146e-06, 1.482686e-05, 
    3.079127e-05, 3.274342e-05, 1.779012e-05, 3.495664e-05, 2.104021e-05, 
    1.400015e-05, 1.727464e-05, 9.904576e-06, 1.018163e-05, 1.919324e-05,
  2.606667e-05, 2.68823e-05, 1.817644e-06, 1.857002e-06, 1.77121e-06, 
    1.353882e-05, 2.942064e-05, 2.857575e-05, 2.739074e-05, 3.901362e-05, 
    3.725239e-05, 2.493515e-05, 8.207585e-06, 2.964937e-06, 3.719889e-06,
  3.521795e-05, 3.942066e-05, 6.060109e-07, 2.197803e-06, 1.26522e-06, 
    5.939077e-07, 9.545411e-07, 5.789221e-06, 1.148539e-05, 2.457951e-05, 
    3.233255e-05, 3.542241e-05, 7.00394e-06, 4.95335e-06, 2.345261e-06,
  5.176008e-05, 8.369964e-05, 1.069882e-05, 6.14873e-07, 1.057847e-06, 
    8.16894e-07, 1.601358e-06, 8.441782e-07, 7.28064e-07, 2.008108e-05, 
    3.364951e-05, 3.480714e-05, 1.51607e-05, 3.124602e-05, 3.878544e-07,
  7.739534e-05, 7.733377e-05, 7.856749e-05, 1.052904e-07, 6.733117e-07, 
    9.107184e-07, 7.183744e-07, 1.213536e-06, 7.599178e-06, 6.319124e-06, 
    2.369621e-05, 3.486456e-05, 3.899396e-05, 2.372849e-05, 1.146652e-05,
  0.0001168446, 0.0001011152, 0.000117045, 6.688495e-05, 1.043609e-07, 
    4.361514e-07, 2.604632e-07, 6.556516e-07, 6.372991e-07, 2.963949e-06, 
    1.03328e-05, 2.627252e-05, 3.031545e-05, 2.171873e-05, 1.292943e-05,
  0.00013861, 0.0001784288, 0.0001672936, 0.0001063731, 1.42044e-08, 
    6.031672e-08, 7.520296e-07, 1.699867e-09, 9.60279e-07, 2.728531e-06, 
    7.748876e-06, 9.570426e-06, 1.664705e-05, 1.035021e-05, 1.397294e-05,
  0.0001969481, 0.0002472312, 0.0002233217, 7.909987e-05, 6.68798e-05, 
    7.513379e-06, 1.25068e-06, 1.549024e-07, 5.856818e-07, 1.662567e-06, 
    1.123501e-05, 1.953973e-05, 1.216644e-05, 1.930896e-05, 1.050082e-05,
  0.0001487313, 0.0002489569, 0.0001610193, 2.423218e-05, 7.157459e-05, 
    5.673747e-05, 4.28281e-09, 1.906975e-06, 8.139933e-07, 3.427703e-06, 
    2.648527e-06, 6.36805e-06, 1.132823e-05, 1.107074e-05, 9.170934e-06,
  4.642545e-06, 5.126722e-06, 5.001518e-06, 2.86674e-05, 3.963496e-05, 
    4.128538e-05, 2.836552e-05, 3.707032e-05, 5.535703e-05, 6.601364e-05, 
    7.541675e-05, 9.986579e-05, 0.0001064921, 0.0001240876, 0.0001717622,
  9.256805e-06, 3.03573e-06, 3.834545e-06, 2.307191e-05, 2.984252e-05, 
    3.923438e-05, 4.373389e-05, 3.422281e-05, 4.765101e-05, 7.634346e-05, 
    8.848825e-05, 0.0001070535, 0.0001229172, 0.0001522618, 0.0001911374,
  1.479828e-05, 1.226199e-05, 2.871325e-06, 1.148051e-05, 3.02459e-05, 
    1.607936e-05, 3.942934e-05, 3.261077e-05, 8.450518e-05, 0.0001031542, 
    7.759851e-05, 9.579715e-05, 0.0001037512, 0.0001136103, 0.0001225433,
  3.244254e-05, 2.118109e-05, 4.647879e-06, 1.774789e-06, 1.602286e-05, 
    2.836042e-05, 6.920614e-05, 5.713663e-05, 2.949841e-05, 8.650465e-05, 
    4.135939e-05, 3.94461e-05, 3.008419e-05, 3.116439e-05, 2.771393e-05,
  3.279785e-05, 4.083054e-05, 9.5553e-06, 3.626983e-06, 1.669938e-06, 
    2.136653e-05, 3.102244e-05, 6.86479e-05, 5.371649e-05, 9.500733e-05, 
    2.772997e-05, 3.6029e-05, 2.466271e-05, 1.864451e-05, 1.711437e-05,
  4.021256e-05, 4.385997e-05, 4.086141e-05, 4.79123e-06, 6.052023e-06, 
    1.048896e-05, 2.839013e-05, 5.538169e-05, 5.768595e-05, 4.392657e-05, 
    7.62694e-05, 2.265424e-06, 6.488107e-06, 4.190518e-06, 8.485603e-06,
  2.810548e-05, 2.207686e-05, 3.580971e-05, 4.323719e-05, 6.670788e-06, 
    4.968314e-06, 1.454764e-05, 4.667788e-05, 4.732024e-05, 2.599126e-05, 
    2.653514e-06, 4.578901e-06, 1.439279e-06, 4.710583e-06, 1.075568e-05,
  1.99815e-05, 3.032411e-05, 3.61866e-05, 4.156875e-05, 1.654767e-05, 
    2.489233e-06, 4.59174e-06, 1.4443e-05, 2.503063e-05, 2.402013e-05, 
    1.389534e-05, 1.917956e-05, 2.521372e-05, 1.599488e-05, 6.838925e-06,
  3.436539e-05, 5.274616e-05, 4.680725e-05, 5.091531e-05, 4.098044e-05, 
    4.426562e-06, 2.816469e-07, 5.839553e-06, 3.115673e-05, 5.108686e-05, 
    3.671242e-05, 2.692184e-05, 1.763426e-05, 2.131716e-05, 3.031837e-05,
  5.974244e-05, 8.604277e-05, 0.0001203491, 8.15777e-05, 4.332381e-05, 
    4.800286e-05, 6.526952e-08, 7.620272e-06, 9.770724e-06, 6.283774e-05, 
    8.588488e-05, 6.238474e-05, 3.649286e-05, 2.940832e-05, 2.871178e-05,
  9.524071e-07, 2.746317e-06, 3.472181e-06, 3.456126e-06, 3.671319e-06, 
    4.222245e-06, 4.916666e-06, 5.08579e-06, 6.109818e-06, 6.903337e-06, 
    8.867441e-06, 1.044296e-05, 2.120486e-05, 2.209397e-05, 4.237209e-05,
  1.29598e-06, 3.260586e-07, 2.009495e-06, 3.204537e-06, 2.12756e-06, 
    1.742941e-06, 3.008888e-06, 3.75746e-06, 4.456477e-06, 4.876081e-06, 
    5.351977e-06, 8.159108e-06, 1.438823e-05, 2.478047e-05, 7.582506e-05,
  2.974416e-07, 1.094585e-06, 1.32892e-06, 2.330135e-06, 1.133835e-06, 
    7.764287e-07, 1.636452e-06, 2.367066e-06, 5.512942e-06, 4.598177e-06, 
    8.91417e-06, 3.101994e-05, 7.318285e-05, 0.0001361911, 0.0002401706,
  1.466863e-07, 6.932192e-07, 1.911607e-06, 2.526602e-06, 2.000679e-06, 
    2.292621e-06, 2.006328e-06, 2.221455e-06, 2.068692e-06, 3.352322e-06, 
    1.017519e-05, 5.461233e-05, 0.0001169833, 0.0001886702, 0.0002618462,
  1.023357e-06, 2.348129e-06, 3.206225e-06, 4.980881e-06, 4.163104e-06, 
    3.176996e-06, 1.942757e-06, 1.70808e-06, 1.637784e-06, 5.033377e-06, 
    2.235711e-05, 6.657189e-05, 0.0001219201, 0.0001702323, 0.0002270255,
  5.096098e-06, 5.712459e-06, 6.680588e-06, 4.410535e-06, 3.606649e-06, 
    3.624395e-06, 3.302986e-06, 5.110546e-06, 9.59909e-06, 3.107766e-05, 
    5.890323e-05, 8.069833e-05, 9.561011e-05, 0.000107062, 0.0001549904,
  5.379793e-06, 8.741678e-06, 1.222411e-05, 9.794778e-06, 7.091412e-06, 
    7.443964e-06, 9.014363e-06, 1.006225e-05, 1.996064e-05, 6.662451e-05, 
    0.0001168545, 0.0001140625, 9.744376e-05, 0.0002126119, 0.0002694618,
  5.082356e-06, 8.453121e-06, 7.947848e-06, 1.800828e-05, 1.690347e-05, 
    1.393915e-05, 9.454532e-06, 2.352814e-05, 5.358185e-05, 4.524873e-05, 
    7.098162e-05, 0.0001099424, 0.0002809414, 0.0003355742, 0.0005332532,
  1.090379e-05, 1.922032e-05, 1.431649e-05, 1.465662e-05, 2.326943e-05, 
    2.558588e-05, 2.492156e-05, 1.690014e-05, 3.052708e-05, 4.377262e-05, 
    7.112967e-05, 0.0001919579, 0.0004790249, 0.0005205508, 0.0006795948,
  8.835093e-06, 1.404524e-05, 3.504573e-05, 5.151451e-05, 3.781761e-05, 
    3.660591e-05, 2.268105e-05, 2.237062e-05, 2.864223e-05, 3.563437e-05, 
    8.419323e-05, 0.0002507705, 0.0004988892, 0.0005642272, 0.0005808607,
  1.975e-09, 3.775485e-09, 1.1807e-07, 9.802262e-07, 3.169576e-06, 
    1.45363e-05, 1.861187e-05, 7.443841e-06, 2.756366e-06, 7.269176e-07, 
    6.666359e-07, 6.417741e-07, 1.831494e-06, 1.70271e-06, 1.8125e-06,
  1.991792e-07, 2.537019e-08, 1.433594e-07, 7.387353e-07, 1.543088e-06, 
    3.664734e-06, 1.332231e-05, 1.032024e-05, 9.122654e-06, 2.427688e-06, 
    6.473909e-07, 1.104972e-06, 1.09003e-06, 1.393122e-06, 1.589943e-06,
  1.466448e-06, 1.810077e-06, 5.456156e-07, 8.166555e-08, 5.930609e-07, 
    2.016059e-06, 4.855896e-06, 6.645218e-06, 5.273802e-06, 6.165005e-06, 
    7.417305e-07, 9.929619e-07, 1.157014e-06, 9.198594e-07, 1.373218e-06,
  2.831367e-06, 1.959728e-06, 1.049147e-06, 1.096366e-06, 7.124677e-07, 
    2.291581e-06, 3.650646e-06, 3.615912e-06, 4.408789e-06, 3.776672e-06, 
    1.802566e-06, 1.740577e-06, 1.212286e-06, 5.591062e-07, 3.945725e-07,
  1.59756e-06, 2.907092e-06, 1.659855e-06, 3.71917e-06, 2.689343e-06, 
    2.792593e-06, 3.616197e-06, 2.686151e-06, 2.927204e-06, 3.679668e-06, 
    1.273959e-06, 4.821903e-07, 4.794393e-07, 4.365888e-07, 3.361325e-07,
  7.669381e-07, 1.944692e-06, 3.376562e-06, 2.195113e-06, 4.572055e-06, 
    3.964419e-06, 4.15938e-06, 3.771075e-06, 3.654606e-06, 4.049246e-06, 
    1.339485e-06, 3.729718e-07, 3.483155e-07, 3.441071e-07, 4.64196e-07,
  1.044581e-06, 2.058484e-06, 4.299523e-06, 6.773619e-06, 4.912357e-06, 
    4.449548e-06, 3.282221e-06, 4.757647e-06, 6.181093e-06, 3.130674e-06, 
    6.966207e-07, 2.71494e-07, 2.004943e-07, 3.521558e-07, 6.053528e-07,
  9.808582e-07, 1.814623e-06, 2.649949e-06, 5.330274e-06, 5.924531e-06, 
    5.000919e-06, 4.877725e-06, 4.569832e-06, 8.622854e-06, 4.150547e-06, 
    3.16532e-06, 1.691567e-06, 1.399816e-06, 1.361965e-06, 5.450732e-07,
  2.92085e-07, 2.111848e-06, 4.204158e-06, 5.302027e-06, 8.195627e-06, 
    7.104033e-06, 7.413651e-06, 5.918587e-06, 8.461467e-06, 4.047224e-06, 
    2.212248e-06, 2.856061e-06, 2.176743e-06, 2.088242e-06, 1.498193e-06,
  3.80277e-09, 1.961452e-07, 2.328627e-06, 9.145429e-06, 8.742403e-06, 
    1.138442e-05, 9.768842e-06, 7.685513e-06, 9.47748e-06, 5.580444e-06, 
    2.301257e-06, 2.44108e-06, 2.076883e-06, 2.739588e-06, 2.703867e-06,
  2.894318e-06, 4.848016e-06, 1.274037e-05, 1.680619e-05, 1.377887e-05, 
    1.22269e-05, 1.007007e-05, 6.089156e-06, 3.467353e-06, 5.395901e-06, 
    4.816106e-06, 6.27408e-06, 7.884333e-06, 7.513795e-06, 9.403221e-06,
  1.580276e-05, 9.531337e-06, 1.696462e-05, 1.58091e-05, 1.27279e-05, 
    9.281489e-06, 1.043614e-05, 6.233077e-06, 3.949424e-06, 4.005447e-06, 
    2.990725e-06, 4.843919e-06, 6.52742e-06, 7.774177e-06, 9.720332e-06,
  1.082155e-05, 1.733224e-05, 1.670947e-05, 1.766255e-05, 1.5123e-05, 
    9.077671e-06, 7.530801e-06, 6.176725e-06, 5.018332e-06, 4.538656e-06, 
    4.006834e-06, 2.698969e-06, 3.679891e-06, 5.147742e-06, 7.588069e-06,
  1.023453e-05, 1.265341e-05, 1.235615e-05, 1.815743e-05, 1.033434e-05, 
    1.294974e-05, 9.366099e-06, 8.146212e-06, 3.401348e-06, 5.248379e-06, 
    4.698769e-06, 2.205361e-06, 2.063494e-06, 1.805969e-06, 2.747249e-06,
  5.572616e-06, 1.063649e-05, 9.19656e-06, 1.291659e-05, 1.578059e-05, 
    1.402085e-05, 1.16439e-05, 8.942859e-06, 7.907612e-06, 5.972983e-06, 
    5.814162e-06, 5.684713e-06, 4.036916e-06, 1.864651e-06, 1.313436e-06,
  4.40883e-06, 7.320954e-06, 1.204666e-05, 7.649608e-06, 1.363084e-05, 
    1.541233e-05, 1.229877e-05, 1.179018e-05, 9.399818e-06, 7.3053e-06, 
    8.448378e-06, 6.170061e-06, 3.101748e-06, 2.677156e-06, 1.710474e-06,
  2.24772e-06, 5.73038e-06, 1.093821e-05, 1.435245e-05, 1.227143e-05, 
    1.477603e-05, 1.249295e-05, 1.119614e-05, 1.402795e-05, 1.073376e-05, 
    7.95803e-06, 8.144891e-06, 6.120749e-06, 5.53277e-06, 2.569769e-06,
  1.327488e-06, 4.199906e-06, 6.316343e-06, 1.278846e-05, 1.002139e-05, 
    1.201331e-05, 1.340768e-05, 1.241444e-05, 1.387676e-05, 1.023683e-05, 
    1.002974e-05, 7.190451e-06, 9.997329e-06, 5.297018e-06, 5.30371e-06,
  1.201729e-06, 4.877065e-06, 6.870614e-06, 8.515612e-06, 1.5218e-05, 
    1.183123e-05, 1.407473e-05, 1.156427e-05, 1.426117e-05, 9.266152e-06, 
    9.225991e-06, 7.956662e-06, 6.90528e-06, 5.825565e-06, 7.274249e-06,
  7.135719e-07, 2.547368e-06, 6.955595e-06, 1.204557e-05, 8.248544e-06, 
    1.712841e-05, 1.744845e-05, 1.700734e-05, 1.387021e-05, 1.558977e-05, 
    1.033435e-05, 1.196842e-05, 1.454027e-05, 2.959727e-06, 3.711571e-06,
  4.21571e-06, 4.741584e-06, 8.642464e-06, 1.208801e-05, 8.301291e-06, 
    7.556623e-06, 6.536583e-06, 6.634095e-06, 5.594877e-06, 5.94883e-06, 
    6.352906e-06, 5.826422e-06, 6.473758e-06, 1.001814e-05, 6.220255e-06,
  2.71828e-05, 1.105801e-05, 1.614063e-05, 1.319172e-05, 8.101051e-06, 
    6.932985e-06, 5.5916e-06, 5.794891e-06, 5.060672e-06, 7.511132e-06, 
    6.614727e-06, 7.169042e-06, 1.05327e-05, 1.403905e-05, 1.390443e-05,
  2.057753e-05, 2.331259e-05, 1.558151e-05, 1.378161e-05, 8.175671e-06, 
    6.363573e-06, 5.927903e-06, 5.739973e-06, 5.939929e-06, 5.135754e-06, 
    4.871467e-06, 5.903368e-06, 7.297229e-06, 1.324491e-05, 1.828946e-05,
  2.225957e-05, 1.90454e-05, 1.207076e-05, 1.427842e-05, 1.07645e-05, 
    7.242516e-06, 7.213333e-06, 6.18177e-06, 5.157604e-06, 5.772799e-06, 
    7.823405e-06, 6.550824e-06, 6.729982e-06, 7.709335e-06, 1.146966e-05,
  1.199914e-05, 1.481474e-05, 1.663342e-05, 1.519196e-05, 1.329371e-05, 
    8.945319e-06, 7.935424e-06, 6.804093e-06, 5.163417e-06, 6.903848e-06, 
    7.85724e-06, 7.735674e-06, 8.251768e-06, 8.043194e-06, 9.140967e-06,
  5.550971e-06, 1.080106e-05, 1.574593e-05, 9.362113e-06, 1.332093e-05, 
    1.08647e-05, 8.088556e-06, 7.13319e-06, 6.17464e-06, 8.291297e-06, 
    7.360381e-06, 9.826089e-06, 1.108648e-05, 1.204784e-05, 1.312906e-05,
  4.066251e-06, 7.437156e-06, 1.423247e-05, 1.696845e-05, 1.358597e-05, 
    1.246961e-05, 7.903279e-06, 6.800758e-06, 1.008858e-05, 8.779446e-06, 
    1.071489e-05, 1.40122e-05, 1.433233e-05, 1.15566e-05, 1.221528e-05,
  1.676667e-06, 5.613657e-06, 9.543155e-06, 1.447675e-05, 9.28377e-06, 
    1.094624e-05, 9.47871e-06, 7.678588e-06, 1.052961e-05, 1.141773e-05, 
    1.581542e-05, 1.478339e-05, 1.177764e-05, 1.577957e-05, 3.849914e-05,
  1.486512e-06, 2.80644e-06, 8.013825e-06, 1.110251e-05, 1.445952e-05, 
    1.049744e-05, 1.101529e-05, 9.889093e-06, 1.421992e-05, 1.801941e-05, 
    2.421722e-05, 2.948541e-05, 7.370381e-05, 0.0002441676, 0.0003051198,
  1.161819e-06, 1.040008e-06, 4.175109e-06, 1.200707e-05, 7.763243e-06, 
    1.877314e-05, 1.105811e-05, 1.411526e-05, 1.296049e-05, 2.356925e-05, 
    3.119344e-05, 6.155712e-05, 0.0002403181, 0.0004543327, 0.0004855225,
  4.209784e-07, 6.602968e-07, 1.342603e-06, 3.604017e-06, 3.861826e-06, 
    3.910408e-06, 3.952023e-06, 3.677107e-06, 4.792792e-06, 6.265662e-06, 
    5.719687e-06, 6.985583e-06, 7.107051e-06, 5.344554e-06, 3.539053e-06,
  4.853966e-06, 1.818738e-06, 3.523499e-06, 4.493577e-06, 3.530065e-06, 
    3.637013e-06, 4.758265e-06, 4.847208e-06, 4.587539e-06, 4.588801e-06, 
    5.855059e-06, 7.282697e-06, 6.985285e-06, 6.647185e-06, 1.197425e-05,
  3.014512e-06, 5.444651e-06, 3.308323e-06, 4.814818e-06, 4.41323e-06, 
    3.949107e-06, 5.056221e-06, 5.286409e-06, 5.544031e-06, 6.222584e-06, 
    7.054867e-06, 9.945644e-06, 1.1825e-05, 4.385312e-05, 0.0001059816,
  3.264523e-06, 4.031321e-06, 2.673345e-06, 4.216696e-06, 6.137413e-06, 
    5.288974e-06, 6.255577e-06, 5.339126e-06, 5.593055e-06, 7.408777e-06, 
    1.295435e-05, 1.792332e-05, 3.098258e-05, 0.000182739, 0.0002825347,
  1.708253e-06, 3.659942e-06, 3.540622e-06, 4.242145e-06, 5.262415e-06, 
    4.495474e-06, 5.263644e-06, 5.005701e-06, 5.771805e-06, 1.161072e-05, 
    1.903036e-05, 2.490895e-05, 9.066885e-05, 0.0003784541, 0.000442816,
  6.394725e-07, 3.146442e-06, 5.692771e-06, 2.718514e-06, 3.730902e-06, 
    4.058359e-06, 2.931828e-06, 4.395854e-06, 7.369919e-06, 1.759758e-05, 
    2.851648e-05, 3.533942e-05, 0.0001680518, 0.0005053282, 0.0005357618,
  4.006765e-07, 2.567807e-06, 5.149053e-06, 6.846385e-06, 3.722521e-06, 
    3.170769e-06, 2.038678e-06, 4.719302e-06, 1.763314e-05, 2.599532e-05, 
    3.344694e-05, 4.827315e-05, 0.000221447, 0.0005348091, 0.0005275332,
  1.673387e-07, 1.902669e-06, 3.052083e-06, 4.342233e-06, 3.824729e-06, 
    1.54757e-06, 2.277546e-06, 7.663219e-06, 3.237382e-05, 4.320034e-05, 
    5.008938e-05, 7.013414e-05, 0.000263813, 0.0005135703, 0.0005312603,
  1.769061e-08, 1.149998e-06, 1.896248e-06, 3.093466e-06, 6.292858e-06, 
    2.491598e-06, 6.785183e-06, 1.978595e-05, 5.104261e-05, 7.652288e-05, 
    6.821274e-05, 0.0001097472, 0.0002731443, 0.00043466, 0.0003865133,
  2.828068e-10, 2.160105e-07, 3.30796e-06, 6.979466e-06, 8.131487e-06, 
    1.640179e-05, 1.416313e-05, 4.233575e-05, 7.330978e-05, 7.496113e-05, 
    7.155984e-05, 0.0001211025, 0.0002300446, 0.000279457, 0.0002397341,
  1.561869e-06, 1.134345e-06, 1.646177e-06, 1.622975e-06, 2.20057e-06, 
    3.026633e-06, 2.629651e-06, 2.183952e-06, 2.801754e-07, 7.619841e-07, 
    3.624741e-06, 6.077624e-06, 9.109465e-06, 8.342066e-06, 1.131868e-05,
  1.008529e-05, 1.318898e-08, 5.910638e-07, 1.092238e-06, 7.090849e-07, 
    1.208459e-06, 2.190032e-06, 1.255329e-06, 4.084355e-07, 1.633088e-06, 
    5.578761e-06, 9.449033e-06, 1.490007e-05, 3.297221e-05, 9.242511e-05,
  4.447107e-06, 7.35373e-06, 2.363799e-07, 9.171457e-07, 3.533421e-07, 
    5.005085e-07, 3.341744e-07, 3.706491e-07, 1.861615e-06, 4.018244e-06, 
    9.279827e-06, 1.726054e-05, 2.994546e-05, 0.0001370302, 0.0001281385,
  4.410797e-06, 5.013354e-06, 6.902147e-07, 8.834535e-07, 2.566699e-07, 
    4.972082e-07, 2.550825e-07, 1.483517e-06, 2.279377e-06, 7.22677e-06, 
    1.54617e-05, 2.012668e-05, 5.156504e-05, 0.0001612223, 7.061826e-05,
  1.695843e-08, 2.138264e-07, 2.144947e-09, 1.279697e-07, 7.111144e-07, 
    2.377662e-07, 4.366847e-07, 1.445987e-06, 3.618259e-06, 8.044474e-06, 
    1.578831e-05, 2.203487e-05, 4.01002e-05, 7.05291e-05, 4.560851e-05,
  2.834876e-10, 1.999216e-08, 1.550144e-07, 2.420469e-07, 4.557532e-07, 
    1.84949e-07, 9.695511e-07, 1.946049e-06, 4.303782e-06, 9.736789e-06, 
    1.459259e-05, 1.977605e-05, 2.022518e-05, 2.177245e-05, 3.227437e-05,
  2.946676e-13, 4.762112e-08, 2.271767e-07, 4.227893e-07, 5.339328e-09, 
    2.62916e-07, 1.425232e-06, 1.700823e-06, 5.046304e-06, 9.069063e-06, 
    1.455882e-05, 2.2505e-05, 1.924453e-05, 1.352757e-05, 2.038017e-05,
  1.703911e-11, 3.650831e-10, 7.958109e-08, 3.646192e-07, 9.986981e-08, 
    1.681799e-07, 5.235872e-07, 1.681809e-06, 6.727443e-06, 9.239e-06, 
    1.49322e-05, 2.591157e-05, 1.803007e-05, 1.571016e-05, 1.984189e-05,
  1.230088e-08, 8.769733e-10, 1.012493e-10, 2.300211e-10, 3.652807e-07, 
    6.037727e-08, 6.09771e-07, 1.839059e-06, 5.850107e-06, 1.077498e-05, 
    1.782232e-05, 2.681925e-05, 1.806021e-05, 1.562529e-05, 1.956016e-05,
  3.400115e-07, 2.085458e-07, 3.32014e-09, 2.380476e-10, 2.593626e-10, 
    7.178821e-07, 7.115308e-07, 2.369459e-06, 5.939205e-06, 8.605761e-06, 
    1.136982e-05, 2.421655e-05, 2.288913e-05, 1.90202e-05, 2.651987e-05,
  3.049609e-06, 2.252629e-06, 7.007061e-06, 5.632988e-05, 4.367945e-05, 
    5.56326e-05, 7.687954e-05, 0.000100811, 0.0002020115, 0.0001460469, 
    0.0001490338, 8.506408e-05, 0.0001520209, 0.0001174527, 7.393198e-05,
  4.244943e-06, 6.509795e-06, 5.057007e-06, 2.131704e-05, 4.394909e-05, 
    4.913957e-05, 6.528412e-05, 5.769488e-05, 0.0001630303, 0.0001884039, 
    0.0001377314, 8.703795e-05, 0.0001258673, 8.923232e-05, 7.427244e-05,
  2.431214e-05, 4.15546e-06, 6.883e-06, 2.465276e-05, 3.345251e-05, 
    5.4869e-05, 7.286374e-05, 7.361604e-05, 7.381719e-05, 0.0001192645, 
    0.0001396146, 8.616887e-05, 4.450488e-05, 2.584593e-05, 2.602192e-05,
  2.718695e-05, 2.863714e-05, 4.321556e-05, 4.691527e-05, 6.12779e-05, 
    4.519136e-05, 4.901772e-05, 5.549657e-05, 3.963235e-05, 4.125871e-05, 
    6.05999e-05, 3.288924e-05, 3.129175e-05, 1.964495e-05, 4.061041e-05,
  2.679845e-05, 4.663317e-05, 2.889496e-05, 3.277351e-05, 5.430253e-05, 
    4.383146e-05, 4.025563e-05, 2.745382e-05, 3.53824e-05, 4.134879e-05, 
    3.687718e-05, 3.13612e-05, 3.387865e-05, 2.990098e-05, 3.234334e-05,
  2.479599e-06, 2.498735e-05, 3.909221e-05, 1.238405e-05, 2.4254e-05, 
    2.607019e-05, 2.8732e-05, 2.087471e-05, 1.731267e-05, 2.202147e-05, 
    2.12259e-05, 2.964885e-05, 2.6923e-05, 1.938548e-05, 1.187143e-05,
  2.809088e-08, 5.954084e-06, 9.818154e-06, 1.043245e-05, 4.010271e-06, 
    4.955584e-06, 1.515549e-05, 1.532503e-05, 1.642765e-05, 2.154965e-05, 
    2.281798e-05, 1.818519e-05, 7.592839e-06, 5.078055e-06, 4.30925e-06,
  2.946158e-10, 7.16309e-10, 5.007047e-08, 6.709524e-08, 4.902026e-10, 
    3.038939e-09, 3.213985e-07, 2.745063e-06, 1.780294e-06, 2.78635e-06, 
    3.26075e-06, 2.872946e-06, 1.449554e-06, 9.701112e-07, 1.231817e-06,
  9.808594e-11, 1.817861e-09, 6.256477e-11, 3.586747e-08, 9.112711e-08, 
    7.293334e-08, 2.792093e-06, 2.929858e-06, 2.787933e-06, 1.931181e-06, 
    1.477654e-06, 1.10624e-06, 4.079012e-06, 3.01247e-06, 3.135955e-06,
  1.440371e-08, 1.131371e-08, 1.456342e-09, 8.513803e-11, 5.673515e-09, 
    1.450434e-07, 4.038675e-06, 3.226543e-06, 5.716695e-06, 2.672848e-06, 
    2.935377e-06, 4.364922e-06, 4.16255e-06, 2.702103e-06, 2.420472e-06,
  3.338845e-08, 1.395053e-06, 6.211282e-08, 5.797066e-07, 3.90915e-07, 
    4.037354e-07, 4.509273e-07, 7.205248e-07, 5.668635e-07, 1.14661e-06, 
    2.993921e-06, 2.943729e-06, 2.927125e-06, 2.231952e-06, 2.161862e-06,
  2.027052e-07, 8.355741e-07, 5.706688e-07, 5.03593e-07, 5.837123e-07, 
    5.159071e-07, 5.937014e-07, 6.154936e-07, 4.065263e-07, 1.975801e-06, 
    1.298829e-06, 3.34014e-06, 2.768604e-06, 2.466267e-06, 2.005901e-06,
  1.041736e-05, 4.486733e-06, 2.769169e-06, 2.003165e-06, 1.902043e-06, 
    1.547601e-06, 7.88003e-07, 5.832114e-07, 4.817368e-07, 1.419711e-06, 
    1.154896e-06, 2.560552e-06, 1.91196e-06, 1.815672e-06, 1.605416e-06,
  2.220339e-05, 9.979773e-06, 6.719958e-06, 4.012075e-06, 1.144451e-06, 
    2.794335e-06, 3.257444e-06, 2.101833e-06, 1.557091e-06, 1.230085e-06, 
    1.868218e-06, 5.881537e-07, 6.655326e-07, 3.507407e-07, 4.170884e-07,
  4.534309e-05, 1.551335e-05, 1.047646e-05, 8.346646e-06, 2.978651e-06, 
    2.146179e-06, 8.944193e-07, 1.450308e-06, 1.222997e-06, 4.093051e-07, 
    9.288761e-07, 1.360989e-06, 2.176335e-06, 3.215843e-06, 2.034949e-06,
  1.044846e-05, 1.52689e-05, 2.01768e-05, 1.068378e-05, 1.381694e-05, 
    6.675566e-06, 2.623412e-06, 1.170061e-06, 5.329345e-07, 5.690541e-07, 
    6.440472e-07, 1.204459e-06, 2.470179e-06, 2.890746e-06, 3.616823e-06,
  1.138517e-08, 1.359759e-05, 2.178864e-05, 2.406333e-05, 2.631318e-05, 
    2.189668e-05, 2.336646e-05, 1.5935e-05, 8.215887e-06, 1.020847e-05, 
    9.323744e-06, 4.584689e-06, 4.145818e-06, 1.072747e-05, 1.380056e-05,
  2.901547e-09, 1.338192e-06, 6.799021e-06, 1.726463e-05, 1.028845e-05, 
    1.892693e-05, 3.009769e-05, 3.275894e-05, 2.985936e-05, 1.790647e-05, 
    1.671476e-05, 1.536344e-05, 1.446619e-05, 1.011467e-05, 8.95793e-06,
  6.353017e-11, 3.703161e-10, 3.894501e-09, 6.465482e-07, 4.713107e-06, 
    1.997493e-06, 9.54929e-06, 1.621141e-05, 2.308531e-05, 1.861917e-05, 
    1.816587e-05, 1.849524e-05, 1.672939e-05, 1.340152e-05, 1.316634e-05,
  3.379585e-10, 5.168428e-09, 1.163605e-08, 2.413904e-08, 2.549312e-09, 
    7.567218e-08, 1.759135e-06, 2.273084e-06, 1.025686e-05, 1.160344e-05, 
    1.106492e-05, 1.344707e-05, 9.595728e-06, 9.940876e-06, 7.418466e-06,
  1.595856e-09, 2.686007e-06, 7.899559e-06, 5.750986e-06, 1.003616e-05, 
    1.041353e-05, 7.514942e-06, 6.030888e-06, 6.195165e-06, 4.881242e-06, 
    3.782948e-06, 2.73991e-06, 3.188458e-06, 2.669376e-06, 2.657614e-06,
  1.963003e-05, 1.348957e-06, 1.097315e-05, 1.188952e-05, 1.615053e-05, 
    7.548983e-06, 4.127871e-06, 4.815771e-06, 7.372227e-06, 7.306581e-06, 
    5.82662e-06, 4.097262e-06, 4.061951e-06, 3.642285e-06, 3.266694e-06,
  8.60683e-06, 1.093896e-05, 1.676342e-05, 2.17244e-05, 2.226641e-05, 
    1.649686e-05, 3.770999e-06, 3.53129e-06, 6.076755e-06, 8.008144e-06, 
    7.72514e-06, 5.355195e-06, 3.89874e-06, 4.294286e-06, 4.357781e-06,
  5.102135e-06, 6.051312e-06, 4.854822e-06, 2.818344e-05, 2.97207e-05, 
    2.037866e-05, 9.366292e-06, 2.720203e-06, 4.37551e-06, 8.245329e-06, 
    8.429756e-06, 6.36473e-06, 7.066172e-06, 5.470427e-06, 3.109215e-06,
  3.956467e-06, 6.267956e-06, 9.741489e-06, 3.036566e-05, 2.342283e-05, 
    2.795779e-05, 1.479032e-05, 3.38003e-06, 3.771995e-06, 4.829458e-06, 
    6.046118e-06, 6.432019e-06, 4.573539e-06, 2.293249e-06, 2.925857e-06,
  1.042503e-06, 6.569367e-06, 1.60877e-06, 1.467344e-05, 1.970946e-05, 
    2.915069e-05, 1.994559e-05, 5.388004e-06, 2.334864e-06, 4.118126e-06, 
    4.759855e-06, 4.735587e-06, 6.371788e-06, 6.608669e-06, 4.255884e-06,
  6.641856e-07, 3.525583e-06, 8.911416e-06, 4.953351e-06, 1.677979e-05, 
    3.494444e-05, 2.810245e-05, 1.901758e-05, 4.507173e-06, 4.682555e-06, 
    5.190925e-06, 5.800821e-06, 8.538922e-06, 9.173807e-06, 4.72495e-06,
  5.832244e-09, 1.333677e-07, 1.395413e-06, 2.369181e-08, 2.02232e-06, 
    1.693606e-05, 2.617075e-05, 2.819837e-05, 1.710931e-05, 8.090105e-06, 
    6.572049e-06, 9.286244e-06, 8.180182e-06, 3.003692e-06, 3.213242e-06,
  2.948811e-07, 3.798976e-07, 2.345239e-07, 1.024374e-08, 2.189499e-08, 
    1.87477e-06, 1.230453e-05, 2.118626e-05, 1.976301e-05, 1.218951e-05, 
    9.57767e-06, 1.082089e-05, 2.062002e-05, 1.202819e-05, 7.919192e-06,
  2.414665e-07, 8.047246e-07, 8.588665e-08, 2.993107e-08, 4.082101e-09, 
    5.057693e-08, 6.111914e-06, 5.852277e-06, 1.254561e-05, 1.480964e-05, 
    1.128169e-05, 1.553716e-05, 8.449315e-05, 0.0001966735, 0.0001877989,
  5.572207e-08, 1.905279e-09, 1.188559e-08, 2.222183e-06, 1.2541e-05, 
    1.238579e-05, 1.229523e-05, 4.783809e-06, 1.074774e-06, 3.435048e-06, 
    4.010055e-06, 5.732451e-06, 3.175948e-06, 2.326239e-05, 0.000262138,
  1.583563e-06, 9.511687e-10, 8.136734e-07, 2.46593e-06, 1.021041e-05, 
    1.346103e-05, 1.207335e-05, 8.939822e-07, 7.094198e-07, 2.158399e-06, 
    3.548854e-06, 2.934356e-06, 1.269227e-05, 0.0001253916, 0.0003876848,
  5.022751e-08, 4.612871e-10, 1.144089e-08, 2.459012e-06, 8.705429e-06, 
    1.346226e-05, 1.198433e-05, 6.715409e-07, 1.329493e-06, 2.669837e-06, 
    4.013093e-06, 7.844815e-06, 5.130985e-05, 0.0002093938, 0.0003651407,
  1.001365e-08, 2.147648e-11, 6.006282e-10, 1.227796e-06, 3.927186e-06, 
    6.877003e-06, 9.757851e-06, 2.813211e-06, 9.013669e-07, 3.990943e-06, 
    5.581466e-06, 2.100886e-05, 6.996711e-05, 0.0001621144, 0.0001746621,
  3.301668e-09, 7.064721e-09, 1.167669e-11, 5.917947e-07, 2.49894e-06, 
    8.367043e-06, 1.200174e-05, 4.34207e-06, 1.589181e-06, 4.618826e-06, 
    1.112776e-05, 2.694895e-05, 6.077694e-05, 0.0001009095, 0.0001322173,
  1.030172e-09, 6.510298e-09, 3.111756e-09, 2.750307e-10, 1.630265e-06, 
    4.045896e-06, 6.072269e-06, 1.136676e-05, 3.930354e-06, 9.649994e-06, 
    9.496067e-06, 1.864687e-05, 4.982658e-05, 8.865548e-05, 0.0001049951,
  5.318116e-09, 1.060554e-08, 2.417445e-08, 1.627334e-09, 8.145398e-07, 
    3.378171e-06, 6.395791e-06, 9.492508e-06, 1.394072e-05, 9.010482e-06, 
    1.48008e-05, 4.916859e-05, 2.89974e-05, 7.187352e-05, 0.0001156373,
  2.368967e-09, 3.371726e-08, 2.154462e-08, 1.398802e-12, 2.194356e-09, 
    1.511085e-06, 1.002986e-05, 9.877999e-06, 2.292266e-05, 1.602566e-05, 
    2.24969e-05, 7.260463e-05, 0.0001034017, 9.364108e-05, 0.0001224032,
  4.448718e-07, 7.614764e-07, 2.675087e-07, 3.497617e-07, 3.763139e-07, 
    1.858726e-09, 5.574815e-06, 1.120336e-05, 1.591088e-05, 1.454604e-05, 
    2.830451e-05, 3.490863e-05, 6.95139e-05, 7.76405e-05, 8.522439e-05,
  1.127973e-06, 5.398999e-06, 3.706593e-06, 3.705401e-06, 1.945674e-06, 
    1.484851e-06, 1.265287e-06, 6.090917e-06, 7.027358e-06, 1.350868e-05, 
    2.467594e-05, 3.182118e-05, 6.368534e-05, 0.0001025503, 6.20432e-05,
  5.139913e-06, 3.332108e-06, 8.447457e-06, 8.890714e-06, 5.192464e-05, 
    8.710541e-05, 0.000101293, 0.0001205778, 0.000127514, 0.000162377, 
    0.0001306838, 0.0001292461, 0.0001277512, 9.394324e-05, 7.701552e-05,
  5.45367e-06, 1.638498e-06, 4.535419e-07, 1.248845e-06, 8.700343e-06, 
    3.509688e-05, 6.936949e-05, 8.53178e-05, 4.645607e-05, 6.716764e-05, 
    7.993203e-05, 0.0001378952, 4.955227e-05, 5.335536e-05, 4.665758e-05,
  5.65749e-06, 5.474616e-06, 3.151355e-06, 1.306872e-06, 1.242053e-06, 
    1.681758e-05, 4.126897e-05, 5.173363e-05, 4.807796e-05, 4.322271e-05, 
    5.462578e-05, 4.135255e-05, 2.511232e-05, 1.13374e-05, 2.552185e-05,
  6.495375e-06, 4.143516e-06, 5.924934e-06, 6.381403e-06, 7.897181e-06, 
    3.459376e-06, 4.97432e-05, 2.946293e-05, 3.481793e-05, 3.266307e-05, 
    4.984623e-05, 5.411446e-05, 2.351782e-05, 2.312623e-05, 1.288126e-05,
  4.158819e-05, 2.151523e-05, 2.683156e-05, 4.132949e-05, 5.529969e-05, 
    4.577068e-05, 3.839776e-05, 6.648461e-06, 1.580097e-05, 3.734112e-05, 
    0.0001138827, 6.76534e-05, 7.265512e-06, 1.742207e-05, 2.623151e-05,
  0.0001416884, 3.499069e-05, 5.137708e-05, 1.480853e-05, 1.872883e-05, 
    1.961047e-05, 1.778527e-05, 8.988043e-06, 1.230205e-05, 9.977978e-05, 
    4.141253e-05, 3.203607e-05, 5.228751e-05, 3.69663e-05, 2.475184e-05,
  0.0001101987, 0.0001273898, 0.000114384, 6.154153e-05, 1.949536e-06, 
    1.850093e-06, 3.037336e-06, 4.693229e-06, 5.776475e-06, 1.834649e-05, 
    2.995405e-05, 5.63123e-05, 3.145569e-05, 3.488476e-05, 1.786109e-05,
  5.887801e-05, 0.0001049149, 8.518043e-05, 7.942739e-05, 9.371625e-07, 
    3.326323e-08, 2.289265e-08, 8.169054e-08, 1.399081e-06, 4.458942e-06, 
    2.773945e-05, 5.286929e-05, 7.57866e-05, 6.528683e-05, 3.674904e-05,
  2.461534e-05, 4.066685e-05, 4.502215e-05, 4.705072e-05, 4.353812e-05, 
    7.110934e-09, 2.426809e-09, 1.761027e-09, 1.788803e-07, 5.033482e-07, 
    6.051245e-06, 2.55071e-05, 3.815844e-05, 1.444778e-05, 4.08702e-05,
  5.456057e-06, 2.239513e-05, 1.73352e-05, 1.733391e-05, 6.214526e-06, 
    8.633338e-06, 3.087049e-09, 7.469326e-10, 3.325217e-07, 6.072298e-07, 
    3.638728e-06, 1.829528e-05, 2.847892e-05, 2.062377e-05, 1.545033e-05,
  2.921035e-05, 1.032088e-05, 2.687818e-07, 2.618813e-08, 7.603509e-08, 
    4.345783e-08, 1.104544e-08, 1.80062e-07, 2.996652e-07, 1.077497e-06, 
    3.489028e-07, 4.863522e-07, 2.120861e-06, 3.582891e-06, 4.247429e-06,
  0.0003985491, 0.0001769959, 3.320269e-05, 5.862306e-06, 1.708602e-07, 
    1.042545e-08, 7.531196e-09, 1.187774e-08, 1.19135e-08, 3.407076e-08, 
    5.192246e-08, 2.285094e-07, 3.555948e-07, 2.863711e-07, 1.33825e-06,
  0.0007051623, 0.0005711641, 0.0002861068, 4.864795e-05, 1.025357e-05, 
    5.725868e-07, 1.831593e-07, 4.454432e-09, 1.624755e-08, 4.543793e-09, 
    1.429112e-08, 7.809011e-08, 4.041478e-08, 1.162549e-07, 1.568943e-07,
  0.0004036948, 0.0004955219, 0.0004579531, 0.0003283878, 9.864359e-05, 
    2.659236e-05, 8.349293e-06, 8.037142e-07, 2.516683e-07, 1.240985e-08, 
    2.453869e-09, 2.49582e-09, 2.823279e-08, 3.839213e-08, 4.881361e-08,
  0.0001754808, 0.0001654442, 0.0003505133, 0.0004809389, 0.0004856627, 
    0.0004083058, 0.0003292172, 0.0001618403, 4.886233e-05, 8.969821e-06, 
    5.148589e-07, 5.309566e-08, 2.540553e-09, 1.005582e-09, 5.144533e-08,
  9.859839e-05, 0.000125073, 6.32168e-05, 3.455895e-05, 0.0001756303, 
    0.0002910943, 0.0004359137, 0.0003839181, 0.000312498, 0.0001808328, 
    7.080819e-05, 1.508886e-05, 2.695261e-06, 1.3877e-07, 1.654917e-08,
  7.934214e-05, 0.0001007688, 9.909261e-05, 9.60829e-05, 6.582351e-06, 
    5.42746e-06, 5.362359e-05, 0.0001654287, 0.0001907961, 0.0001211615, 
    0.0002434839, 0.0001326224, 9.560146e-05, 4.56417e-05, 1.894067e-05,
  4.224948e-05, 6.731212e-05, 7.592519e-05, 8.333997e-05, 1.461758e-06, 
    9.945032e-07, 1.24461e-06, 1.83819e-05, 9.590139e-05, 0.0001292495, 
    0.0001242831, 0.0001660026, 0.0001117634, 8.958956e-05, 7.369825e-05,
  9.963164e-05, 6.401383e-05, 4.480294e-05, 1.431934e-05, 2.136175e-05, 
    5.729197e-09, 6.565751e-08, 6.502105e-07, 2.859428e-06, 4.315802e-05, 
    6.718024e-05, 9.466901e-05, 9.543134e-05, 0.0001193392, 9.610421e-05,
  0.0001129511, 0.0001232384, 0.0001044466, 4.152342e-05, 6.558382e-09, 
    1.049778e-06, 2.03968e-08, 4.144054e-07, 1.798548e-06, 1.179194e-05, 
    3.017045e-05, 4.001173e-05, 4.352552e-05, 8.338488e-05, 7.696428e-05,
  2.542852e-07, 8.349029e-08, 3.374457e-08, 6.172069e-07, 3.258767e-08, 
    7.606732e-08, 5.956098e-08, 1.199166e-08, 1.492275e-08, 1.374401e-08, 
    4.045257e-07, 1.305556e-06, 3.507985e-06, 3.678388e-06, 3.280262e-06,
  4.981294e-05, 1.753503e-05, 1.615516e-06, 6.94936e-06, 7.430973e-06, 
    6.264779e-06, 6.427235e-06, 2.455791e-07, 1.306771e-07, 1.785108e-07, 
    6.573629e-08, 6.089722e-08, 1.941435e-08, 4.790361e-07, 2.914635e-06,
  0.000185583, 5.330797e-05, 3.93069e-05, 2.509706e-05, 1.969532e-05, 
    1.939092e-05, 2.754086e-05, 1.138383e-05, 1.043136e-05, 3.319465e-06, 
    2.827244e-06, 3.234673e-06, 9.479804e-08, 1.355203e-08, 1.255979e-08,
  0.000140862, 6.444608e-05, 3.212181e-05, 5.074723e-05, 5.613104e-05, 
    5.986194e-05, 0.0001135888, 0.0001494848, 0.000116379, 0.0001276409, 
    5.744401e-05, 1.03649e-05, 4.55095e-06, 2.222631e-06, 6.190372e-08,
  0.0001845454, 0.0001700769, 5.876916e-06, 1.024996e-06, 1.116604e-05, 
    5.127344e-05, 4.958705e-05, 2.415745e-05, 6.210061e-05, 0.0001298301, 
    0.0002053248, 0.0001477845, 9.675926e-05, 1.316617e-05, 4.93467e-06,
  0.000180679, 0.0001879508, 0.0001573574, 5.088824e-07, 4.959211e-07, 
    1.059006e-06, 4.765539e-05, 9.904492e-06, 1.089384e-05, 6.275419e-05, 
    7.599395e-05, 0.0001098022, 0.0001933112, 0.0001875374, 0.0001780934,
  8.593162e-05, 0.0001393503, 0.0001689203, 0.0001156517, 2.160461e-07, 
    2.46814e-07, 3.986227e-06, 3.899417e-05, 2.740825e-05, 4.010113e-05, 
    2.072217e-05, 1.641184e-05, 1.416722e-05, 6.548716e-05, 0.0002390099,
  5.187425e-05, 7.525866e-05, 0.0001118404, 0.0001338769, 1.86565e-06, 
    1.674711e-07, 4.780658e-07, 8.626683e-06, 8.476657e-06, 1.994414e-05, 
    2.464603e-05, 3.625761e-05, 4.260354e-05, 4.682443e-05, 5.575328e-05,
  6.505662e-05, 4.944927e-05, 8.884422e-05, 0.0001445201, 0.0001065979, 
    6.436411e-06, 2.560604e-06, 2.09996e-06, 1.305064e-06, 3.361939e-06, 
    7.440755e-06, 1.688826e-05, 2.883439e-05, 3.265893e-05, 5.599053e-05,
  5.342515e-05, 7.895583e-05, 8.967316e-05, 0.0001465585, 0.0001829239, 
    0.0001689892, 3.060117e-06, 2.049298e-06, 1.059005e-06, 1.085046e-06, 
    2.306149e-06, 5.562952e-06, 1.294878e-05, 1.934468e-05, 3.181424e-05,
  0.0005724921, 0.0004991345, 0.0004084253, 0.0004953382, 0.000234628, 
    0.000151633, 5.285362e-05, 2.729453e-06, 9.11719e-06, 4.608687e-06, 
    4.736654e-06, 3.50508e-06, 2.894473e-07, 2.518166e-07, 1.577648e-06,
  0.0002354302, 0.0001407784, 0.0001010268, 0.000166327, 0.0004256957, 
    0.0002644942, 0.0002380626, 0.0001068229, 1.553751e-05, 1.395587e-05, 
    1.945777e-05, 1.895339e-05, 3.765532e-06, 6.832904e-07, 7.536763e-08,
  0.0002007643, 0.0001924638, 6.158341e-05, 4.759829e-05, 4.965936e-05, 
    0.000328933, 0.0002945204, 0.0002353104, 6.388531e-05, 4.349456e-05, 
    3.286897e-05, 1.114155e-05, 1.041183e-05, 1.116494e-05, 3.303594e-06,
  0.0001602822, 0.0001516652, 6.297281e-06, 2.657822e-06, 2.20226e-05, 
    0.0001334653, 0.000514942, 0.0003918709, 0.0001544755, 0.0001048343, 
    7.994464e-05, 5.399631e-05, 3.025788e-05, 2.435084e-05, 3.49667e-05,
  0.0001407832, 0.0001202029, 3.199834e-06, 1.306163e-06, 4.049531e-07, 
    3.276838e-06, 0.000230981, 0.0001937411, 8.244145e-05, 5.22862e-05, 
    6.474537e-05, 5.246212e-05, 8.690725e-05, 6.232892e-05, 2.060977e-05,
  8.19184e-05, 9.977935e-05, 9.268984e-05, 5.924259e-06, 8.555545e-07, 
    1.215765e-06, 1.615786e-05, 4.473359e-05, 4.832146e-05, 9.239052e-05, 
    2.482453e-05, 2.816401e-05, 3.807573e-05, 6.954695e-05, 3.079711e-05,
  0.0001056665, 0.0001030669, 0.0001345056, 8.909928e-05, 3.949334e-06, 
    3.624597e-06, 1.50429e-05, 4.692681e-05, 7.689917e-05, 5.301357e-05, 
    4.843226e-05, 4.343014e-05, 3.977355e-05, 3.114429e-05, 2.919191e-05,
  0.0001198561, 0.0001017422, 0.0001241486, 0.0001107875, 2.020442e-05, 
    1.549352e-05, 1.710537e-05, 2.560982e-05, 3.527782e-05, 3.806497e-05, 
    4.253949e-05, 4.975999e-05, 6.270347e-05, 5.299068e-05, 3.753572e-05,
  0.0001198217, 0.0001284642, 0.0001500398, 0.0001111194, 7.154796e-05, 
    3.100522e-05, 2.713083e-05, 1.315187e-05, 2.674125e-05, 2.911151e-05, 
    2.963425e-05, 3.028734e-05, 4.206216e-05, 5.191676e-05, 4.970513e-05,
  0.0001043946, 0.0001193307, 0.0001276282, 0.0001450311, 6.997376e-05, 
    4.743157e-05, 3.487059e-05, 1.602168e-05, 1.537243e-05, 1.451303e-05, 
    1.885696e-05, 1.983336e-05, 2.739602e-05, 3.377676e-05, 3.338173e-05,
  0.0001576495, 0.0003456098, 0.0005832039, 0.0007387983, 0.0009269112, 
    0.001031487, 0.001088443, 0.0009945682, 0.000897034, 0.0008686339, 
    0.000830691, 0.0007361749, 0.0006492223, 0.0005197102, 0.0004662889,
  4.543833e-05, 8.14351e-05, 0.0001666317, 0.0002358792, 0.0002698166, 
    0.0003403638, 0.0004765223, 0.0005592598, 0.0004714791, 0.000439465, 
    0.0004518589, 0.000464773, 0.0004572427, 0.0004682489, 0.0004368995,
  1.90052e-05, 1.378266e-05, 1.515227e-05, 1.104303e-05, 9.959203e-06, 
    1.49077e-05, 0.0001115112, 0.0001472407, 0.0001802779, 0.0001817857, 
    0.0002094895, 0.0002388825, 0.0003066691, 0.0003648958, 0.0003643697,
  1.221502e-05, 8.721432e-06, 1.24372e-05, 9.261018e-06, 7.300816e-06, 
    9.47979e-06, 3.445074e-05, 3.175638e-05, 3.675252e-05, 6.837145e-05, 
    6.807626e-05, 0.000110151, 0.0001182566, 0.0001641736, 0.0001853979,
  1.881126e-05, 1.657055e-05, 8.986452e-06, 7.458952e-06, 2.218679e-06, 
    4.972318e-06, 4.304511e-06, 5.096939e-06, 6.08703e-06, 3.552812e-05, 
    4.414563e-05, 5.91413e-05, 7.124737e-05, 7.080966e-05, 7.407788e-05,
  4.493149e-05, 3.894321e-05, 2.575727e-05, 3.631735e-06, 4.37086e-06, 
    3.146555e-06, 2.167603e-06, 2.205593e-06, 2.984846e-06, 1.704671e-05, 
    1.082677e-05, 1.570113e-05, 3.381888e-05, 5.220791e-05, 7.703451e-05,
  9.63584e-05, 9.136662e-05, 6.26192e-05, 2.887374e-05, 1.031011e-06, 
    2.528084e-06, 8.019189e-07, 8.97642e-07, 2.328984e-05, 3.114372e-05, 
    8.138174e-06, 1.117641e-05, 1.787193e-05, 3.116338e-05, 4.283784e-05,
  0.000205431, 0.0002421841, 0.0001644716, 3.834041e-05, 6.269825e-06, 
    2.049903e-06, 4.609432e-07, 7.402475e-07, 3.305708e-06, 9.508601e-06, 
    2.034986e-05, 1.264737e-05, 2.363625e-05, 6.201777e-05, 5.731178e-05,
  0.0002454856, 0.0002011185, 0.0001965626, 0.0002094369, 0.0001318573, 
    1.338702e-05, 3.220887e-06, 2.447427e-06, 2.599718e-06, 6.534877e-06, 
    1.263637e-05, 1.760659e-05, 3.947789e-05, 4.404105e-05, 5.961181e-05,
  0.0001421373, 0.0001498504, 0.0001386099, 0.0001191103, 0.0002044329, 
    0.0001520321, 1.829418e-05, 1.061676e-05, 4.615817e-06, 5.405414e-06, 
    4.538455e-05, 3.334419e-05, 8.23799e-05, 8.720903e-05, 6.449544e-05,
  4.120194e-17, 1.301956e-16, 7.288856e-14, 7.417895e-12, 9.045665e-09, 
    8.741256e-07, 9.787699e-07, 9.056819e-07, 7.890185e-07, 1.498862e-06, 
    9.531373e-06, 3.483328e-05, 4.510199e-05, 4.926997e-05, 4.814273e-05,
  3.756936e-10, 2.697136e-15, 6.986972e-18, 4.259555e-12, 4.7289e-08, 
    8.137771e-07, 6.46699e-07, 1.625714e-06, 1.753129e-06, 2.177923e-06, 
    8.479077e-06, 3.816465e-05, 4.136769e-05, 3.144859e-05, 2.926585e-05,
  2.304886e-08, 2.721013e-12, 8.344639e-23, 1.440072e-23, 2.240582e-09, 
    3.217511e-07, 5.130304e-07, 1.458841e-06, 2.674293e-06, 3.081535e-06, 
    1.116705e-05, 2.84014e-05, 3.62739e-05, 3.216124e-05, 2.520148e-05,
  6.512162e-08, 8.483043e-12, 1.664119e-12, 5.611171e-13, 5.005064e-12, 
    3.416188e-09, 1.705068e-07, 1.154189e-06, 1.437286e-06, 3.490384e-06, 
    5.698202e-06, 2.459926e-05, 3.581672e-05, 3.320152e-05, 2.943707e-05,
  2.808869e-07, 3.345976e-08, 1.082477e-10, 3.147108e-12, 7.699644e-13, 
    3.214084e-12, 3.221848e-09, 5.619327e-07, 1.224891e-06, 1.35445e-06, 
    5.20568e-06, 1.719457e-05, 2.735807e-05, 2.482514e-05, 3.163536e-05,
  2.1304e-06, 7.936412e-08, 1.574219e-08, 1.833879e-11, 3.953748e-12, 
    3.586143e-13, 1.043572e-10, 1.015149e-07, 6.810319e-07, 7.155728e-07, 
    2.124425e-06, 3.979812e-06, 7.900912e-06, 2.01799e-05, 2.082604e-05,
  6.279623e-06, 2.497135e-06, 8.921527e-07, 5.468501e-08, 4.772273e-11, 
    1.953422e-12, 4.512176e-11, 2.823305e-08, 4.118809e-07, 6.900735e-07, 
    1.468889e-06, 2.118996e-06, 4.3186e-06, 7.471246e-06, 1.5332e-05,
  6.649519e-06, 6.504847e-06, 5.445617e-06, 2.978137e-07, 2.729201e-09, 
    1.6525e-10, 7.205928e-09, 6.079492e-09, 1.647774e-08, 5.926487e-07, 
    9.325003e-07, 1.653937e-06, 2.625101e-06, 4.421154e-06, 7.080351e-06,
  6.666876e-05, 4.166006e-06, 2.039215e-05, 1.993631e-05, 2.763368e-06, 
    4.898351e-09, 8.034366e-11, 1.10899e-07, 3.063178e-07, 6.278702e-07, 
    5.751803e-07, 7.34866e-07, 1.674707e-06, 2.538829e-06, 4.610209e-06,
  9.538439e-05, 0.0001131611, 2.343048e-05, 2.451324e-05, 2.282253e-05, 
    4.366018e-06, 9.200862e-09, 5.686224e-08, 9.358874e-08, 2.358391e-07, 
    1.018437e-07, 5.633871e-07, 6.221629e-07, 2.120243e-06, 1.009436e-05,
  0.0003908153, 0.0003433988, 0.0002137004, 5.89314e-05, 3.522327e-06, 
    4.855622e-06, 5.267501e-06, 4.06842e-06, 3.831508e-06, 2.114934e-07, 
    2.239402e-08, 6.284719e-09, 9.919916e-11, 5.408027e-11, 5.574214e-11,
  0.0001517735, 0.000193628, 0.0002357255, 0.0001422495, 3.729518e-05, 
    2.67148e-06, 6.526532e-06, 8.158038e-06, 1.606687e-06, 3.489536e-07, 
    3.67852e-08, 8.224561e-09, 5.196813e-10, 1.131824e-10, 1.218225e-11,
  9.266785e-05, 5.602981e-05, 9.942309e-05, 0.0001278678, 6.14567e-05, 
    3.417155e-06, 5.440229e-06, 7.726967e-06, 3.583897e-06, 1.076553e-06, 
    1.262381e-07, 6.451827e-09, 1.18109e-10, 7.780959e-11, 7.793668e-11,
  9.816929e-05, 3.979501e-05, 3.116972e-05, 6.745006e-05, 7.490109e-05, 
    2.00143e-05, 6.689575e-06, 8.618601e-06, 6.871521e-06, 2.632426e-06, 
    2.76952e-08, 5.191827e-08, 9.492813e-11, 2.566008e-11, 4.975665e-11,
  5.322802e-05, 2.11417e-05, 1.090496e-05, 2.241425e-05, 4.132322e-05, 
    4.36931e-05, 2.892016e-06, 5.681739e-06, 8.353527e-06, 5.892818e-06, 
    2.423631e-07, 4.38655e-09, 4.348492e-10, 2.215581e-11, 1.081703e-09,
  2.375287e-05, 9.766757e-06, 2.45729e-06, 1.043246e-06, 5.499516e-06, 
    1.852201e-05, 6.499246e-06, 4.28102e-06, 8.387328e-06, 7.34198e-06, 
    1.577267e-07, 2.059368e-08, 1.834544e-09, 3.923796e-09, 4.478751e-08,
  3.064098e-05, 3.098389e-05, 3.1039e-05, 2.211679e-06, 3.826866e-07, 
    1.044782e-06, 5.390391e-06, 5.384112e-06, 7.201684e-06, 6.098024e-06, 
    2.590736e-07, 7.316057e-09, 2.17419e-08, 8.447086e-08, 6.008104e-08,
  2.418267e-05, 2.782251e-05, 3.974546e-05, 3.421541e-05, 1.405342e-08, 
    4.130916e-07, 1.624007e-06, 1.411821e-06, 5.968539e-06, 3.093834e-06, 
    9.809143e-07, 4.841309e-08, 5.297706e-08, 2.888828e-07, 3.408062e-07,
  2.645262e-05, 3.157761e-05, 4.555726e-05, 2.993183e-05, 8.743054e-06, 
    2.737416e-07, 1.767971e-06, 5.603018e-07, 1.779719e-06, 1.035281e-06, 
    2.644759e-08, 2.065976e-07, 1.119003e-07, 6.520153e-08, 7.915316e-07,
  3.498129e-05, 2.619221e-05, 4.862316e-05, 5.445388e-05, 1.973037e-05, 
    2.936647e-06, 1.289459e-06, 1.405121e-06, 1.067367e-06, 7.813112e-07, 
    1.16657e-07, 1.157632e-07, 4.034536e-07, 9.3997e-08, 1.475453e-07,
  3.030099e-05, 0.0001748816, 0.0003867477, 0.0005850227, 0.0005733176, 
    0.0005405114, 0.0005048173, 0.000543827, 0.0006076199, 0.0005516854, 
    0.0003073371, 9.80464e-05, 4.547471e-05, 2.861537e-05, 1.000873e-05,
  5.180507e-05, 3.43334e-05, 0.0001631887, 0.0003599623, 0.0004900793, 
    0.0005254495, 0.0004804912, 0.0004594623, 0.0005497266, 0.0006274749, 
    0.0005824305, 0.0003093773, 0.000150377, 9.533772e-05, 5.273177e-05,
  6.339824e-05, 3.134065e-05, 1.185901e-05, 5.427862e-05, 0.0001699472, 
    0.0002422038, 0.0002715043, 0.0002831711, 0.0003447938, 0.000464905, 
    0.0005301033, 0.0004108407, 0.000198689, 0.0001298556, 0.0001462214,
  0.0003230439, 0.0001574838, 0.0001568998, 4.358924e-06, 6.88809e-06, 
    2.539369e-05, 8.453299e-05, 0.000103617, 9.693582e-05, 0.0001840207, 
    0.0003202634, 0.0003357249, 0.0002097595, 0.0001053569, 0.0001085648,
  0.0001843778, 0.0001654185, 3.467472e-05, 3.746562e-06, 3.783382e-06, 
    4.487303e-06, 1.584295e-05, 2.366496e-05, 3.594457e-05, 4.006932e-05, 
    7.153674e-05, 0.0001606429, 0.0001590575, 5.995176e-05, 3.092049e-05,
  0.0001459859, 0.0001677189, 0.0001496266, 4.96737e-07, 7.537136e-07, 
    1.552439e-06, 7.177173e-06, 8.413702e-06, 1.114955e-05, 1.464679e-05, 
    3.074026e-05, 4.446362e-05, 7.811878e-05, 3.692705e-05, 7.934322e-06,
  6.683715e-05, 0.0001017941, 0.0001022618, 6.795473e-05, 6.025199e-09, 
    1.942135e-07, 3.964967e-06, 3.495297e-06, 4.437637e-06, 6.285648e-06, 
    1.108223e-05, 1.830762e-05, 2.773791e-05, 2.211664e-05, 5.024608e-06,
  4.052271e-05, 6.373158e-05, 4.789945e-05, 6.844228e-05, 1.993553e-09, 
    6.562501e-09, 3.094626e-06, 2.880399e-06, 2.279004e-06, 2.997629e-06, 
    6.19388e-06, 9.592647e-06, 1.136272e-05, 7.100225e-06, 2.473017e-06,
  4.605252e-05, 5.988699e-05, 6.485086e-05, 8.841199e-05, 7.595381e-05, 
    6.196421e-09, 1.113002e-06, 3.060269e-06, 2.05932e-06, 2.211309e-06, 
    5.604057e-06, 5.444426e-06, 5.761417e-06, 4.030926e-06, 9.807001e-07,
  7.802813e-05, 8.224534e-05, 9.613245e-05, 9.206658e-05, 8.213644e-05, 
    8.817686e-05, 7.738104e-09, 2.673487e-06, 1.133545e-06, 2.431478e-06, 
    4.453894e-06, 4.859155e-06, 6.193877e-06, 4.257973e-06, 2.24905e-06,
  7.893491e-07, 3.161827e-07, 1.34483e-06, 5.297388e-06, 6.091537e-06, 
    8.165011e-06, 6.087936e-06, 6.371884e-06, 1.524254e-05, 4.354806e-05, 
    6.460331e-05, 6.040674e-05, 5.851221e-05, 8.291614e-05, 9.978656e-05,
  1.122339e-06, 3.244953e-07, 9.902668e-07, 2.008868e-06, 2.169098e-06, 
    4.863453e-06, 5.552039e-06, 5.178175e-06, 4.990228e-06, 2.566659e-05, 
    7.813581e-05, 0.0001133077, 6.239348e-05, 5.634562e-05, 6.753712e-05,
  3.021579e-07, 4.304234e-07, 3.037952e-07, 6.701775e-07, 1.521421e-06, 
    2.692708e-06, 4.521292e-06, 3.686113e-06, 3.87196e-06, 7.730231e-06, 
    6.95701e-05, 0.0001873275, 0.0001799492, 7.150257e-05, 6.543061e-05,
  6.199778e-07, 2.212878e-07, 8.582118e-08, 4.862914e-07, 9.344241e-07, 
    1.868895e-06, 1.858171e-06, 1.723107e-06, 2.064635e-06, 5.459254e-06, 
    6.092675e-05, 0.0001951524, 0.0003014537, 0.0002207981, 8.492934e-05,
  1.442389e-06, 1.629299e-06, 1.382313e-06, 7.62309e-07, 8.708564e-07, 
    9.246187e-07, 1.479223e-06, 1.908719e-06, 1.996651e-06, 6.883761e-06, 
    4.522152e-05, 0.0001637711, 0.000331565, 0.0003775374, 0.000273936,
  5.322595e-05, 4.883611e-05, 6.055017e-05, 1.072807e-05, 3.203637e-06, 
    8.469118e-07, 8.285454e-07, 2.296761e-06, 4.903025e-06, 7.658036e-06, 
    2.012049e-05, 7.59663e-05, 0.0002351052, 0.0004245441, 0.0004413129,
  6.047037e-05, 3.641692e-05, 7.974465e-05, 8.878873e-05, 2.618537e-05, 
    1.076275e-05, 6.727935e-06, 7.276184e-06, 1.280502e-05, 2.295023e-05, 
    3.152535e-05, 4.669181e-05, 0.0001155385, 0.0003201654, 0.0004437202,
  0.0001420879, 8.622307e-05, 5.137353e-05, 4.298027e-05, 3.330484e-05, 
    2.105992e-05, 9.048363e-06, 5.517092e-06, 1.146865e-05, 3.082033e-05, 
    5.523261e-05, 8.253884e-05, 0.000124962, 0.0002192921, 0.0003274421,
  0.0001840332, 0.000143452, 9.540822e-05, 8.7897e-05, 2.903112e-05, 
    1.289705e-05, 3.424587e-06, 7.687738e-07, 1.106371e-06, 3.455835e-06, 
    1.507703e-05, 4.558602e-05, 9.162408e-05, 0.0001369676, 0.0001859644,
  9.910134e-05, 9.711321e-05, 0.0001258624, 0.0001156772, 7.345655e-05, 
    6.758088e-05, 1.726187e-06, 3.863908e-07, 1.12121e-07, 2.887956e-07, 
    6.419269e-07, 4.631594e-06, 1.70275e-05, 6.122791e-05, 7.734589e-05,
  2.714557e-09, 2.197106e-09, 1.978481e-08, 7.211727e-08, 4.290548e-07, 
    3.214121e-06, 6.075953e-06, 1.482569e-05, 1.627727e-05, 1.594169e-05, 
    1.519423e-05, 1.50857e-05, 1.026709e-05, 9.391571e-06, 9.099565e-06,
  2.848904e-09, 2.325803e-09, 2.415086e-09, 2.461343e-08, 8.813895e-08, 
    1.00712e-06, 3.407567e-06, 8.226297e-06, 1.210645e-05, 1.554063e-05, 
    1.732372e-05, 1.237278e-05, 7.853345e-06, 1.02875e-05, 1.251274e-05,
  1.286319e-07, 4.678785e-08, 3.85771e-09, 3.605227e-09, 9.004272e-08, 
    3.258492e-07, 9.682351e-07, 4.178587e-06, 8.23656e-06, 1.439616e-05, 
    1.25224e-05, 1.224832e-05, 1.371102e-05, 1.281472e-05, 1.685303e-05,
  1.00169e-05, 8.537268e-08, 5.372675e-08, 1.174039e-08, 2.059959e-09, 
    1.374817e-08, 9.402086e-07, 2.08029e-06, 4.446502e-06, 9.464181e-06, 
    1.066445e-05, 1.990856e-05, 1.564762e-05, 1.146127e-05, 1.125197e-05,
  0.0001253728, 4.766162e-05, 8.438458e-06, 6.198965e-07, 1.250461e-07, 
    2.808165e-09, 9.121751e-08, 7.98975e-07, 2.415181e-06, 3.960798e-06, 
    9.679981e-06, 1.36638e-05, 1.392113e-05, 1.591064e-05, 1.080912e-05,
  0.0002875039, 0.000219391, 0.0001374136, 5.258419e-05, 1.356617e-05, 
    1.200422e-06, 3.264422e-09, 3.983405e-08, 2.785697e-07, 2.115251e-06, 
    3.698069e-06, 7.276877e-06, 9.809227e-06, 1.497564e-05, 1.453633e-05,
  0.000291621, 0.0002432147, 0.0001644158, 8.012188e-05, 2.366085e-05, 
    3.355152e-06, 1.28396e-09, 1.619353e-09, 1.483312e-08, 9.329692e-08, 
    1.973092e-06, 3.588614e-06, 6.084746e-06, 1.025173e-05, 1.196933e-05,
  0.0001926856, 0.0001117426, 7.058487e-05, 2.463864e-05, 3.901567e-06, 
    5.514784e-08, 2.517144e-09, 3.851008e-10, 1.330524e-09, 1.080491e-08, 
    9.855548e-08, 8.557874e-07, 3.358695e-06, 5.729572e-06, 8.255931e-06,
  0.0002867253, 0.0001794006, 0.0001026452, 3.230028e-05, 5.969506e-06, 
    1.178697e-07, 4.552645e-09, 1.658119e-09, 2.514153e-10, 1.216387e-09, 
    2.276709e-09, 2.971044e-09, 9.379287e-08, 1.259122e-06, 6.486478e-06,
  0.0002108877, 0.0001872717, 0.0001793396, 7.839291e-05, 4.026512e-05, 
    5.267241e-06, 8.115081e-08, 2.794583e-08, 1.063698e-09, 1.812644e-10, 
    1.626878e-10, 1.558708e-09, 2.542665e-09, 8.523838e-08, 4.426481e-07,
  2.193381e-06, 5.318793e-10, 3.294022e-09, 6.323031e-07, 2.17157e-06, 
    7.924586e-06, 6.110165e-06, 7.740937e-06, 9.989097e-06, 1.845789e-05, 
    2.688097e-05, 4.863597e-05, 2.24383e-05, 1.778016e-05, 5.623661e-06,
  2.651605e-05, 1.095842e-06, 4.086306e-07, 6.766732e-07, 9.665182e-07, 
    2.144666e-06, 3.996086e-06, 4.470499e-06, 6.624711e-06, 1.008673e-05, 
    2.039579e-05, 2.799731e-05, 4.126579e-05, 1.343998e-05, 9.198548e-06,
  2.256594e-05, 1.264152e-05, 1.519051e-06, 7.767219e-07, 4.600025e-07, 
    1.139418e-06, 4.186277e-06, 5.732763e-06, 5.592567e-06, 6.840238e-06, 
    1.07413e-05, 1.94051e-05, 2.386946e-05, 3.484137e-05, 1.771004e-05,
  4.661924e-05, 3.771297e-05, 1.138552e-05, 4.051692e-06, 6.360143e-07, 
    4.780983e-07, 1.188323e-06, 2.820912e-06, 4.817551e-06, 6.683948e-06, 
    9.457926e-06, 1.215515e-05, 2.161218e-05, 2.338142e-05, 4.717211e-05,
  5.140449e-05, 4.332597e-05, 3.298771e-05, 1.970609e-05, 6.830318e-06, 
    1.856445e-06, 1.423058e-06, 1.331668e-06, 1.940087e-06, 6.622524e-06, 
    1.002124e-05, 1.411565e-05, 1.614983e-05, 1.598098e-05, 2.660197e-05,
  5.901715e-05, 0.0001135747, 0.0001852507, 0.0001467641, 0.0001289973, 
    0.0001023724, 6.204688e-05, 3.792227e-05, 2.522498e-05, 2.678772e-05, 
    3.843867e-05, 4.419143e-05, 4.599043e-05, 3.778342e-05, 5.181306e-05,
  0.0001197618, 0.0001748654, 0.0003201608, 0.0004310295, 0.0004931514, 
    0.0005645478, 0.0006139373, 0.0006552897, 0.0006012511, 0.0005148898, 
    0.0004427765, 0.0003442877, 0.0002779494, 0.0002333466, 0.0001994091,
  9.408516e-05, 0.0001984842, 0.0002120036, 0.0003146531, 0.000361946, 
    0.0005538846, 0.0008200892, 0.001026748, 0.001135373, 0.001067966, 
    0.0009465618, 0.0007628363, 0.0006112205, 0.0004923457, 0.0003285091,
  0.0002544709, 0.0003333557, 0.0002310152, 8.347534e-05, 0.0001028159, 
    8.477832e-05, 0.0002473838, 0.0004312046, 0.0008174945, 0.0006458108, 
    0.0007438699, 0.0007590698, 0.0007271442, 0.0006194954, 0.0004043549,
  0.0002104946, 0.0001857267, 0.0002853836, 0.0002987912, 0.0002842737, 
    0.0001944985, 2.123377e-06, 3.194299e-06, 1.487558e-05, 0.0001177438, 
    0.0002482434, 0.0003165785, 0.000384194, 0.0003594684, 0.0002557873,
  9.652078e-10, 1.496724e-11, 3.155343e-12, 2.414836e-11, 2.064226e-07, 
    6.830742e-07, 8.218504e-07, 4.05975e-06, 3.059005e-06, 1.409933e-06, 
    2.226855e-06, 4.977479e-06, 6.473325e-06, 8.361762e-06, 1.119975e-05,
  3.572325e-07, 1.113567e-09, 7.3503e-09, 7.549321e-10, 4.18431e-07, 
    5.384861e-07, 5.364393e-06, 6.227758e-06, 3.662068e-06, 2.554272e-06, 
    3.300861e-06, 5.118346e-06, 7.881067e-06, 7.538874e-06, 5.518814e-06,
  1.63686e-06, 2.205496e-06, 4.731342e-07, 8.522189e-07, 5.497639e-07, 
    3.403314e-06, 4.90209e-06, 3.578325e-06, 2.9803e-06, 3.429501e-06, 
    3.798597e-06, 4.756348e-06, 7.605892e-06, 6.20445e-06, 1.00691e-05,
  3.69775e-06, 3.071036e-06, 1.410164e-06, 1.96267e-06, 2.915778e-06, 
    3.887227e-06, 6.788876e-06, 3.535606e-06, 2.481834e-06, 4.194741e-06, 
    5.474272e-06, 7.007536e-06, 7.269684e-06, 8.176681e-06, 1.046354e-05,
  4.753587e-06, 5.947696e-06, 4.621956e-06, 4.775386e-06, 5.809139e-06, 
    6.91198e-06, 7.129798e-06, 2.791387e-06, 2.404408e-06, 3.07863e-06, 
    3.881408e-06, 6.685679e-06, 8.20294e-06, 1.033241e-05, 1.321203e-05,
  1.196905e-05, 7.126813e-06, 1.059588e-05, 4.924815e-06, 5.866349e-06, 
    5.433472e-06, 4.533386e-06, 2.846544e-06, 3.119343e-06, 3.580321e-06, 
    5.24097e-06, 7.804215e-06, 8.29416e-06, 9.992984e-06, 1.511829e-05,
  2.789678e-05, 1.765338e-05, 2.056689e-05, 1.138922e-05, 4.348079e-06, 
    3.540708e-06, 2.895593e-06, 2.390239e-06, 4.406397e-06, 6.01273e-06, 
    7.034112e-06, 9.68232e-06, 9.349845e-06, 6.105971e-06, 2.398471e-05,
  1.109666e-05, 1.659563e-05, 1.158932e-05, 8.862994e-06, 5.214531e-06, 
    3.073404e-06, 3.264014e-06, 2.043862e-06, 2.826159e-06, 4.480483e-06, 
    9.005874e-06, 7.97456e-06, 9.273083e-06, 1.428332e-05, 7.896998e-05,
  4.895304e-06, 4.677943e-06, 2.534395e-06, 3.592147e-06, 6.706364e-06, 
    2.513697e-06, 3.851861e-06, 2.803069e-06, 3.932108e-06, 6.897567e-06, 
    1.044847e-05, 1.045097e-05, 3.495397e-05, 0.0001319396, 0.0002938482,
  1.028808e-05, 9.861876e-06, 1.156389e-05, 1.074358e-05, 8.750237e-06, 
    7.829843e-06, 5.061111e-06, 6.476214e-06, 5.607041e-06, 7.000675e-06, 
    6.785433e-06, 1.218958e-05, 4.664489e-05, 0.0001739462, 0.0003820077,
  2.388355e-11, 4.478527e-10, 2.422363e-09, 6.087614e-10, 3.9797e-10, 
    1.560666e-10, 3.181061e-10, 4.365027e-08, 3.227528e-06, 1.922071e-06, 
    2.231853e-06, 2.801168e-06, 1.456693e-06, 3.83829e-06, 2.030617e-06,
  1.787288e-08, 2.22083e-10, 2.1231e-10, 3.730234e-10, 1.354355e-09, 
    1.500105e-09, 1.323226e-09, 1.582563e-07, 3.277915e-06, 7.70764e-07, 
    1.973585e-06, 7.475066e-07, 7.109795e-07, 9.847333e-07, 8.485861e-07,
  1.303469e-08, 1.243472e-07, 2.774166e-10, 5.183085e-09, 5.71988e-10, 
    1.284528e-09, 1.908061e-09, 5.014832e-07, 1.222368e-06, 1.131208e-06, 
    1.321263e-06, 4.509455e-07, 1.79398e-06, 8.92835e-07, 1.893863e-06,
  6.344905e-07, 3.170174e-07, 3.329972e-09, 6.824427e-08, 6.97321e-09, 
    6.854833e-10, 7.435766e-08, 5.038644e-07, 1.111692e-06, 2.061435e-06, 
    1.560567e-06, 2.052501e-06, 1.756671e-06, 4.772639e-06, 4.235525e-06,
  2.081145e-07, 1.295004e-06, 6.618613e-07, 5.053842e-07, 3.843886e-07, 
    7.407984e-08, 2.523177e-07, 4.733956e-07, 1.230252e-06, 2.882226e-06, 
    3.45944e-06, 3.254019e-06, 2.974519e-06, 5.403673e-06, 8.108813e-06,
  2.579748e-07, 6.459731e-07, 2.325368e-06, 4.367663e-07, 7.722082e-07, 
    8.488284e-07, 5.1366e-07, 8.086438e-07, 1.773024e-06, 2.501305e-06, 
    4.799976e-06, 4.845355e-06, 3.657168e-06, 6.081089e-06, 9.015756e-06,
  8.398554e-07, 3.219116e-07, 1.74197e-06, 3.222713e-06, 1.284101e-06, 
    8.30167e-07, 6.963654e-07, 7.947299e-07, 1.445178e-06, 2.696383e-06, 
    4.032465e-06, 5.22082e-06, 4.766551e-06, 5.044664e-06, 1.001573e-05,
  2.196299e-06, 8.359429e-08, 5.101186e-07, 1.760145e-06, 1.191559e-06, 
    1.482602e-06, 1.024939e-06, 1.522515e-06, 2.054564e-06, 3.03649e-06, 
    3.643941e-06, 4.288823e-06, 4.790907e-06, 5.389238e-06, 1.061943e-05,
  7.498927e-06, 1.992113e-06, 1.0963e-06, 1.316722e-07, 2.567843e-06, 
    1.099126e-06, 1.713751e-06, 2.096563e-06, 2.289224e-06, 1.484048e-06, 
    2.926122e-06, 4.265937e-06, 5.897154e-06, 9.134118e-06, 1.164142e-05,
  3.892662e-05, 1.760797e-05, 5.385639e-06, 9.475955e-07, 3.372574e-07, 
    1.155856e-06, 9.278422e-07, 1.465832e-06, 2.176949e-06, 2.478165e-06, 
    1.971904e-06, 4.371086e-06, 7.448751e-06, 1.069245e-05, 1.076761e-05,
  2.353981e-09, 6.77785e-08, 8.047009e-09, 2.390506e-07, 1.020589e-06, 
    1.576953e-06, 5.695425e-06, 1.12374e-05, 8.914006e-06, 2.047625e-05, 
    1.715534e-05, 1.950637e-05, 1.612705e-05, 1.314874e-05, 6.2881e-06,
  2.02132e-06, 2.119674e-07, 8.874227e-07, 8.508125e-07, 2.3958e-06, 
    1.211457e-06, 8.512385e-06, 1.510165e-06, 3.16444e-06, 1.334844e-06, 
    7.048227e-07, 1.193966e-06, 3.088091e-06, 7.020518e-06, 9.074058e-06,
  5.996853e-06, 1.717934e-06, 9.841499e-07, 1.258376e-06, 3.533447e-07, 
    1.985905e-07, 1.913912e-07, 3.851048e-07, 5.23126e-08, 6.696287e-07, 
    6.267204e-08, 8.670406e-08, 5.386696e-07, 1.04873e-06, 1.337207e-06,
  9.97697e-06, 1.056565e-05, 5.177026e-06, 4.712431e-06, 2.350592e-06, 
    2.944497e-07, 6.54356e-08, 2.205861e-07, 4.652939e-08, 3.706449e-08, 
    1.581324e-08, 5.091407e-09, 3.03899e-08, 3.374308e-07, 1.345672e-06,
  1.018288e-05, 1.525321e-05, 8.215558e-06, 6.962342e-06, 4.389098e-06, 
    3.063726e-06, 2.896496e-06, 1.611626e-06, 4.276873e-07, 2.355331e-07, 
    6.518687e-08, 9.71648e-09, 1.064766e-07, 7.722757e-07, 5.523935e-07,
  1.224129e-05, 1.489571e-05, 2.48678e-05, 4.354624e-05, 4.698412e-05, 
    3.258903e-05, 1.001354e-05, 3.757645e-06, 3.315198e-06, 7.7098e-07, 
    4.879583e-07, 3.898201e-08, 4.063459e-08, 1.192874e-07, 2.019378e-07,
  7.076513e-05, 0.0001921591, 0.0003985678, 0.0005667903, 0.0005820887, 
    0.0003929639, 0.0001355913, 4.500726e-05, 1.554506e-05, 1.950488e-06, 
    1.104373e-06, 9.67103e-09, 2.856602e-08, 3.368227e-08, 4.847447e-07,
  0.000166512, 0.0003913423, 0.0006385936, 0.0008092962, 0.0008584361, 
    0.0007469355, 0.0003384714, 6.175364e-05, 1.986847e-05, 8.661948e-06, 
    2.874783e-06, 8.207447e-07, 4.080199e-07, 8.610091e-07, 1.747416e-06,
  0.0002799222, 0.0004159422, 0.0004749636, 0.0005013401, 0.0006851836, 
    0.0007144601, 0.0003685027, 8.022877e-05, 1.861672e-05, 9.391894e-06, 
    5.016962e-06, 3.866414e-06, 4.172409e-06, 4.681887e-06, 6.543796e-06,
  0.0003802578, 0.0004311817, 0.0003299367, 0.000295976, 0.0003825445, 
    0.0003749353, 0.0002115831, 4.187248e-05, 9.72224e-06, 8.269028e-06, 
    5.859174e-06, 5.152478e-06, 6.052248e-06, 5.761474e-06, 6.165898e-06,
  1.14808e-05, 6.27453e-05, 4.104587e-05, 5.990851e-06, 3.450523e-06, 
    3.526951e-06, 4.640582e-06, 4.343671e-06, 7.343281e-06, 1.177542e-05, 
    1.335632e-05, 1.070085e-05, 7.340232e-06, 5.302123e-06, 2.625185e-06,
  0.0001097794, 0.0001563343, 9.355469e-05, 1.607661e-05, 4.61196e-06, 
    4.419941e-06, 1.80222e-06, 1.12773e-06, 1.245835e-06, 2.304971e-06, 
    3.543559e-06, 7.633402e-06, 9.18715e-06, 1.58177e-05, 9.561639e-06,
  8.649721e-05, 0.0001548038, 7.265233e-05, 9.809922e-06, 5.607905e-06, 
    5.565396e-06, 2.062582e-06, 1.094215e-06, 7.033449e-07, 8.707232e-07, 
    3.642667e-07, 5.217059e-07, 1.242529e-06, 3.514836e-06, 5.626935e-06,
  4.839036e-05, 9.038855e-05, 5.324209e-05, 2.428885e-05, 2.162495e-05, 
    1.84221e-05, 1.448983e-05, 4.120996e-06, 1.838375e-06, 9.214445e-07, 
    9.807605e-07, 1.695108e-07, 8.224722e-08, 1.050122e-07, 2.049959e-07,
  2.019728e-05, 6.65934e-05, 7.671096e-05, 6.302153e-05, 5.694475e-05, 
    6.752301e-05, 4.251055e-05, 1.694144e-05, 4.420257e-06, 1.735514e-06, 
    2.240834e-07, 6.65747e-07, 9.674909e-07, 3.086331e-07, 8.036032e-08,
  1.415106e-05, 4.562666e-05, 7.954023e-05, 9.698276e-05, 0.0001095339, 
    0.0001010674, 7.766141e-05, 3.772947e-05, 1.494701e-05, 6.63634e-06, 
    4.072476e-06, 2.593991e-06, 3.007831e-06, 2.223454e-06, 2.103794e-07,
  5.162871e-06, 1.974914e-05, 6.085276e-05, 9.702341e-05, 0.0001196651, 
    0.0001364005, 0.0001186483, 7.068837e-05, 4.200533e-05, 1.360802e-05, 
    7.729891e-06, 6.884385e-06, 4.45144e-06, 3.025991e-06, 7.888656e-07,
  5.780376e-06, 1.295343e-05, 2.952013e-05, 6.580137e-05, 9.667216e-05, 
    0.0001289583, 0.0001347602, 0.0001106493, 6.115766e-05, 2.32435e-05, 
    7.69375e-06, 5.642315e-06, 3.242687e-06, 1.974063e-06, 4.157606e-06,
  8.581061e-06, 1.455611e-05, 1.807713e-05, 2.697448e-05, 5.440107e-05, 
    0.0001122291, 0.000165685, 0.0001190192, 6.996369e-05, 3.923661e-05, 
    1.210142e-05, 5.834986e-06, 4.617295e-06, 4.914371e-06, 3.315259e-06,
  6.440586e-06, 1.062305e-05, 1.206656e-05, 1.046576e-05, 1.005594e-05, 
    6.747404e-05, 0.0002200059, 0.000194043, 0.0001115175, 6.119531e-05, 
    2.658499e-05, 8.902966e-06, 5.016814e-06, 4.355901e-06, 3.847546e-06,
  1.962107e-05, 7.887809e-05, 0.0002246438, 0.0001672057, 3.351721e-05, 
    1.694115e-05, 1.072563e-05, 7.78205e-06, 1.297484e-05, 3.39053e-05, 
    8.188033e-05, 0.0001531622, 0.000161487, 8.081417e-05, 1.999493e-06,
  3.769011e-05, 5.225662e-05, 8.498099e-05, 5.431738e-05, 2.419337e-05, 
    2.438211e-05, 1.62773e-05, 1.072105e-05, 2.677382e-05, 7.593928e-05, 
    0.0001391884, 0.0001776574, 0.0001634113, 7.276454e-05, 3.699546e-06,
  2.443369e-05, 3.033407e-05, 2.007272e-05, 2.941113e-05, 2.007333e-05, 
    2.080479e-05, 3.660894e-05, 5.889349e-05, 0.00012839, 0.0002231581, 
    0.0002709522, 0.0002062805, 8.634543e-05, 1.855874e-05, 4.586261e-06,
  2.80823e-05, 1.802802e-05, 1.914329e-05, 2.210125e-05, 3.55927e-05, 
    5.481683e-05, 0.0001075653, 0.0001590463, 0.0002538613, 0.0003661156, 
    0.0003678489, 0.0002257793, 7.82639e-05, 1.3715e-05, 3.975243e-06,
  2.502361e-05, 1.895409e-05, 1.110084e-05, 1.534152e-05, 3.55599e-05, 
    6.650627e-05, 0.0001236246, 0.0001843518, 0.000240658, 0.0003036961, 
    0.0002769669, 0.0001567896, 7.568576e-05, 2.937051e-05, 1.510339e-05,
  9.525945e-06, 7.810894e-06, 3.5559e-06, 4.072715e-06, 8.371453e-06, 
    4.36728e-05, 7.241908e-05, 0.000106652, 0.0001423664, 0.0001724912, 
    0.0001013398, 4.637623e-05, 2.09409e-05, 1.258004e-05, 7.021988e-06,
  1.420216e-06, 4.218581e-06, 3.558847e-06, 1.096645e-06, 1.371892e-06, 
    1.085593e-05, 3.666132e-05, 5.538817e-05, 7.006267e-05, 6.200831e-05, 
    4.027971e-05, 1.520335e-05, 8.069446e-06, 3.156415e-06, 2.965786e-06,
  1.647017e-07, 1.169345e-06, 5.857524e-07, 3.548545e-07, 4.054817e-08, 
    1.479804e-06, 7.823554e-06, 3.61592e-05, 3.761742e-05, 2.871593e-05, 
    2.911494e-05, 2.217803e-05, 5.54691e-06, 5.428722e-06, 3.27573e-06,
  5.37074e-07, 1.156768e-07, 1.326924e-07, 1.582641e-07, 4.488887e-07, 
    2.443308e-08, 6.338643e-07, 2.078274e-05, 2.648056e-05, 2.273769e-05, 
    2.340957e-05, 7.695761e-06, 4.805549e-06, 5.588267e-06, 3.726283e-06,
  1.426815e-06, 2.096025e-06, 3.959253e-06, 1.795835e-06, 1.639141e-06, 
    2.606382e-06, 8.589844e-08, 6.211341e-07, 1.947017e-05, 1.904444e-05, 
    1.152887e-05, 3.949671e-06, 3.379988e-06, 5.428538e-06, 3.792387e-06,
  1.578375e-05, 9.825753e-06, 1.786219e-05, 4.246783e-05, 5.058848e-05, 
    6.046528e-05, 6.231292e-05, 6.970791e-05, 6.723971e-05, 3.189226e-05, 
    2.534563e-05, 3.118177e-05, 0.0001096521, 0.000237176, 0.0003039556,
  2.278139e-05, 1.229402e-05, 1.236679e-05, 2.382141e-05, 2.717365e-05, 
    4.023846e-05, 3.808748e-05, 4.209427e-05, 3.700955e-05, 3.165647e-05, 
    2.371612e-05, 3.929686e-05, 7.61207e-05, 0.0001392564, 0.0001156514,
  5.097077e-05, 3.57677e-05, 3.076452e-05, 3.275807e-05, 3.604448e-05, 
    3.705423e-05, 3.457838e-05, 2.41806e-05, 3.06833e-05, 2.54544e-05, 
    3.058432e-05, 3.289097e-05, 2.908405e-05, 2.173187e-05, 1.687498e-05,
  0.0001115479, 8.690375e-05, 4.839717e-05, 4.143355e-05, 2.538662e-05, 
    2.10107e-05, 2.09311e-05, 2.435351e-05, 2.012084e-05, 2.114144e-05, 
    2.179499e-05, 2.909045e-05, 2.25473e-05, 1.512184e-05, 2.177569e-05,
  0.0001131495, 9.094696e-05, 5.545321e-05, 3.205362e-05, 2.392465e-05, 
    1.736703e-05, 1.571053e-05, 1.538594e-05, 1.672244e-05, 2.130149e-05, 
    2.242414e-05, 3.129866e-05, 2.188508e-05, 1.827535e-05, 3.001852e-05,
  0.0001377628, 0.0001317373, 0.0001045122, 6.354759e-05, 4.560215e-05, 
    3.320465e-05, 2.328205e-05, 2.092028e-05, 2.325564e-05, 2.621359e-05, 
    2.602716e-05, 2.204272e-05, 2.629041e-05, 3.924543e-05, 5.119501e-05,
  0.0001793456, 0.0001827275, 0.0001907173, 0.0001696632, 0.00014402, 
    0.000123056, 8.848454e-05, 7.555861e-05, 5.89056e-05, 5.534697e-05, 
    6.457853e-05, 6.743556e-05, 7.564246e-05, 8.178477e-05, 8.536929e-05,
  0.000222765, 0.0002481084, 0.0002254394, 0.0002084294, 0.0002049011, 
    0.0001733464, 0.0001526347, 0.0001407941, 0.0001401785, 0.000134651, 
    0.0001178752, 0.0001346027, 0.0001289123, 0.0001286338, 0.0001403636,
  0.0002167218, 0.0002551146, 0.0002282848, 0.0002039903, 0.0001979379, 
    0.0001671308, 0.0001408974, 0.0001200229, 0.000115961, 0.0001157227, 
    0.0001429147, 0.0001618699, 0.0001727052, 0.0001804348, 0.0001882967,
  0.0001062806, 0.0001641684, 0.0001981683, 0.0002133769, 0.0002141718, 
    0.0002052687, 0.0001590633, 0.0001121065, 0.0001049862, 0.0001159713, 
    0.0001396218, 0.0001658338, 0.0001719198, 0.0001962546, 0.0002297608,
  7.311959e-06, 3.834831e-06, 5.011252e-06, 2.470787e-05, 2.452831e-05, 
    2.248352e-05, 2.880025e-05, 5.109047e-05, 5.86989e-05, 8.759512e-05, 
    9.036643e-05, 7.965221e-05, 7.194175e-05, 5.383972e-05, 5.985448e-05,
  6.676185e-06, 5.64472e-06, 8.683652e-06, 2.043398e-05, 1.947773e-05, 
    2.451715e-05, 2.892818e-05, 2.926094e-05, 5.153801e-05, 6.307845e-05, 
    8.305912e-05, 8.333941e-05, 6.787913e-05, 6.486541e-05, 6.106011e-05,
  4.565785e-06, 3.423959e-06, 1.811241e-05, 2.162574e-05, 2.331457e-05, 
    2.832055e-05, 2.666379e-05, 3.402814e-05, 4.471456e-05, 4.621956e-05, 
    6.364552e-05, 6.402666e-05, 6.522284e-05, 7.022054e-05, 4.946957e-05,
  2.605769e-06, 2.421644e-06, 1.040735e-05, 2.215041e-05, 2.529437e-05, 
    2.604606e-05, 2.969771e-05, 2.880554e-05, 2.995168e-05, 3.548549e-05, 
    4.925333e-05, 5.44515e-05, 6.321693e-05, 5.826378e-05, 4.578682e-05,
  1.12539e-06, 1.662746e-06, 4.446641e-06, 1.666397e-05, 2.79306e-05, 
    2.411455e-05, 2.09513e-05, 2.315416e-05, 2.201443e-05, 2.694559e-05, 
    3.246126e-05, 4.065734e-05, 4.292614e-05, 4.216267e-05, 3.789591e-05,
  1.120362e-07, 9.903439e-07, 2.886105e-06, 5.638579e-06, 2.837099e-05, 
    2.615817e-05, 1.900109e-05, 1.750017e-05, 1.796114e-05, 1.957552e-05, 
    2.003724e-05, 2.135178e-05, 2.831974e-05, 2.661835e-05, 3.472789e-05,
  4.662063e-09, 9.939672e-09, 9.637718e-07, 4.921647e-06, 1.797952e-05, 
    2.364585e-05, 2.143672e-05, 1.543545e-05, 1.447404e-05, 1.20314e-05, 
    1.201488e-05, 1.625685e-05, 1.704115e-05, 2.098458e-05, 2.433164e-05,
  3.824026e-09, 3.692625e-08, 7.093897e-07, 3.421608e-06, 8.544331e-06, 
    1.784625e-05, 2.219552e-05, 1.63527e-05, 1.270317e-05, 1.026937e-05, 
    1.065227e-05, 9.515039e-06, 1.179563e-05, 1.53552e-05, 1.706449e-05,
  6.443584e-08, 1.365635e-07, 3.516835e-07, 2.276643e-06, 7.596332e-06, 
    1.182827e-05, 2.024596e-05, 2.056788e-05, 1.442212e-05, 1.05499e-05, 
    8.88011e-06, 8.4425e-06, 9.802268e-06, 1.094193e-05, 3.07321e-05,
  2.255664e-08, 1.940071e-08, 2.282264e-07, 6.33575e-07, 5.803928e-06, 
    1.11896e-05, 1.30112e-05, 2.266286e-05, 1.870188e-05, 1.253486e-05, 
    8.381833e-06, 8.312352e-06, 1.106622e-05, 1.960376e-05, 5.271997e-05,
  1.684483e-08, 3.820791e-10, 4.014137e-07, 2.694163e-06, 3.255519e-06, 
    5.149718e-06, 4.496786e-06, 5.959388e-06, 6.605631e-06, 9.826515e-06, 
    9.615532e-06, 1.162374e-05, 1.435914e-05, 1.645891e-05, 4.057149e-05,
  1.161384e-06, 2.60747e-07, 4.140487e-08, 4.067807e-06, 3.424471e-06, 
    4.287487e-06, 4.98724e-06, 5.339209e-06, 6.712861e-06, 8.604642e-06, 
    9.199888e-06, 1.085963e-05, 1.38966e-05, 1.847501e-05, 3.255907e-05,
  2.24567e-06, 2.694599e-06, 2.00879e-06, 2.819001e-06, 3.268123e-06, 
    2.52541e-06, 3.261437e-06, 4.945647e-06, 4.081662e-06, 6.643355e-06, 
    8.061316e-06, 1.070954e-05, 1.313784e-05, 1.863552e-05, 1.893924e-05,
  2.581906e-06, 3.628593e-06, 3.314924e-06, 3.561241e-06, 3.273342e-06, 
    3.431654e-06, 2.204856e-06, 2.75738e-06, 3.272311e-06, 4.079932e-06, 
    8.096226e-06, 9.457293e-06, 1.408809e-05, 1.746713e-05, 2.861998e-05,
  2.740709e-06, 3.618076e-06, 2.796352e-06, 3.37996e-06, 2.928121e-06, 
    3.139843e-06, 1.193743e-06, 1.850723e-06, 2.952577e-06, 3.986217e-06, 
    4.373341e-06, 7.352167e-06, 1.074639e-05, 1.82322e-05, 2.28665e-05,
  1.561234e-06, 2.790545e-06, 2.815947e-06, 2.402634e-06, 3.269959e-06, 
    4.068154e-06, 1.812164e-06, 1.758217e-06, 1.614503e-06, 2.347215e-06, 
    3.4124e-06, 4.928462e-06, 7.908533e-06, 1.118907e-05, 1.813109e-05,
  5.764087e-07, 1.597312e-06, 3.126331e-06, 2.85323e-06, 2.725632e-06, 
    2.715472e-06, 2.145751e-06, 1.937758e-06, 2.401772e-06, 1.747973e-06, 
    3.826351e-06, 4.868113e-06, 7.907607e-06, 9.42286e-06, 1.320283e-05,
  4.314972e-09, 1.14475e-06, 1.578642e-06, 3.469814e-06, 1.656053e-06, 
    1.254169e-06, 2.762655e-06, 1.605802e-06, 2.020114e-06, 1.763197e-06, 
    1.949e-06, 4.246996e-06, 5.297557e-06, 8.106219e-06, 9.682132e-06,
  4.531873e-07, 5.682901e-07, 9.666419e-07, 1.83408e-06, 2.058227e-06, 
    2.297043e-06, 2.163282e-06, 2.189742e-06, 2.318048e-06, 1.836145e-06, 
    1.704516e-06, 3.113633e-06, 4.207635e-06, 4.614039e-06, 7.977584e-06,
  3.457271e-06, 9.402557e-07, 6.527734e-07, 2.324982e-06, 1.83982e-06, 
    2.285737e-06, 1.245952e-06, 3.089633e-06, 2.776667e-06, 1.931418e-06, 
    1.578239e-06, 1.629744e-06, 2.156884e-06, 5.210484e-06, 6.146636e-06,
  5.003338e-06, 5.533388e-06, 4.44243e-06, 2.64182e-05, 3.063469e-05, 
    1.970104e-05, 1.184457e-05, 7.096382e-06, 5.046727e-06, 5.323835e-06, 
    5.626931e-06, 7.187889e-06, 5.803607e-06, 4.573116e-06, 5.567956e-06,
  1.724835e-05, 1.161973e-05, 5.393683e-06, 4.329412e-05, 4.117877e-05, 
    2.069166e-05, 1.16486e-05, 9.176383e-06, 3.119818e-06, 2.47409e-06, 
    4.225193e-06, 5.304135e-06, 7.676534e-06, 4.882089e-06, 4.64311e-06,
  1.29653e-05, 2.196396e-05, 2.068675e-05, 5.171169e-05, 5.572937e-05, 
    3.053708e-05, 1.28202e-05, 4.390336e-06, 2.616987e-06, 3.39954e-06, 
    4.47402e-06, 6.121707e-06, 6.066294e-06, 6.481741e-06, 6.446066e-06,
  1.149643e-05, 1.714641e-05, 2.570164e-05, 4.622601e-05, 5.15733e-05, 
    2.546678e-05, 9.41836e-06, 4.877847e-06, 2.200837e-06, 1.727046e-06, 
    1.356494e-06, 3.639936e-06, 3.763011e-06, 4.103165e-06, 5.64857e-06,
  9.91856e-06, 1.217526e-05, 9.878851e-06, 2.92046e-05, 3.429287e-05, 
    1.847148e-05, 8.095927e-06, 5.893322e-06, 4.20374e-06, 3.142881e-06, 
    3.236341e-06, 2.520413e-06, 2.541881e-06, 2.996784e-06, 4.644388e-06,
  3.853307e-06, 7.731428e-06, 8.143174e-06, 1.044138e-05, 2.061414e-05, 
    2.230165e-05, 1.426432e-05, 7.593845e-06, 6.045184e-06, 5.726085e-06, 
    5.115774e-06, 3.64272e-06, 2.861915e-06, 1.655615e-06, 1.832327e-06,
  9.082662e-06, 9.583303e-06, 1.128606e-05, 7.36945e-06, 1.136572e-05, 
    1.680636e-05, 1.855115e-05, 1.278732e-05, 6.476532e-06, 4.855311e-06, 
    4.718615e-06, 4.761712e-06, 3.813546e-06, 3.276022e-06, 4.672076e-06,
  2.664727e-05, 1.395794e-05, 4.428187e-06, 6.127297e-06, 2.154899e-06, 
    1.01293e-05, 2.034072e-05, 1.591708e-05, 9.965711e-06, 6.939674e-06, 
    4.85605e-06, 4.176374e-06, 3.877084e-06, 3.646265e-06, 2.609404e-06,
  4.752413e-05, 2.967255e-05, 9.011885e-06, 2.797758e-06, 3.122047e-06, 
    5.307043e-06, 1.467658e-05, 1.458222e-05, 1.262071e-05, 7.585203e-06, 
    5.835336e-06, 3.835964e-06, 3.707983e-06, 4.238136e-06, 2.433403e-06,
  4.619571e-05, 4.861266e-05, 1.851375e-05, 5.056681e-06, 2.578708e-06, 
    3.873956e-06, 1.272138e-05, 1.034951e-05, 1.353229e-05, 8.365321e-06, 
    6.81863e-06, 7.168444e-06, 5.687597e-06, 3.924592e-06, 2.548036e-06,
  1.010511e-05, 5.265053e-06, 3.344956e-05, 0.0004126913, 0.0006233438, 
    0.0003633042, 3.888679e-05, 1.511625e-05, 3.515523e-06, 1.730316e-06, 
    2.412096e-06, 1.292035e-05, 1.039336e-05, 3.108363e-06, 3.820323e-06,
  2.504414e-05, 2.815859e-06, 1.380784e-05, 0.0002754412, 0.000472641, 
    0.0001881958, 2.772609e-05, 8.015617e-06, 3.787294e-06, 2.080927e-06, 
    1.558461e-06, 5.840518e-06, 1.333397e-05, 9.961151e-06, 3.259685e-06,
  1.95297e-05, 3.515881e-05, 4.893432e-05, 0.0001794183, 0.0002812622, 
    0.0001001406, 2.164464e-05, 6.587828e-06, 4.376529e-06, 2.072285e-06, 
    1.750733e-06, 1.358295e-06, 4.505203e-06, 5.867412e-06, 3.587511e-06,
  1.231001e-05, 3.681207e-05, 3.941394e-05, 7.336969e-05, 0.0001182233, 
    6.438652e-05, 2.181279e-05, 9.217136e-06, 6.209353e-06, 4.045826e-06, 
    2.470751e-06, 1.813631e-06, 1.466765e-06, 2.076128e-06, 3.021554e-06,
  1.216839e-05, 6.72245e-06, 9.821195e-06, 5.389801e-05, 6.847047e-05, 
    6.475028e-05, 3.323268e-05, 1.378039e-05, 1.08101e-05, 9.016168e-06, 
    5.181963e-06, 2.977031e-06, 3.221576e-06, 1.611486e-06, 2.483503e-06,
  2.18725e-05, 9.62623e-06, 5.986755e-06, 4.666223e-06, 3.575991e-05, 
    6.07188e-05, 4.678592e-05, 2.520314e-05, 1.505559e-05, 1.097425e-05, 
    9.563119e-06, 5.135103e-06, 2.734102e-06, 3.01062e-06, 1.91997e-06,
  3.179467e-05, 1.931379e-05, 2.834308e-05, 1.299996e-05, 1.509585e-05, 
    3.376889e-05, 4.703368e-05, 3.997847e-05, 2.531131e-05, 1.651538e-05, 
    1.257411e-05, 7.797174e-06, 5.184093e-06, 2.964301e-06, 2.410738e-06,
  7.777425e-05, 6.716155e-05, 6.960836e-05, 5.045845e-05, 1.880433e-05, 
    2.795534e-05, 4.262256e-05, 5.089012e-05, 3.778866e-05, 2.41923e-05, 
    1.67935e-05, 1.340637e-05, 7.958253e-06, 4.949145e-06, 3.067657e-06,
  0.0001126213, 0.0001073977, 8.338322e-05, 0.0001007254, 8.678444e-05, 
    4.280694e-05, 5.014194e-05, 5.345439e-05, 4.007131e-05, 2.766353e-05, 
    1.928773e-05, 1.709888e-05, 1.075298e-05, 5.821365e-06, 3.487632e-06,
  4.346263e-05, 7.215331e-05, 8.963753e-05, 7.82425e-05, 9.981186e-05, 
    5.567789e-05, 5.714586e-05, 4.256159e-05, 3.619424e-05, 2.565118e-05, 
    1.907162e-05, 1.508315e-05, 1.433265e-05, 1.159453e-05, 5.981453e-06,
  9.820388e-07, 2.288119e-06, 1.746013e-06, 2.33779e-05, 6.67841e-05, 
    0.0002571627, 0.0003602159, 0.0002336823, 0.0002542485, 0.0002763578, 
    0.0002578889, 0.000199993, 9.076291e-05, 1.142852e-05, 3.396012e-06,
  8.668909e-06, 1.764222e-06, 3.711864e-07, 3.075514e-05, 4.568594e-05, 
    0.0002278626, 0.0003060797, 0.0002933142, 0.0002884255, 0.0003140378, 
    0.0003656072, 0.000347367, 0.0001849951, 4.172873e-05, 4.91911e-06,
  8.062892e-06, 5.808907e-06, 9.636124e-06, 1.946805e-05, 4.859289e-05, 
    0.0001252037, 0.000276503, 0.0002375425, 0.0003390417, 0.000343799, 
    0.0003973183, 0.0004030529, 0.000262903, 7.810551e-05, 5.27098e-06,
  9.172087e-06, 7.491493e-06, 6.438464e-06, 1.929837e-05, 3.079052e-05, 
    9.036709e-05, 0.0002520055, 0.0003415912, 0.0004162915, 0.0003437238, 
    0.0003639823, 0.0003788695, 0.0002640315, 9.532918e-05, 8.316471e-06,
  1.00115e-05, 5.954655e-06, 1.378057e-06, 7.870184e-06, 2.430796e-05, 
    6.44604e-05, 0.0002219114, 0.0004769863, 0.0004286154, 0.000308157, 
    0.0001923834, 0.0001468703, 9.718332e-05, 3.530828e-05, 5.848941e-06,
  1.79438e-05, 1.71487e-05, 9.714478e-06, 3.403066e-06, 1.359929e-05, 
    5.787997e-05, 0.0001378305, 0.0002926448, 0.000249569, 0.0001697057, 
    7.927399e-05, 3.807027e-05, 1.824284e-05, 6.349579e-06, 5.307117e-06,
  1.962593e-05, 2.702445e-05, 2.781599e-05, 2.156025e-05, 1.315741e-05, 
    6.384515e-05, 0.0001010547, 0.0001511014, 0.0001304459, 8.803626e-05, 
    7.612139e-05, 2.844424e-05, 8.603795e-06, 4.39618e-06, 8.741396e-06,
  2.786744e-05, 2.846401e-05, 4.459959e-05, 4.35612e-05, 3.07662e-06, 
    1.911342e-05, 7.598419e-05, 9.026084e-05, 9.920231e-05, 5.843718e-05, 
    4.423459e-05, 2.978071e-05, 1.540899e-05, 7.245288e-06, 7.699537e-06,
  6.516595e-05, 4.165837e-05, 7.008488e-05, 3.724774e-05, 2.351538e-05, 
    3.892355e-06, 2.57418e-05, 7.767089e-05, 4.413553e-05, 3.097211e-05, 
    3.837797e-05, 2.137107e-05, 2.610608e-05, 2.19961e-05, 8.164897e-06,
  7.888653e-05, 5.84077e-05, 3.478393e-05, 4.635186e-05, 2.003156e-05, 
    2.181409e-05, 2.42181e-05, 7.539096e-05, 4.967611e-05, 3.538863e-05, 
    2.827653e-05, 1.840632e-05, 2.398556e-05, 2.121399e-05, 9.519879e-06,
  4.978704e-06, 1.759227e-06, 1.67285e-06, 1.10177e-05, 6.976152e-06, 
    6.000755e-06, 3.734915e-06, 4.795313e-06, 5.768029e-06, 8.783072e-06, 
    1.077976e-05, 2.963994e-05, 2.687008e-05, 2.772716e-05, 3.747433e-05,
  1.421249e-05, 1.26606e-06, 1.59369e-07, 4.230227e-07, 4.716081e-06, 
    1.031543e-05, 1.27381e-05, 1.79388e-05, 1.797678e-05, 8.885769e-06, 
    2.830611e-05, 8.261864e-05, 0.0001458393, 0.0001732177, 0.0002045369,
  1.28394e-05, 1.392092e-05, 9.573603e-06, 6.500863e-06, 1.701978e-05, 
    4.635954e-05, 7.346174e-05, 6.330858e-05, 1.940113e-05, 5.744909e-05, 
    8.488999e-05, 0.0001459509, 0.0002547601, 0.0002895985, 0.0002412652,
  3.448243e-05, 5.470843e-05, 5.888152e-05, 6.192501e-05, 8.133106e-05, 
    6.193468e-05, 0.0001764489, 0.0001571627, 2.106462e-05, 3.711859e-05, 
    4.919952e-05, 9.22784e-05, 0.0001856361, 0.0002413477, 0.0001746938,
  0.0001081109, 0.0001468624, 6.870245e-05, 3.834778e-05, 2.618314e-05, 
    7.667603e-06, 1.294422e-05, 7.420932e-05, 6.040136e-06, 2.073921e-05, 
    4.328848e-05, 6.766112e-05, 7.980235e-05, 9.110268e-05, 7.571896e-05,
  0.0001867315, 0.0001975168, 0.0001956295, 3.634739e-08, 9.710585e-08, 
    8.918079e-08, 8.951299e-08, 1.637972e-05, 1.603199e-05, 6.690836e-06, 
    3.737998e-05, 5.508687e-05, 4.891106e-05, 1.362016e-05, 9.740642e-06,
  0.0002090515, 0.0001818316, 0.0001948524, 0.000114359, 2.07509e-08, 
    2.468765e-08, 1.582879e-08, 5.645765e-08, 4.660296e-06, 2.477497e-05, 
    3.589998e-05, 2.196022e-05, 1.07165e-05, 1.001237e-05, 9.019422e-06,
  0.0001518771, 0.0001428593, 0.0001211881, 9.02005e-05, 2.037223e-08, 
    4.189693e-09, 9.083018e-10, 7.169808e-09, 1.485755e-06, 7.014616e-06, 
    2.469422e-05, 2.2861e-05, 1.230947e-05, 8.193795e-06, 5.475955e-06,
  6.84561e-05, 6.981008e-05, 6.722563e-05, 5.119656e-05, 3.034293e-05, 
    2.99945e-09, 7.839583e-10, 6.932797e-10, 3.283862e-07, 1.502237e-06, 
    6.185639e-06, 7.123242e-06, 8.062571e-06, 4.845698e-06, 1.345968e-06,
  5.413259e-05, 5.432315e-05, 3.735846e-05, 2.296302e-05, 2.386882e-05, 
    2.101327e-05, 2.664983e-10, 1.215184e-10, 7.946706e-08, 5.789404e-07, 
    3.01956e-06, 4.827045e-06, 7.039161e-06, 3.533742e-06, 1.469423e-06,
  1.373538e-09, 5.434843e-10, 1.278015e-10, 6.916707e-11, 1.07187e-10, 
    1.334238e-10, 4.550796e-10, 1.583817e-08, 3.561109e-07, 1.239393e-06, 
    1.69597e-08, 2.085409e-09, 2.055037e-08, 8.646544e-08, 3.873634e-07,
  1.712697e-08, 6.332281e-10, 1.115431e-10, 1.832143e-10, 1.592918e-10, 
    1.094714e-10, 9.380564e-11, 9.729469e-11, 2.55715e-10, 3.51467e-10, 
    3.481643e-06, 8.576521e-06, 1.351618e-05, 5.946001e-05, 0.0001493283,
  2.414056e-05, 9.508875e-09, 1.052145e-09, 1.839849e-09, 2.031836e-08, 
    4.689583e-08, 2.428286e-06, 5.764392e-06, 2.358949e-05, 4.606745e-05, 
    0.0001134253, 0.0002084638, 0.0003012626, 0.0004164746, 0.000500321,
  3.332467e-05, 1.630217e-05, 3.687499e-06, 2.687585e-05, 7.603551e-05, 
    0.0001172142, 0.0001510327, 0.0003039039, 0.0002476352, 0.0003542472, 
    0.0004627672, 0.0005416155, 0.0005715387, 0.0005599312, 0.0004779736,
  0.0001015763, 6.720748e-05, 1.614267e-05, 3.827789e-05, 6.71454e-05, 
    0.0001069416, 0.0001387252, 0.0002210231, 0.0003488752, 0.0003600781, 
    0.0004020994, 0.0004269908, 0.0004502448, 0.0004744678, 0.0004681368,
  0.0001391363, 8.406249e-05, 9.633925e-05, 6.162482e-06, 9.294331e-07, 
    1.444933e-06, 9.477572e-06, 5.271825e-05, 0.0001019683, 0.0001209187, 
    0.0001626051, 0.0002029025, 0.0002439899, 0.0002909973, 0.0003110768,
  0.0001758997, 0.0001996531, 0.0002375502, 0.0001358628, 1.02871e-06, 
    4.251706e-07, 4.485738e-07, 2.37151e-06, 5.615726e-05, 6.083939e-05, 
    7.092136e-05, 7.329119e-05, 8.2812e-05, 0.0001227628, 0.0001741275,
  0.0001157304, 0.0001700507, 0.0002275588, 0.000236191, 4.668535e-07, 
    6.024064e-08, 2.141119e-08, 3.791986e-08, 1.422381e-06, 5.237227e-05, 
    7.425342e-05, 7.117193e-05, 6.894036e-05, 8.433167e-05, 4.760167e-05,
  8.763354e-05, 8.058258e-05, 8.724222e-05, 0.0001470871, 9.588431e-05, 
    7.051702e-08, 7.561291e-09, 5.977048e-09, 3.485682e-07, 5.443289e-07, 
    3.46622e-05, 4.412554e-05, 4.561227e-05, 3.065634e-05, 3.042918e-07,
  5.749825e-05, 8.767299e-05, 9.337591e-05, 8.739685e-05, 7.011242e-05, 
    6.175665e-05, 1.933772e-09, 5.242156e-10, 2.463232e-07, 2.891373e-08, 
    3.774566e-06, 1.554929e-05, 2.979865e-05, 2.429882e-05, 2.361387e-05,
  2.960703e-08, 2.139218e-08, 1.206459e-08, 9.884357e-10, 2.624808e-09, 
    1.224487e-09, 4.645513e-10, 9.663086e-11, 1.726759e-10, 5.505617e-11, 
    2.553766e-10, 3.77109e-08, 3.360515e-07, 7.960984e-07, 1.939486e-06,
  8.491861e-06, 7.696664e-07, 1.313993e-06, 6.506465e-08, 1.334859e-08, 
    2.076223e-09, 4.040564e-09, 1.150827e-09, 9.778259e-10, 5.815449e-10, 
    7.219987e-11, 2.564738e-11, 1.2433e-10, 1.647913e-08, 9.961627e-08,
  3.970419e-05, 7.888041e-06, 2.917543e-06, 1.957115e-06, 5.059935e-08, 
    1.577291e-08, 2.454672e-09, 1.860273e-09, 6.110906e-10, 2.026291e-09, 
    1.815317e-09, 8.726434e-10, 1.765646e-09, 1.794279e-10, 2.380361e-10,
  0.0001454098, 6.349355e-05, 8.311702e-07, 9.149432e-08, 5.166261e-08, 
    4.485116e-09, 2.560746e-10, 2.168448e-10, 2.528029e-09, 2.040552e-09, 
    2.898101e-10, 2.460429e-10, 9.14499e-11, 9.540321e-11, 1.454305e-09,
  0.0001493932, 5.015797e-05, 1.404879e-05, 1.631118e-07, 6.734166e-08, 
    3.510137e-07, 1.110129e-08, 1.289593e-09, 7.356766e-10, 8.654428e-10, 
    1.901351e-09, 3.447857e-09, 5.158368e-09, 3.537421e-09, 1.944072e-09,
  0.000336759, 0.0001845613, 2.356743e-05, 6.458789e-06, 3.171175e-06, 
    9.311273e-07, 1.799347e-07, 1.533653e-07, 1.520733e-08, 1.630251e-08, 
    6.44785e-09, 7.174742e-10, 5.617534e-10, 2.166688e-09, 2.385483e-09,
  0.0003137198, 0.0003250976, 9.348661e-05, 5.378188e-05, 3.121395e-05, 
    2.254556e-05, 7.501723e-05, 1.565254e-05, 8.619426e-06, 9.978591e-06, 
    6.973639e-06, 1.786047e-06, 3.277596e-07, 8.132761e-07, 2.34923e-06,
  0.0001883733, 0.000213298, 0.0002982367, 0.0003608025, 0.0001432862, 
    8.364745e-07, 3.071424e-05, 5.708841e-05, 7.3984e-05, 0.0001811291, 
    0.0002240628, 0.0001859108, 8.675003e-05, 6.724062e-05, 8.034168e-05,
  8.202199e-05, 0.0001223023, 0.0001650199, 0.0002472467, 0.0003053711, 
    6.178564e-06, 8.135731e-07, 2.68109e-05, 5.103007e-05, 0.0002781443, 
    0.0002959826, 0.0001902857, 0.0002427406, 0.0001935095, 0.0001321466,
  9.192547e-05, 9.85939e-05, 0.0001098327, 0.0001792354, 0.0002340767, 
    0.0001374923, 1.074898e-07, 2.003181e-07, 3.110288e-06, 8.616113e-05, 
    0.0001262502, 0.0001431799, 0.0001279887, 0.0001699835, 0.0001406584,
  3.011573e-06, 1.897637e-07, 1.729864e-09, 2.8435e-13, 2.738337e-14, 
    1.933457e-13, 9.366046e-11, 1.212205e-10, 9.353309e-10, 2.397587e-08, 
    2.093525e-08, 8.48686e-08, 8.360683e-07, 2.296248e-06, 1.639125e-06,
  1.753642e-05, 2.06609e-06, 3.775257e-08, 2.416916e-10, 1.550716e-11, 
    2.855359e-14, 4.535506e-13, 3.036646e-11, 7.045923e-11, 1.522601e-10, 
    6.093748e-10, 1.549166e-07, 1.922648e-07, 3.919961e-07, 1.554924e-06,
  1.653782e-05, 1.002088e-05, 4.725584e-07, 5.877971e-09, 5.073216e-12, 
    8.511536e-12, 2.729405e-12, 1.679826e-11, 2.403466e-11, 1.808856e-11, 
    2.879498e-11, 1.828675e-10, 1.919077e-10, 1.60375e-07, 3.901173e-07,
  2.941709e-05, 1.437531e-05, 1.211974e-06, 3.510265e-08, 1.084394e-10, 
    1.97696e-11, 1.531175e-09, 2.256497e-09, 5.302838e-10, 2.633555e-11, 
    4.222239e-11, 3.40142e-10, 1.487815e-12, 5.784876e-11, 4.48456e-10,
  3.888884e-05, 2.759616e-05, 2.101803e-06, 1.710489e-07, 1.018852e-07, 
    4.325455e-08, 4.683923e-08, 6.14818e-07, 2.962961e-07, 2.170897e-07, 
    8.332578e-08, 1.799351e-09, 8.394267e-11, 4.112335e-12, 3.424779e-12,
  6.995413e-05, 3.858575e-05, 2.884053e-05, 4.253865e-06, 6.738284e-06, 
    1.792347e-06, 1.287358e-06, 1.51704e-06, 2.507969e-06, 3.355822e-06, 
    3.011096e-06, 9.501134e-07, 3.886908e-08, 1.333455e-10, 1.891278e-12,
  8.348507e-05, 0.0001017112, 3.067441e-05, 2.382007e-05, 4.142555e-06, 
    5.104387e-06, 1.341143e-05, 1.573968e-05, 1.933742e-05, 2.20484e-05, 
    9.847778e-06, 4.588342e-06, 1.452031e-06, 1.065041e-08, 1.635916e-08,
  9.591059e-05, 0.0001123218, 0.0001120375, 8.736997e-05, 5.858183e-06, 
    1.02795e-05, 2.937824e-05, 5.591579e-05, 7.231519e-05, 5.166527e-05, 
    3.689839e-05, 3.40484e-05, 2.662809e-05, 1.1388e-05, 5.852206e-06,
  5.811355e-05, 8.588179e-05, 0.0001383962, 0.0001901417, 0.0002109002, 
    2.692792e-05, 5.687831e-05, 7.748604e-05, 0.0001915441, 0.0001063639, 
    6.851608e-05, 5.122064e-05, 5.200815e-05, 5.495794e-05, 3.872624e-05,
  2.027726e-05, 3.298101e-05, 7.77532e-05, 0.0002231656, 0.0002794518, 
    0.0002337962, 6.020027e-06, 5.072775e-07, 0.0001653882, 9.689512e-05, 
    5.462697e-05, 3.586812e-05, 5.65093e-05, 5.410691e-05, 5.888689e-05,
  3.078074e-07, 1.973296e-08, 7.180607e-10, 2.301905e-08, 2.007417e-06, 
    2.778088e-06, 3.91674e-06, 2.965994e-06, 1.002126e-06, 4.051838e-08, 
    3.531804e-09, 5.470339e-09, 3.594441e-07, 7.275632e-07, 1.62916e-06,
  4.839349e-06, 3.265446e-07, 4.473377e-09, 7.142152e-08, 2.21233e-06, 
    2.736286e-06, 6.737109e-06, 4.515137e-06, 3.904298e-06, 7.785182e-07, 
    1.15138e-07, 8.51267e-11, 3.881414e-09, 4.18799e-07, 2.349095e-06,
  4.438705e-06, 3.22621e-06, 9.55183e-08, 4.533798e-07, 3.649102e-06, 
    4.540206e-06, 7.711963e-06, 6.180561e-06, 4.272853e-06, 4.022878e-06, 
    2.232212e-06, 3.296811e-09, 4.529738e-10, 9.494045e-09, 9.123987e-07,
  5.665499e-06, 5.536661e-06, 1.456496e-06, 5.172615e-07, 2.556464e-06, 
    4.067231e-06, 5.874741e-06, 5.996423e-06, 6.375963e-06, 4.971671e-06, 
    1.749522e-06, 4.431101e-07, 1.292652e-08, 1.354195e-09, 2.960688e-10,
  5.116861e-06, 9.391223e-06, 1.965921e-06, 3.489561e-06, 4.716465e-06, 
    3.856745e-06, 8.840913e-06, 9.89573e-06, 1.18386e-05, 1.304655e-05, 
    6.178115e-06, 4.420644e-06, 2.038221e-06, 1.510169e-08, 1.864945e-08,
  4.348825e-06, 4.75113e-06, 6.833132e-06, 1.183235e-06, 5.030248e-06, 
    8.651064e-06, 8.436953e-06, 1.283551e-05, 1.615592e-05, 1.739741e-05, 
    3.181074e-05, 2.760693e-05, 5.153182e-06, 1.965609e-06, 1.82207e-07,
  3.407937e-06, 7.038211e-06, 1.566649e-05, 9.841493e-06, 5.303317e-06, 
    4.026869e-06, 1.30427e-05, 1.322128e-05, 1.358973e-05, 2.223843e-05, 
    2.309203e-05, 3.792789e-05, 3.650879e-05, 1.090347e-05, 4.670448e-06,
  2.187551e-06, 5.017685e-06, 2.661991e-05, 1.866407e-05, 2.359166e-07, 
    3.009823e-06, 6.89219e-06, 4.875168e-06, 4.771361e-06, 1.215493e-05, 
    1.239237e-05, 3.259625e-05, 8.660185e-05, 4.605584e-05, 1.589601e-05,
  2.433167e-06, 5.058786e-06, 1.084257e-05, 1.491649e-05, 1.867874e-05, 
    1.709282e-06, 9.796749e-06, 4.428223e-06, 7.397782e-06, 1.935612e-05, 
    2.498009e-05, 4.566426e-05, 8.796119e-05, 8.352681e-05, 6.706822e-05,
  2.623485e-06, 3.496656e-06, 9.025009e-06, 2.095454e-05, 3.066348e-05, 
    1.419441e-05, 2.099752e-05, 1.78516e-05, 1.565762e-05, 2.743271e-05, 
    5.453697e-05, 8.658721e-05, 7.459972e-05, 7.595004e-05, 5.757356e-05,
  9.784681e-06, 1.509699e-05, 2.303278e-05, 2.162773e-05, 4.077524e-06, 
    1.512695e-05, 5.884114e-06, 8.505438e-06, 1.049556e-05, 7.163304e-06, 
    1.386796e-06, 5.309534e-07, 2.173452e-06, 3.269036e-06, 4.655038e-06,
  0.0001000943, 8.131285e-06, 1.627561e-05, 1.534446e-05, 8.024845e-06, 
    6.951665e-06, 5.31926e-06, 5.974463e-06, 8.181948e-06, 4.928553e-06, 
    2.527251e-07, 2.221462e-07, 6.902093e-07, 1.56491e-06, 3.160188e-06,
  0.0001201873, 0.0001223729, 1.108756e-05, 1.165889e-05, 1.283887e-05, 
    6.055406e-06, 5.4496e-06, 5.457047e-06, 6.064968e-06, 1.648312e-06, 
    5.109692e-06, 5.511802e-07, 6.30576e-07, 1.287852e-06, 3.047631e-06,
  0.0001081666, 0.0001054857, 5.09794e-06, 6.266619e-06, 5.14225e-06, 
    5.618689e-06, 4.730992e-06, 4.342928e-06, 4.475129e-06, 4.941453e-06, 
    4.710163e-06, 8.76133e-07, 2.086333e-06, 8.09887e-07, 3.266044e-06,
  7.874288e-05, 7.449045e-05, 1.696564e-06, 2.494303e-06, 3.588924e-06, 
    6.279662e-06, 4.240054e-06, 4.043246e-06, 3.365273e-06, 2.909748e-06, 
    5.076754e-06, 6.937923e-06, 3.656523e-06, 1.844362e-06, 2.337935e-06,
  4.249538e-05, 4.901116e-05, 6.290308e-05, 1.368114e-06, 2.813062e-06, 
    9.579096e-07, 4.008223e-06, 4.209931e-06, 2.072345e-06, 2.394066e-06, 
    6.453266e-06, 5.924491e-06, 6.287365e-06, 4.827132e-06, 4.778964e-06,
  2.052188e-05, 3.173003e-05, 3.616492e-05, 3.672919e-05, 5.439957e-07, 
    1.613968e-07, 1.761375e-06, 3.488481e-06, 3.701428e-06, 1.788598e-06, 
    2.981142e-06, 5.903139e-06, 1.212665e-05, 9.103586e-06, 3.593106e-06,
  1.060418e-05, 1.402085e-05, 2.915178e-05, 4.982784e-05, 2.405569e-08, 
    7.049139e-09, 5.133837e-06, 1.243348e-06, 4.842115e-06, 3.59882e-06, 
    1.720269e-06, 3.893872e-06, 1.198422e-05, 1.582962e-05, 2.347271e-05,
  7.602375e-06, 1.167381e-05, 3.00761e-05, 4.676462e-05, 3.043281e-05, 
    2.51325e-08, 2.107705e-06, 1.888886e-06, 2.866763e-06, 4.622661e-06, 
    2.696769e-06, 4.537043e-06, 5.054212e-06, 3.016892e-06, 2.039771e-05,
  2.591221e-06, 6.138464e-06, 1.953355e-05, 4.208419e-05, 9.148712e-05, 
    3.95973e-05, 4.767206e-07, 3.826893e-06, 7.165893e-06, 4.355214e-06, 
    4.626232e-06, 5.488277e-06, 4.183712e-06, 3.836688e-06, 1.266633e-05,
  1.029474e-05, 3.232403e-06, 1.576366e-08, 1.601499e-08, 2.152072e-08, 
    4.886468e-08, 1.913412e-06, 3.53843e-06, 3.758639e-06, 2.806861e-06, 
    1.995497e-06, 3.718072e-07, 1.29022e-06, 2.489865e-06, 8.688773e-06,
  0.0001238425, 1.07399e-05, 8.923018e-07, 2.980378e-09, 5.375087e-09, 
    1.279684e-08, 2.659767e-06, 2.643376e-06, 4.01952e-06, 5.068642e-06, 
    8.0577e-07, 5.275948e-07, 4.689135e-07, 1.812252e-06, 6.820517e-06,
  0.0001526307, 7.246881e-05, 3.238606e-06, 5.007019e-09, 1.429761e-07, 
    1.638817e-06, 1.772533e-06, 1.844396e-06, 3.107531e-06, 1.888934e-06, 
    1.467134e-06, 1.145111e-06, 1.376761e-06, 3.023904e-06, 5.447309e-06,
  0.0001382299, 9.045643e-05, 2.687871e-06, 7.841338e-09, 3.48756e-09, 
    1.519984e-06, 2.002229e-06, 2.603969e-06, 1.445249e-06, 1.209201e-06, 
    1.034705e-06, 9.593605e-07, 2.629099e-06, 3.162831e-06, 4.183278e-06,
  8.392978e-05, 7.352674e-05, 6.633682e-07, 1.914154e-09, 1.424948e-07, 
    2.922383e-07, 1.106268e-06, 2.263032e-06, 1.472723e-06, 2.092198e-06, 
    2.065788e-06, 2.259633e-06, 2.197526e-06, 2.744532e-06, 4.760414e-06,
  4.861261e-05, 4.583286e-05, 2.962384e-05, 3.135607e-09, 2.672533e-08, 
    4.570957e-08, 9.872834e-08, 3.622687e-07, 2.227658e-06, 1.959814e-06, 
    3.050071e-06, 2.637179e-06, 2.69781e-06, 2.356004e-06, 4.061488e-06,
  1.906901e-05, 3.209869e-05, 2.329787e-05, 1.18974e-05, 4.707796e-10, 
    3.868965e-09, 1.096508e-06, 5.302122e-07, 1.423747e-06, 2.592901e-06, 
    2.303824e-06, 3.988912e-06, 2.568657e-06, 2.01199e-06, 4.300178e-06,
  1.150363e-05, 1.479777e-05, 1.415398e-05, 1.90777e-05, 1.552871e-09, 
    2.047103e-10, 6.6836e-07, 6.246771e-07, 1.909807e-06, 3.417966e-06, 
    2.441797e-06, 4.304786e-06, 3.086896e-06, 3.590315e-06, 2.205462e-06,
  7.297701e-06, 6.227008e-06, 9.95658e-06, 1.35908e-05, 1.688392e-05, 
    2.12058e-09, 2.143474e-07, 1.015755e-06, 1.181599e-06, 2.366402e-06, 
    4.588832e-06, 4.764403e-06, 3.70708e-06, 3.970705e-06, 3.175926e-06,
  5.973694e-06, 3.060639e-06, 4.379454e-06, 1.132064e-05, 2.452721e-05, 
    1.635933e-05, 1.336483e-09, 1.61415e-06, 8.950811e-07, 1.496132e-06, 
    3.542866e-06, 3.65644e-06, 3.809861e-06, 4.200204e-06, 3.651431e-06,
  0.0002742502, 0.0002817186, 0.0002850501, 0.0002932379, 0.0002560768, 
    0.000191492, 0.0001427487, 0.0001123317, 8.401432e-05, 5.966451e-05, 
    2.961244e-05, 5.792607e-06, 5.691105e-06, 9.093851e-06, 9.89316e-06,
  0.0004097987, 0.0003238733, 0.0002562864, 0.0001463986, 5.041358e-05, 
    2.295548e-05, 2.143004e-05, 2.66462e-05, 2.22525e-05, 2.355129e-05, 
    1.509224e-05, 2.296328e-06, 6.063256e-06, 8.014171e-06, 1.030772e-05,
  0.0003674445, 0.0002712502, 0.0001277483, 5.749163e-05, 5.119681e-05, 
    3.150647e-05, 2.455918e-05, 2.334432e-05, 2.936258e-05, 1.69954e-05, 
    4.148352e-06, 2.292598e-06, 7.481426e-06, 7.581578e-06, 9.831017e-06,
  0.0002498321, 0.0001626095, 0.0001002149, 7.859558e-05, 5.671886e-05, 
    2.384411e-05, 1.907684e-05, 1.403521e-05, 1.142826e-05, 3.330862e-06, 
    1.130916e-06, 3.427834e-06, 3.688791e-06, 6.008603e-06, 1.195469e-05,
  0.000105992, 0.0001178519, 0.0001173532, 7.205331e-05, 3.446177e-05, 
    5.424083e-06, 2.015268e-06, 8.467138e-07, 2.072049e-07, 5.035788e-07, 
    2.099411e-06, 5.277289e-06, 7.616004e-06, 5.572767e-06, 1.08928e-05,
  2.996035e-05, 6.084132e-05, 8.42126e-05, 0.0001259093, 1.001424e-05, 
    1.36888e-07, 1.365331e-07, 1.994806e-07, 2.667011e-07, 6.469767e-07, 
    2.799082e-06, 3.922382e-06, 5.40933e-06, 4.805956e-06, 6.685063e-06,
  0.0002329576, 0.0001624196, 0.0002107422, 8.406065e-05, 8.636256e-06, 
    2.709045e-06, 1.50353e-06, 2.617593e-07, 5.360959e-07, 1.034061e-06, 
    1.881453e-06, 2.950723e-06, 2.684629e-06, 5.770367e-06, 9.263244e-06,
  0.0005286231, 0.0004438155, 0.0002588223, 9.427239e-05, 8.676909e-06, 
    5.010626e-06, 1.684461e-06, 9.020746e-07, 1.269743e-06, 1.062061e-06, 
    1.298118e-06, 3.102233e-06, 4.139466e-06, 3.870597e-06, 6.174751e-06,
  0.0006327017, 0.0004703996, 0.0002572717, 9.034057e-05, 5.063668e-05, 
    6.389474e-06, 1.6335e-06, 1.79776e-06, 9.56907e-07, 1.86278e-06, 
    2.397115e-06, 2.371149e-06, 2.685289e-06, 4.97345e-06, 6.172847e-06,
  0.000451602, 0.0003591307, 0.0002221833, 0.0001187109, 4.757595e-05, 
    2.014197e-05, 1.224258e-06, 6.590298e-07, 7.013766e-07, 8.925765e-07, 
    2.522296e-06, 2.582475e-06, 3.164409e-06, 3.497023e-06, 4.42639e-06,
  5.173121e-13, 3.354839e-13, 5.751935e-13, 7.269979e-13, 1.148274e-10, 
    2.741703e-08, 1.384591e-06, 6.303138e-06, 1.338363e-05, 2.730174e-05, 
    6.045819e-05, 9.886125e-05, 0.0001130673, 0.0001337119, 0.0001412799,
  3.657905e-12, 1.370465e-12, 3.54245e-12, 1.12807e-09, 4.797375e-07, 
    3.293362e-06, 1.307828e-05, 3.206735e-05, 5.863243e-05, 0.0001043477, 
    0.0001531476, 0.000207274, 0.0002382402, 0.0002741382, 0.000293307,
  3.948934e-09, 5.195001e-11, 5.083324e-09, 3.539289e-07, 7.305058e-06, 
    4.850358e-05, 9.796697e-05, 0.00015258, 0.0002126965, 0.000277244, 
    0.0003300674, 0.0003356898, 0.0003479767, 0.0003548713, 0.0003687138,
  2.138356e-07, 2.240423e-08, 2.22748e-07, 7.067579e-06, 5.07654e-05, 
    0.0001240043, 0.0001845101, 0.0002194584, 0.0002370486, 0.0002544812, 
    0.0002577358, 0.0002515488, 0.0002554481, 0.000263598, 0.0002521033,
  4.143959e-06, 6.006497e-07, 1.398697e-06, 1.578547e-05, 6.385627e-05, 
    0.0001183504, 0.0001275447, 0.0001257888, 0.0001314991, 0.0001400279, 
    0.0001408655, 0.0001342015, 0.0001308097, 0.0001190827, 0.0001090151,
  5.201277e-06, 6.350912e-06, 9.252229e-06, 2.174009e-05, 4.18255e-05, 
    3.527988e-05, 2.485321e-05, 2.301323e-05, 3.026542e-05, 3.38888e-05, 
    4.516694e-05, 4.874558e-05, 4.717626e-05, 4.105349e-05, 4.646324e-05,
  2.668579e-06, 1.266436e-05, 3.092003e-05, 5.025489e-05, 4.945294e-05, 
    2.324868e-05, 1.371044e-05, 2.816224e-05, 3.626143e-06, 9.305432e-06, 
    2.976493e-05, 3.980314e-05, 4.548977e-05, 4.843199e-05, 4.905386e-05,
  1.451148e-05, 5.566137e-05, 0.0001441863, 0.0001856046, 0.0001356511, 
    0.0001259964, 9.468839e-05, 6.603892e-05, 6.680098e-05, 1.937606e-05, 
    2.417127e-05, 3.253444e-05, 4.514051e-05, 4.666981e-05, 3.793457e-05,
  6.592268e-05, 0.0002201103, 0.0003103819, 0.0003502734, 0.0003179392, 
    0.000223102, 0.0001549852, 0.0001257764, 0.0001198409, 0.0001357586, 
    0.0001151278, 9.379286e-05, 0.0001116256, 7.903903e-05, 1.26831e-05,
  9.549136e-05, 0.000287052, 0.0004263275, 0.0005108345, 0.0004821155, 
    0.000366614, 0.0002361376, 0.0001581627, 0.0001768691, 0.0001811751, 
    0.0001457943, 8.901595e-05, 7.616931e-05, 7.035527e-05, 8.982443e-06,
  2.936943e-07, 1.243646e-06, 6.862076e-07, 7.628011e-07, 2.977777e-07, 
    1.342416e-06, 5.064106e-06, 9.936761e-06, 1.002915e-05, 1.259335e-05, 
    1.308835e-05, 1.065637e-05, 9.574821e-06, 1.453634e-05, 1.079548e-05,
  1.130709e-06, 4.091913e-08, 2.832802e-08, 1.841588e-07, 7.269416e-07, 
    9.522533e-07, 3.270975e-06, 3.748487e-06, 6.329085e-06, 8.649707e-06, 
    9.697013e-06, 1.046146e-05, 1.180596e-05, 1.123984e-05, 8.972734e-06,
  1.024753e-07, 4.407611e-07, 2.365562e-08, 9.456696e-09, 4.8508e-08, 
    5.464417e-07, 1.282155e-06, 2.48755e-06, 2.585814e-06, 3.76551e-06, 
    6.911426e-06, 7.707343e-06, 7.510222e-06, 9.545508e-06, 9.712182e-06,
  5.883792e-09, 4.656489e-08, 9.193948e-08, 5.665428e-08, 8.173836e-07, 
    1.872565e-06, 1.773355e-06, 2.690378e-06, 2.832166e-06, 3.851026e-06, 
    4.230765e-06, 6.321506e-06, 7.920782e-06, 7.302361e-06, 7.129061e-06,
  8.166936e-09, 1.995868e-08, 2.15943e-06, 1.634795e-06, 3.41925e-06, 
    3.395197e-06, 3.033381e-06, 4.889342e-06, 6.764017e-06, 5.157287e-06, 
    4.656316e-06, 6.386438e-06, 4.878923e-06, 4.543844e-06, 4.372435e-06,
  2.049911e-07, 3.778162e-07, 1.742442e-06, 4.617429e-06, 6.164592e-06, 
    4.16526e-06, 2.736648e-06, 3.579902e-06, 3.920098e-06, 3.366362e-06, 
    3.36563e-06, 4.520897e-06, 2.84889e-06, 2.270438e-06, 2.900784e-06,
  2.024238e-06, 2.920805e-07, 1.156717e-06, 4.796041e-06, 5.423709e-06, 
    2.637427e-06, 2.806443e-06, 1.320501e-06, 2.040096e-06, 2.491651e-06, 
    3.822604e-06, 2.799354e-06, 4.153769e-07, 7.97108e-07, 8.215172e-07,
  7.584596e-06, 3.868689e-06, 7.168793e-07, 5.856069e-06, 7.933564e-06, 
    4.210528e-06, 2.734232e-06, 2.179557e-06, 2.424307e-06, 1.370671e-06, 
    1.109736e-06, 1.033943e-06, 2.74878e-06, 5.220401e-06, 1.027929e-05,
  1.154692e-05, 1.519265e-05, 7.905423e-06, 2.999988e-06, 5.633918e-06, 
    3.737033e-06, 9.469304e-06, 6.454714e-06, 1.008153e-05, 1.04513e-05, 
    8.222978e-06, 7.515136e-06, 9.841568e-06, 1.366156e-05, 2.620691e-05,
  7.068134e-06, 1.463815e-05, 2.912857e-05, 3.089003e-05, 2.63019e-05, 
    2.958225e-05, 1.630055e-05, 3.188683e-05, 4.485335e-05, 7.341585e-05, 
    0.0001080686, 9.689209e-05, 0.0001044374, 8.642285e-05, 7.827932e-05,
  8.241964e-06, 8.54759e-07, 9.27664e-07, 9.927235e-06, 1.960947e-05, 
    2.111757e-05, 1.928611e-05, 1.802349e-05, 2.175106e-05, 1.915759e-05, 
    2.114314e-05, 1.605977e-05, 1.746864e-05, 1.551636e-05, 1.412308e-05,
  1.917315e-05, 4.655012e-06, 3.404488e-07, 3.468039e-06, 1.358113e-05, 
    2.078349e-05, 2.17954e-05, 2.065437e-05, 1.558506e-05, 1.398293e-05, 
    1.299214e-05, 1.376094e-05, 1.191275e-05, 1.839517e-05, 1.162347e-05,
  1.199313e-05, 1.057735e-05, 1.525458e-06, 3.12651e-06, 1.110084e-05, 
    1.889997e-05, 2.2494e-05, 2.029973e-05, 1.380188e-05, 1.075761e-05, 
    1.027086e-05, 9.34574e-06, 8.136651e-06, 9.296459e-06, 1.019718e-05,
  2.77178e-06, 3.644631e-06, 2.338575e-07, 2.352108e-06, 8.624176e-06, 
    1.523351e-05, 1.892033e-05, 1.882702e-05, 1.378622e-05, 1.252884e-05, 
    9.360021e-06, 7.45836e-06, 8.059295e-06, 8.89627e-06, 9.530371e-06,
  2.132487e-06, 2.112971e-06, 2.94704e-06, 3.230398e-06, 6.020558e-06, 
    1.086158e-05, 1.221209e-05, 1.363603e-05, 1.296579e-05, 1.048143e-05, 
    8.777912e-06, 8.542004e-06, 8.236789e-06, 7.095849e-06, 5.94892e-06,
  2.2234e-07, 2.587316e-06, 3.293075e-06, 4.216658e-06, 5.345727e-06, 
    8.04222e-06, 1.044831e-05, 1.080298e-05, 1.146575e-05, 1.09627e-05, 
    1.069514e-05, 9.534499e-06, 8.010532e-06, 7.272968e-06, 7.348459e-06,
  1.382397e-07, 1.054755e-06, 6.586703e-06, 4.668907e-06, 4.302562e-06, 
    8.05055e-06, 1.041308e-05, 9.738867e-06, 1.093199e-05, 9.642105e-06, 
    9.283688e-06, 9.028587e-06, 8.03972e-06, 7.745748e-06, 6.64035e-06,
  2.668672e-07, 4.920539e-07, 3.314588e-06, 4.958535e-06, 6.370773e-06, 
    6.576688e-06, 1.093099e-05, 1.036195e-05, 9.771337e-06, 7.386857e-06, 
    8.574702e-06, 8.426283e-06, 7.428909e-06, 6.441283e-06, 5.539395e-06,
  2.286726e-07, 1.015733e-06, 1.233541e-06, 3.219117e-06, 1.035268e-05, 
    7.787174e-06, 8.878091e-06, 1.378275e-05, 9.683816e-06, 7.577781e-06, 
    7.029294e-06, 6.610122e-06, 6.313136e-06, 6.369862e-06, 6.883887e-06,
  6.973031e-08, 2.953159e-07, 1.53838e-06, 3.933587e-06, 5.928885e-06, 
    1.153142e-05, 9.171666e-06, 1.266321e-05, 1.064774e-05, 6.742396e-06, 
    5.85727e-06, 5.190127e-06, 6.071849e-06, 6.450444e-06, 7.721042e-06,
  3.084182e-07, 1.65318e-06, 1.248615e-06, 3.035955e-06, 4.069297e-06, 
    5.889552e-06, 9.968385e-06, 1.54017e-05, 2.551062e-05, 3.24111e-05, 
    2.744532e-05, 4.261797e-05, 5.116962e-05, 7.121728e-05, 6.876772e-05,
  8.301815e-07, 6.39209e-07, 1.436641e-06, 4.607495e-06, 5.11856e-06, 
    5.435656e-06, 7.690759e-06, 1.253654e-05, 1.887588e-05, 2.634842e-05, 
    3.278935e-05, 3.33616e-05, 5.732126e-05, 6.467181e-05, 5.758929e-05,
  2.879947e-07, 1.150512e-06, 1.579146e-06, 5.256548e-06, 9.73746e-06, 
    8.209527e-06, 5.985172e-06, 8.57892e-06, 1.283271e-05, 2.086863e-05, 
    2.697053e-05, 2.855297e-05, 4.035142e-05, 4.901251e-05, 4.982082e-05,
  1.894876e-07, 6.230877e-07, 2.749378e-06, 4.803266e-06, 1.118003e-05, 
    1.242882e-05, 9.031195e-06, 8.117677e-06, 9.380718e-06, 1.602021e-05, 
    2.524266e-05, 3.10311e-05, 3.318471e-05, 3.669604e-05, 3.982942e-05,
  1.1201e-06, 9.239521e-07, 3.113903e-07, 5.3313e-06, 1.161327e-05, 
    1.529521e-05, 1.356658e-05, 9.536537e-06, 7.058065e-06, 9.182268e-06, 
    1.497298e-05, 2.14747e-05, 4.621077e-05, 5.20781e-05, 3.906123e-05,
  2.727741e-06, 8.7042e-07, 8.966064e-07, 1.673067e-06, 1.079831e-05, 
    1.59471e-05, 1.703842e-05, 1.309012e-05, 9.914262e-06, 7.716544e-06, 
    9.69e-06, 1.573346e-05, 2.0714e-05, 4.100734e-05, 5.413292e-05,
  2.120215e-06, 1.848032e-06, 6.225071e-07, 1.56189e-06, 7.103934e-06, 
    1.54568e-05, 1.934658e-05, 1.673851e-05, 1.420038e-05, 1.031592e-05, 
    9.393771e-06, 9.772828e-06, 1.351072e-05, 2.246192e-05, 3.53271e-05,
  8.883501e-08, 1.07415e-06, 4.565233e-07, 1.158301e-06, 3.286707e-06, 
    1.117067e-05, 1.968074e-05, 2.118985e-05, 1.854609e-05, 1.374741e-05, 
    1.143534e-05, 1.202416e-05, 1.425395e-05, 1.576184e-05, 1.992362e-05,
  4.337365e-11, 1.000544e-07, 4.579739e-07, 3.554129e-07, 2.47523e-06, 
    3.814233e-06, 1.579207e-05, 2.012632e-05, 1.767113e-05, 2.03842e-05, 
    1.447857e-05, 1.313218e-05, 1.568538e-05, 1.546671e-05, 1.80404e-05,
  2.363384e-15, 2.694906e-12, 7.082409e-08, 1.450625e-07, 8.169904e-07, 
    4.171881e-06, 5.757729e-06, 1.879106e-05, 1.867172e-05, 1.863255e-05, 
    2.142998e-05, 1.95334e-05, 1.658785e-05, 2.232775e-05, 1.677895e-05,
  3.642736e-09, 9.045133e-09, 3.753086e-09, 1.965828e-07, 1.078644e-06, 
    1.652455e-06, 2.228407e-06, 2.675584e-06, 4.784356e-06, 1.033413e-05, 
    1.699909e-05, 2.614568e-05, 5.045116e-05, 4.649447e-05, 3.465313e-05,
  1.488776e-07, 7.14189e-09, 6.191069e-09, 1.623193e-07, 3.484575e-06, 
    3.464399e-06, 3.575606e-06, 3.296902e-06, 4.009308e-06, 5.538792e-06, 
    8.74098e-06, 1.511765e-05, 3.546411e-05, 4.195965e-05, 4.525938e-05,
  1.777078e-07, 3.000057e-07, 5.741425e-08, 2.202317e-08, 4.030217e-06, 
    2.980485e-06, 4.089345e-06, 4.870962e-06, 2.862527e-06, 3.840428e-06, 
    5.827489e-06, 8.373992e-06, 2.176481e-05, 4.00651e-05, 5.014201e-05,
  1.24794e-07, 2.870385e-07, 2.562309e-07, 2.358025e-08, 1.710991e-06, 
    3.356603e-06, 6.04375e-06, 4.784498e-06, 4.538058e-06, 3.252337e-06, 
    4.44174e-06, 6.675857e-06, 1.41123e-05, 3.035219e-05, 5.293306e-05,
  5.789367e-08, 8.484329e-08, 4.668512e-08, 3.275939e-07, 1.194655e-06, 
    2.437649e-06, 5.021349e-06, 4.47054e-06, 4.261332e-06, 4.10686e-06, 
    3.293458e-06, 5.583874e-06, 8.542125e-06, 1.776898e-05, 4.258087e-05,
  4.856243e-09, 1.27618e-07, 2.442721e-07, 1.016982e-07, 1.808524e-06, 
    1.63769e-06, 3.083719e-06, 4.379465e-06, 4.934276e-06, 3.818826e-06, 
    3.127618e-06, 4.107837e-06, 7.49753e-06, 9.607857e-06, 2.275042e-05,
  5.239588e-09, 6.035074e-08, 5.457443e-07, 7.598223e-07, 4.373087e-07, 
    4.385436e-07, 1.941969e-06, 3.482778e-06, 4.473412e-06, 3.78938e-06, 
    3.732078e-06, 2.855763e-06, 5.476691e-06, 7.111538e-06, 1.215381e-05,
  1.367745e-10, 3.564127e-09, 1.788706e-07, 1.276503e-06, 5.149737e-07, 
    3.988135e-07, 6.909845e-07, 2.437413e-06, 3.04199e-06, 3.69501e-06, 
    4.313958e-06, 2.842336e-06, 3.54569e-06, 3.802579e-06, 6.603874e-06,
  2.691826e-08, 9.039985e-08, 6.37526e-09, 2.825741e-07, 1.344639e-06, 
    8.656072e-07, 3.045528e-07, 8.537146e-07, 1.873315e-06, 3.437579e-06, 
    4.283383e-06, 4.652992e-06, 3.842984e-06, 3.099457e-06, 3.306886e-06,
  5.807295e-07, 8.976388e-07, 4.275233e-07, 5.487969e-09, 5.725355e-09, 
    7.709911e-07, 1.612e-06, 4.516926e-07, 7.491997e-07, 1.276983e-06, 
    3.35754e-06, 4.199158e-06, 3.868666e-06, 3.068139e-06, 3.350733e-06,
  4.736588e-08, 3.339232e-08, 7.591839e-07, 1.600102e-06, 5.351702e-06, 
    6.288804e-06, 2.190284e-07, 1.019953e-06, 2.98515e-06, 1.566616e-05, 
    2.182337e-05, 1.243605e-05, 3.044685e-06, 2.909629e-07, 1.814793e-06,
  1.529789e-07, 5.74339e-08, 1.420411e-07, 6.880987e-07, 5.421602e-06, 
    5.493952e-06, 1.952233e-07, 8.943603e-08, 2.333832e-06, 7.268803e-06, 
    2.473457e-05, 2.115475e-05, 6.114132e-06, 1.989956e-06, 2.075219e-06,
  2.795765e-07, 2.01444e-07, 1.076941e-07, 9.4124e-07, 5.189351e-06, 
    6.718624e-06, 1.768932e-06, 1.925682e-07, 4.402085e-07, 2.675512e-06, 
    1.24863e-05, 1.978376e-05, 1.077676e-05, 4.385014e-06, 2.903473e-05,
  4.206041e-07, 1.750948e-07, 8.185292e-08, 2.193679e-07, 4.56024e-06, 
    1.643589e-06, 1.46531e-06, 3.921601e-07, 1.512697e-07, 1.333678e-07, 
    6.357016e-06, 1.468231e-05, 1.83136e-05, 1.660558e-05, 4.031731e-06,
  3.973131e-07, 1.805656e-07, 3.126717e-08, 4.775491e-08, 7.837381e-07, 
    2.335628e-06, 3.26482e-06, 3.365289e-07, 3.744734e-07, 7.846622e-07, 
    4.454989e-06, 1.027373e-05, 2.441036e-05, 1.942958e-05, 1.134234e-05,
  1.474494e-07, 2.699159e-07, 2.468621e-08, 3.749422e-08, 5.433747e-07, 
    3.156487e-06, 1.226646e-06, 4.817996e-07, 8.57903e-07, 4.244725e-07, 
    1.771548e-07, 5.812621e-06, 1.472107e-05, 2.100304e-05, 1.54869e-05,
  3.305724e-07, 2.471752e-07, 3.150983e-07, 5.180132e-08, 1.663524e-07, 
    1.420313e-06, 3.198012e-06, 2.222363e-06, 7.387516e-07, 7.953359e-07, 
    1.124883e-06, 2.85554e-06, 1.060407e-05, 2.270921e-05, 1.911305e-05,
  1.601494e-07, 1.726287e-07, 1.970375e-07, 1.808624e-07, 3.890891e-08, 
    8.833666e-07, 2.254766e-06, 2.508692e-06, 1.837776e-06, 3.726294e-07, 
    6.736532e-07, 7.123014e-07, 3.537133e-06, 1.431138e-05, 2.216523e-05,
  4.147504e-07, 1.837546e-07, 4.124176e-08, 6.884004e-08, 1.570676e-07, 
    5.754786e-07, 2.427246e-06, 2.756183e-06, 1.71555e-06, 7.138479e-07, 
    4.19308e-07, 6.796276e-07, 1.706829e-06, 8.188294e-06, 1.43277e-05,
  2.218871e-07, 2.111061e-07, 1.188845e-07, 1.104558e-08, 4.114181e-09, 
    5.888171e-09, 1.583078e-06, 1.793136e-06, 2.886252e-06, 1.180514e-06, 
    7.060249e-07, 6.237208e-07, 1.543104e-06, 2.048317e-06, 8.582913e-06,
  3.679109e-05, 8.875751e-06, 3.631096e-07, 1.16984e-07, 7.20142e-06, 
    2.281915e-05, 3.527052e-05, 1.928497e-05, 4.926149e-06, 9.573257e-06, 
    2.041068e-05, 1.788957e-05, 1.166029e-06, 1.903566e-07, 7.05153e-07,
  5.57731e-06, 4.590189e-09, 2.707526e-09, 2.646447e-08, 5.681279e-06, 
    1.351546e-05, 2.756564e-05, 1.656899e-05, 6.846192e-07, 4.027954e-06, 
    1.656927e-05, 3.156157e-05, 5.235263e-06, 4.226387e-08, 9.000065e-09,
  5.660137e-07, 9.753539e-09, 1.955338e-09, 5.861655e-08, 8.181883e-06, 
    1.432598e-05, 2.491116e-05, 1.838319e-05, 1.535374e-06, 2.371993e-06, 
    9.995959e-06, 2.746438e-05, 7.451471e-06, 8.83664e-08, 3.72403e-09,
  3.882679e-07, 3.650394e-07, 2.485677e-09, 2.386012e-07, 9.186109e-06, 
    8.622578e-06, 1.800173e-05, 2.038097e-05, 5.94784e-06, 9.467295e-07, 
    5.855108e-06, 2.298279e-05, 1.53866e-05, 4.60376e-07, 1.988096e-09,
  4.503992e-07, 1.316789e-07, 8.032014e-10, 7.190699e-08, 4.07673e-06, 
    7.423253e-06, 1.41359e-05, 1.939421e-05, 8.582331e-06, 8.277338e-07, 
    3.598859e-06, 1.873575e-05, 2.950676e-05, 1.330901e-06, 1.839733e-09,
  5.07181e-07, 3.978957e-07, 2.018049e-07, 6.901473e-09, 1.027991e-06, 
    4.225434e-06, 8.211739e-06, 1.375253e-05, 1.145719e-05, 2.93074e-06, 
    1.760835e-06, 7.534406e-06, 2.718634e-05, 5.208958e-06, 1.826042e-08,
  8.95929e-07, 1.245778e-06, 5.919625e-07, 1.376933e-07, 2.996514e-07, 
    1.145039e-06, 7.286799e-06, 1.274271e-05, 9.963491e-06, 3.987796e-06, 
    1.761518e-07, 3.512576e-06, 2.181891e-05, 2.020132e-05, 2.809624e-10,
  1.227026e-06, 1.229483e-06, 4.925428e-07, 3.478862e-07, 1.075273e-09, 
    2.587707e-07, 6.300277e-06, 1.042838e-05, 9.504096e-06, 6.290014e-06, 
    5.427704e-07, 1.276556e-06, 1.059255e-05, 2.537402e-05, 4.341574e-06,
  1.858811e-06, 9.569344e-07, 2.969655e-07, 1.237488e-07, 4.510969e-08, 
    1.458863e-08, 4.876974e-06, 8.071649e-06, 8.063492e-06, 5.56944e-06, 
    6.524691e-07, 1.903197e-07, 4.542787e-06, 1.658324e-05, 1.208056e-05,
  1.423851e-06, 8.220873e-07, 4.442022e-07, 5.95415e-08, 1.90325e-10, 
    3.389721e-09, 2.143991e-06, 8.534279e-06, 5.738672e-06, 4.13717e-06, 
    1.286801e-06, 1.055718e-08, 5.984301e-07, 6.464064e-06, 1.280573e-05,
  0.0001175348, 0.0001834469, 0.000239265, 0.0002493258, 0.0002248004, 
    0.000218102, 0.0001728491, 0.0002099642, 0.0002710887, 0.0003055545, 
    0.0002356097, 0.0002428536, 0.0001709187, 0.0002093773, 7.362204e-05,
  0.0001221192, 0.0001564145, 0.0001549096, 0.0001695871, 0.0002003913, 
    0.0001607402, 0.0001764927, 0.0001726213, 0.0001872466, 0.0002159193, 
    0.0002572017, 0.000274634, 0.0002581298, 0.0002778413, 8.254854e-05,
  7.989485e-05, 8.128184e-05, 9.034265e-05, 0.0001110769, 0.0001915711, 
    0.0001503164, 0.0001685384, 0.0001468904, 0.0001412158, 0.000149321, 
    0.0001128138, 0.000199621, 0.0001880992, 0.0001739012, 7.089583e-05,
  2.166057e-05, 1.688248e-05, 3.795082e-05, 4.957603e-05, 0.0001047668, 
    9.728084e-05, 0.0001335108, 0.0001127645, 0.0001254841, 0.000121068, 
    0.0001218071, 9.279473e-05, 0.0001898192, 0.0001246495, 6.141709e-05,
  1.416751e-05, 1.688368e-05, 2.216896e-05, 2.541773e-05, 6.308931e-05, 
    6.041662e-05, 6.69943e-05, 0.0001212499, 0.0001178976, 0.0001370965, 
    0.0001250952, 0.0001699272, 0.0001071493, 0.0001095274, 6.447045e-05,
  1.471582e-05, 1.787505e-05, 1.648645e-05, 1.285358e-05, 4.301254e-05, 
    5.553048e-05, 8.406665e-05, 0.0001037066, 0.0001272207, 0.0001656504, 
    0.0001966852, 0.0002168224, 9.227692e-05, 7.341077e-05, 6.118129e-05,
  8.998641e-06, 3.561685e-05, 4.813679e-05, 4.191466e-05, 2.140705e-05, 
    4.359083e-05, 6.448843e-05, 0.0001058211, 9.416844e-05, 0.0001443625, 
    0.0001026159, 0.0001188717, 8.671448e-05, 7.931113e-05, 4.708523e-05,
  1.723972e-05, 2.588902e-05, 2.781892e-05, 3.224939e-05, 3.43608e-05, 
    8.155014e-05, 7.58541e-05, 5.767677e-05, 5.404208e-05, 3.146568e-05, 
    4.853537e-05, 5.016144e-05, 6.876739e-05, 5.77082e-05, 4.08852e-05,
  2.963619e-05, 2.694548e-05, 1.335493e-05, 1.135356e-05, 1.975603e-05, 
    3.200491e-05, 3.853827e-05, 4.14673e-05, 1.96615e-05, 2.120027e-05, 
    1.868743e-05, 3.176162e-05, 3.480751e-05, 3.586967e-05, 3.746e-05,
  1.385828e-05, 1.45293e-05, 1.056957e-05, 8.416459e-06, 4.975886e-06, 
    4.837183e-06, 2.102922e-07, 7.273453e-06, 1.592549e-05, 1.788355e-05, 
    1.855414e-05, 1.38619e-05, 1.876965e-05, 2.186517e-05, 3.188883e-05,
  1.657342e-05, 3.061951e-05, 1.834999e-05, 3.939237e-05, 3.678708e-05, 
    2.987538e-05, 5.675096e-05, 7.72342e-05, 0.0001552473, 0.0002173136, 
    0.0001915387, 0.0001152356, 8.607864e-05, 5.405576e-05, 0.0001324689,
  2.264268e-06, 5.988689e-06, 2.860823e-05, 5.539045e-05, 4.516073e-05, 
    3.828447e-05, 5.049972e-05, 4.165914e-05, 4.870239e-05, 7.016997e-05, 
    0.0001106287, 0.0001171067, 0.000121545, 8.741851e-05, 0.0001245672,
  8.239181e-07, 8.498979e-07, 1.311713e-05, 3.960207e-05, 5.336387e-05, 
    5.580124e-05, 3.88273e-05, 3.114603e-05, 3.012474e-05, 2.918376e-05, 
    3.055645e-05, 3.774567e-05, 7.903085e-05, 8.52254e-05, 0.0001459584,
  5.268e-07, 5.996507e-07, 2.146158e-06, 2.064467e-05, 3.631414e-05, 
    4.220313e-05, 3.308422e-05, 2.640776e-05, 2.763292e-05, 2.805499e-05, 
    1.773579e-05, 1.851954e-05, 2.575738e-05, 0.0001297511, 0.0002338178,
  3.274975e-07, 3.86952e-07, 1.074777e-07, 5.931233e-06, 1.706983e-05, 
    2.551218e-05, 2.249982e-05, 2.066175e-05, 1.803509e-05, 2.092957e-05, 
    2.547572e-05, 1.477381e-05, 7.640717e-05, 0.0001942376, 0.0002328837,
  5.594535e-11, 7.920607e-11, 2.631382e-09, 2.302912e-08, 4.522542e-06, 
    1.070616e-05, 1.223292e-05, 1.214455e-05, 1.31372e-05, 1.213906e-05, 
    2.370073e-05, 5.740835e-05, 0.0001830813, 0.0001950187, 0.0002887436,
  2.941801e-24, 1.073057e-18, 2.075494e-14, 9.169299e-12, 2.148543e-10, 
    1.042608e-06, 7.424529e-06, 1.061438e-05, 2.475297e-05, 4.236789e-05, 
    9.285455e-05, 0.0001997877, 0.0003221059, 0.0002603504, 0.0003660402,
  4.573976e-12, 1.751995e-13, 5.475721e-16, 4.768212e-09, 1.349569e-11, 
    1.572283e-06, 2.294148e-05, 3.773242e-05, 8.172719e-05, 0.000118343, 
    0.0002139395, 0.0002001273, 0.0002355185, 0.0003185888, 0.0003731356,
  2.268213e-08, 2.338945e-07, 3.807089e-07, 2.376126e-06, 5.782511e-06, 
    2.040807e-05, 3.318112e-05, 6.849451e-05, 0.0001288781, 0.0001558022, 
    0.0001190734, 0.000171835, 0.0002464189, 0.0002326044, 0.000319476,
  1.397321e-06, 5.228627e-06, 7.480073e-06, 1.60383e-05, 1.099392e-05, 
    4.666216e-06, 2.681727e-05, 5.025756e-05, 4.820412e-05, 0.0001241823, 
    0.000158393, 0.0002020738, 0.0001934774, 0.0001702736, 0.0002019425,
  0.000274716, 0.0002427627, 0.0002435248, 0.0002349844, 0.0001357288, 
    4.417905e-05, 2.545663e-05, 1.4543e-05, 2.835853e-05, 3.150467e-05, 
    1.706233e-05, 7.369695e-06, 9.276469e-06, 1.030883e-05, 1.440762e-05,
  0.0003799445, 0.0004000826, 0.0004923826, 0.0004942964, 0.0003786027, 
    0.0001919437, 6.052949e-05, 9.184084e-06, 9.255439e-06, 1.156092e-05, 
    2.405704e-05, 2.020634e-05, 2.427183e-05, 3.460955e-05, 4.731932e-05,
  0.0003892358, 0.0005197804, 0.0006029956, 0.0006249125, 0.0005572964, 
    0.0004352949, 0.0003487761, 0.0001724618, 1.222915e-05, 6.373746e-06, 
    5.108398e-06, 1.498746e-05, 2.231389e-05, 5.402364e-05, 5.166998e-05,
  0.0003869972, 0.0005334595, 0.0006416752, 0.0005734863, 0.0004436671, 
    0.0003606172, 0.0003011415, 0.0002047323, 7.435945e-05, 2.130384e-06, 
    3.681788e-06, 3.972017e-06, 1.038768e-05, 2.854607e-05, 3.9363e-05,
  0.0003735496, 0.0005122285, 0.0005316788, 0.0003679938, 0.0002628174, 
    0.000406799, 0.0004620241, 0.0002632319, 2.578518e-05, 5.517204e-06, 
    4.061302e-06, 4.488495e-06, 5.831823e-06, 5.570468e-06, 1.102004e-05,
  0.0003574473, 0.0003796528, 0.000256514, 0.0001150815, 0.0001130769, 
    0.0001970676, 0.0002858846, 0.0001387033, 3.410574e-05, 5.563633e-06, 
    3.795456e-06, 2.665825e-06, 2.810334e-06, 3.706567e-06, 3.616821e-06,
  0.0002200164, 0.0001826326, 0.0001113176, 0.0001293192, 0.0001084693, 
    0.0001501463, 0.0001250003, 7.225758e-05, 3.824438e-05, 2.564877e-05, 
    1.297272e-06, 2.425689e-06, 2.18051e-06, 3.065567e-06, 3.357284e-06,
  0.0001113291, 0.000114857, 0.0001868255, 0.0002121205, 0.0001563355, 
    0.0001446238, 6.921049e-05, 0.0001222877, 4.339761e-05, 3.114706e-05, 
    1.933693e-05, 2.836922e-06, 1.836031e-06, 2.619361e-06, 3.902364e-06,
  0.0002052777, 0.0002207023, 0.0002047133, 0.0002011315, 0.0002532681, 
    0.0001682333, 7.675758e-05, 7.052018e-06, 2.77897e-06, 1.682508e-05, 
    4.469904e-06, 3.286814e-06, 2.656523e-06, 2.372943e-06, 2.938202e-06,
  0.0002501621, 0.0003303512, 0.0003030834, 0.0003755081, 0.0003525422, 
    0.0002208707, 7.21175e-05, 3.828584e-06, 1.11366e-06, 4.689376e-07, 
    9.416138e-06, 4.292439e-06, 2.247056e-06, 1.617552e-06, 1.352257e-06,
  0.001082655, 0.001032621, 0.0008594766, 0.000749319, 0.0005221789, 
    0.0004215491, 0.0004157215, 0.0003156935, 0.0001708341, 7.448552e-05, 
    3.450625e-05, 7.091401e-06, 2.31707e-06, 2.864135e-06, 1.30523e-06,
  0.0008575927, 0.0007233248, 0.0005318873, 0.0005771238, 0.0005439061, 
    0.0005652663, 0.0007142414, 0.0008260411, 0.0005798707, 0.0002408373, 
    8.197067e-05, 4.06588e-05, 2.040804e-05, 4.73193e-06, 1.007487e-06,
  0.0005287395, 0.0003485497, 0.0001580801, 0.0001132054, 0.0002403166, 
    0.0003459104, 0.0007139541, 0.001172701, 0.001113118, 0.0005828026, 
    0.0001901933, 6.548239e-05, 3.627112e-05, 1.313096e-05, 5.828231e-06,
  0.000348014, 0.0002305058, 0.0001220284, 2.270457e-05, 1.473523e-05, 
    0.0001058735, 0.0005013609, 0.0007599054, 0.0009666905, 0.0008710348, 
    0.0004560211, 0.0002359114, 0.0001361632, 8.361954e-05, 5.057496e-05,
  0.0002498711, 0.0001074415, 6.456252e-05, 4.270509e-05, 1.464694e-05, 
    4.746795e-05, 0.000264345, 0.0004786608, 0.0008111558, 0.0007741643, 
    0.000596009, 0.0004226769, 0.0003057402, 0.0001937083, 0.0001152998,
  0.0002688594, 0.0001096431, 3.853759e-05, 3.27236e-05, 4.245855e-05, 
    7.460045e-05, 0.0001740677, 0.0004094253, 0.0003782035, 0.0003600239, 
    0.0004894665, 0.0005094332, 0.0003864171, 0.0002780056, 0.0001670234,
  0.0003105694, 0.0001887777, 8.007792e-05, 6.08041e-05, 8.227407e-05, 
    0.00010674, 0.0001696008, 0.0001848043, 0.0002825647, 0.0002284877, 
    0.0004081272, 0.0005556575, 0.0004981011, 0.0003209104, 0.0001771796,
  0.0003049031, 0.0002547087, 0.0001424314, 9.291812e-05, 7.529504e-05, 
    0.0001603496, 0.000180431, 0.0001870707, 0.0001799454, 0.0001877909, 
    0.0003457757, 0.0005368321, 0.00048995, 0.0003507849, 0.0001806459,
  0.0002833956, 0.0002155705, 0.0001198169, 9.235147e-05, 0.0001051305, 
    0.0001803097, 0.0002271595, 0.0002603703, 0.0001817692, 0.0002103535, 
    0.0003704752, 0.0005058128, 0.0004811661, 0.0003568237, 0.0001915285,
  0.0001465361, 0.0001526755, 0.0001007, 5.183049e-05, 8.797477e-05, 
    0.0001869148, 0.0002675042, 0.0002481323, 0.0002317886, 0.0003505494, 
    0.000476651, 0.0004880552, 0.0004089726, 0.0003602059, 0.0002383944,
  0.0001631722, 0.0001821804, 0.0002077503, 0.0002749269, 0.0003124181, 
    0.0003224613, 0.0003243135, 0.0003185988, 0.0003038297, 0.0002930393, 
    0.0003092717, 0.000361728, 0.0003483632, 0.0002732633, 0.000191158,
  0.000206825, 0.0002177096, 0.0002123624, 0.000243473, 0.0002476945, 
    0.0002654431, 0.0002488303, 0.0002348835, 0.0003006353, 0.0003899689, 
    0.0004914908, 0.0005029695, 0.000406939, 0.0003286027, 0.0002585081,
  0.0001642467, 0.0001565418, 0.0001559308, 0.0001606623, 0.0001173236, 
    4.934323e-05, 2.620822e-05, 4.130189e-05, 7.754584e-05, 9.238142e-05, 
    0.0001269108, 0.0002048552, 0.0003071044, 0.0003429673, 0.0003347642,
  0.0001066362, 7.65046e-05, 0.000122034, 0.000103654, 2.104286e-05, 
    1.492586e-05, 2.516006e-05, 1.414082e-05, 4.966691e-06, 1.100448e-05, 
    2.782021e-05, 5.753325e-05, 0.0001737333, 0.000290182, 0.0003026418,
  5.440546e-05, 4.948207e-05, 9.033662e-05, 5.897645e-05, 3.173415e-05, 
    3.479473e-05, 1.211571e-05, 5.239887e-07, 8.615484e-07, 7.363944e-07, 
    1.041889e-06, 5.681586e-06, 6.285425e-05, 0.00020596, 0.0003035348,
  3.505131e-05, 4.889938e-05, 6.486307e-05, 3.977148e-05, 5.921314e-05, 
    3.709723e-05, 7.077245e-06, 3.665373e-06, 3.360102e-06, 2.955135e-06, 
    2.651261e-06, 3.74661e-06, 1.650651e-05, 0.0001387128, 0.0003112645,
  2.955439e-05, 4.394948e-05, 5.54551e-05, 4.745817e-05, 0.0001257009, 
    0.0001137461, 4.22898e-05, 2.003496e-05, 1.593691e-05, 9.574069e-06, 
    5.48395e-06, 6.79526e-06, 7.463874e-06, 0.0001030824, 0.0003121265,
  4.818426e-05, 5.154456e-05, 3.301074e-05, 4.449336e-05, 0.0001197887, 
    0.0001522569, 0.0001113265, 4.957542e-05, 3.039903e-05, 1.924389e-05, 
    1.46261e-05, 1.222126e-05, 1.016866e-05, 7.769018e-05, 0.0002717578,
  0.0001063417, 8.647795e-05, 5.97625e-05, 5.437749e-05, 7.74088e-05, 
    0.0001663975, 0.0001341053, 0.0001055626, 4.284437e-05, 4.736408e-05, 
    3.747086e-05, 3.269989e-05, 2.21899e-05, 5.560524e-05, 0.0001857481,
  9.866057e-05, 0.0001266495, 0.0001231925, 0.0001081392, 5.936715e-05, 
    3.416667e-05, 0.0001730346, 0.0001213237, 0.0001077424, 0.0001017714, 
    5.911156e-05, 4.262732e-05, 2.812152e-05, 4.080478e-05, 0.0001176022,
  1.484246e-10, 6.546504e-10, 8.732621e-10, 1.47525e-09, 2.918002e-09, 
    5.263628e-10, 5.619821e-10, 6.096442e-10, 3.021604e-07, 5.939902e-07, 
    4.002758e-06, 3.116972e-06, 2.532909e-06, 1.258631e-06, 8.364557e-07,
  5.484387e-11, 5.019767e-11, 2.92132e-10, 3.805188e-10, 1.994057e-10, 
    6.388603e-10, 5.887208e-11, 2.185262e-10, 6.538089e-08, 5.482023e-07, 
    1.032968e-06, 1.780371e-06, 2.416807e-06, 1.978464e-06, 1.514085e-06,
  1.484064e-11, 2.496927e-11, 2.9498e-11, 1.300669e-10, 6.337685e-11, 
    6.820318e-11, 9.653366e-10, 8.999059e-09, 9.422274e-09, 4.481037e-08, 
    1.83108e-06, 2.000261e-06, 2.81972e-06, 1.759946e-06, 1.064521e-06,
  5.763436e-11, 1.608046e-11, 2.625889e-11, 4.680531e-11, 1.004546e-10, 
    4.031961e-10, 4.375903e-08, 1.129759e-06, 1.246209e-06, 9.237449e-07, 
    1.319719e-06, 2.257078e-06, 1.146249e-06, 3.913693e-06, 6.682254e-06,
  8.855824e-12, 2.271552e-11, 3.967922e-11, 3.763463e-11, 4.18983e-11, 
    6.327654e-07, 3.585748e-06, 3.394851e-06, 1.814975e-06, 1.648613e-06, 
    2.690109e-06, 3.693315e-06, 3.844789e-06, 3.71038e-06, 7.52927e-06,
  2.08223e-25, 1.216686e-11, 1.808912e-11, 1.350402e-11, 2.721582e-08, 
    3.814937e-06, 9.052681e-06, 1.801609e-06, 2.022733e-06, 4.484458e-06, 
    5.577717e-06, 6.390505e-06, 6.048367e-06, 4.395606e-06, 4.749552e-06,
  5.269467e-26, 8.59141e-12, 3.752525e-10, 4.931464e-09, 1.393513e-06, 
    1.109519e-05, 1.54238e-05, 4.339361e-06, 6.128522e-06, 7.883228e-06, 
    6.023904e-06, 6.752205e-06, 6.001809e-06, 5.120332e-06, 6.389515e-06,
  1.919358e-26, 1.326991e-09, 1.844871e-08, 4.955095e-08, 1.953078e-06, 
    1.423431e-05, 3.370578e-05, 1.524532e-05, 1.115158e-05, 5.613475e-06, 
    5.496111e-06, 6.19111e-06, 7.055611e-06, 7.291591e-06, 7.034636e-06,
  9.875537e-10, 1.52752e-08, 1.139608e-07, 6.175073e-07, 2.087097e-06, 
    8.05735e-06, 1.166879e-05, 4.285927e-05, 1.716208e-05, 7.555182e-06, 
    1.473841e-05, 1.527938e-05, 2.263033e-05, 2.149467e-05, 1.59525e-05,
  1.346531e-09, 5.44901e-08, 6.910029e-07, 1.974797e-06, 3.591924e-07, 
    7.189074e-07, 1.576662e-05, 3.579363e-05, 5.496744e-05, 2.162361e-05, 
    2.152635e-05, 3.431498e-05, 4.206268e-05, 2.613715e-05, 1.893006e-05,
  7.304925e-15, 3.806518e-11, 6.793239e-11, 6.42714e-10, 2.488516e-09, 
    4.786939e-08, 3.305575e-08, 2.994868e-08, 8.411343e-07, 1.588596e-06, 
    1.934096e-06, 3.578999e-06, 2.192132e-06, 5.947868e-06, 5.197985e-06,
  3.593889e-15, 1.17122e-11, 1.115904e-21, 5.956316e-15, 4.01339e-11, 
    5.613748e-10, 1.298611e-09, 1.667606e-09, 1.992976e-09, 2.861569e-08, 
    1.503849e-07, 7.117141e-07, 1.858518e-06, 1.819104e-06, 4.78126e-06,
  4.06728e-12, 5.79274e-12, 7.387593e-22, 4.466925e-22, 6.837684e-16, 
    1.7155e-10, 8.129832e-11, 4.801188e-10, 6.649634e-10, 1.993006e-08, 
    1.865457e-07, 6.365085e-07, 9.82571e-07, 1.855091e-06, 2.563836e-06,
  1.502878e-11, 6.869473e-15, 7.22909e-22, 6.046716e-22, 6.786722e-22, 
    6.150724e-22, 5.11884e-22, 3.617439e-11, 3.861205e-12, 1.430645e-08, 
    4.762674e-08, 4.126344e-07, 2.05799e-06, 3.182096e-06, 2.810702e-06,
  1.118992e-10, 7.216293e-14, 5.666961e-15, 4.29739e-22, 3.422352e-22, 
    4.037609e-22, 3.010287e-22, 4.365208e-22, 2.418658e-12, 3.00004e-11, 
    2.376342e-09, 7.937211e-07, 1.595151e-06, 2.351497e-06, 5.891264e-06,
  1.667907e-12, 3.295222e-19, 8.794289e-18, 5.45787e-22, 4.683483e-22, 
    3.45554e-22, 2.445009e-22, 1.850018e-22, 3.46962e-12, 9.09731e-12, 
    1.993118e-10, 1.050653e-07, 6.53456e-07, 3.097315e-06, 7.43767e-06,
  2.485666e-12, 3.041987e-15, 8.789928e-22, 5.407367e-22, 5.605145e-22, 
    3.365298e-22, 3.03868e-22, 3.234958e-22, 1.69926e-12, 3.88172e-13, 
    3.649725e-10, 2.755776e-07, 6.942074e-07, 2.577902e-06, 3.220204e-06,
  1.222608e-11, 1.553276e-13, 1.325517e-15, 1.178696e-17, 5.389253e-22, 
    3.176866e-22, 2.579548e-22, 1.859974e-22, 1.540742e-14, 1.091964e-13, 
    4.122586e-09, 5.709629e-07, 9.794973e-07, 1.808066e-06, 3.997071e-06,
  2.555695e-11, 5.502484e-10, 3.681104e-12, 4.155292e-15, 2.852686e-16, 
    5.049349e-22, 2.588656e-22, 2.452074e-22, 7.326733e-16, 1.113838e-13, 
    1.211964e-08, 6.553823e-07, 1.322164e-06, 1.255316e-06, 3.192907e-06,
  2.135191e-10, 5.380787e-12, 2.526274e-13, 3.020864e-13, 4.235379e-12, 
    6.215153e-11, 3.475299e-22, 2.390922e-13, 8.120342e-13, 1.891493e-12, 
    5.13615e-07, 1.356987e-07, 1.512561e-06, 2.691848e-06, 2.523379e-06,
  1.769825e-06, 7.397301e-08, 1.880483e-07, 5.281346e-08, 2.893566e-06, 
    2.162788e-06, 2.900656e-06, 4.054541e-06, 4.787462e-06, 8.27595e-06, 
    6.580361e-06, 2.844296e-06, 3.604921e-06, 1.159049e-05, 1.607427e-05,
  7.912874e-06, 1.512787e-06, 5.085256e-07, 2.896755e-07, 3.198651e-06, 
    1.578235e-06, 1.845915e-06, 2.227914e-06, 1.877355e-06, 4.012886e-06, 
    4.75228e-06, 5.967311e-06, 4.468187e-06, 9.379677e-06, 1.122934e-05,
  6.932858e-06, 6.023226e-06, 9.599642e-07, 4.256414e-07, 3.884759e-06, 
    2.584384e-06, 2.89767e-06, 2.36807e-06, 1.754524e-06, 1.806314e-06, 
    3.353524e-06, 4.548503e-06, 4.888062e-06, 6.499587e-06, 9.986526e-06,
  7.870282e-06, 5.174812e-06, 3.759456e-06, 7.100202e-07, 4.256115e-06, 
    3.848789e-06, 2.522782e-06, 1.647108e-06, 1.861944e-06, 2.194803e-06, 
    3.873611e-06, 3.191678e-06, 4.755881e-06, 4.345391e-06, 5.058026e-06,
  6.921916e-06, 6.518444e-06, 2.408931e-06, 1.371061e-06, 1.813488e-06, 
    3.753e-06, 2.192876e-06, 1.796061e-06, 1.511032e-06, 1.312879e-06, 
    2.031548e-06, 2.617664e-06, 2.988316e-06, 4.387623e-06, 3.115637e-06,
  7.071468e-06, 3.473444e-06, 5.888583e-06, 6.965089e-07, 4.549113e-07, 
    1.943315e-06, 2.649343e-06, 2.682778e-06, 2.635699e-06, 3.301868e-06, 
    3.842137e-06, 3.418062e-06, 3.250281e-06, 4.238702e-06, 4.878912e-06,
  6.765106e-06, 6.270364e-06, 9.042237e-06, 5.39649e-06, 3.024034e-07, 
    1.618806e-06, 1.605678e-06, 2.424426e-06, 3.19812e-06, 3.011674e-06, 
    2.829318e-06, 3.000322e-06, 4.517506e-06, 1.246898e-05, 1.571648e-05,
  5.238102e-06, 5.235855e-06, 4.513574e-06, 3.4006e-06, 1.19929e-07, 
    1.093362e-06, 1.416276e-06, 2.15306e-06, 2.81906e-06, 2.691243e-06, 
    3.943361e-06, 6.863368e-06, 1.396386e-05, 1.615952e-05, 1.692551e-05,
  3.178058e-06, 2.602209e-06, 1.443507e-06, 1.962714e-06, 5.185313e-07, 
    6.677811e-09, 5.229134e-07, 7.658857e-07, 4.663741e-06, 4.990306e-06, 
    5.085299e-06, 7.094849e-06, 7.418328e-06, 6.848763e-06, 7.763872e-06,
  9.033619e-07, 1.327039e-06, 1.910434e-06, 1.27346e-06, 8.496291e-07, 
    5.181612e-07, 2.49392e-09, 4.288445e-08, 1.880172e-06, 3.44914e-06, 
    4.875932e-06, 5.622483e-06, 5.188977e-06, 5.342909e-06, 5.999629e-06,
  4.217915e-07, 3.914025e-09, 2.66565e-10, 7.304656e-11, 7.24257e-11, 
    2.731133e-10, 1.573736e-09, 2.949311e-10, 2.212013e-10, 4.634359e-08, 
    6.743189e-07, 6.463387e-07, 5.647149e-07, 1.425143e-06, 2.27192e-06,
  7.780407e-06, 4.283986e-08, 5.238037e-10, 3.97735e-11, 2.852071e-09, 
    3.507112e-10, 1.06818e-09, 1.67414e-09, 1.703938e-10, 2.947821e-10, 
    4.885412e-09, 2.058061e-08, 2.148653e-08, 5.03071e-07, 1.484599e-06,
  3.840842e-06, 5.740457e-07, 1.336704e-08, 6.938203e-10, 2.082671e-08, 
    2.299931e-09, 1.724171e-09, 9.139933e-09, 1.806994e-09, 2.887695e-08, 
    3.873816e-08, 4.421882e-08, 8.25557e-08, 4.791812e-07, 7.902212e-07,
  5.344951e-06, 1.718976e-06, 3.77457e-07, 2.850246e-08, 7.306153e-07, 
    4.115877e-07, 1.885025e-07, 2.323298e-07, 7.74858e-08, 3.091018e-08, 
    1.706731e-08, 2.514506e-07, 4.849394e-07, 8.45146e-07, 1.062707e-06,
  7.547399e-06, 5.29067e-06, 7.779009e-07, 7.629593e-07, 1.546571e-06, 
    2.064215e-06, 1.459759e-06, 1.27652e-06, 8.612103e-07, 5.344556e-07, 
    1.116414e-06, 1.096773e-06, 1.3782e-06, 1.578896e-06, 2.003045e-06,
  6.305218e-06, 6.395515e-06, 1.896152e-06, 3.470881e-06, 1.393973e-06, 
    3.533645e-06, 3.211528e-06, 1.893215e-06, 1.712654e-06, 1.036027e-06, 
    1.270487e-06, 1.783466e-06, 2.314056e-06, 2.596031e-06, 2.562861e-06,
  7.789909e-06, 7.65546e-06, 9.282696e-06, 2.727778e-06, 1.84982e-06, 
    2.76254e-06, 4.658135e-06, 3.484539e-06, 2.358974e-06, 1.541225e-06, 
    1.749697e-06, 2.072594e-06, 1.98777e-06, 2.568825e-06, 3.965089e-06,
  5.175299e-06, 9.026789e-06, 1.303437e-05, 1.263383e-05, 1.738124e-06, 
    3.28326e-06, 5.501888e-06, 5.335668e-06, 3.0321e-06, 3.253494e-06, 
    3.032578e-06, 2.349109e-06, 3.217488e-06, 5.762507e-06, 6.490808e-06,
  2.396327e-06, 6.539483e-06, 7.19234e-06, 9.745364e-06, 1.120537e-05, 
    4.2724e-06, 5.888078e-06, 6.975767e-06, 5.084565e-06, 4.499635e-06, 
    5.64692e-06, 6.096967e-06, 5.937435e-06, 7.565917e-06, 5.560269e-06,
  2.306403e-07, 7.636264e-07, 1.727802e-06, 6.386257e-06, 4.147075e-06, 
    1.259173e-05, 6.664093e-06, 7.166133e-06, 5.902855e-06, 4.886679e-06, 
    6.548039e-06, 8.034365e-06, 9.489469e-06, 7.832463e-06, 7.766173e-06,
  4.488375e-09, 1.113975e-06, 1.848482e-06, 1.313336e-07, 1.181617e-06, 
    2.12746e-06, 3.925099e-07, 2.135447e-07, 5.307903e-07, 4.170862e-07, 
    3.534381e-07, 3.592985e-07, 5.637849e-08, 7.100093e-08, 3.886877e-06,
  1.180617e-06, 6.016971e-08, 5.531254e-07, 4.622826e-09, 2.924316e-06, 
    4.401082e-06, 1.684393e-06, 5.189713e-07, 4.833443e-07, 2.104576e-07, 
    2.031207e-08, 4.089372e-09, 4.559226e-08, 3.546848e-07, 1.201039e-06,
  1.293132e-06, 1.339778e-06, 8.508357e-07, 1.785684e-08, 4.446295e-06, 
    4.27184e-06, 4.076675e-06, 1.386876e-06, 1.154479e-06, 2.169016e-07, 
    4.543514e-08, 6.01491e-10, 1.260287e-09, 4.067734e-08, 5.1665e-07,
  3.63299e-06, 7.081725e-07, 4.431657e-07, 6.407604e-08, 5.164784e-06, 
    3.150755e-06, 4.448305e-06, 4.490655e-06, 2.081366e-06, 1.244774e-06, 
    7.738702e-08, 1.264875e-08, 1.284951e-08, 4.212764e-09, 2.421995e-08,
  1.023012e-06, 1.915625e-06, 4.893853e-07, 1.518999e-07, 2.266272e-06, 
    5.147027e-06, 2.775654e-06, 1.737202e-06, 1.31406e-07, 1.06174e-07, 
    8.418674e-08, 4.385666e-08, 1.552893e-08, 1.158467e-10, 1.420258e-08,
  1.296441e-06, 2.119971e-06, 1.618297e-06, 3.099596e-07, 2.811843e-07, 
    4.38632e-06, 3.441619e-06, 3.150565e-06, 1.478612e-07, 4.458131e-08, 
    1.150198e-07, 7.079403e-07, 4.680521e-08, 2.402774e-09, 3.286732e-08,
  1.187009e-06, 2.770461e-06, 4.340831e-06, 2.907e-06, 8.295278e-07, 
    3.323399e-06, 4.603893e-06, 3.133627e-06, 2.234434e-06, 3.484735e-08, 
    2.48803e-08, 2.742744e-09, 1.495677e-10, 2.214265e-09, 1.145117e-09,
  2.201413e-07, 8.713317e-07, 1.915226e-06, 4.817328e-06, 1.485201e-06, 
    3.756956e-06, 6.474699e-06, 3.687485e-06, 3.158716e-06, 3.025056e-07, 
    5.295364e-07, 5.762199e-08, 2.394156e-10, 3.559301e-12, 3.678925e-11,
  1.332157e-08, 3.032756e-08, 8.667099e-08, 1.566723e-06, 3.24262e-06, 
    4.732387e-06, 4.911026e-06, 7.733804e-06, 5.62272e-06, 3.813996e-06, 
    2.045327e-06, 1.061692e-07, 1.191411e-10, 1.79391e-12, 5.524282e-11,
  2.094503e-08, 1.657801e-08, 7.244218e-09, 3.937287e-08, 1.627743e-07, 
    1.966672e-06, 3.246835e-06, 7.073473e-06, 7.195875e-06, 6.542457e-06, 
    5.531084e-06, 3.257286e-06, 1.558724e-06, 3.667465e-08, 1.299094e-11,
  4.384825e-09, 3.341275e-08, 1.182626e-06, 5.965377e-08, 6.495603e-06, 
    4.312536e-06, 2.813755e-06, 8.884653e-06, 6.124595e-06, 5.792579e-06, 
    2.509175e-06, 1.377091e-06, 1.410285e-06, 5.466904e-07, 2.146556e-06,
  1.482044e-06, 2.437078e-08, 6.358344e-08, 1.132449e-08, 5.950444e-06, 
    4.407077e-06, 2.931857e-06, 2.590987e-06, 4.695257e-06, 2.467701e-06, 
    2.013127e-06, 1.725417e-06, 1.354031e-06, 2.225108e-06, 3.020037e-06,
  4.555494e-07, 6.978567e-08, 5.394544e-09, 2.910775e-08, 1.121078e-06, 
    4.226838e-06, 4.503528e-06, 2.570755e-06, 4.010314e-06, 1.11499e-06, 
    8.447761e-07, 3.569768e-07, 1.738353e-06, 4.151895e-06, 6.543867e-06,
  5.614483e-07, 2.452374e-09, 3.283107e-11, 5.17172e-08, 2.786083e-07, 
    5.375198e-06, 3.566416e-06, 2.197006e-06, 2.291575e-06, 1.714084e-06, 
    1.873595e-06, 1.237493e-06, 1.587214e-06, 2.166281e-06, 4.302573e-06,
  1.225733e-07, 3.80248e-09, 9.009669e-11, 3.774026e-08, 1.462656e-07, 
    1.943137e-06, 5.520981e-06, 4.88565e-06, 2.229002e-06, 1.596909e-06, 
    3.36084e-06, 3.260571e-06, 5.816285e-06, 3.662426e-06, 4.181947e-06,
  1.666645e-08, 7.037428e-09, 1.394688e-09, 1.053556e-11, 1.120434e-09, 
    6.320007e-09, 2.617336e-06, 4.165979e-06, 2.160827e-06, 1.816073e-06, 
    2.938867e-06, 4.77298e-06, 6.304407e-06, 6.33124e-06, 4.499868e-06,
  5.117691e-10, 2.946903e-09, 6.850344e-09, 9.803877e-12, 4.842307e-10, 
    9.069153e-08, 2.699711e-06, 2.42402e-06, 5.123608e-06, 1.040197e-06, 
    2.202e-06, 6.02028e-06, 5.965604e-06, 4.296101e-06, 4.659566e-06,
  8.546665e-13, 2.915922e-15, 4.727149e-14, 1.188685e-11, 9.502601e-10, 
    2.511541e-07, 3.17657e-06, 3.820392e-06, 3.655437e-06, 1.814299e-06, 
    4.791177e-07, 3.87431e-06, 5.10783e-06, 3.476701e-06, 1.817973e-06,
  0, 1.797449e-15, 1.174375e-14, 7.939665e-08, 1.25707e-09, 6.860765e-08, 
    2.015087e-06, 3.182818e-06, 3.42202e-06, 3.196762e-06, 1.820881e-06, 
    7.41224e-07, 2.293326e-06, 2.176814e-06, 2.014032e-06,
  9.072301e-16, 3.549756e-16, 7.633409e-12, 1.434216e-11, 2.162927e-09, 
    2.598053e-09, 1.500979e-07, 3.484696e-06, 3.051095e-06, 4.037102e-06, 
    2.140167e-06, 1.851537e-06, 1.802319e-06, 2.418455e-06, 1.942714e-06,
  3.447916e-07, 5.048026e-07, 1.845359e-06, 3.734476e-06, 3.982597e-06, 
    6.112206e-06, 1.234044e-05, 1.274345e-05, 3.231608e-06, 8.995018e-06, 
    8.830105e-06, 6.171115e-06, 9.950089e-06, 1.230758e-05, 1.488429e-05,
  3.074041e-06, 3.623558e-08, 3.322323e-08, 2.177047e-07, 6.430069e-08, 
    2.377463e-06, 4.323368e-06, 2.173185e-06, 1.94515e-06, 1.075508e-05, 
    9.977e-06, 7.82717e-06, 7.841018e-06, 7.302108e-06, 7.496279e-06,
  1.93399e-06, 1.333685e-06, 1.340746e-08, 1.019885e-08, 1.766649e-08, 
    2.021932e-06, 5.126049e-06, 4.571491e-06, 4.261457e-06, 6.295974e-07, 
    5.704161e-06, 5.007907e-06, 4.281419e-06, 3.731554e-06, 2.651981e-06,
  1.245781e-06, 2.165763e-07, 2.188349e-09, 2.079375e-09, 7.039139e-09, 
    7.458023e-07, 4.052964e-06, 4.271684e-06, 3.353044e-06, 3.223102e-07, 
    2.574127e-06, 4.099388e-06, 3.704459e-06, 3.464427e-06, 3.981496e-06,
  4.642665e-07, 3.127983e-07, 2.707915e-10, 3.749133e-12, 1.769926e-10, 
    2.285305e-08, 1.433565e-06, 4.881088e-06, 3.892079e-06, 3.757534e-07, 
    2.108796e-07, 5.821608e-07, 1.355078e-06, 1.942468e-06, 3.010954e-06,
  2.04399e-08, 2.199601e-07, 1.089113e-09, 1.093007e-12, 3.004888e-10, 
    1.539138e-07, 1.869159e-06, 5.033462e-06, 4.660292e-06, 1.572228e-06, 
    7.869655e-07, 1.222774e-06, 2.670313e-06, 2.415095e-06, 2.503885e-06,
  5.553545e-08, 3.235131e-07, 2.880558e-07, 1.341697e-09, 2.031919e-09, 
    1.414409e-07, 3.338024e-06, 3.953662e-06, 2.066247e-06, 9.72043e-07, 
    9.881434e-07, 1.661785e-06, 3.567897e-06, 4.428934e-06, 5.43584e-06,
  1.4569e-07, 1.212688e-07, 4.401438e-09, 5.31119e-09, 3.523401e-09, 
    7.477374e-08, 5.191127e-06, 7.755088e-06, 1.215044e-06, 4.242855e-07, 
    5.378703e-07, 3.051591e-06, 4.136217e-06, 7.302669e-06, 6.137638e-06,
  1.796638e-07, 9.26641e-08, 3.669042e-08, 3.420535e-10, 5.545657e-09, 
    1.848239e-07, 1.187058e-05, 1.771523e-05, 2.97054e-06, 7.122255e-07, 
    6.136892e-07, 1.394454e-06, 3.189897e-06, 5.794775e-06, 5.142866e-06,
  1.918201e-07, 3.361485e-07, 9.909968e-08, 5.481008e-08, 3.884628e-07, 
    4.554457e-06, 1.860066e-06, 7.401294e-05, 5.694659e-07, 2.897148e-07, 
    8.191972e-07, 6.780964e-07, 2.462016e-06, 6.530326e-06, 6.465642e-06,
  4.280616e-11, 3.178596e-08, 1.342633e-06, 4.071611e-06, 1.892128e-06, 
    2.451343e-06, 5.756419e-06, 1.206327e-05, 1.890361e-05, 2.784743e-05, 
    1.954628e-05, 1.458809e-05, 1.420606e-05, 1.662647e-05, 1.665871e-05,
  1.01488e-10, 6.44565e-08, 1.85413e-06, 5.954109e-06, 6.8565e-06, 
    7.580313e-06, 9.732661e-06, 1.390844e-05, 1.594427e-05, 1.727297e-05, 
    9.305823e-06, 7.949172e-06, 1.112679e-05, 1.330178e-05, 1.286877e-05,
  3.240185e-10, 1.102607e-10, 2.597478e-07, 5.486922e-06, 6.252482e-06, 
    4.513984e-06, 9.93174e-06, 7.797631e-06, 7.612181e-06, 3.335633e-06, 
    1.9408e-06, 5.545356e-06, 9.030755e-06, 1.155401e-05, 1.269945e-05,
  1.823358e-07, 4.435285e-11, 2.257361e-07, 3.642055e-06, 4.254442e-06, 
    8.570922e-06, 1.031551e-05, 6.948374e-06, 2.730686e-06, 6.707576e-07, 
    1.858206e-06, 4.418985e-06, 5.697375e-06, 7.770058e-06, 9.568466e-06,
  7.590896e-08, 6.453192e-09, 1.449781e-07, 1.186389e-06, 1.514478e-06, 
    3.254334e-06, 1.176987e-05, 1.621708e-05, 4.556728e-06, 1.155816e-06, 
    1.830517e-07, 2.047458e-06, 1.104857e-06, 3.447476e-06, 4.713175e-06,
  1.105802e-07, 4.297177e-08, 1.988731e-07, 4.074638e-08, 5.098709e-08, 
    7.439584e-07, 1.237784e-05, 6.637682e-06, 3.395674e-06, 2.650362e-06, 
    6.326203e-07, 3.274749e-07, 2.79812e-07, 6.194185e-08, 1.501772e-07,
  1.297035e-07, 5.300787e-07, 3.36901e-06, 8.099319e-07, 1.436087e-08, 
    3.219536e-07, 1.195776e-05, 1.23272e-05, 1.327939e-06, 3.978319e-07, 
    1.2478e-06, 5.583881e-07, 1.217635e-07, 2.206115e-07, 4.814108e-07,
  4.644477e-08, 4.162134e-07, 3.284132e-06, 3.673858e-06, 1.1557e-08, 
    7.141728e-09, 8.557937e-06, 1.090741e-05, 1.544459e-06, 1.717995e-06, 
    5.393205e-07, 2.87308e-07, 5.750339e-07, 1.164285e-06, 1.408859e-06,
  1.137081e-07, 3.377939e-07, 7.022368e-07, 2.576952e-06, 5.52036e-06, 
    2.802722e-09, 5.76302e-06, 5.050255e-06, 1.258365e-06, 2.384347e-06, 
    1.092567e-06, 6.177715e-07, 1.225583e-06, 1.420552e-06, 2.160504e-06,
  3.289545e-08, 1.143341e-07, 2.27727e-07, 4.429873e-07, 5.204317e-06, 
    1.10014e-05, 2.682489e-09, 4.720857e-06, 5.445669e-07, 9.365134e-07, 
    1.480856e-06, 1.187063e-06, 1.844843e-06, 1.450775e-06, 1.712837e-06,
  6.8578e-10, 1.344403e-07, 8.713576e-06, 1.267918e-05, 6.420429e-06, 
    5.584364e-06, 5.839804e-06, 9.600907e-06, 1.269282e-05, 1.280561e-05, 
    1.259455e-05, 1.34162e-05, 1.442425e-05, 1.310606e-05, 1.549552e-05,
  2.894988e-06, 7.286981e-08, 2.639336e-06, 1.160207e-05, 3.975322e-06, 
    7.167785e-06, 5.805641e-06, 6.845916e-06, 7.889081e-06, 9.043129e-06, 
    9.919367e-06, 9.001084e-06, 6.500042e-06, 6.724705e-06, 6.864675e-06,
  2.968256e-06, 5.418973e-06, 1.01145e-07, 1.594275e-06, 3.241838e-07, 
    5.201868e-07, 1.198623e-06, 1.499681e-06, 1.876069e-06, 1.961106e-06, 
    2.714464e-06, 2.676198e-06, 2.24015e-06, 2.358287e-06, 1.873672e-06,
  3.224314e-06, 5.605263e-06, 4.892229e-09, 2.521305e-08, 1.042436e-08, 
    9.314516e-08, 1.708414e-07, 9.462233e-08, 1.002921e-08, 2.157282e-09, 
    1.508887e-09, 1.530338e-08, 2.447474e-08, 3.98292e-08, 6.28169e-08,
  3.223009e-06, 7.60681e-06, 1.290492e-09, 4.387836e-10, 5.059109e-10, 
    1.50537e-09, 1.616012e-10, 4.614631e-09, 1.451257e-06, 2.046235e-09, 
    1.323865e-08, 1.158562e-08, 1.390169e-08, 1.604806e-08, 2.202852e-08,
  1.076512e-05, 1.037543e-05, 1.754556e-05, 8.750912e-10, 1.140758e-10, 
    8.154313e-11, 1.975743e-10, 4.744841e-09, 4.619501e-07, 4.384179e-07, 
    3.851437e-07, 4.459167e-07, 1.414568e-08, 1.007726e-08, 1.763632e-08,
  9.917209e-06, 3.448369e-05, 4.445979e-05, 3.068901e-05, 1.125899e-10, 
    6.414976e-11, 1.489195e-10, 3.43182e-07, 8.386489e-07, 7.941942e-07, 
    2.285802e-06, 3.800494e-06, 9.627732e-07, 3.050275e-07, 6.924749e-07,
  1.117337e-05, 1.802186e-05, 3.93927e-05, 4.129826e-05, 3.936454e-10, 
    7.679896e-11, 1.076925e-10, 3.463161e-08, 4.776951e-07, 2.06907e-06, 
    3.856861e-06, 4.727186e-06, 3.983855e-06, 1.554654e-06, 7.855654e-07,
  1.553356e-05, 1.8275e-05, 3.569289e-05, 3.992235e-05, 1.458142e-05, 
    2.517374e-11, 1.794418e-10, 1.579983e-07, 1.85383e-07, 4.306632e-06, 
    1.152565e-05, 6.279852e-06, 3.807732e-06, 1.565403e-06, 1.287521e-06,
  2.988065e-05, 3.270739e-05, 2.69982e-05, 2.437537e-05, 1.447049e-05, 
    1.594698e-06, 2.101891e-10, 7.313024e-07, 7.958521e-07, 6.566042e-06, 
    1.599263e-05, 7.782104e-06, 4.525703e-06, 3.198629e-06, 1.661948e-06,
  4.337198e-06, 1.186324e-06, 3.549808e-06, 6.068107e-06, 4.215764e-06, 
    8.003716e-06, 8.803629e-06, 1.836303e-05, 1.613185e-05, 2.026915e-05, 
    1.97204e-05, 2.514684e-05, 2.822576e-05, 3.041807e-05, 3.44447e-05,
  2.697333e-05, 1.203275e-06, 2.150153e-06, 4.448216e-06, 1.665432e-06, 
    2.173688e-06, 6.138139e-06, 8.871427e-06, 8.785108e-06, 1.395933e-05, 
    1.214016e-05, 1.461235e-05, 2.008883e-05, 2.166409e-05, 2.252846e-05,
  6.574469e-06, 1.086711e-05, 2.971264e-07, 3.771931e-07, 2.521579e-07, 
    4.216967e-07, 9.556179e-07, 8.082356e-07, 1.938213e-06, 3.197218e-06, 
    5.220338e-06, 6.672342e-06, 7.135908e-06, 1.127271e-05, 1.755486e-05,
  2.827841e-06, 4.604476e-06, 2.876508e-09, 3.477037e-09, 8.291914e-09, 
    1.362202e-07, 1.363933e-07, 9.118452e-08, 1.810006e-07, 2.228558e-07, 
    4.765591e-07, 1.695817e-06, 2.547607e-06, 4.815388e-06, 7.601519e-06,
  5.071844e-06, 1.04285e-05, 2.857626e-06, 7.571247e-10, 8.8905e-10, 
    4.591948e-10, 7.794015e-06, 1.42993e-05, 1.281855e-05, 6.317611e-07, 
    9.820488e-07, 5.29866e-07, 1.638802e-07, 2.474028e-07, 6.045871e-06,
  4.889007e-06, 3.058006e-06, 3.841598e-06, 5.826699e-10, 1.055462e-09, 
    6.883127e-10, 4.417592e-07, 2.112998e-05, 1.686736e-05, 8.396843e-06, 
    4.813462e-06, 5.512878e-06, 6.793033e-06, 2.427867e-06, 2.813018e-06,
  4.827379e-06, 2.97131e-06, 5.064857e-06, 6.579781e-06, 6.629489e-10, 
    1.273734e-09, 5.42567e-07, 2.785058e-07, 1.610185e-05, 1.587505e-05, 
    1.182362e-05, 1.84197e-05, 1.492922e-05, 1.220342e-05, 7.081314e-06,
  3.537272e-06, 5.318771e-06, 8.660239e-06, 1.533018e-05, 6.531239e-10, 
    1.421286e-09, 1.316789e-07, 5.436888e-07, 4.477883e-06, 1.874931e-05, 
    2.552229e-05, 2.905021e-05, 2.125346e-05, 1.108235e-05, 5.717803e-06,
  5.716315e-06, 6.405635e-06, 1.231144e-05, 2.095389e-05, 9.752896e-06, 
    7.063116e-10, 1.130156e-09, 4.611575e-06, 2.535875e-06, 1.416253e-05, 
    3.19881e-05, 2.661748e-05, 1.540645e-05, 4.48293e-06, 7.343224e-07,
  6.024184e-06, 9.293305e-06, 1.179073e-05, 2.193592e-05, 1.994791e-05, 
    1.696595e-05, 8.705293e-10, 1.258916e-06, 2.592844e-06, 1.905981e-05, 
    3.4414e-05, 1.234679e-05, 3.616782e-06, 1.38147e-06, 3.243862e-07,
  1.954069e-06, 8.224431e-06, 1.489102e-05, 8.657564e-06, 6.275706e-07, 
    1.305232e-06, 3.556929e-07, 2.069758e-07, 3.076999e-07, 4.68605e-07, 
    4.705994e-07, 7.511208e-07, 1.397518e-06, 2.830788e-06, 6.474053e-06,
  1.575937e-05, 8.864141e-06, 6.203261e-06, 1.119656e-05, 1.133413e-05, 
    3.124015e-06, 2.197535e-06, 2.008827e-06, 2.991925e-06, 2.60861e-06, 
    4.419418e-06, 5.396003e-06, 7.195922e-06, 1.156332e-05, 1.472183e-05,
  1.670787e-05, 1.023216e-05, 5.763642e-06, 3.996108e-06, 1.283815e-05, 
    8.468278e-06, 7.654371e-06, 3.923838e-06, 6.211289e-06, 7.994874e-06, 
    8.387273e-06, 1.005329e-05, 1.16008e-05, 1.384037e-05, 1.751634e-05,
  1.01374e-05, 1.077741e-05, 3.21194e-06, 6.796926e-06, 5.34173e-06, 
    1.379881e-05, 1.0869e-05, 1.023463e-05, 1.766082e-05, 9.203892e-06, 
    6.984912e-06, 1.089739e-05, 1.161378e-05, 1.491217e-05, 1.492557e-05,
  4.361794e-06, 6.989368e-06, 3.440803e-06, 3.715821e-06, 5.475424e-06, 
    5.618542e-06, 9.614517e-06, 1.720318e-05, 1.166721e-05, 1.558661e-05, 
    1.563635e-05, 1.924441e-05, 2.581333e-05, 2.40079e-05, 1.574465e-05,
  2.392218e-06, 1.803837e-06, 5.985272e-06, 7.594662e-07, 2.129648e-06, 
    4.294281e-06, 6.426869e-06, 8.490738e-06, 1.619107e-05, 4.61822e-05, 
    4.040814e-05, 4.467811e-05, 4.933168e-05, 2.567627e-05, 3.33248e-05,
  2.296587e-06, 2.314214e-06, 5.435697e-06, 5.113449e-06, 3.731644e-08, 
    8.498748e-07, 3.217099e-06, 2.87567e-06, 7.74915e-06, 5.319588e-05, 
    5.090213e-05, 5.586176e-05, 4.063407e-05, 4.956792e-05, 4.179282e-05,
  2.222854e-06, 2.935751e-06, 3.797675e-06, 4.218994e-06, 3.143316e-10, 
    5.28039e-09, 7.174602e-08, 1.402992e-06, 4.841454e-06, 2.048996e-05, 
    6.159307e-05, 5.494628e-05, 5.376486e-05, 5.000832e-05, 5.580198e-05,
  1.693805e-06, 2.37967e-06, 2.849445e-06, 6.839937e-06, 3.993519e-06, 
    7.447229e-10, 8.752199e-10, 5.925699e-07, 1.413291e-05, 2.314884e-05, 
    2.405767e-05, 3.610429e-05, 7.497789e-05, 5.970494e-05, 6.143671e-05,
  1.305754e-06, 2.114597e-06, 2.660192e-06, 6.898264e-06, 6.952449e-06, 
    6.265736e-06, 9.20809e-10, 8.347093e-10, 8.922826e-06, 1.818272e-05, 
    1.591909e-05, 5.159697e-05, 3.88907e-05, 3.650342e-05, 4.475833e-05,
  7.513822e-07, 2.771823e-06, 4.211037e-06, 1.320799e-06, 2.567357e-06, 
    4.378996e-06, 5.737866e-06, 1.356963e-06, 1.943941e-08, 8.32879e-10, 
    2.479774e-09, 1.475161e-07, 2.658698e-07, 2.103297e-06, 2.972654e-06,
  1.502601e-05, 3.483568e-06, 3.027598e-06, 3.231864e-06, 3.72528e-06, 
    6.853965e-06, 5.525005e-06, 1.041424e-06, 5.723373e-08, 6.162433e-10, 
    1.164387e-08, 3.126891e-08, 1.279501e-08, 4.644705e-07, 2.780957e-06,
  1.71185e-05, 1.481798e-05, 1.847586e-06, 2.059e-06, 3.802276e-06, 
    9.604373e-06, 9.001281e-06, 1.417896e-06, 1.233969e-07, 3.423692e-10, 
    1.631169e-09, 2.677106e-08, 1.569002e-08, 8.942095e-08, 7.048299e-07,
  1.936779e-05, 1.398307e-05, 4.527364e-06, 3.047961e-06, 3.396201e-06, 
    1.505265e-05, 1.505616e-05, 2.005459e-06, 1.526956e-07, 1.14753e-09, 
    6.684909e-11, 1.852524e-09, 6.989693e-08, 4.225697e-07, 4.722331e-07,
  7.949474e-06, 1.22602e-05, 5.157771e-07, 4.412414e-06, 3.557864e-06, 
    7.485022e-06, 1.485374e-05, 1.39831e-05, 3.502798e-06, 2.576481e-07, 
    1.357499e-08, 2.171018e-11, 2.071446e-09, 2.912179e-07, 5.760928e-08,
  5.2894e-06, 6.730096e-06, 4.474987e-06, 3.163132e-07, 3.834283e-06, 
    3.188293e-06, 9.209098e-06, 1.005871e-05, 5.807343e-06, 6.814804e-06, 
    8.756953e-07, 1.335662e-09, 5.988464e-10, 1.749569e-08, 4.585499e-08,
  5.615895e-06, 5.959624e-06, 1.115974e-05, 5.840738e-06, 1.074965e-06, 
    2.687474e-06, 5.888881e-06, 6.766348e-06, 1.181504e-05, 4.488484e-06, 
    5.254426e-06, 2.285902e-06, 4.358142e-07, 4.20024e-09, 7.994666e-09,
  1.495224e-06, 5.523484e-06, 7.608261e-06, 9.74249e-06, 1.318857e-07, 
    1.583816e-06, 1.82915e-06, 5.291301e-06, 7.960514e-06, 9.309642e-06, 
    9.932603e-06, 8.878746e-06, 6.686027e-06, 1.422219e-06, 6.217873e-07,
  8.428471e-07, 1.652447e-06, 5.483211e-06, 4.35532e-06, 7.153157e-06, 
    2.547071e-07, 9.295566e-07, 1.582727e-06, 3.792892e-06, 6.220428e-06, 
    1.153318e-05, 1.540347e-05, 8.980957e-06, 5.995523e-06, 5.559709e-06,
  4.352418e-07, 6.14391e-07, 1.338458e-06, 2.487766e-06, 3.540864e-06, 
    3.768678e-06, 2.098229e-07, 8.745492e-07, 4.499409e-06, 5.183825e-06, 
    4.14455e-06, 1.041729e-05, 1.340055e-05, 1.445639e-05, 8.201713e-06,
  5.696139e-06, 3.632661e-06, 1.729162e-06, 2.15045e-06, 2.849018e-06, 
    3.119195e-06, 1.24927e-05, 3.382913e-05, 6.222614e-05, 7.006071e-05, 
    2.464884e-05, 1.833118e-05, 1.032725e-05, 1.810141e-06, 8.792568e-07,
  5.831502e-05, 1.978923e-06, 3.78189e-07, 3.815616e-07, 2.620842e-07, 
    7.108568e-07, 1.643062e-05, 4.830481e-05, 3.879523e-05, 0.0001024448, 
    2.657167e-05, 3.381384e-06, 2.364797e-06, 2.929999e-06, 2.751518e-06,
  2.308228e-05, 1.609227e-05, 8.347106e-08, 3.040053e-07, 9.877933e-08, 
    1.123418e-06, 1.10427e-05, 4.736183e-05, 2.972927e-05, 1.426701e-06, 
    9.518191e-07, 9.791233e-07, 1.66759e-06, 2.7059e-06, 1.410579e-06,
  6.192638e-06, 5.771037e-06, 1.58085e-08, 4.023938e-08, 3.161406e-08, 
    1.504489e-06, 1.761283e-06, 3.080526e-05, 1.624215e-05, 2.185531e-06, 
    9.741404e-07, 6.946393e-07, 9.290646e-07, 6.518317e-07, 8.927025e-07,
  4.579765e-06, 5.055725e-06, 2.939133e-09, 7.946848e-09, 1.870266e-08, 
    6.281743e-07, 1.50675e-06, 1.587508e-05, 1.103003e-05, 1.36436e-05, 
    6.954442e-06, 2.930704e-06, 8.454218e-07, 9.92786e-07, 4.709624e-07,
  1.147711e-06, 2.755821e-06, 4.442472e-06, 5.172283e-09, 4.196799e-08, 
    1.510824e-07, 1.563952e-06, 8.589937e-06, 1.31858e-05, 7.739109e-06, 
    6.68078e-06, 7.088961e-06, 3.061679e-06, 5.624947e-07, 2.168507e-07,
  1.959386e-06, 1.393182e-06, 3.131913e-06, 6.630797e-06, 6.765013e-09, 
    1.613147e-07, 2.289956e-06, 1.753203e-06, 9.072654e-06, 9.233967e-06, 
    1.041127e-05, 7.779762e-06, 4.143762e-06, 1.231472e-06, 5.674055e-08,
  1.254445e-06, 7.30302e-07, 1.428093e-06, 3.326661e-06, 6.059496e-09, 
    1.807536e-07, 9.206022e-07, 2.369188e-06, 2.734658e-06, 5.273731e-06, 
    6.059994e-06, 9.264991e-06, 5.527959e-06, 7.550062e-07, 5.142703e-08,
  9.491316e-07, 1.53739e-07, 4.182499e-07, 2.178112e-06, 2.720756e-06, 
    2.258473e-09, 8.441545e-07, 2.755322e-06, 2.761411e-06, 3.064511e-06, 
    8.156827e-06, 9.876869e-06, 7.053641e-06, 2.239613e-06, 1.538876e-07,
  5.622937e-07, 1.982701e-07, 3.347851e-08, 3.451893e-08, 1.944104e-07, 
    6.164857e-07, 5.133046e-08, 2.556024e-06, 2.888064e-06, 4.586958e-06, 
    8.803306e-06, 9.166305e-06, 8.880671e-06, 7.539486e-06, 8.918157e-07,
  2.985872e-06, 1.266297e-06, 1.607016e-06, 3.358781e-06, 3.907774e-06, 
    3.938637e-06, 3.840618e-06, 5.301702e-06, 4.107947e-06, 8.741427e-06, 
    2.45061e-05, 4.087491e-05, 5.494544e-05, 6.899104e-05, 7.766289e-05,
  1.219013e-05, 6.173247e-06, 2.889637e-06, 1.804638e-06, 3.274984e-06, 
    4.934862e-06, 5.844307e-06, 5.984576e-06, 9.111163e-06, 2.369098e-05, 
    0.0001076207, 6.177574e-05, 7.457524e-05, 7.820022e-05, 8.571062e-05,
  9.645831e-06, 7.084812e-06, 1.732945e-06, 6.481303e-07, 5.612999e-07, 
    1.369056e-06, 1.707407e-06, 5.900122e-06, 3.120307e-05, 6.306407e-05, 
    4.944869e-05, 4.494385e-05, 6.025678e-05, 6.946673e-05, 8.267382e-05,
  1.000965e-05, 5.5001e-06, 1.214508e-06, 1.127414e-06, 7.604629e-07, 
    1.706343e-06, 1.788142e-05, 3.194272e-05, 4.299193e-05, 2.890638e-05, 
    1.360655e-05, 1.931398e-05, 2.925838e-05, 3.822767e-05, 5.258555e-05,
  4.651772e-05, 9.499806e-06, 7.856407e-06, 3.531686e-06, 2.367568e-06, 
    5.487647e-06, 1.360575e-05, 3.32285e-05, 6.248932e-05, 2.683886e-05, 
    5.346441e-05, 6.921961e-05, 1.256066e-05, 0.0001254124, 7.582964e-05,
  4.584319e-05, 6.24677e-05, 1.387084e-05, 5.117044e-06, 3.685346e-06, 
    1.396745e-05, 1.889772e-05, 3.716203e-05, 5.086476e-05, 6.358547e-05, 
    6.042575e-05, 8.599181e-05, 5.709289e-05, 5.597268e-05, 5.93903e-05,
  3.144944e-05, 4.505655e-05, 6.310317e-05, 2.233283e-05, 2.740613e-06, 
    1.75901e-05, 1.063895e-05, 2.170004e-05, 4.22241e-05, 6.014791e-05, 
    6.656162e-05, 6.977037e-05, 7.914478e-05, 8.740847e-05, 9.830758e-05,
  1.536744e-05, 2.820781e-05, 3.866366e-05, 5.231766e-05, 2.34291e-05, 
    2.162476e-05, 2.550535e-05, 1.130156e-05, 4.205059e-05, 4.82207e-05, 
    3.805991e-05, 6.593797e-05, 7.864768e-05, 8.296676e-05, 7.36642e-05,
  1.075771e-05, 9.675374e-06, 1.303516e-05, 2.446361e-05, 2.842011e-05, 
    5.433997e-06, 6.764612e-06, 9.002246e-06, 1.482652e-05, 4.765996e-05, 
    5.832979e-05, 6.05755e-05, 7.238216e-05, 6.504413e-05, 6.322854e-05,
  3.242706e-06, 2.544209e-06, 1.426698e-06, 2.796882e-06, 4.813309e-06, 
    7.709865e-06, 6.928357e-09, 1.817061e-06, 4.987272e-06, 1.289337e-05, 
    2.56841e-05, 2.371785e-05, 3.486505e-05, 2.432471e-05, 3.147882e-05,
  0.0001029991, 4.594694e-05, 3.990547e-06, 5.353112e-07, 1.040375e-06, 
    3.079867e-06, 8.106298e-06, 1.190838e-05, 1.57842e-05, 2.661891e-05, 
    3.589934e-05, 4.633328e-05, 6.342426e-05, 5.504876e-05, 5.741135e-05,
  5.1845e-05, 6.526824e-05, 3.353536e-05, 3.976056e-06, 9.260073e-07, 
    1.450765e-06, 2.365472e-06, 4.056308e-06, 7.080762e-06, 1.381442e-05, 
    1.844191e-05, 2.384231e-05, 2.929019e-05, 4.330486e-05, 6.409032e-05,
  2.9109e-05, 3.047922e-05, 5.270075e-05, 2.913565e-05, 6.772094e-06, 
    1.073622e-06, 1.082567e-06, 2.570092e-06, 5.033306e-06, 8.008185e-06, 
    1.279825e-05, 1.759841e-05, 2.209554e-05, 3.037846e-05, 5.570576e-05,
  4.88915e-05, 1.635477e-05, 2.556805e-05, 4.00754e-05, 2.834502e-05, 
    7.747905e-06, 6.67588e-07, 4.038665e-07, 1.769693e-06, 3.672062e-06, 
    6.770425e-06, 1.015362e-05, 1.508444e-05, 2.267943e-05, 2.992468e-05,
  1.530054e-05, 1.406315e-05, 1.664414e-05, 2.307277e-05, 3.497647e-05, 
    2.547578e-05, 6.374011e-06, 1.29233e-06, 4.414424e-07, 1.295622e-06, 
    5.387878e-06, 7.624354e-06, 8.687682e-06, 1.260267e-05, 1.599686e-05,
  3.027539e-05, 1.413318e-05, 1.525886e-05, 1.259721e-05, 2.659057e-05, 
    3.63558e-05, 2.300204e-05, 3.625645e-06, 1.84896e-06, 1.546756e-06, 
    1.8934e-06, 4.310295e-06, 5.73157e-06, 6.222868e-06, 7.900864e-06,
  7.352958e-05, 7.406743e-05, 2.439413e-05, 1.526958e-05, 1.103785e-05, 
    2.194036e-05, 2.777544e-05, 1.708753e-05, 4.960288e-06, 2.285541e-06, 
    1.756216e-06, 2.949903e-06, 2.459797e-06, 3.608729e-06, 4.733915e-06,
  4.244089e-05, 0.0001021187, 8.29999e-05, 4.296445e-05, 2.475517e-05, 
    1.23425e-05, 4.872013e-05, 1.823751e-05, 9.431797e-06, 4.276058e-06, 
    3.602111e-06, 3.935926e-06, 2.828828e-06, 2.894977e-06, 2.476967e-06,
  4.720877e-06, 3.256868e-05, 6.820863e-05, 9.030027e-05, 9.145159e-05, 
    7.536147e-05, 4.609175e-05, 3.319271e-05, 7.454503e-06, 6.09357e-06, 
    5.062336e-06, 4.264644e-06, 4.165921e-06, 3.064981e-06, 3.332487e-06,
  4.39799e-06, 5.297778e-06, 1.064302e-05, 4.149831e-05, 8.049993e-05, 
    5.434361e-05, 7.154806e-05, 8.166847e-05, 3.135188e-05, 1.094654e-05, 
    1.288804e-05, 8.91692e-06, 9.766776e-06, 2.47747e-05, 2.487671e-05,
  3.557744e-05, 1.548652e-05, 5.005176e-06, 6.223357e-06, 5.847477e-06, 
    6.796613e-06, 1.634084e-05, 2.985802e-05, 3.02923e-05, 5.203628e-05, 
    5.362673e-05, 7.268137e-05, 5.114529e-05, 7.256066e-05, 0.0001193907,
  4.58392e-05, 3.730124e-05, 2.448306e-05, 7.274254e-06, 7.806508e-06, 
    6.66033e-06, 1.038792e-05, 1.604381e-05, 2.172375e-05, 3.317659e-05, 
    4.460053e-05, 4.837276e-05, 4.663834e-05, 5.772826e-05, 0.0001027407,
  4.061206e-05, 5.020656e-05, 5.485632e-05, 3.642396e-05, 1.349671e-05, 
    1.037612e-05, 8.456673e-06, 1.350366e-05, 1.999036e-05, 2.719964e-05, 
    3.274662e-05, 4.020918e-05, 4.454036e-05, 7.158091e-05, 5.6804e-05,
  2.184709e-05, 3.920042e-05, 6.635368e-05, 7.029264e-05, 5.868083e-05, 
    3.659634e-05, 2.348627e-05, 1.728359e-05, 1.563906e-05, 2.083592e-05, 
    3.009142e-05, 3.129983e-05, 4.385146e-05, 3.691183e-05, 3.57274e-05,
  1.204862e-05, 7.121948e-06, 3.395952e-05, 6.884415e-05, 7.866218e-05, 
    8.375572e-05, 7.056122e-05, 4.973683e-05, 3.762131e-05, 2.591751e-05, 
    2.581068e-05, 3.09563e-05, 3.420303e-05, 3.296359e-05, 2.754578e-05,
  3.980979e-05, 3.010113e-05, 9.216776e-06, 2.715833e-05, 6.309699e-05, 
    9.185576e-05, 0.0001087067, 0.0001033872, 8.86604e-05, 6.068798e-05, 
    4.651131e-05, 3.786191e-05, 3.683952e-05, 3.234322e-05, 2.130046e-05,
  7.045291e-05, 6.771032e-05, 6.466685e-05, 2.540931e-05, 2.296949e-05, 
    5.643968e-05, 9.766701e-05, 0.000120947, 0.0001316882, 0.0001152921, 
    8.801209e-05, 6.226599e-05, 4.114378e-05, 2.365667e-05, 1.514741e-05,
  4.702557e-05, 6.077188e-05, 3.761033e-05, 6.149957e-05, 1.029207e-06, 
    2.691701e-05, 4.550856e-05, 0.0001067888, 0.0001321531, 0.0001378096, 
    0.0001103784, 7.087796e-05, 2.529608e-05, 1.407006e-05, 7.702709e-06,
  2.878414e-05, 4.144707e-05, 3.751867e-05, 4.217648e-05, 4.76299e-05, 
    5.884051e-06, 4.611809e-05, 9.702152e-05, 0.0001618781, 9.727885e-05, 
    6.541557e-05, 4.269371e-05, 9.714371e-06, 2.609979e-06, 2.97543e-06,
  8.678675e-06, 1.068147e-05, 1.35826e-05, 3.206008e-05, 2.707432e-05, 
    3.097924e-05, 1.406458e-05, 3.098269e-05, 7.342876e-05, 3.196395e-05, 
    1.799236e-05, 4.612884e-06, 9.582446e-07, 1.299093e-06, 1.49835e-06,
  2.872753e-07, 7.986044e-08, 1.163104e-09, 7.448244e-13, 3.334007e-13, 
    1.209575e-13, 1.281205e-12, 1.872973e-08, 4.550208e-07, 2.679463e-06, 
    3.804439e-06, 6.416304e-06, 1.242806e-05, 2.068757e-05, 3.710404e-05,
  9.89139e-08, 9.801521e-08, 1.644499e-07, 2.758979e-08, 5.601623e-09, 
    9.321528e-09, 2.799632e-24, 7.496823e-08, 9.997155e-08, 5.483677e-07, 
    4.440559e-06, 8.939551e-06, 1.461071e-05, 2.196526e-05, 2.399882e-05,
  4.819093e-08, 3.416874e-08, 2.999903e-07, 1.783193e-07, 2.298055e-07, 
    3.544163e-08, 1.287836e-07, 1.0401e-07, 1.541541e-07, 4.561169e-07, 
    1.028384e-06, 4.418882e-06, 8.562339e-06, 1.996618e-05, 4.179875e-05,
  1.05781e-07, 1.271843e-07, 6.424874e-08, 4.563701e-07, 2.904053e-07, 
    2.145213e-07, 2.660811e-07, 3.299635e-07, 4.347667e-12, 3.469121e-07, 
    1.004329e-06, 2.754621e-06, 5.949639e-06, 1.353268e-05, 5.62106e-05,
  7.898867e-07, 1.063676e-06, 3.673306e-08, 2.690692e-07, 1.492376e-07, 
    3.837352e-07, 3.720924e-07, 3.505338e-07, 3.918381e-07, 9.28507e-07, 
    1.564704e-06, 2.59211e-06, 6.420859e-06, 1.288296e-05, 4.475039e-05,
  1.278467e-06, 1.633177e-06, 1.137285e-06, 1.996576e-06, 6.880056e-07, 
    5.664732e-07, 2.983685e-07, 2.31092e-07, 6.859698e-07, 5.253681e-07, 
    6.57383e-07, 3.063865e-06, 6.515118e-06, 2.827937e-05, 3.735004e-05,
  3.031489e-06, 2.493339e-06, 6.598797e-06, 2.352087e-06, 2.393718e-06, 
    1.247955e-06, 8.096134e-07, 4.878615e-07, 6.395946e-07, 1.401563e-06, 
    2.222269e-06, 5.371734e-06, 2.103742e-05, 3.759397e-05, 4.597757e-05,
  1.488195e-05, 6.781666e-06, 2.307206e-06, 4.914592e-06, 9.107659e-07, 
    3.475465e-06, 6.746444e-06, 3.594421e-06, 2.609656e-06, 8.822717e-06, 
    2.690344e-05, 4.716507e-05, 5.828537e-05, 5.029244e-05, 5.670773e-05,
  6.29312e-06, 1.15738e-05, 3.6903e-06, 3.662271e-06, 4.960507e-06, 
    1.240921e-05, 5.916253e-06, 6.273065e-06, 2.31669e-05, 3.78029e-05, 
    8.980349e-05, 0.0001280425, 0.0001398745, 0.0001064027, 7.509705e-05,
  2.249167e-06, 6.349401e-06, 1.588692e-05, 1.515654e-05, 1.50567e-05, 
    1.168569e-05, 1.139998e-05, 3.101968e-05, 5.002665e-05, 9.785244e-05, 
    0.0001139106, 0.0001743421, 0.0001919187, 0.0001938623, 0.0001419773,
  7.304575e-07, 3.902008e-06, 1.097651e-05, 1.873328e-05, 2.58723e-05, 
    4.392953e-05, 6.970004e-05, 9.14605e-05, 9.778547e-05, 6.720488e-05, 
    3.883899e-05, 2.280574e-05, 2.426666e-05, 1.003392e-05, 1.180223e-05,
  2.865638e-05, 1.274738e-08, 2.762746e-08, 4.58283e-07, 1.005306e-05, 
    2.229025e-05, 3.704309e-05, 5.485771e-05, 7.356988e-05, 9.876295e-05, 
    9.70784e-05, 6.961566e-05, 3.738984e-05, 2.348771e-05, 2.085194e-05,
  2.037388e-05, 1.273904e-05, 4.26333e-09, 1.645799e-08, 3.436855e-08, 
    1.045627e-05, 2.60945e-05, 3.357769e-05, 2.512111e-05, 6.279371e-05, 
    4.33958e-05, 7.139473e-05, 8.095298e-05, 7.555367e-05, 5.551911e-05,
  1.84913e-05, 1.374465e-05, 1.765235e-09, 3.697032e-09, 4.5833e-09, 
    4.392621e-08, 5.577817e-07, 6.834475e-06, 1.487758e-05, 3.626324e-05, 
    3.887737e-05, 5.325883e-05, 0.0001078442, 6.254729e-05, 8.756432e-05,
  1.928793e-05, 1.206689e-05, 3.339401e-10, 1.104669e-09, 4.974384e-09, 
    3.187396e-07, 8.581599e-07, 1.125516e-06, 1.17609e-06, 2.085299e-06, 
    1.179319e-05, 3.428465e-05, 3.413231e-05, 4.071379e-05, 9.883138e-05,
  1.578503e-05, 6.181176e-06, 6.310382e-08, 4.155954e-10, 1.123861e-07, 
    1.178396e-06, 1.554755e-06, 1.089726e-06, 7.147948e-07, 1.271237e-06, 
    8.407714e-07, 1.21914e-06, 1.155948e-06, 3.910572e-07, 8.70008e-06,
  4.874653e-06, 6.80986e-06, 9.535319e-07, 1.336804e-08, 6.343097e-08, 
    3.370126e-07, 1.709927e-06, 1.374912e-06, 1.044585e-06, 6.384792e-07, 
    7.679158e-07, 4.667428e-07, 6.271469e-07, 7.810885e-07, 6.875557e-07,
  2.310778e-06, 3.187407e-06, 1.217464e-06, 1.43188e-07, 2.41638e-09, 
    3.863038e-09, 7.854496e-07, 1.592416e-06, 1.81756e-06, 1.049465e-06, 
    1.451651e-06, 1.103279e-06, 1.429877e-06, 1.046629e-06, 6.024423e-07,
  2.015737e-06, 1.476164e-06, 1.191091e-06, 1.117207e-06, 1.00628e-09, 
    4.891359e-12, 3.860818e-08, 1.508486e-06, 1.640023e-06, 2.765403e-06, 
    2.145323e-06, 2.697317e-06, 1.673342e-06, 1.221564e-06, 5.72211e-07,
  7.619204e-07, 1.543266e-06, 1.685395e-06, 2.08363e-06, 4.393256e-07, 
    1.433724e-07, 3.232118e-09, 9.884257e-07, 1.249997e-06, 3.048391e-06, 
    2.573121e-06, 1.887351e-06, 2.443982e-06, 3.127331e-06, 9.392818e-07,
  1.371267e-05, 8.220039e-06, 5.051212e-06, 2.619822e-06, 2.664214e-06, 
    3.136006e-06, 3.703162e-06, 3.934131e-06, 2.164111e-06, 3.332249e-06, 
    4.741299e-06, 6.482569e-06, 7.471961e-06, 6.837563e-06, 8.99e-06,
  8.63539e-06, 6.126653e-06, 6.209616e-06, 8.424086e-06, 9.186353e-06, 
    7.048825e-06, 5.098992e-06, 4.936953e-06, 4.178093e-06, 3.573515e-06, 
    3.373032e-06, 3.406037e-06, 3.406428e-06, 3.884669e-06, 2.900837e-06,
  8.634112e-06, 4.313356e-06, 3.161344e-06, 2.237596e-06, 4.267587e-06, 
    6.388932e-06, 3.517992e-06, 2.461342e-06, 4.645776e-06, 7.90706e-06, 
    6.887297e-06, 7.653434e-06, 7.175934e-06, 5.474945e-06, 3.874668e-06,
  1.08384e-05, 6.56598e-06, 2.018602e-06, 1.545201e-06, 1.107851e-06, 
    3.910427e-06, 2.273478e-05, 1.963849e-05, 1.998388e-05, 8.099953e-06, 
    6.979362e-06, 1.25897e-05, 1.873158e-05, 2.213482e-05, 2.357313e-05,
  1.181579e-05, 8.955021e-06, 4.709267e-06, 1.35305e-06, 1.434893e-06, 
    2.475489e-06, 7.923625e-06, 1.729736e-05, 2.055093e-05, 2.543134e-05, 
    3.792869e-05, 3.704302e-05, 4.291777e-05, 0.0001036622, 5.765189e-05,
  4.870003e-05, 2.409819e-05, 9.962352e-06, 4.60839e-06, 3.180913e-06, 
    3.916044e-06, 5.200277e-06, 2.338681e-05, 2.950732e-05, 4.595249e-05, 
    4.027338e-05, 3.608376e-05, 5.608614e-05, 0.0001231711, 7.463119e-05,
  6.837657e-05, 6.416501e-05, 3.397921e-05, 2.665278e-05, 3.45084e-06, 
    2.886399e-06, 5.179777e-06, 2.817963e-05, 3.665553e-05, 3.866828e-05, 
    3.797871e-05, 3.671754e-05, 2.8186e-05, 4.417897e-05, 9.421192e-05,
  4.115135e-05, 6.803474e-05, 6.421711e-05, 7.685989e-05, 1.029705e-05, 
    4.7719e-06, 1.39356e-05, 2.667328e-05, 3.538522e-05, 4.572552e-05, 
    3.041431e-05, 2.649866e-05, 3.160291e-05, 2.965636e-05, 5.94192e-05,
  1.617325e-05, 1.619102e-05, 3.422892e-05, 5.244149e-05, 6.10534e-05, 
    1.487146e-05, 1.820861e-05, 1.893468e-05, 2.390308e-05, 2.814406e-05, 
    3.082299e-05, 2.401469e-05, 3.362988e-05, 4.820993e-05, 4.0487e-05,
  1.207588e-05, 7.97465e-06, 9.403558e-06, 9.427427e-06, 3.065541e-05, 
    4.905481e-05, 4.372746e-06, 1.57222e-05, 2.90623e-05, 3.545526e-05, 
    4.284941e-05, 4.026731e-05, 4.20908e-05, 4.759577e-05, 4.375514e-05,
  3.477425e-08, 5.14121e-09, 2.106582e-09, 1.194218e-09, 3.501275e-09, 
    1.241607e-10, 4.145109e-07, 1.175295e-06, 3.963137e-06, 5.459352e-06, 
    6.982124e-06, 5.617922e-06, 5.452738e-06, 6.435783e-06, 6.627894e-06,
  8.100028e-06, 1.466554e-08, 2.346157e-09, 2.126943e-10, 2.263731e-08, 
    3.027867e-08, 1.224598e-07, 9.249513e-07, 2.601117e-06, 5.773884e-06, 
    5.687291e-06, 6.059763e-06, 5.568242e-06, 6.891992e-06, 8.569739e-06,
  1.342326e-05, 2.157416e-06, 2.421735e-07, 4.584398e-10, 2.757193e-08, 
    4.304803e-07, 1.483714e-08, 1.667734e-07, 1.966675e-06, 4.45056e-06, 
    5.721619e-06, 5.661837e-06, 5.524868e-06, 5.702388e-06, 6.452914e-06,
  5.057862e-05, 1.873371e-05, 1.304079e-06, 4.578206e-09, 1.22554e-07, 
    6.048713e-07, 2.430213e-08, 1.506006e-09, 9.522672e-08, 2.28887e-06, 
    3.492642e-06, 4.120795e-06, 4.459342e-06, 5.613914e-06, 4.731558e-06,
  8.408697e-05, 6.24958e-05, 2.496457e-06, 1.732583e-07, 4.906144e-09, 
    2.086849e-07, 5.420157e-09, 2.264322e-09, 4.610075e-09, 2.618552e-08, 
    1.68145e-07, 8.165098e-07, 2.518455e-06, 2.254115e-06, 4.261206e-06,
  0.0001057003, 7.776383e-05, 5.332154e-05, 2.296244e-06, 3.372489e-06, 
    1.000269e-06, 1.506164e-06, 7.024948e-08, 5.241983e-10, 3.903929e-10, 
    2.393241e-08, 1.008737e-07, 1.073061e-07, 5.179015e-07, 1.433202e-06,
  9.486966e-05, 0.0001035246, 6.382668e-05, 3.860674e-05, 2.697415e-06, 
    7.318095e-06, 4.081158e-06, 3.777415e-06, 1.717894e-07, 8.508371e-09, 
    1.034445e-09, 1.475829e-08, 1.122857e-07, 1.795933e-07, 1.077558e-06,
  5.814989e-05, 6.421137e-05, 4.704416e-05, 5.358371e-05, 1.065981e-05, 
    9.653384e-06, 1.76606e-05, 6.524122e-06, 1.977135e-06, 1.13046e-06, 
    7.983105e-07, 2.912247e-08, 3.950552e-08, 1.557195e-07, 4.209888e-07,
  2.947164e-05, 3.46546e-05, 2.831343e-05, 3.185077e-05, 3.464836e-05, 
    3.943484e-05, 2.202784e-05, 1.010969e-05, 6.876772e-06, 7.98305e-06, 
    3.318773e-06, 2.540858e-07, 4.15883e-08, 1.099271e-08, 8.341363e-08,
  1.881366e-05, 2.175152e-05, 9.462259e-06, 1.789857e-05, 6.231708e-06, 
    1.386121e-05, 3.411769e-05, 4.831258e-05, 5.184022e-05, 1.537365e-05, 
    1.406004e-05, 6.795933e-06, 5.666786e-06, 1.929475e-07, 1.705771e-07,
  1.403792e-07, 7.666263e-07, 1.408059e-07, 4.024596e-07, 2.01983e-06, 
    2.055025e-06, 1.148466e-05, 2.64303e-05, 2.613779e-05, 1.916063e-05, 
    2.839367e-05, 1.357338e-05, 5.762665e-06, 1.861526e-06, 2.290289e-06,
  4.767301e-05, 3.520311e-08, 1.32898e-08, 8.714922e-08, 3.399319e-06, 
    4.021915e-06, 4.286315e-06, 1.26852e-05, 1.780378e-05, 2.459549e-05, 
    2.51988e-05, 1.595321e-05, 8.918217e-06, 4.690228e-06, 1.487596e-05,
  6.720251e-05, 4.546028e-05, 2.344693e-07, 1.643976e-07, 1.952757e-06, 
    1.812916e-06, 7.505227e-06, 7.31508e-06, 1.112314e-05, 1.411843e-05, 
    1.492631e-05, 1.282787e-05, 4.484886e-06, 9.806703e-06, 2.328676e-05,
  8.608361e-05, 0.0001027309, 1.321032e-06, 6.691405e-08, 1.240326e-07, 
    3.703371e-05, 2.268999e-05, 1.415026e-05, 5.349515e-06, 6.018132e-06, 
    6.496537e-06, 7.795098e-06, 9.650597e-06, 1.51286e-05, 7.395104e-06,
  7.105627e-05, 9.461889e-05, 2.388703e-06, 6.987295e-08, 9.689558e-08, 
    2.845435e-05, 6.405091e-05, 4.496186e-05, 1.077192e-05, 1.257057e-06, 
    1.58971e-06, 2.430902e-06, 3.361774e-06, 3.869978e-06, 2.988836e-06,
  4.60463e-05, 5.075007e-05, 7.77302e-05, 1.635902e-08, 6.26412e-06, 
    3.925653e-05, 5.130546e-05, 8.665563e-05, 2.839562e-05, 7.83282e-07, 
    1.852107e-06, 3.864755e-07, 5.421577e-08, 3.522287e-07, 1.022992e-06,
  2.227794e-05, 4.182124e-05, 3.920348e-05, 6.679435e-05, 8.639779e-09, 
    1.398013e-05, 6.239241e-05, 7.631454e-05, 6.975821e-05, 3.687959e-05, 
    4.344738e-06, 6.426105e-06, 1.35844e-06, 2.070901e-06, 2.331346e-06,
  6.328819e-05, 6.69336e-05, 5.510487e-05, 5.612591e-05, 4.796739e-08, 
    5.101674e-06, 1.577238e-05, 5.210045e-05, 7.315444e-05, 6.588399e-05, 
    4.744131e-05, 5.900306e-05, 5.626982e-05, 3.705387e-05, 9.066422e-06,
  0.0001392742, 0.0001190655, 6.922512e-05, 4.330033e-05, 3.110091e-05, 
    9.0201e-08, 5.186687e-06, 3.659585e-05, 6.98068e-05, 5.981057e-05, 
    7.897789e-05, 0.0001146431, 8.629954e-05, 9.703503e-05, 5.043163e-05,
  0.0001331233, 0.0001214622, 6.508278e-05, 5.034224e-05, 5.245237e-05, 
    2.781819e-05, 4.89913e-08, 1.843675e-06, 4.971704e-05, 5.838197e-05, 
    4.009343e-05, 5.472599e-05, 9.445911e-05, 9.389241e-05, 7.266612e-05,
  3.961058e-06, 7.38366e-06, 3.95084e-06, 5.456321e-06, 6.670577e-06, 
    6.217411e-06, 3.688821e-06, 3.613818e-06, 4.063787e-06, 8.200744e-07, 
    8.870611e-08, 2.195688e-10, 6.27382e-11, 8.158282e-11, 1.397702e-10,
  7.356957e-06, 6.12632e-06, 2.626312e-06, 1.688666e-06, 3.8719e-06, 
    3.183849e-06, 4.703562e-06, 9.745633e-06, 4.817559e-06, 1.81128e-06, 
    2.694351e-07, 1.421515e-08, 9.161177e-11, 1.403979e-10, 1.671689e-10,
  9.644629e-06, 1.10778e-05, 5.860385e-06, 3.295021e-07, 5.288468e-07, 
    2.057062e-06, 3.79547e-06, 3.67925e-06, 6.934046e-06, 8.120236e-06, 
    8.17212e-07, 3.439848e-07, 1.211629e-07, 4.719646e-10, 1.128523e-10,
  8.172108e-06, 6.811416e-06, 5.844152e-06, 4.237729e-06, 3.750693e-06, 
    4.91316e-06, 3.683168e-06, 3.533333e-06, 5.237085e-06, 8.014106e-06, 
    7.550096e-06, 4.257569e-06, 1.957549e-06, 4.0067e-07, 1.306225e-07,
  5.570087e-06, 5.461954e-06, 2.137712e-06, 2.205397e-06, 7.872753e-07, 
    6.646661e-06, 5.283932e-06, 3.876346e-06, 3.309998e-06, 4.779368e-06, 
    6.98134e-06, 9.148314e-06, 9.761241e-06, 6.757182e-06, 5.332594e-06,
  2.480302e-06, 8.158515e-06, 5.621064e-06, 3.628415e-07, 4.365762e-06, 
    2.787255e-06, 1.136266e-05, 1.544674e-05, 6.733618e-06, 3.274191e-06, 
    2.415081e-06, 5.55828e-06, 7.911212e-06, 1.027579e-05, 8.025466e-06,
  1.264238e-06, 3.102749e-06, 8.178326e-06, 5.451958e-06, 2.950807e-06, 
    4.387794e-06, 5.549738e-06, 1.184509e-05, 2.517543e-05, 1.229561e-05, 
    2.432594e-06, 1.379068e-06, 2.385374e-06, 4.644525e-06, 7.096796e-06,
  2.015749e-06, 3.655816e-06, 7.885509e-06, 1.136597e-05, 1.390994e-06, 
    1.856393e-05, 5.475435e-06, 5.624239e-06, 1.251308e-05, 1.642579e-05, 
    1.833894e-05, 3.553182e-06, 1.687967e-06, 2.194496e-06, 1.757199e-06,
  6.368444e-06, 3.281579e-06, 2.646961e-06, 3.54251e-06, 1.160582e-05, 
    1.09131e-05, 1.421561e-05, 2.764959e-05, 2.849514e-05, 3.05765e-05, 
    2.186557e-05, 1.508993e-05, 1.653787e-05, 1.185592e-05, 2.6023e-06,
  1.304102e-05, 7.473309e-06, 4.334831e-06, 1.111309e-06, 1.763826e-06, 
    1.481214e-05, 1.815846e-05, 6.356001e-05, 8.232857e-05, 6.456337e-05, 
    1.501283e-05, 1.122942e-05, 2.395282e-05, 1.261854e-05, 3.396551e-05,
  4.009171e-06, 9.806599e-06, 9.666647e-06, 9.690059e-07, 2.656227e-06, 
    9.489011e-07, 3.357787e-06, 6.032612e-06, 4.639951e-06, 3.743855e-06, 
    3.584419e-06, 5.74525e-07, 8.915757e-08, 8.344293e-08, 3.827502e-08,
  6.039369e-06, 5.508863e-06, 3.665507e-06, 4.906934e-08, 5.695364e-07, 
    9.898624e-07, 4.477895e-06, 3.068983e-06, 2.389573e-06, 3.194488e-06, 
    3.872065e-06, 1.796651e-06, 4.00626e-07, 1.82043e-07, 5.644439e-07,
  3.40494e-06, 3.852376e-06, 1.056492e-06, 1.971294e-08, 1.966452e-08, 
    2.500273e-06, 2.962473e-06, 5.23816e-06, 4.582701e-06, 2.323325e-06, 
    3.791831e-06, 2.769184e-06, 6.880297e-07, 6.534174e-08, 3.509145e-07,
  3.071541e-06, 1.049517e-06, 2.966284e-07, 1.845691e-08, 7.133464e-09, 
    8.958586e-07, 1.656115e-06, 2.252903e-06, 4.857621e-06, 4.303567e-06, 
    3.157818e-06, 3.85309e-06, 1.658185e-06, 5.563778e-07, 4.936405e-07,
  1.205018e-06, 2.931662e-06, 5.587387e-07, 3.591816e-10, 2.958231e-09, 
    6.206193e-07, 3.559177e-06, 2.179421e-06, 5.449244e-06, 3.562691e-06, 
    4.840176e-06, 3.932882e-06, 4.114161e-06, 1.33165e-06, 1.714654e-07,
  1.280672e-07, 1.202845e-06, 1.771671e-06, 4.120843e-07, 6.581661e-10, 
    4.926872e-08, 9.078616e-07, 2.045376e-06, 1.932573e-06, 3.511281e-06, 
    2.760935e-06, 3.351648e-06, 4.327281e-06, 2.679267e-06, 1.939708e-06,
  5.388165e-08, 1.179875e-06, 3.253832e-06, 2.35119e-06, 1.546204e-07, 
    1.686082e-07, 8.377447e-07, 1.795496e-06, 3.434832e-06, 3.038543e-06, 
    2.013153e-06, 4.690069e-06, 3.150939e-06, 3.93817e-06, 3.837161e-06,
  1.287092e-09, 1.085598e-07, 2.941281e-06, 2.917262e-06, 1.290621e-09, 
    6.749918e-07, 1.320394e-06, 1.309033e-06, 1.278431e-06, 2.523653e-06, 
    3.628328e-06, 3.124803e-06, 3.026033e-06, 3.563763e-06, 3.374953e-06,
  2.776414e-11, 1.325679e-10, 6.07385e-10, 9.038712e-07, 2.182542e-06, 
    2.882176e-07, 2.4654e-06, 1.107659e-06, 1.468854e-06, 1.990431e-06, 
    3.299501e-06, 3.539408e-06, 3.404525e-06, 5.137686e-06, 5.408137e-06,
  1.318778e-10, 1.048353e-07, 4.83231e-07, 1.541472e-06, 4.426971e-07, 
    4.035533e-06, 4.01291e-06, 2.606048e-06, 2.042478e-06, 1.681518e-06, 
    1.865605e-06, 2.310831e-06, 3.482777e-06, 4.813765e-06, 3.779922e-06,
  9.948543e-07, 2.273288e-06, 4.3525e-06, 3.637069e-07, 4.318874e-07, 
    5.302738e-07, 2.651508e-06, 8.207637e-07, 6.716851e-07, 2.677668e-06, 
    5.13757e-06, 6.828604e-07, 4.662652e-06, 1.049981e-05, 9.869347e-06,
  1.935633e-06, 5.100721e-07, 2.431071e-06, 4.736398e-08, 4.250999e-08, 
    2.642528e-07, 2.839407e-06, 5.622639e-07, 6.549346e-08, 4.137257e-07, 
    1.874406e-06, 4.218352e-06, 2.537071e-06, 6.22228e-06, 3.534584e-06,
  5.970985e-07, 8.446554e-07, 1.572747e-07, 4.472981e-10, 3.055999e-09, 
    5.090184e-07, 1.316145e-06, 6.897484e-07, 8.660089e-07, 6.725943e-07, 
    5.579179e-07, 2.159036e-06, 1.65396e-07, 2.499515e-06, 2.109866e-07,
  2.557533e-06, 4.023539e-07, 2.81835e-09, 1.132633e-10, 1.006025e-09, 
    4.772739e-08, 8.09327e-07, 6.784333e-07, 9.309669e-07, 1.755591e-06, 
    2.499027e-07, 1.538988e-07, 4.870602e-07, 1.814828e-06, 1.705166e-06,
  1.023499e-06, 3.433242e-07, 2.715563e-09, 7.298034e-11, 1.097427e-10, 
    5.530754e-08, 4.58439e-07, 1.074607e-06, 8.423715e-07, 2.072953e-06, 
    1.995749e-06, 1.116464e-06, 8.694183e-07, 1.598664e-06, 4.189954e-06,
  1.112119e-06, 3.447134e-07, 7.220652e-08, 1.536971e-08, 3.980046e-11, 
    7.541221e-10, 4.016827e-07, 1.296869e-06, 1.574677e-06, 1.288904e-06, 
    2.42239e-06, 3.049023e-06, 1.5196e-06, 3.479196e-06, 4.913273e-06,
  9.588938e-07, 1.093992e-06, 1.001405e-06, 2.111284e-07, 3.043771e-10, 
    1.556182e-09, 4.581064e-07, 2.153439e-06, 2.750365e-06, 1.423164e-06, 
    1.99942e-06, 3.55135e-06, 2.796287e-06, 1.515509e-06, 5.81048e-06,
  2.230055e-08, 6.707697e-07, 4.74373e-07, 1.964876e-07, 6.646171e-08, 
    3.893166e-08, 1.874449e-06, 7.097768e-07, 3.086151e-06, 3.665173e-06, 
    1.739537e-06, 4.915932e-06, 5.536036e-06, 3.084039e-06, 5.709351e-06,
  7.29456e-07, 2.477996e-07, 5.410567e-08, 2.182172e-07, 3.061558e-07, 
    3.071267e-07, 4.054631e-06, 7.48232e-07, 2.36634e-06, 3.584828e-06, 
    2.383322e-06, 2.983914e-06, 4.822452e-06, 2.746614e-06, 3.663605e-06,
  2.279848e-06, 1.136174e-06, 1.713968e-06, 1.314183e-06, 4.222837e-07, 
    3.27262e-07, 7.34935e-07, 7.373555e-06, 2.393417e-06, 1.252834e-06, 
    1.008968e-06, 1.670893e-06, 2.138211e-06, 6.544522e-06, 3.62487e-06,
  1.676144e-09, 2.596261e-08, 1.092973e-06, 2.898953e-06, 5.786327e-06, 
    1.09546e-05, 1.684222e-05, 2.36808e-05, 2.723646e-05, 2.327188e-05, 
    2.94536e-05, 3.726589e-05, 4.951183e-05, 6.784807e-05, 8.112574e-05,
  6.791142e-06, 3.721793e-09, 6.144621e-09, 2.907204e-07, 2.534252e-06, 
    6.547739e-06, 1.269389e-05, 1.405321e-05, 1.396691e-05, 1.946383e-05, 
    2.289283e-05, 2.800771e-05, 4.098739e-05, 6.151081e-05, 8.027817e-05,
  2.953618e-06, 6.583841e-06, 5.122342e-09, 4.551654e-08, 1.867441e-06, 
    4.149081e-06, 9.143779e-06, 9.488734e-06, 1.370547e-05, 1.460064e-05, 
    1.616342e-05, 2.255915e-05, 3.545624e-05, 4.933372e-05, 7.065392e-05,
  1.586644e-07, 2.946625e-07, 3.580771e-09, 4.792037e-09, 5.689056e-08, 
    1.118896e-06, 2.827742e-06, 6.439186e-06, 6.727259e-06, 5.669251e-06, 
    7.579807e-06, 7.838968e-06, 1.249136e-05, 2.512564e-05, 3.777019e-05,
  7.788381e-09, 1.470911e-08, 1.709579e-09, 7.769181e-10, 2.726238e-09, 
    2.527889e-08, 3.972126e-07, 1.459105e-06, 3.884375e-06, 6.05704e-06, 
    7.862844e-06, 6.884753e-06, 8.444879e-06, 1.005912e-05, 1.235108e-05,
  2.541607e-09, 3.492635e-10, 2.221266e-09, 2.303319e-10, 2.055578e-10, 
    1.909497e-09, 1.004512e-08, 3.595005e-07, 1.014323e-06, 1.249325e-06, 
    8.945204e-06, 1.19197e-05, 9.119107e-06, 3.918909e-06, 5.497078e-06,
  3.801703e-10, 9.343091e-11, 9.931308e-11, 8.436806e-11, 3.250671e-13, 
    2.605179e-10, 1.798745e-08, 8.385724e-08, 1.767854e-06, 3.27618e-06, 
    5.629959e-06, 9.900285e-06, 1.352108e-05, 1.197872e-06, 6.21478e-06,
  3.929411e-15, 9.735247e-10, 4.256473e-13, 3.453128e-13, 8.604347e-13, 
    1.436325e-10, 2.528629e-07, 3.766348e-09, 6.185224e-07, 2.734543e-06, 
    6.530749e-06, 9.068599e-06, 6.802704e-06, 4.752713e-06, 8.11706e-06,
  1.533622e-16, 1.850922e-10, 5.660953e-13, 1.232607e-13, 2.429855e-15, 
    4.762648e-13, 1.111828e-09, 4.77489e-07, 1.641751e-07, 3.721877e-06, 
    5.843486e-06, 7.218424e-06, 9.979927e-06, 7.123952e-06, 4.842728e-06,
  1.059691e-16, 2.047422e-13, 6.406578e-13, 1.123737e-12, 2.621378e-14, 
    1.99567e-17, 3.867493e-10, 2.959456e-07, 1.139011e-06, 4.796141e-06, 
    6.927116e-06, 1.106962e-05, 1.222936e-05, 1.074093e-05, 7.840951e-06,
  1.489997e-06, 4.514135e-06, 4.383766e-06, 7.561296e-06, 1.006237e-05, 
    9.897686e-06, 5.937816e-06, 2.981258e-06, 1.655562e-06, 3.193614e-07, 
    1.157416e-07, 2.639831e-07, 7.030043e-07, 2.149132e-06, 5.183274e-06,
  1.547945e-05, 7.130677e-06, 6.138659e-06, 5.155791e-06, 7.434398e-06, 
    1.033244e-05, 1.20034e-05, 1.142774e-05, 9.749772e-06, 4.67367e-06, 
    1.756572e-06, 6.814393e-07, 7.27359e-07, 2.199485e-06, 2.532245e-06,
  2.211921e-05, 1.024001e-05, 5.176349e-06, 4.878523e-06, 7.951573e-06, 
    8.013243e-06, 1.250859e-05, 1.553329e-05, 1.327286e-05, 1.302304e-05, 
    9.737925e-06, 6.110822e-06, 3.119462e-06, 3.654696e-06, 3.919929e-06,
  1.156752e-05, 1.460176e-05, 3.119179e-06, 3.194504e-06, 4.393857e-06, 
    1.039848e-05, 9.763237e-06, 1.164886e-05, 1.43471e-05, 2.116091e-05, 
    1.606784e-05, 1.576657e-05, 1.398852e-05, 1.438191e-05, 1.180114e-05,
  7.55794e-06, 1.107404e-05, 1.264796e-05, 4.087851e-06, 3.001186e-06, 
    1.089699e-05, 8.572462e-06, 7.099963e-06, 1.094778e-05, 1.471477e-05, 
    1.819148e-05, 2.429387e-05, 2.390531e-05, 2.122348e-05, 2.708416e-05,
  1.457639e-06, 3.788425e-06, 9.30806e-06, 9.210639e-06, 3.947967e-06, 
    5.477115e-06, 7.482701e-06, 6.891586e-06, 7.462937e-06, 1.025255e-05, 
    1.458747e-05, 1.761824e-05, 2.284843e-05, 2.688562e-05, 2.978145e-05,
  4.055529e-08, 3.294214e-07, 4.515129e-06, 1.100651e-05, 1.489897e-05, 
    8.482762e-06, 7.205421e-06, 5.176179e-06, 1.005102e-05, 1.02455e-05, 
    1.024997e-05, 1.600806e-05, 2.681129e-05, 3.242578e-05, 3.135025e-05,
  1.383732e-09, 1.341618e-07, 9.853011e-07, 4.697494e-06, 6.900163e-06, 
    9.388275e-06, 7.412606e-06, 5.020026e-06, 3.743084e-06, 7.406257e-06, 
    1.792846e-05, 2.323962e-05, 2.342165e-05, 3.800554e-05, 4.010351e-05,
  3.735094e-09, 2.252424e-09, 1.4345e-07, 1.603319e-06, 5.248144e-06, 
    9.655661e-06, 1.334926e-05, 8.445571e-06, 4.862127e-06, 5.206624e-06, 
    1.094029e-05, 2.822217e-05, 3.098146e-05, 3.166883e-05, 3.466473e-05,
  6.521342e-09, 5.287478e-08, 5.577806e-08, 6.821915e-07, 1.499305e-06, 
    2.935705e-06, 8.879201e-06, 8.370478e-06, 8.403087e-06, 7.873669e-06, 
    1.28059e-05, 2.55955e-05, 1.870669e-05, 2.532968e-05, 3.903388e-05,
  2.224326e-07, 2.754562e-07, 6.26927e-07, 1.361353e-06, 2.578793e-06, 
    9.75999e-06, 1.198618e-05, 1.063307e-05, 1.007227e-05, 4.413481e-06, 
    2.158524e-06, 8.025085e-07, 6.695497e-07, 1.676605e-06, 3.57863e-06,
  1.090214e-05, 1.35485e-06, 3.179856e-06, 1.990087e-06, 7.878783e-06, 
    5.076785e-06, 1.046091e-05, 1.218567e-05, 9.022941e-06, 4.999923e-06, 
    2.954345e-06, 2.141571e-06, 1.649701e-06, 2.02057e-06, 3.117474e-06,
  9.561373e-06, 8.041168e-06, 1.826962e-06, 3.313448e-06, 1.108823e-05, 
    4.83708e-06, 8.129829e-06, 1.04664e-05, 8.918791e-06, 5.704865e-06, 
    4.79501e-06, 2.638907e-06, 1.954321e-06, 3.112616e-06, 3.708791e-06,
  7.215926e-06, 8.492488e-06, 3.485098e-06, 4.855267e-06, 9.090565e-06, 
    1.16901e-05, 6.689364e-06, 1.04508e-05, 8.267495e-06, 9.07459e-06, 
    7.076415e-06, 5.876586e-06, 5.135495e-06, 3.963633e-06, 5.207906e-06,
  8.329116e-06, 7.559709e-06, 9.689737e-06, 9.861029e-06, 8.680263e-06, 
    1.187814e-05, 7.836064e-06, 1.027201e-05, 1.071368e-05, 1.020764e-05, 
    8.06327e-06, 8.048747e-06, 6.435557e-06, 6.913132e-06, 6.49724e-06,
  4.300178e-06, 8.240974e-06, 1.214094e-05, 1.257479e-05, 8.568497e-06, 
    1.270012e-05, 7.865285e-06, 3.985177e-06, 1.102364e-05, 1.075385e-05, 
    6.922583e-06, 7.526353e-06, 8.189725e-06, 7.780694e-06, 9.794393e-06,
  8.367463e-07, 4.156944e-06, 1.615594e-05, 1.542207e-05, 1.111745e-05, 
    7.45322e-06, 1.716795e-05, 5.379796e-06, 9.991871e-06, 1.130289e-05, 
    9.735484e-06, 8.374888e-06, 9.506721e-06, 7.552828e-06, 9.273153e-06,
  2.548952e-07, 2.65809e-06, 1.703002e-05, 1.082212e-05, 7.565457e-06, 
    8.305437e-06, 1.677262e-05, 4.001614e-06, 5.029671e-06, 6.386656e-06, 
    1.051156e-05, 9.5945e-06, 8.484123e-06, 5.033181e-06, 5.032559e-06,
  2.853817e-07, 5.594394e-07, 4.271614e-06, 1.059367e-05, 1.371097e-05, 
    1.816486e-05, 8.575152e-06, 1.540146e-05, 1.868822e-06, 7.950309e-06, 
    8.692122e-06, 1.250191e-05, 1.174761e-05, 9.936452e-06, 5.343833e-06,
  4.871112e-08, 6.068311e-07, 2.187968e-06, 3.151701e-06, 5.578022e-06, 
    6.617618e-06, 2.823479e-05, 9.343465e-06, 1.513796e-05, 5.130151e-06, 
    6.470284e-06, 9.412156e-06, 1.126882e-05, 1.064961e-05, 1.113209e-05,
  0.0003064697, 0.0002088509, 0.000135624, 8.988516e-05, 7.258751e-05, 
    7.497791e-05, 7.495357e-05, 4.366304e-05, 1.300799e-05, 1.022704e-05, 
    1.247804e-05, 1.02898e-05, 4.888323e-06, 4.655041e-06, 1.827862e-06,
  0.0001911641, 0.0001003405, 6.850536e-05, 5.308726e-05, 5.571735e-05, 
    0.000158644, 0.0001816669, 2.480637e-05, 1.140992e-05, 1.045028e-05, 
    1.140218e-05, 1.044173e-05, 6.011885e-06, 3.647777e-06, 3.483888e-06,
  0.0001084426, 6.461777e-05, 6.116492e-05, 6.449082e-05, 7.339718e-05, 
    0.0002247779, 0.0001962022, 3.154086e-05, 1.535847e-05, 9.898683e-06, 
    1.063555e-05, 7.81136e-06, 5.138334e-06, 2.118853e-06, 3.06448e-06,
  7.181142e-05, 6.54526e-05, 6.513258e-05, 8.714068e-05, 0.0001795972, 
    0.0002167645, 0.0001182738, 3.83074e-05, 1.311706e-05, 1.14296e-05, 
    9.299862e-06, 8.237662e-06, 7.52323e-06, 3.701155e-06, 4.514338e-06,
  6.151692e-05, 6.313335e-05, 7.27351e-05, 0.0001167619, 0.0001395954, 
    0.0002926222, 9.70674e-05, 2.336553e-05, 1.643199e-05, 9.174551e-06, 
    9.546335e-06, 8.514796e-06, 9.0297e-06, 6.148945e-06, 5.008349e-06,
  5.319869e-05, 0.0001317409, 7.4009e-05, 7.690272e-05, 0.0001043427, 
    9.831778e-05, 2.512974e-05, 2.152647e-05, 1.129406e-05, 8.797697e-06, 
    6.810221e-06, 8.085669e-06, 9.078155e-06, 8.849725e-06, 5.915922e-06,
  5.847976e-05, 8.18471e-05, 0.0001063879, 9.63598e-05, 3.642982e-05, 
    8.668549e-06, 1.106996e-05, 1.490492e-05, 8.054642e-06, 8.411163e-06, 
    7.782442e-06, 1.322408e-05, 1.050748e-05, 6.516281e-06, 6.154158e-06,
  7.455658e-05, 8.175607e-05, 8.670423e-05, 2.295507e-05, 1.607579e-06, 
    3.253695e-06, 1.251801e-05, 5.568325e-06, 3.409844e-06, 6.044317e-06, 
    9.239899e-06, 7.80144e-06, 1.029424e-05, 8.677947e-06, 7.103016e-06,
  4.253919e-05, 3.703761e-05, 1.492875e-05, 3.385016e-08, 2.176878e-07, 
    1.010248e-07, 8.978638e-06, 2.591627e-06, 8.454449e-07, 4.423699e-06, 
    8.22231e-06, 9.027817e-06, 1.222104e-05, 8.086515e-06, 7.531174e-06,
  3.029267e-05, 1.200872e-05, 4.545442e-08, 1.280841e-07, 7.65446e-09, 
    4.907927e-07, 2.469055e-06, 8.743819e-06, 5.215532e-07, 1.568234e-06, 
    9.549024e-06, 7.783981e-06, 7.107313e-06, 9.525632e-06, 9.269425e-06,
  1.629743e-12, 7.024085e-12, 2.105014e-11, 2.866691e-12, 2.570702e-13, 
    1.141128e-06, 2.439813e-05, 6.248306e-05, 0.0001665842, 9.271129e-05, 
    0.0001006674, 0.0001011, 9.288952e-05, 8.304748e-05, 7.018029e-05,
  7.039654e-12, 9.96147e-13, 8.01266e-14, 6.110448e-12, 4.896266e-11, 
    1.428167e-06, 2.067811e-05, 0.000128837, 7.062248e-05, 0.0001730972, 
    9.683528e-05, 9.895842e-05, 0.0001039562, 6.833667e-05, 6.860923e-05,
  2.688218e-11, 1.256891e-10, 1.769708e-10, 4.272107e-11, 1.775255e-07, 
    5.607503e-07, 1.660956e-05, 0.0001721967, 0.0001654782, 0.0002019815, 
    0.0001053938, 0.0001493034, 7.868205e-05, 9.289248e-05, 8.758369e-05,
  2.29281e-12, 1.29891e-10, 4.805539e-08, 1.613838e-07, 4.904998e-07, 
    3.088454e-06, 3.534339e-05, 0.0002180096, 0.0002129539, 0.0001924149, 
    0.0001476663, 0.0001233005, 0.0001163625, 0.0001217166, 0.0001226431,
  3.191787e-10, 2.177259e-11, 1.695815e-07, 1.70304e-06, 7.787677e-07, 
    2.742596e-05, 9.176767e-05, 0.0001530353, 0.0001838691, 0.0001813083, 
    0.0002032343, 0.0001476487, 0.0001570999, 0.0001497824, 0.000135694,
  1.51203e-07, 1.107399e-07, 3.625444e-07, 1.673664e-06, 1.453975e-05, 
    6.077008e-05, 0.0001530856, 0.0002667466, 0.0002439389, 0.0001854344, 
    0.000219189, 0.0001911216, 0.0001832168, 0.0001655869, 0.0001303963,
  3.11472e-07, 8.141745e-07, 3.124923e-06, 1.309032e-05, 5.280007e-05, 
    9.867836e-05, 0.0001271462, 0.0001631858, 0.0001816985, 0.0002353936, 
    0.0002141117, 0.000225293, 0.0002010032, 0.0001799335, 0.0001320664,
  3.841987e-06, 9.603104e-06, 2.085999e-05, 5.215526e-05, 5.160238e-05, 
    7.025368e-05, 8.107371e-05, 0.0001066515, 0.0001467985, 0.0001888666, 
    0.0002051935, 0.0002184609, 0.0002576929, 0.0002124665, 0.0001672226,
  4.717106e-05, 5.685268e-05, 8.239004e-05, 5.380241e-05, 4.286907e-05, 
    3.472454e-05, 3.430037e-05, 3.641229e-05, 8.146677e-05, 0.0001045633, 
    0.0001630049, 0.0001494637, 0.0002570971, 0.0002419007, 0.0001597409,
  5.42762e-05, 4.687633e-05, 3.801281e-05, 3.608365e-05, 2.750378e-05, 
    3.025929e-05, 1.986882e-05, 1.797186e-05, 3.139587e-05, 6.97399e-05, 
    9.115991e-05, 0.0001296579, 0.0001709191, 0.0001499212, 0.0001449045,
  0.0001398458, 8.065227e-05, 3.620528e-05, 1.396783e-05, 4.577812e-06, 
    8.821408e-07, 5.837012e-07, 3.251051e-06, 3.403607e-06, 2.815451e-06, 
    2.688947e-06, 2.309265e-06, 2.419172e-06, 9.09076e-07, 6.237502e-07,
  9.378554e-05, 1.221862e-06, 7.685867e-07, 5.015163e-07, 6.041066e-07, 
    3.601632e-06, 4.201181e-06, 4.164201e-06, 3.509016e-06, 3.248757e-06, 
    2.557571e-06, 3.159759e-06, 4.261883e-06, 4.645288e-06, 2.160934e-06,
  4.908244e-05, 2.185146e-05, 3.418808e-07, 1.823685e-07, 1.199509e-06, 
    5.385726e-06, 2.930556e-06, 2.669428e-06, 2.456893e-06, 2.656725e-06, 
    3.351555e-06, 4.837859e-06, 5.415406e-06, 3.558668e-06, 3.310982e-06,
  4.296114e-05, 3.879897e-05, 1.219822e-07, 2.205186e-07, 1.010259e-06, 
    8.609789e-06, 9.218645e-06, 1.551262e-06, 2.500704e-06, 2.028729e-06, 
    7.26316e-07, 1.071976e-06, 4.369113e-06, 5.394821e-06, 4.395738e-06,
  2.842738e-05, 1.97509e-05, 1.485611e-08, 2.594259e-08, 5.39433e-07, 
    1.469221e-06, 3.254629e-06, 1.04228e-06, 1.999133e-06, 9.853773e-07, 
    9.495716e-07, 3.408002e-07, 3.036519e-07, 1.236509e-06, 3.61714e-06,
  1.454337e-05, 1.309174e-05, 1.185612e-05, 8.45121e-10, 4.938676e-07, 
    3.276291e-07, 4.714996e-06, 6.501516e-07, 6.297106e-07, 2.662654e-07, 
    4.297655e-08, 1.112706e-07, 7.259029e-08, 2.219662e-07, 1.031155e-06,
  4.335248e-06, 7.499951e-06, 9.409105e-06, 1.130617e-05, 2.648772e-08, 
    2.066268e-08, 7.013894e-07, 1.137239e-07, 2.708747e-07, 1.037984e-08, 
    1.559292e-07, 2.522673e-08, 7.867785e-09, 4.096492e-07, 3.337182e-07,
  6.565515e-07, 1.662259e-06, 3.666918e-06, 9.780545e-06, 5.302408e-08, 
    1.218239e-09, 8.076466e-07, 1.329207e-07, 3.010746e-07, 8.229277e-08, 
    2.051733e-08, 1.025173e-08, 1.318684e-08, 3.276801e-07, 1.171076e-07,
  8.946447e-07, 5.207455e-07, 1.047777e-06, 2.572649e-06, 7.867427e-06, 
    8.072409e-09, 4.294837e-07, 1.302319e-06, 2.013797e-07, 5.241678e-07, 
    1.014014e-08, 8.779382e-09, 4.656079e-09, 1.452349e-07, 3.822112e-07,
  6.239541e-07, 4.971791e-07, 9.604548e-09, 1.452138e-07, 3.136535e-08, 
    4.688045e-07, 4.411675e-09, 1.930754e-06, 9.4935e-07, 7.189339e-07, 
    7.382347e-08, 1.650195e-10, 3.113632e-09, 3.834695e-08, 3.271808e-07,
  0.0002035308, 0.0002249651, 0.0002524981, 0.0002482051, 0.0002635643, 
    0.0002676965, 0.0002644054, 0.0002628555, 0.0002798667, 0.0002131203, 
    0.0002280232, 0.0002020265, 0.0002044079, 0.0001928923, 0.000180897,
  0.0003008758, 0.000279963, 0.0002536839, 0.0002331524, 0.0002123725, 
    0.0002023948, 0.0001947022, 0.000206818, 0.0001729607, 0.0001780175, 
    0.0001762648, 0.0001738248, 0.0001534106, 0.0001505209, 0.0001387717,
  0.000489458, 0.0003692089, 0.0002288824, 0.0001745485, 0.0001532717, 
    0.0001393759, 0.000168532, 0.0001342711, 0.0001969565, 0.0001331945, 
    0.0001367532, 0.0001190344, 0.0001052304, 8.756966e-05, 7.543939e-05,
  0.0005393392, 0.0005103852, 0.0004080996, 0.0002861079, 0.0001789812, 
    0.0001352623, 9.305742e-05, 0.0001094691, 0.0001835976, 0.000134987, 
    0.0001098483, 0.0001035697, 8.255473e-05, 6.390813e-05, 5.173939e-05,
  0.0003702616, 0.0003296584, 0.0002623235, 0.0001947424, 0.000151982, 
    0.0001177184, 0.0001011935, 5.847148e-05, 7.653853e-05, 0.0001521215, 
    7.365453e-05, 7.763578e-05, 6.472921e-05, 5.050351e-05, 4.195466e-05,
  0.0001529757, 0.0001101162, 6.147574e-05, 4.903134e-05, 6.271155e-05, 
    5.827858e-05, 4.81083e-05, 4.083367e-05, 5.500857e-05, 5.077087e-05, 
    5.166847e-05, 6.522045e-05, 2.885261e-05, 2.98277e-05, 2.625206e-05,
  2.192259e-05, 1.345416e-05, 2.744263e-05, 2.737253e-05, 2.519567e-05, 
    2.07486e-05, 1.461622e-05, 1.923635e-05, 2.305527e-05, 1.212065e-05, 
    2.379703e-05, 2.058246e-05, 2.465329e-05, 1.593471e-05, 1.494443e-05,
  1.14961e-05, 1.380184e-05, 1.215449e-05, 4.012999e-05, 9.192801e-08, 
    6.759051e-07, 1.773479e-06, 2.773185e-06, 2.073538e-06, 4.101233e-06, 
    1.434712e-05, 1.685698e-05, 1.494588e-05, 1.466648e-06, 2.158961e-06,
  3.063302e-06, 3.147519e-06, 1.152013e-05, 2.807112e-05, 2.276501e-05, 
    2.230297e-08, 2.172944e-08, 3.21051e-08, 4.824532e-07, 2.087123e-06, 
    4.396797e-06, 1.303977e-05, 1.925858e-05, 1.603133e-06, 6.053795e-07,
  6.425328e-07, 2.072221e-06, 1.030536e-06, 5.916784e-07, 6.513118e-08, 
    4.561974e-07, 1.57983e-10, 8.893229e-10, 2.479227e-09, 9.403296e-07, 
    4.361195e-06, 1.343813e-05, 2.578588e-05, 2.183025e-05, 1.10945e-05,
  4.127835e-05, 5.660453e-05, 6.599343e-05, 7.675806e-05, 7.4178e-05, 
    7.052117e-05, 7.69929e-05, 8.763478e-05, 0.0001005478, 0.0001130026, 
    0.0001224536, 0.0001274835, 0.0001320317, 0.0001341219, 0.0001290819,
  7.749857e-05, 0.0001377915, 0.0001986359, 0.0002125205, 0.0002312296, 
    0.0002081301, 0.000183426, 0.0001661181, 0.0001503539, 0.000142083, 
    0.0001395798, 0.0001447804, 0.0001506115, 0.0001600415, 0.0001734856,
  0.0001089307, 0.0002226642, 0.0003342627, 0.0003748548, 0.000355847, 
    0.0002988627, 0.0002519482, 0.0002214681, 0.0002062343, 0.0002159595, 
    0.0002172451, 0.0002255568, 0.0002608154, 0.000326111, 0.0003793176,
  6.29731e-05, 0.0001726785, 0.000315213, 0.0004199132, 0.0004533841, 
    0.0005075387, 0.0004972015, 0.0004966025, 0.0004294915, 0.0003979295, 
    0.0004143892, 0.0003972295, 0.0004107127, 0.0004304734, 0.0004475363,
  5.107609e-05, 0.0001371478, 0.0002522569, 0.0003404447, 0.000439796, 
    0.0004890517, 0.0005608723, 0.0005050782, 0.0006301412, 0.0005512742, 
    0.0004764115, 0.0004786414, 0.0003587346, 0.0002730924, 0.0001714863,
  6.897152e-05, 0.0001362985, 0.0001747767, 0.0001550031, 0.0001615335, 
    0.0001888086, 0.0002163899, 0.0002251687, 0.000221465, 0.000203487, 
    0.0002454382, 0.0002684099, 0.0002343576, 0.0002272752, 0.0001963216,
  0.0002134282, 0.0002734207, 0.0002775378, 0.0002594691, 0.0002334123, 
    0.0002547111, 0.0002971619, 0.0003258119, 0.0003375916, 0.0003251897, 
    0.0003040679, 0.0002862739, 0.0002495203, 0.0002376594, 0.0002123686,
  0.0003024897, 0.0003994084, 0.0004160923, 0.0004207571, 0.0003904562, 
    0.0003916011, 0.0004135374, 0.0003947701, 0.0003959765, 0.0003653195, 
    0.0003285902, 0.0002685327, 0.0002284105, 0.0001880197, 0.0001246772,
  0.0002998832, 0.0003782023, 0.0003982851, 0.000404482, 0.0003947232, 
    0.0003399264, 0.0002869866, 0.0002714157, 0.0002520009, 0.0002337041, 
    0.0001912246, 0.0001600687, 0.0001578602, 9.139685e-05, 2.986753e-05,
  0.0001708631, 0.0002470832, 0.0002371181, 0.0002102701, 0.0001962296, 
    0.0001861584, 0.000133434, 0.0001170011, 0.0001127702, 0.0001014565, 
    7.907661e-05, 5.665245e-05, 3.416909e-05, 3.360447e-05, 8.079016e-06,
  0.0001078555, 0.0001308755, 6.541357e-05, 3.894544e-05, 4.801761e-05, 
    8.21517e-05, 0.0001290624, 0.0001276835, 9.53534e-05, 0.0001090076, 
    0.0001530324, 0.0001651624, 0.0001729283, 0.0001713936, 0.0001899976,
  1.035135e-05, 6.355774e-05, 0.0001032713, 6.450755e-05, 8.99434e-05, 
    9.664486e-05, 9.49568e-05, 0.0001069659, 8.681838e-05, 8.725721e-05, 
    9.082681e-05, 9.078361e-05, 9.442757e-05, 7.681162e-05, 0.000117667,
  1.763044e-06, 6.673088e-06, 4.773196e-05, 9.094206e-05, 0.0001137621, 
    8.723719e-05, 7.729633e-05, 7.75696e-05, 9.067527e-05, 7.563767e-05, 
    6.888328e-05, 5.901793e-05, 6.041975e-05, 6.382706e-05, 7.470912e-05,
  1.143662e-06, 1.507906e-06, 1.498255e-05, 5.059145e-05, 9.324839e-05, 
    9.642283e-05, 9.167971e-05, 9.274858e-05, 9.561512e-05, 7.660131e-05, 
    7.567032e-05, 6.896709e-05, 7.388461e-05, 7.343916e-05, 6.497763e-05,
  1.469273e-06, 2.539502e-06, 6.081851e-06, 3.941374e-05, 7.373067e-05, 
    9.017972e-05, 9.673629e-05, 8.883367e-05, 8.335819e-05, 8.492335e-05, 
    8.129352e-05, 0.0001004218, 0.0001158531, 0.0001073238, 8.73188e-05,
  4.310533e-07, 6.301393e-07, 2.04206e-06, 1.221287e-05, 4.411916e-05, 
    6.509903e-05, 8.231189e-05, 8.72488e-05, 0.0001022028, 9.805949e-05, 
    0.0001033344, 0.0001080856, 9.791205e-05, 9.007444e-05, 8.724368e-05,
  8.461924e-07, 3.86816e-07, 1.316663e-06, 1.555186e-06, 2.021694e-05, 
    4.95179e-05, 7.457077e-05, 8.856197e-05, 0.0001112915, 0.0001133328, 
    0.00010184, 9.490002e-05, 6.92683e-05, 6.550701e-05, 7.422312e-05,
  1.325119e-06, 4.889314e-07, 1.595868e-06, 3.467924e-06, 9.148013e-06, 
    3.425822e-05, 6.818354e-05, 7.608932e-05, 6.820755e-05, 6.639977e-05, 
    5.744795e-05, 6.400787e-05, 6.103714e-05, 6.904953e-05, 9.095034e-05,
  5.19206e-06, 6.670174e-06, 1.929644e-06, 1.413187e-05, 3.945417e-05, 
    6.180984e-05, 7.488317e-05, 7.565539e-05, 7.282395e-05, 7.802179e-05, 
    9.273062e-05, 9.940696e-05, 0.0001238608, 0.0001745434, 0.0002839374,
  5.622836e-06, 3.607791e-05, 8.482803e-05, 0.0001104397, 0.0001253466, 
    0.0001581117, 0.0001710805, 0.0001777387, 0.0001733577, 0.0001849924, 
    0.000193625, 0.0002381966, 0.0003069407, 0.0004277139, 0.0005455489,
  4.345548e-05, 3.466299e-05, 5.518058e-06, 9.750121e-06, 4.187342e-05, 
    6.499855e-05, 0.0001043737, 0.0001034431, 0.0001063229, 8.964108e-05, 
    0.0001019882, 0.0001034804, 7.622194e-05, 7.8676e-05, 7.547124e-05,
  2.112803e-06, 2.889423e-05, 2.18153e-05, 2.253242e-05, 4.8987e-05, 
    6.444997e-05, 0.0001014168, 0.0001248987, 0.0001100734, 9.503397e-05, 
    9.911044e-05, 0.000110642, 0.0001108119, 8.513354e-05, 7.849625e-05,
  2.323828e-07, 7.690062e-07, 3.806254e-05, 4.127889e-05, 5.458435e-05, 
    5.583374e-05, 5.564361e-05, 0.0001398112, 0.000103714, 0.0001156467, 
    9.92514e-05, 9.53983e-05, 9.473602e-05, 8.803332e-05, 7.725909e-05,
  4.995333e-08, 9.155418e-08, 1.283751e-05, 3.414298e-05, 6.885009e-05, 
    5.564161e-05, 5.175491e-05, 7.155329e-05, 9.646e-05, 0.0001391604, 
    9.642045e-05, 7.459176e-05, 7.54225e-05, 7.256043e-05, 7.321851e-05,
  1.097189e-08, 3.170086e-08, 3.832241e-06, 3.606018e-05, 7.587689e-05, 
    7.169547e-05, 5.421162e-05, 4.455166e-05, 8.155638e-05, 0.0001225237, 
    0.0001074785, 8.023906e-05, 6.971847e-05, 6.82099e-05, 7.214891e-05,
  3.88319e-13, 1.700287e-10, 4.153774e-09, 5.834809e-06, 7.582211e-05, 
    8.164351e-05, 6.430577e-05, 4.363333e-05, 5.799356e-05, 9.474307e-05, 
    0.0001060142, 9.620139e-05, 7.673597e-05, 6.38666e-05, 6.613538e-05,
  2.508353e-11, 5.001113e-12, 1.852354e-10, 7.781479e-10, 2.729406e-05, 
    8.451678e-05, 8.981008e-05, 6.362054e-05, 5.759391e-05, 6.392683e-05, 
    8.989449e-05, 9.959071e-05, 8.484477e-05, 6.726047e-05, 6.61555e-05,
  1.187675e-10, 9.190214e-11, 1.020075e-11, 1.263707e-10, 9.447981e-10, 
    5.34694e-05, 9.134682e-05, 8.744028e-05, 6.915547e-05, 6.077302e-05, 
    8.115102e-05, 8.421615e-05, 0.0001101452, 8.403889e-05, 6.450044e-05,
  4.861453e-10, 5.254597e-10, 5.983375e-11, 1.461721e-11, 1.496442e-10, 
    2.021567e-07, 6.727416e-05, 9.672296e-05, 8.708614e-05, 6.621555e-05, 
    5.992196e-05, 7.261759e-05, 8.695626e-05, 8.048538e-05, 6.242257e-05,
  3.912701e-10, 2.061221e-09, 1.080279e-09, 1.767754e-10, 1.802519e-11, 
    1.264245e-10, 1.027466e-05, 7.114772e-05, 9.762784e-05, 7.82469e-05, 
    5.876645e-05, 5.223864e-05, 6.492035e-05, 6.684764e-05, 6.759161e-05,
  2.61486e-06, 1.348975e-05, 5.273933e-06, 1.218965e-05, 5.262665e-05, 
    7.138996e-05, 8.698717e-05, 7.683667e-05, 0.000128911, 0.0001526739, 
    0.0002149796, 0.0002791083, 0.0001105839, 8.95158e-05, 4.806196e-05,
  7.272732e-08, 9.589675e-07, 7.606484e-06, 1.669682e-05, 5.767722e-05, 
    7.739067e-05, 8.672423e-05, 8.758928e-05, 8.725872e-05, 0.0001181983, 
    0.0001696048, 0.0001956703, 0.0002389916, 0.0001543069, 8.495509e-05,
  8.536865e-09, 4.813672e-09, 1.854589e-06, 1.9148e-05, 5.324574e-05, 
    5.999758e-05, 7.401522e-05, 8.360438e-05, 9.840191e-05, 0.0001036361, 
    0.0001150597, 0.0001453012, 0.0002107827, 0.0001901107, 0.0001448871,
  6.509322e-12, 1.200912e-10, 3.423454e-08, 2.163222e-06, 3.880512e-05, 
    6.372613e-05, 6.654237e-05, 7.612474e-05, 8.562514e-05, 9.215836e-05, 
    0.0001021887, 0.0001168126, 0.0001787743, 0.0001621035, 0.0001612365,
  3.416157e-14, 2.726096e-11, 2.403587e-09, 5.033482e-07, 1.512553e-05, 
    4.503752e-05, 6.420304e-05, 6.131008e-05, 6.877346e-05, 7.67785e-05, 
    9.061734e-05, 0.0001174717, 0.0001425242, 0.000160322, 0.0001571419,
  5.626644e-23, 4.534639e-12, 1.164059e-11, 8.772022e-10, 6.147284e-06, 
    3.109626e-05, 5.115776e-05, 5.754485e-05, 6.249973e-05, 5.937394e-05, 
    7.616053e-05, 9.182814e-05, 0.000114079, 0.0001293605, 0.0001393494,
  1.571262e-11, 6.328264e-13, 2.8233e-12, 3.043458e-12, 1.479883e-07, 
    1.277464e-05, 4.599459e-05, 5.520008e-05, 6.120954e-05, 5.674914e-05, 
    6.439246e-05, 7.007862e-05, 8.927299e-05, 0.0001009001, 0.0001020499,
  3.877962e-11, 5.886942e-11, 3.51755e-12, 1.818732e-13, 1.229695e-10, 
    3.311062e-06, 2.576685e-05, 4.695974e-05, 5.938935e-05, 6.050154e-05, 
    5.548259e-05, 5.744678e-05, 7.039158e-05, 8.489787e-05, 0.0001058648,
  1.41774e-10, 3.864246e-10, 9.681562e-11, 3.054798e-11, 1.570661e-13, 
    1.72339e-09, 9.220845e-06, 2.950278e-05, 4.692702e-05, 5.266331e-05, 
    5.687738e-05, 5.205369e-05, 5.739213e-05, 6.002577e-05, 7.54616e-05,
  2.672562e-12, 3.689987e-10, 7.552635e-10, 4.084117e-10, 4.329924e-11, 
    4.801036e-14, 1.649444e-06, 1.779365e-05, 4.275969e-05, 5.475364e-05, 
    5.667259e-05, 5.288848e-05, 5.294414e-05, 5.055507e-05, 5.751798e-05,
  2.335737e-05, 9.633674e-06, 3.225038e-09, 1.443846e-06, 1.08519e-05, 
    1.565468e-05, 1.76926e-05, 2.507967e-05, 4.28842e-05, 6.157783e-05, 
    9.564962e-05, 9.782146e-05, 4.070833e-05, 2.509785e-05, 2.870799e-05,
  2.336109e-06, 1.076511e-05, 2.808493e-06, 5.177749e-06, 1.548262e-05, 
    2.0752e-05, 1.931579e-05, 2.042211e-05, 1.782113e-05, 5.021593e-05, 
    9.390464e-05, 9.337613e-05, 8.385163e-05, 4.236702e-05, 2.868724e-05,
  3.559332e-07, 7.855783e-07, 4.666097e-06, 1.196749e-05, 2.377015e-05, 
    2.319203e-05, 2.369211e-05, 1.900903e-05, 2.745074e-05, 4.552848e-05, 
    6.216203e-05, 6.646873e-05, 9.668225e-05, 8.695632e-05, 5.065127e-05,
  8.959021e-08, 7.57586e-07, 2.589741e-06, 4.467905e-06, 2.485033e-05, 
    2.704388e-05, 2.451434e-05, 1.995117e-05, 2.403511e-05, 2.394748e-05, 
    3.154238e-05, 5.805869e-05, 6.406214e-05, 9.269505e-05, 9.857259e-05,
  6.064673e-10, 1.678556e-07, 4.931409e-08, 3.849447e-07, 2.035845e-05, 
    3.564384e-05, 2.904005e-05, 2.018768e-05, 2.574001e-05, 2.018837e-05, 
    2.609618e-05, 3.659545e-05, 5.350205e-05, 6.180178e-05, 8.191752e-05,
  9.050985e-14, 1.751854e-09, 1.367344e-08, 7.569383e-07, 1.047104e-05, 
    3.605965e-05, 3.475162e-05, 2.596412e-05, 2.63544e-05, 1.935572e-05, 
    2.787999e-05, 2.946622e-05, 3.808451e-05, 4.537408e-05, 6.407723e-05,
  1.426517e-22, 2.507317e-14, 1.151808e-10, 4.060537e-11, 2.647676e-06, 
    3.074831e-05, 3.941315e-05, 3.579546e-05, 3.200986e-05, 2.706952e-05, 
    2.510149e-05, 2.224158e-05, 2.834537e-05, 3.989058e-05, 4.64124e-05,
  2.629398e-22, 1.936644e-22, 8.412566e-14, 6.776523e-13, 5.600531e-11, 
    7.838382e-06, 3.455774e-05, 4.266714e-05, 3.667032e-05, 2.990765e-05, 
    2.460738e-05, 2.059807e-05, 2.260086e-05, 2.809882e-05, 3.5963e-05,
  1.700549e-22, 2.123453e-22, 3.223423e-16, 1.923117e-15, 5.351583e-12, 
    4.311385e-08, 1.606483e-05, 4.054926e-05, 3.466791e-05, 3.574819e-05, 
    3.203854e-05, 2.457658e-05, 2.644045e-05, 3.10816e-05, 2.676016e-05,
  1.931022e-22, 2.915675e-22, 2.346308e-22, 2.632253e-22, 4.504425e-14, 
    7.020006e-10, 3.153029e-07, 2.32786e-05, 4.704362e-05, 3.897394e-05, 
    3.769452e-05, 3.160568e-05, 3.00604e-05, 3.306823e-05, 3.277115e-05,
  3.51544e-06, 5.61461e-06, 9.283026e-09, 2.679484e-08, 9.641438e-06, 
    2.165827e-05, 2.325911e-05, 1.442101e-05, 1.226422e-05, 1.539471e-05, 
    2.538571e-05, 2.514609e-05, 1.151133e-05, 6.188198e-06, 8.732482e-06,
  1.995427e-07, 1.626282e-06, 1.188411e-08, 6.65621e-08, 6.959024e-06, 
    1.614849e-05, 1.904873e-05, 1.201349e-05, 9.123775e-06, 1.315179e-05, 
    2.048849e-05, 2.801555e-05, 2.181887e-05, 8.352212e-06, 7.234335e-06,
  1.541743e-08, 3.500342e-09, 5.133065e-07, 2.954049e-07, 7.500907e-06, 
    1.127153e-05, 1.158177e-05, 1.17963e-05, 9.023335e-06, 1.163384e-05, 
    1.276171e-05, 1.956273e-05, 2.096219e-05, 1.562929e-05, 7.733191e-06,
  7.156737e-10, 1.504864e-07, 4.054857e-07, 6.653669e-07, 4.328872e-06, 
    1.101413e-05, 1.159044e-05, 1.381154e-05, 1.266313e-05, 1.152549e-05, 
    9.603483e-06, 1.170123e-05, 1.243311e-05, 1.867303e-05, 1.581402e-05,
  2.416773e-11, 1.768771e-09, 1.267025e-06, 2.383515e-07, 1.203407e-06, 
    8.744601e-06, 1.262003e-05, 1.66533e-05, 1.696833e-05, 1.552469e-05, 
    1.245618e-05, 1.204962e-05, 1.224549e-05, 1.274376e-05, 1.908887e-05,
  5.172775e-11, 2.890643e-10, 8.952647e-09, 4.619692e-07, 1.703356e-06, 
    7.795978e-06, 1.287849e-05, 1.635013e-05, 1.967312e-05, 1.849632e-05, 
    1.595482e-05, 1.348573e-05, 1.320703e-05, 1.21334e-05, 1.352884e-05,
  4.107302e-11, 1.980524e-11, 2.392944e-09, 1.415387e-07, 1.924574e-06, 
    5.849813e-06, 1.287959e-05, 1.843778e-05, 1.884063e-05, 1.713606e-05, 
    1.397156e-05, 1.480245e-05, 1.239231e-05, 1.984741e-05, 3.041649e-05,
  1.915394e-10, 6.139945e-11, 1.940524e-10, 1.174392e-10, 1.107929e-07, 
    4.611329e-06, 1.094581e-05, 1.815707e-05, 2.076022e-05, 2.101062e-05, 
    1.674251e-05, 1.436427e-05, 1.101013e-05, 1.472738e-05, 1.561885e-05,
  4.816039e-10, 2.51445e-10, 1.496484e-10, 1.922111e-11, 1.596676e-12, 
    1.561975e-07, 7.22207e-06, 1.480851e-05, 2.35917e-05, 2.297109e-05, 
    1.869969e-05, 1.11367e-05, 1.019111e-05, 1.266086e-05, 1.251429e-05,
  3.406712e-09, 5.349074e-10, 3.937344e-10, 1.874371e-10, 8.294954e-11, 
    1.100672e-11, 1.611765e-07, 9.136756e-06, 2.057515e-05, 2.545111e-05, 
    2.071799e-05, 1.401046e-05, 1.105456e-05, 8.382625e-06, 7.095871e-06,
  2.321502e-06, 3.374104e-06, 4.254734e-07, 8.305751e-07, 1.587689e-05, 
    4.680305e-05, 3.882794e-05, 5.389149e-05, 7.476859e-05, 0.0001004492, 
    0.0001094755, 0.0001192, 0.0001011701, 9.042882e-05, 8.729212e-05,
  4.423356e-07, 3.054872e-06, 8.265619e-07, 1.807878e-07, 9.763561e-06, 
    2.567552e-05, 4.015998e-05, 4.729035e-05, 5.829973e-05, 7.277776e-05, 
    8.31932e-05, 0.0001167147, 0.0001069482, 9.156248e-05, 9.901547e-05,
  6.05781e-08, 2.388107e-07, 1.636033e-06, 1.951134e-06, 1.230187e-05, 
    1.508868e-05, 2.765066e-05, 3.913713e-05, 5.063e-05, 5.936869e-05, 
    6.657141e-05, 8.205795e-05, 9.582716e-05, 9.939439e-05, 9.992865e-05,
  7.151811e-08, 2.67398e-07, 5.407761e-07, 5.137433e-07, 2.404143e-06, 
    7.364803e-06, 1.862919e-05, 2.617128e-05, 3.305938e-05, 3.979098e-05, 
    4.685259e-05, 5.931349e-05, 6.482493e-05, 7.225958e-05, 8.862364e-05,
  6.236694e-09, 1.690285e-07, 5.580246e-07, 1.983451e-07, 1.442013e-07, 
    5.368233e-06, 1.215466e-05, 1.325318e-05, 1.751645e-05, 2.271836e-05, 
    3.176676e-05, 4.332679e-05, 5.24201e-05, 6.042697e-05, 6.322769e-05,
  2.58794e-09, 5.149779e-09, 2.050119e-07, 1.680019e-07, 3.678107e-08, 
    2.674527e-06, 5.74766e-06, 6.995607e-06, 1.024191e-05, 1.240411e-05, 
    1.892623e-05, 2.653014e-05, 3.772003e-05, 4.071695e-05, 6.3785e-05,
  1.110961e-08, 4.432052e-09, 5.586978e-08, 4.48879e-07, 3.281828e-07, 
    4.163854e-06, 4.056483e-06, 4.424028e-06, 7.146677e-06, 9.952792e-06, 
    1.278695e-05, 1.533161e-05, 2.111736e-05, 2.734849e-05, 3.391196e-05,
  7.19143e-08, 2.962939e-08, 9.112704e-09, 1.477942e-08, 7.868592e-07, 
    1.110358e-06, 1.345901e-06, 3.34383e-06, 4.340744e-06, 6.581091e-06, 
    9.542998e-06, 1.18906e-05, 1.389279e-05, 1.445678e-05, 1.520282e-05,
  1.042462e-07, 5.535051e-08, 5.010963e-08, 8.534454e-09, 2.613108e-09, 
    3.652322e-07, 4.085902e-07, 5.728556e-07, 1.386358e-06, 3.911151e-06, 
    6.87657e-06, 8.184908e-06, 9.068125e-06, 1.074535e-05, 1.061047e-05,
  1.029115e-06, 6.041011e-07, 6.64034e-08, 1.19889e-07, 4.431363e-08, 
    3.65696e-09, 3.990045e-10, 9.249024e-08, 1.508516e-06, 2.812107e-06, 
    4.682406e-06, 6.048197e-06, 7.747794e-06, 9.949908e-06, 1.235262e-05,
  6.641246e-09, 6.896527e-09, 8.462415e-08, 1.317328e-07, 5.604507e-07, 
    3.003404e-06, 1.496491e-05, 2.193753e-05, 3.164546e-05, 3.781695e-05, 
    4.565838e-05, 4.779606e-05, 3.318845e-05, 2.910682e-05, 3.307495e-05,
  7.554537e-08, 1.781525e-07, 2.635477e-08, 8.916777e-09, 6.426228e-07, 
    3.347846e-06, 7.272657e-06, 1.62439e-05, 2.129611e-05, 2.588064e-05, 
    3.253642e-05, 3.790504e-05, 3.793019e-05, 3.301606e-05, 3.460248e-05,
  1.453881e-07, 1.134984e-08, 3.885861e-07, 2.366839e-08, 1.870216e-06, 
    3.649008e-06, 5.329433e-06, 1.033997e-05, 1.640322e-05, 2.079458e-05, 
    2.125267e-05, 2.431746e-05, 2.621454e-05, 2.226783e-05, 1.91616e-05,
  4.059589e-08, 2.745908e-07, 8.089817e-07, 3.571048e-07, 1.594763e-06, 
    6.36491e-06, 1.015901e-05, 1.423264e-05, 2.504881e-05, 2.079547e-05, 
    2.141454e-05, 2.180518e-05, 2.261652e-05, 2.084293e-05, 1.86062e-05,
  9.656226e-08, 5.550576e-07, 2.78627e-07, 7.838689e-07, 2.330934e-07, 
    4.858381e-06, 8.891714e-06, 1.375274e-05, 2.191972e-05, 2.528395e-05, 
    2.609355e-05, 3.392524e-05, 3.820748e-05, 3.243805e-05, 2.736352e-05,
  3.270063e-07, 1.843424e-06, 4.253975e-07, 1.949916e-06, 8.722452e-07, 
    1.43157e-06, 5.530494e-06, 1.018388e-05, 1.751955e-05, 2.053866e-05, 
    2.619182e-05, 3.360838e-05, 3.865816e-05, 3.808568e-05, 3.98296e-05,
  6.553211e-07, 2.037486e-06, 3.77634e-06, 2.097042e-06, 3.049733e-06, 
    6.515988e-06, 5.974476e-06, 7.66808e-06, 1.077799e-05, 1.265639e-05, 
    1.780498e-05, 2.49138e-05, 3.102062e-05, 4.079908e-05, 4.763422e-05,
  1.324866e-07, 7.898831e-07, 1.8672e-06, 3.207532e-06, 6.641883e-06, 
    8.334039e-06, 7.921604e-06, 6.893379e-06, 8.82366e-06, 1.242471e-05, 
    1.662331e-05, 1.986668e-05, 2.510044e-05, 3.111358e-05, 3.951107e-05,
  1.967001e-06, 4.574415e-06, 8.609926e-07, 1.594905e-06, 4.01323e-06, 
    4.366447e-06, 7.922635e-06, 9.745623e-06, 9.260022e-06, 1.005478e-05, 
    1.323374e-05, 1.531167e-05, 2.157724e-05, 2.458317e-05, 3.079391e-05,
  1.497759e-06, 4.521922e-06, 9.198184e-06, 1.230712e-05, 9.84328e-06, 
    4.911598e-06, 9.263853e-06, 1.180748e-05, 8.681042e-06, 8.349571e-06, 
    9.671909e-06, 1.192262e-05, 1.580363e-05, 2.105225e-05, 2.264173e-05,
  1.35333e-06, 8.966848e-07, 4.519037e-07, 2.901429e-07, 1.106119e-06, 
    5.940603e-06, 1.200653e-05, 3.387395e-05, 4.623068e-05, 5.234963e-05, 
    5.989429e-05, 5.324331e-05, 3.701323e-05, 3.208299e-05, 2.675591e-05,
  7.808922e-07, 1.265518e-06, 2.429437e-06, 1.327891e-06, 2.300684e-06, 
    3.251075e-06, 2.938774e-06, 1.184581e-05, 2.727574e-05, 3.740377e-05, 
    5.372737e-05, 5.804809e-05, 6.116747e-05, 4.840294e-05, 4.726387e-05,
  1.119006e-06, 4.988115e-07, 2.945954e-06, 2.162928e-06, 7.336376e-06, 
    3.159056e-06, 3.951955e-06, 6.134143e-06, 2.025823e-05, 2.745819e-05, 
    3.080461e-05, 3.795886e-05, 4.296681e-05, 5.761276e-05, 4.33712e-05,
  1.151785e-06, 2.553868e-07, 1.820881e-06, 2.438109e-06, 7.961548e-06, 
    9.218847e-06, 7.441474e-06, 6.907111e-06, 1.236783e-05, 2.306849e-05, 
    2.623626e-05, 2.915099e-05, 2.57255e-05, 2.43559e-05, 3.557906e-05,
  1.068224e-06, 1.843734e-06, 1.15325e-06, 1.396599e-06, 5.431976e-06, 
    8.784215e-06, 1.247368e-05, 8.813756e-06, 1.445963e-05, 2.008985e-05, 
    2.585729e-05, 2.913357e-05, 3.078105e-05, 3.320468e-05, 3.052891e-05,
  3.196801e-07, 1.622967e-07, 7.793558e-07, 1.484667e-07, 8.435414e-07, 
    1.815117e-06, 1.450008e-05, 1.316735e-05, 1.275186e-05, 1.960602e-05, 
    2.082555e-05, 2.865522e-05, 3.355608e-05, 3.243479e-05, 3.115626e-05,
  2.167267e-06, 1.35005e-07, 2.040128e-08, 6.313361e-08, 5.645891e-08, 
    1.164036e-06, 7.032823e-06, 1.206742e-05, 1.602189e-05, 1.768983e-05, 
    1.472121e-05, 2.355816e-05, 2.679004e-05, 3.132396e-05, 3.239428e-05,
  6.067724e-07, 2.891521e-06, 1.288338e-06, 2.594085e-07, 7.460199e-09, 
    1.58607e-06, 2.913303e-06, 5.531154e-06, 1.11982e-05, 1.513877e-05, 
    1.357262e-05, 1.992279e-05, 2.413602e-05, 2.916593e-05, 3.38948e-05,
  5.031825e-06, 1.876426e-06, 8.020926e-07, 1.374762e-06, 2.937221e-07, 
    2.502283e-06, 1.576143e-06, 3.750571e-06, 6.256692e-06, 1.101837e-05, 
    1.13365e-05, 1.302168e-05, 1.904484e-05, 2.285239e-05, 2.736371e-05,
  6.807256e-07, 2.328841e-07, 3.003661e-06, 3.279037e-06, 4.810332e-06, 
    4.721857e-06, 6.028542e-06, 7.649932e-06, 6.892902e-06, 8.401616e-06, 
    7.44517e-06, 9.146269e-06, 1.338498e-05, 1.716268e-05, 2.200727e-05,
  1.674318e-06, 3.88232e-06, 9.72088e-08, 1.598723e-06, 2.584946e-05, 
    3.836134e-05, 3.400595e-05, 3.29261e-05, 1.950543e-05, 1.081007e-05, 
    1.358606e-05, 1.580182e-05, 1.277192e-05, 1.460076e-05, 1.356539e-05,
  5.893498e-07, 3.866996e-07, 1.02747e-06, 5.705235e-07, 2.016276e-05, 
    3.257993e-05, 3.996747e-05, 3.460035e-05, 3.42283e-05, 2.998546e-05, 
    3.003808e-05, 1.737031e-05, 1.353772e-05, 1.264182e-05, 1.031101e-05,
  1.822705e-07, 7.932491e-07, 1.737973e-06, 1.472441e-06, 1.818519e-05, 
    2.467568e-05, 3.010772e-05, 3.909431e-05, 4.316582e-05, 3.841384e-05, 
    4.475713e-05, 4.453251e-05, 4.500174e-05, 2.526134e-05, 1.831573e-05,
  2.324612e-07, 6.110797e-07, 1.610987e-06, 2.620625e-06, 9.700711e-06, 
    1.872509e-05, 2.288071e-05, 2.955895e-05, 3.824437e-05, 3.766614e-05, 
    3.669243e-05, 4.632769e-05, 5.2658e-05, 6.335331e-05, 4.307195e-05,
  2.058345e-07, 4.215399e-07, 1.124957e-06, 4.064856e-06, 6.29996e-06, 
    1.198211e-05, 1.771586e-05, 1.969346e-05, 2.719912e-05, 3.111563e-05, 
    3.546877e-05, 3.814023e-05, 4.100605e-05, 4.915628e-05, 5.342599e-05,
  6.189224e-08, 9.56793e-08, 2.81834e-07, 9.036037e-07, 2.446626e-06, 
    7.434713e-06, 1.35603e-05, 1.418375e-05, 1.890573e-05, 2.253078e-05, 
    2.693087e-05, 3.081347e-05, 3.345029e-05, 3.646147e-05, 3.930684e-05,
  2.240083e-08, 3.700908e-08, 4.075241e-08, 2.754503e-08, 2.052076e-06, 
    3.399445e-06, 1.193918e-05, 1.318056e-05, 1.327174e-05, 1.714527e-05, 
    2.043479e-05, 2.124939e-05, 2.337606e-05, 2.982266e-05, 3.165258e-05,
  1.516891e-10, 1.892842e-08, 4.539459e-10, 1.106327e-08, 1.588441e-07, 
    4.275728e-07, 8.449137e-06, 1.270446e-05, 9.402032e-06, 1.145953e-05, 
    1.398308e-05, 1.700587e-05, 1.977541e-05, 2.202175e-05, 2.659988e-05,
  1.150227e-08, 1.219241e-08, 1.761807e-08, 3.587141e-10, 1.142201e-06, 
    6.249043e-08, 3.313543e-06, 3.927581e-06, 6.244445e-06, 6.257247e-06, 
    1.227012e-05, 1.000384e-05, 1.347374e-05, 1.774468e-05, 1.642654e-05,
  5.367911e-08, 7.356439e-08, 5.171343e-09, 8.981897e-09, 4.949937e-09, 
    1.438269e-08, 8.115679e-07, 3.207586e-06, 1.818093e-06, 4.58959e-06, 
    6.828816e-06, 1.335772e-05, 7.855624e-06, 1.002676e-05, 1.335774e-05,
  9.211347e-08, 5.416429e-08, 7.193189e-08, 3.055962e-07, 9.980722e-06, 
    1.806962e-05, 1.354266e-05, 2.791332e-05, 3.474539e-05, 3.424969e-05, 
    3.493888e-05, 3.793436e-05, 3.205035e-05, 2.944058e-05, 3.192246e-05,
  1.983947e-07, 2.24966e-07, 3.672884e-08, 7.838499e-08, 7.150487e-06, 
    1.100946e-05, 1.17212e-05, 2.13779e-05, 2.82296e-05, 3.251066e-05, 
    3.814117e-05, 4.007503e-05, 3.31991e-05, 2.984847e-05, 3.255821e-05,
  4.614712e-09, 4.242886e-08, 6.616657e-09, 5.738028e-09, 7.799824e-06, 
    1.318038e-05, 1.501133e-05, 1.507561e-05, 2.263785e-05, 2.760582e-05, 
    3.383191e-05, 3.866859e-05, 4.863284e-05, 4.386532e-05, 3.522333e-05,
  5.593816e-09, 2.432892e-09, 1.115754e-08, 2.76891e-08, 4.901284e-06, 
    9.342442e-06, 9.397671e-06, 1.276276e-05, 1.502625e-05, 1.969943e-05, 
    2.314482e-05, 2.637629e-05, 3.465973e-05, 3.885714e-05, 4.519189e-05,
  1.270909e-08, 1.528067e-08, 1.218051e-09, 9.90924e-10, 2.251609e-07, 
    3.57729e-06, 1.099257e-05, 1.047833e-05, 1.255245e-05, 1.388545e-05, 
    1.692078e-05, 2.129645e-05, 2.48644e-05, 2.892745e-05, 3.876888e-05,
  4.734819e-10, 1.685705e-09, 1.538752e-08, 2.824229e-09, 4.776427e-08, 
    1.222047e-06, 5.310194e-06, 9.823435e-06, 8.9225e-06, 1.087464e-05, 
    1.467229e-05, 1.321726e-05, 2.19518e-05, 2.603777e-05, 3.054761e-05,
  5.78075e-10, 3.105303e-10, 1.261554e-10, 2.246928e-10, 2.833116e-07, 
    1.450076e-06, 4.085204e-06, 7.763902e-06, 1.218221e-05, 8.882685e-06, 
    1.086821e-05, 1.489719e-05, 1.666555e-05, 1.778637e-05, 2.07534e-05,
  4.316235e-10, 9.619611e-10, 3.381088e-10, 5.573634e-12, 2.318619e-09, 
    4.781061e-07, 1.855133e-07, 5.383183e-06, 1.174928e-05, 1.391902e-05, 
    8.954229e-06, 1.185872e-05, 1.316102e-05, 1.445912e-05, 1.624417e-05,
  3.641747e-11, 1.879693e-08, 4.67319e-10, 7.774505e-11, 3.414356e-11, 
    8.112272e-09, 5.817539e-09, 1.090431e-06, 1.410437e-06, 7.987763e-06, 
    9.246491e-06, 9.753003e-06, 1.193759e-05, 1.303817e-05, 1.450345e-05,
  1.41858e-09, 6.131801e-08, 2.134742e-08, 1.725731e-09, 3.013035e-10, 
    2.706237e-11, 2.716771e-09, 1.346851e-07, 5.357504e-07, 1.496215e-06, 
    1.493871e-06, 7.590049e-06, 1.119056e-05, 9.817754e-06, 1.442846e-05,
  8.863674e-13, 7.470014e-11, 2.837711e-09, 1.330291e-11, 6.278086e-17, 
    1.584087e-09, 1.728898e-08, 1.035845e-07, 4.401236e-07, 5.032235e-07, 
    1.03349e-06, 2.21208e-06, 2.361674e-06, 3.025077e-06, 2.542036e-06,
  3.126075e-09, 1.426466e-10, 8.852863e-09, 7.17708e-09, 7.691207e-12, 
    6.851914e-12, 7.010555e-09, 1.153219e-07, 2.759596e-07, 6.404883e-07, 
    1.147704e-06, 1.617347e-06, 4.047641e-06, 3.405984e-06, 3.077338e-06,
  3.18741e-09, 1.521772e-07, 9.633055e-08, 3.096602e-08, 4.522386e-08, 
    4.444539e-10, 1.036863e-10, 2.619269e-08, 1.658904e-07, 4.394853e-07, 
    8.650936e-07, 1.293562e-06, 2.464369e-06, 3.93786e-06, 4.257693e-06,
  1.300515e-08, 1.687716e-09, 2.331062e-07, 1.391748e-07, 2.421941e-07, 
    1.27283e-08, 2.56038e-08, 1.631177e-08, 3.880814e-08, 2.727874e-07, 
    2.482303e-07, 8.417681e-07, 1.475965e-06, 2.367242e-06, 3.883722e-06,
  4.056074e-07, 1.597445e-08, 6.78458e-08, 2.278761e-07, 1.818746e-07, 
    5.070112e-08, 1.704952e-07, 1.159698e-09, 8.965092e-09, 5.242153e-08, 
    3.743816e-07, 5.263591e-07, 1.345606e-06, 2.17042e-06, 4.433256e-06,
  9.907969e-07, 5.855803e-07, 3.003942e-08, 1.501943e-07, 4.797317e-07, 
    7.321934e-07, 3.358828e-07, 2.017302e-07, 2.913566e-09, 1.633868e-07, 
    2.438777e-07, 5.184079e-07, 9.854516e-07, 2.078864e-06, 3.47757e-06,
  8.341643e-07, 5.866945e-07, 6.173159e-07, 5.330236e-08, 1.020487e-07, 
    9.293859e-07, 7.383168e-07, 4.545974e-07, 8.277664e-07, 1.768345e-07, 
    2.552493e-07, 4.094436e-07, 4.678433e-07, 1.156646e-06, 1.955269e-06,
  2.569503e-08, 2.621264e-07, 6.43772e-07, 4.722805e-07, 2.286553e-07, 
    9.930957e-07, 1.944485e-06, 2.789071e-06, 1.347697e-06, 3.664016e-07, 
    4.576072e-07, 4.737388e-07, 4.440248e-07, 6.827715e-07, 1.282408e-06,
  8.455842e-11, 1.845546e-08, 4.428555e-07, 3.514282e-07, 3.582292e-07, 
    8.937417e-07, 5.698449e-07, 4.479914e-06, 9.557104e-07, 9.692791e-07, 
    6.339706e-07, 7.887385e-07, 6.646695e-07, 4.603946e-07, 4.922562e-07,
  2.276661e-12, 7.2807e-08, 1.588664e-07, 1.769199e-07, 1.442765e-07, 
    4.980592e-07, 4.484203e-07, 1.011878e-06, 1.893859e-06, 1.085924e-06, 
    5.595556e-07, 1.054469e-06, 9.944637e-07, 1.056162e-06, 7.886104e-07,
  6.441658e-08, 1.128905e-08, 7.026704e-09, 2.262604e-07, 2.417719e-08, 
    2.614937e-07, 2.605604e-06, 5.487806e-06, 1.037845e-05, 9.328257e-06, 
    7.013181e-06, 1.396572e-05, 9.728733e-07, 2.928208e-06, 4.124292e-06,
  1.049604e-06, 5.496924e-09, 1.026755e-08, 3.278686e-07, 1.807619e-07, 
    1.417297e-08, 2.717574e-06, 1.080926e-05, 8.634706e-06, 6.47856e-06, 
    5.695846e-06, 6.590713e-06, 1.842302e-06, 1.195966e-06, 3.13857e-06,
  1.147378e-06, 2.978053e-07, 1.030205e-08, 1.051914e-07, 1.503726e-07, 
    2.217283e-08, 1.529098e-06, 9.707835e-06, 8.623801e-06, 5.601876e-06, 
    5.585684e-06, 5.718806e-06, 3.966936e-06, 1.806912e-06, 5.914923e-07,
  7.866994e-07, 1.593802e-08, 2.017549e-09, 7.372043e-09, 3.330492e-09, 
    6.97063e-08, 2.477176e-06, 9.00442e-06, 9.73881e-06, 4.633134e-06, 
    3.0282e-06, 1.21161e-06, 5.009726e-07, 4.700584e-07, 5.04807e-07,
  1.129047e-06, 1.056799e-09, 1.555919e-09, 6.903459e-09, 7.218556e-09, 
    2.777831e-09, 9.155436e-07, 5.094347e-06, 6.245655e-06, 3.129379e-06, 
    1.566126e-06, 9.340756e-07, 2.159628e-07, 1.221207e-06, 1.200093e-06,
  4.802944e-07, 3.69186e-10, 1.207802e-10, 2.530486e-09, 5.310238e-10, 
    5.742047e-09, 7.024152e-07, 2.409781e-06, 3.851548e-06, 2.14593e-06, 
    1.757034e-06, 1.125441e-06, 9.298931e-07, 1.891986e-06, 1.66286e-06,
  7.92821e-07, 2.576131e-07, 1.87628e-10, 4.513573e-11, 2.885373e-10, 
    1.157566e-08, 1.562015e-06, 2.491448e-06, 3.205023e-06, 4.199701e-06, 
    1.733127e-06, 1.075642e-06, 7.709747e-07, 1.803236e-06, 1.683035e-06,
  4.733113e-08, 8.901119e-10, 8.031551e-11, 1.078853e-11, 4.770297e-10, 
    1.649828e-08, 1.180622e-06, 2.58182e-06, 2.310901e-06, 2.343856e-06, 
    1.78035e-06, 3.536098e-07, 4.171957e-07, 1.215267e-06, 1.288355e-06,
  1.33496e-10, 1.793547e-12, 2.871221e-18, 1.289753e-12, 1.155693e-09, 
    2.474699e-08, 7.781782e-07, 2.74944e-06, 1.49589e-06, 1.52294e-06, 
    1.005895e-06, 3.728839e-08, 2.460639e-07, 3.761612e-07, 3.549125e-07,
  1.119719e-07, 3.535933e-12, 4.07148e-15, 2.153651e-14, 2.269595e-13, 
    1.166181e-10, 1.295968e-08, 6.242113e-06, 2.318173e-06, 2.701284e-06, 
    9.174553e-07, 1.159899e-07, 2.563551e-07, 5.449957e-07, 2.031773e-07,
  2.090288e-06, 3.911854e-06, 5.057042e-06, 6.96325e-06, 9.745887e-06, 
    1.731129e-05, 6.291982e-05, 3.247053e-05, 5.616517e-05, 3.694466e-05, 
    3.902128e-05, 4.780755e-05, 4.248351e-05, 5.806254e-05, 7.166033e-05,
  7.424795e-06, 1.184759e-06, 2.057416e-06, 3.285972e-06, 4.358604e-06, 
    5.946875e-06, 2.124355e-05, 1.653234e-05, 1.893977e-05, 1.035947e-05, 
    1.219451e-05, 1.872564e-05, 7.900527e-06, 1.455184e-05, 1.785774e-05,
  4.137189e-06, 1.900806e-06, 1.246707e-07, 6.35106e-08, 7.552229e-08, 
    4.0235e-07, 2.344726e-06, 2.811889e-06, 2.406727e-06, 2.539413e-06, 
    2.277955e-06, 3.123563e-06, 4.185567e-06, 4.184846e-06, 1.897877e-06,
  3.095079e-06, 3.292218e-07, 1.386337e-08, 8.913215e-07, 1.16178e-06, 
    1.402992e-06, 7.209121e-07, 1.343054e-06, 2.945837e-06, 1.009957e-06, 
    7.950325e-07, 5.189755e-07, 1.441986e-07, 6.254473e-07, 5.815398e-07,
  8.695387e-07, 2.253953e-08, 3.847775e-08, 7.54036e-06, 9.43094e-06, 
    3.833322e-06, 6.401362e-07, 1.405311e-06, 4.563985e-07, 3.852824e-07, 
    1.334904e-06, 6.246628e-07, 3.294135e-07, 6.024888e-08, 2.408999e-07,
  2.043011e-06, 2.873173e-07, 1.85339e-06, 1.580535e-05, 1.034618e-05, 
    2.395319e-06, 1.036597e-07, 9.455176e-07, 5.527255e-07, 6.877095e-07, 
    1.283616e-06, 9.324173e-07, 1.733305e-06, 9.345125e-07, 3.153005e-07,
  1.606888e-06, 3.218637e-06, 5.146676e-06, 1.489755e-05, 5.694524e-06, 
    9.362474e-07, 4.050833e-08, 1.37703e-06, 5.998423e-07, 6.642161e-07, 
    2.084638e-06, 1.871239e-06, 1.112792e-06, 1.712794e-06, 1.614366e-06,
  2.371777e-06, 3.688542e-06, 1.046707e-05, 1.161632e-05, 2.683682e-06, 
    5.619635e-09, 8.34067e-09, 1.613391e-06, 8.260898e-07, 2.720004e-06, 
    4.267037e-06, 2.220902e-06, 1.614792e-06, 1.606968e-06, 3.366271e-06,
  1.111262e-06, 2.150602e-06, 2.076492e-06, 7.6662e-07, 6.919848e-09, 
    4.012887e-10, 2.475022e-09, 1.283052e-06, 1.714374e-06, 2.691535e-06, 
    5.046475e-06, 2.685071e-06, 2.484965e-06, 2.380801e-06, 2.956263e-06,
  8.756174e-08, 1.153959e-08, 4.734529e-09, 2.304431e-09, 9.549181e-09, 
    3.773715e-09, 1.44089e-09, 1.538909e-06, 1.204589e-06, 1.801325e-06, 
    3.671717e-06, 2.137609e-06, 4.973802e-06, 3.753523e-06, 2.90871e-06,
  1.559307e-11, 1.46846e-12, 4.957084e-10, 1.515682e-08, 2.553562e-07, 
    4.610324e-06, 2.198709e-05, 2.405198e-05, 3.441027e-05, 3.294256e-05, 
    2.242614e-05, 2.528673e-05, 1.894947e-05, 1.526907e-05, 7.950344e-06,
  8.599289e-09, 1.729801e-09, 1.309077e-08, 3.864857e-08, 6.097681e-08, 
    1.128631e-06, 3.41962e-05, 2.265777e-05, 3.341006e-05, 3.25334e-05, 
    3.915343e-05, 3.379742e-05, 1.82568e-05, 1.663064e-05, 1.259649e-05,
  2.063118e-06, 5.414391e-06, 4.154433e-07, 1.999304e-07, 1.183385e-07, 
    6.344061e-06, 2.69738e-05, 5.096265e-05, 2.439933e-05, 4.807676e-05, 
    2.887332e-05, 3.0197e-05, 2.686561e-05, 2.51068e-05, 2.28068e-05,
  3.385991e-06, 3.716466e-06, 1.539793e-06, 1.710942e-06, 1.703019e-06, 
    4.834872e-06, 2.8009e-05, 4.401921e-05, 3.846867e-05, 4.705253e-05, 
    3.920747e-05, 3.417295e-05, 4.090603e-05, 4.393969e-05, 4.950542e-05,
  5.78515e-06, 8.479323e-06, 2.921579e-06, 2.027044e-06, 2.388281e-06, 
    3.943397e-06, 2.082272e-05, 3.550642e-05, 3.580004e-05, 6.031895e-05, 
    5.071746e-05, 4.306811e-05, 4.556035e-05, 6.040505e-05, 6.912144e-05,
  1.024878e-05, 9.887772e-06, 2.513564e-06, 7.106193e-08, 2.169972e-07, 
    3.287063e-06, 1.136985e-05, 2.683286e-05, 5.17521e-05, 3.958199e-05, 
    7.484339e-05, 5.720378e-05, 5.037125e-05, 6.023082e-05, 6.477726e-05,
  1.955759e-05, 1.504972e-05, 1.033748e-05, 2.01635e-06, 1.043787e-07, 
    2.26218e-06, 1.046268e-05, 5.128865e-05, 3.494718e-05, 4.582345e-05, 
    3.728595e-05, 0.0001044813, 4.014993e-05, 3.717862e-05, 4.206819e-05,
  6.933216e-05, 4.599166e-05, 1.782167e-05, 8.887343e-06, 2.753378e-06, 
    5.706868e-06, 2.049669e-05, 1.750623e-05, 1.840228e-05, 5.583584e-05, 
    1.376294e-05, 1.903049e-05, 3.224577e-05, 2.222363e-05, 2.652057e-05,
  8.78846e-05, 9.979967e-05, 8.179369e-05, 6.656769e-05, 2.84068e-05, 
    8.812743e-06, 3.693295e-06, 2.179379e-06, 4.566069e-06, 6.545906e-06, 
    5.615807e-06, 1.148567e-05, 7.585193e-06, 1.198125e-05, 9.074955e-06,
  2.515477e-05, 3.174255e-05, 2.675693e-05, 2.050694e-05, 2.237444e-05, 
    2.378519e-05, 6.802817e-06, 3.826817e-06, 2.452961e-06, 1.708659e-06, 
    2.408587e-06, 1.150723e-05, 2.543862e-05, 5.164791e-05, 2.689206e-05,
  1.478644e-08, 2.403175e-08, 2.410649e-08, 3.668728e-08, 6.96498e-08, 
    6.906016e-08, 6.334801e-09, 1.211194e-06, 2.502653e-06, 4.33046e-06, 
    4.084876e-06, 5.889308e-06, 5.550474e-06, 3.341644e-06, 4.121241e-06,
  8.765929e-08, 1.131675e-08, 2.332808e-08, 7.316063e-09, 2.455476e-08, 
    8.369588e-09, 4.756392e-08, 1.675178e-08, 5.661584e-07, 1.550092e-06, 
    3.061518e-06, 4.040719e-06, 5.624206e-06, 4.693735e-06, 3.98443e-06,
  4.037956e-07, 2.190501e-08, 3.816693e-09, 6.242423e-10, 3.814162e-09, 
    1.559247e-08, 5.537026e-08, 2.4532e-08, 3.028152e-08, 2.145676e-07, 
    5.418789e-07, 2.178521e-06, 3.738533e-06, 4.476979e-06, 3.002246e-06,
  1.542536e-06, 4.633909e-08, 2.959548e-09, 1.361297e-09, 7.829012e-10, 
    1.237476e-09, 8.407217e-09, 1.808481e-08, 7.793457e-09, 1.089549e-08, 
    6.523109e-09, 3.150944e-07, 6.405292e-07, 6.750273e-07, 1.371477e-06,
  3.13391e-06, 3.83481e-07, 6.198452e-09, 1.931718e-09, 1.865842e-09, 
    1.528672e-09, 3.675534e-09, 1.511199e-09, 1.357123e-09, 2.669049e-09, 
    5.131582e-09, 5.647013e-09, 1.193925e-08, 3.444072e-07, 1.167338e-06,
  6.509851e-06, 2.578978e-06, 2.967213e-07, 1.613208e-07, 5.730022e-09, 
    4.655615e-09, 9.259266e-08, 4.216814e-08, 1.394634e-08, 4.23466e-09, 
    1.060953e-09, 3.940293e-09, 6.149248e-09, 9.61962e-09, 5.499756e-08,
  5.104015e-05, 2.5967e-05, 8.661348e-06, 2.773141e-06, 2.088508e-07, 
    2.283057e-07, 1.358935e-06, 5.376945e-07, 4.729772e-07, 1.981032e-08, 
    2.002333e-09, 7.334041e-09, 1.951919e-09, 1.212072e-08, 5.164869e-09,
  7.36627e-05, 0.0001020237, 0.0001026849, 0.0001361918, 0.0001332087, 
    0.0001201338, 4.622913e-05, 5.836423e-06, 3.627013e-06, 3.928784e-06, 
    5.889982e-09, 1.406425e-09, 2.122957e-09, 2.952066e-09, 1.483788e-08,
  2.674933e-05, 7.866306e-05, 9.643537e-05, 0.0001480792, 0.0002183684, 
    0.0002480592, 0.0003000369, 0.0003244108, 0.0002537445, 5.523478e-05, 
    2.469866e-06, 1.79342e-09, 6.894361e-10, 2.361353e-09, 3.414569e-09,
  1.282102e-05, 2.131929e-05, 2.296666e-05, 1.796733e-05, 4.384786e-05, 
    7.578715e-05, 0.0001411715, 0.0002596169, 0.0002904238, 0.0001900225, 
    7.164406e-05, 3.527932e-05, 2.909017e-05, 2.210768e-05, 1.565536e-05,
  1.6772e-05, 1.683032e-05, 1.829249e-05, 1.90653e-05, 2.260885e-05, 
    2.006176e-05, 1.991945e-05, 2.507047e-05, 1.991601e-05, 1.919679e-05, 
    1.663724e-05, 4.282814e-05, 4.235261e-06, 5.446358e-06, 6.902511e-06,
  1.8407e-05, 3.683138e-06, 8.395282e-06, 1.423485e-05, 1.462624e-05, 
    2.353414e-05, 3.273801e-05, 2.021217e-05, 2.260603e-05, 2.201279e-05, 
    2.288906e-05, 2.049051e-05, 2.032793e-05, 7.166933e-06, 9.90285e-06,
  1.306932e-05, 1.050536e-05, 4.691114e-06, 5.53499e-06, 8.006262e-06, 
    1.657338e-05, 2.737177e-05, 1.589843e-05, 2.548852e-05, 1.632322e-05, 
    6.551128e-06, 5.747962e-06, 1.360797e-05, 5.603571e-06, 9.860914e-06,
  1.776917e-05, 8.363194e-06, 3.052859e-06, 3.441598e-06, 1.905848e-06, 
    2.295128e-06, 1.15333e-05, 1.353197e-05, 1.510072e-05, 5.872413e-06, 
    3.706307e-06, 2.304913e-06, 1.760953e-06, 9.316587e-07, 5.173461e-07,
  4.581322e-06, 5.654242e-06, 3.347745e-07, 1.707389e-07, 1.336548e-06, 
    2.445153e-06, 3.506541e-06, 6.052551e-06, 7.01391e-06, 4.988717e-06, 
    3.126879e-06, 2.378953e-06, 3.011544e-07, 1.534561e-06, 2.276658e-06,
  4.923026e-06, 5.828591e-06, 3.159804e-06, 2.451617e-07, 6.662662e-07, 
    2.849725e-07, 1.480883e-06, 4.633196e-06, 8.867564e-06, 8.233163e-06, 
    8.280957e-06, 5.049787e-06, 1.351731e-06, 2.136956e-06, 1.713047e-06,
  8.014069e-06, 5.476852e-06, 5.634909e-06, 3.374805e-06, 8.482833e-09, 
    2.315585e-08, 2.798409e-06, 3.197856e-06, 1.199252e-05, 9.598207e-06, 
    7.835042e-06, 6.329718e-06, 1.804759e-06, 1.241645e-06, 2.079672e-07,
  2.485066e-06, 4.492326e-06, 5.744962e-06, 4.678623e-06, 1.430994e-08, 
    1.342338e-08, 4.864247e-07, 3.838025e-06, 1.094695e-05, 1.936574e-05, 
    1.211945e-05, 4.706802e-06, 2.618451e-06, 1.599828e-06, 7.317679e-07,
  4.449426e-06, 1.850616e-06, 4.946073e-06, 3.998655e-06, 7.882518e-07, 
    1.877135e-07, 8.758523e-08, 6.236561e-07, 5.568357e-06, 1.408428e-05, 
    1.433349e-05, 4.453901e-06, 3.408848e-06, 1.823778e-06, 1.498634e-06,
  3.15064e-06, 4.707953e-06, 3.087162e-06, 9.083441e-07, 7.555565e-07, 
    1.89144e-06, 7.224869e-08, 4.82413e-08, 7.162969e-07, 6.15718e-06, 
    1.237366e-05, 1.070014e-05, 3.032576e-06, 2.563854e-06, 2.812171e-06,
  0.0004583704, 0.0004882106, 0.0004828577, 0.0004050686, 0.0003114747, 
    0.0001911369, 0.0001465466, 8.5579e-05, 8.904017e-05, 0.0001149211, 
    0.0001138451, 0.0001810586, 0.0002331596, 0.0002338676, 0.0001977627,
  0.0004501847, 0.000431144, 0.0003307052, 0.0001805089, 7.350583e-05, 
    5.022719e-05, 4.748075e-05, 3.557884e-05, 3.690795e-05, 5.329894e-05, 
    8.871782e-05, 9.758465e-05, 0.0001104625, 0.00012129, 0.0001490495,
  0.0003268967, 0.0002553064, 0.0001155927, 3.815583e-05, 3.832497e-06, 
    3.067068e-06, 6.193688e-06, 7.936133e-06, 2.414981e-05, 2.35347e-05, 
    4.278345e-05, 4.543387e-05, 0.0001098988, 5.816715e-05, 9.570675e-05,
  0.0001505837, 5.391466e-05, 1.130087e-05, 2.028241e-06, 2.981537e-06, 
    1.10928e-06, 6.540287e-07, 6.012765e-06, 1.162682e-05, 1.17295e-05, 
    7.215722e-06, 3.301357e-06, 4.118524e-06, 8.966704e-06, 2.560525e-05,
  6.173345e-05, 5.095534e-05, 5.799064e-06, 1.202425e-06, 2.686799e-06, 
    2.836553e-06, 2.582279e-06, 2.814048e-06, 3.773396e-06, 4.888117e-06, 
    2.244885e-06, 2.977716e-06, 6.840888e-06, 4.620018e-07, 2.529884e-06,
  5.97603e-05, 6.548852e-05, 4.120125e-05, 3.10158e-06, 6.573396e-06, 
    1.111138e-05, 7.973799e-06, 1.673157e-06, 2.317868e-06, 9.081906e-06, 
    1.362047e-05, 1.482414e-05, 8.760993e-06, 5.650219e-06, 1.362593e-05,
  7.902408e-05, 7.259786e-05, 6.655128e-05, 5.200489e-05, 7.922982e-06, 
    1.81171e-05, 1.164034e-05, 2.60384e-06, 4.566416e-06, 7.938476e-06, 
    1.25798e-05, 1.176524e-05, 1.189166e-05, 3.79649e-06, 3.579228e-06,
  9.205846e-05, 9.816667e-05, 8.532598e-05, 4.604866e-05, 1.260869e-05, 
    1.361153e-05, 7.921553e-06, 2.169541e-06, 1.140779e-07, 6.403886e-06, 
    9.902489e-06, 8.044902e-06, 1.068191e-05, 1.055739e-05, 5.993572e-06,
  0.0001007473, 7.860526e-05, 4.124532e-05, 2.670142e-05, 9.528065e-06, 
    6.857537e-06, 3.354343e-06, 7.338543e-07, 1.823256e-07, 4.393444e-06, 
    9.392326e-06, 1.168341e-05, 1.086353e-05, 1.038837e-05, 1.351161e-05,
  5.34629e-05, 6.577936e-05, 3.717291e-05, 9.474758e-06, 1.718665e-06, 
    1.546049e-06, 9.589556e-07, 3.001959e-07, 2.747063e-07, 2.549464e-06, 
    8.081383e-06, 1.345117e-05, 1.358452e-05, 1.422943e-05, 9.369173e-06,
  3.209923e-05, 7.47637e-05, 0.0001334329, 0.0002285221, 0.0002827841, 
    0.0003064586, 0.0002569702, 0.0002246215, 0.0001688407, 0.000138972, 
    7.739071e-05, 7.222512e-05, 9.286713e-05, 0.0001368595, 0.0001461728,
  1.584687e-05, 3.630841e-05, 9.479793e-05, 0.0001388292, 0.0001803401, 
    0.0001591445, 0.0001525793, 0.000116836, 0.000145008, 0.0001281211, 
    0.0001327446, 0.0001502016, 0.0001181033, 0.000129019, 0.0001052771,
  5.936822e-06, 1.445478e-05, 4.065603e-05, 5.602123e-05, 0.0001009786, 
    0.0001035863, 0.0001118698, 8.530189e-05, 0.0001010659, 0.0001131522, 
    0.0001286791, 0.0001151051, 0.0001051559, 9.853196e-05, 6.500147e-05,
  8.838453e-06, 1.498911e-05, 2.124777e-05, 2.783652e-05, 5.935339e-05, 
    7.339653e-05, 8.704057e-05, 0.0001012085, 0.0001141763, 9.984957e-05, 
    7.802376e-05, 6.975173e-05, 6.161955e-05, 5.859633e-05, 3.845973e-05,
  9.030535e-06, 1.101517e-05, 1.785011e-05, 1.590179e-05, 3.072838e-05, 
    5.279032e-05, 7.641477e-05, 0.0001098045, 0.0001069681, 8.857928e-05, 
    5.735201e-05, 4.512084e-05, 3.726824e-05, 3.923677e-05, 3.649827e-05,
  1.264318e-05, 1.165875e-05, 1.380592e-05, 9.226009e-06, 1.586262e-05, 
    3.457766e-05, 6.976716e-05, 0.0001082372, 0.0001364979, 7.896475e-05, 
    5.073585e-05, 5.284882e-05, 3.591129e-05, 3.636442e-05, 3.608691e-05,
  7.842048e-06, 1.176689e-05, 1.695702e-05, 2.263727e-05, 1.768531e-05, 
    3.336483e-05, 6.875998e-05, 9.359187e-05, 8.297913e-05, 5.856947e-05, 
    4.143536e-05, 4.696937e-05, 5.30873e-05, 3.354558e-05, 4.063803e-05,
  2.568663e-06, 1.094741e-05, 1.777072e-05, 2.008513e-05, 3.041526e-06, 
    2.338296e-05, 5.580453e-05, 4.157679e-05, 4.991091e-05, 4.594149e-05, 
    4.532604e-05, 2.964861e-05, 4.342193e-05, 3.143307e-05, 3.774012e-05,
  6.475385e-06, 2.104399e-05, 2.800042e-05, 3.507222e-05, 4.291766e-05, 
    5.166952e-06, 2.379894e-05, 2.990461e-05, 4.000239e-05, 3.687908e-05, 
    2.937035e-05, 3.466775e-05, 5.442595e-05, 3.944571e-05, 6.530141e-05,
  1.666317e-05, 1.526056e-05, 2.653499e-05, 4.78438e-05, 4.722148e-05, 
    3.496049e-05, 6.588507e-06, 1.161896e-05, 1.817656e-05, 3.151911e-05, 
    3.702251e-05, 2.66287e-05, 2.260771e-05, 7.901905e-05, 2.747024e-05,
  6.91841e-05, 5.30745e-05, 3.089752e-05, 8.586486e-05, 2.669748e-05, 
    9.673752e-05, 0.0001291489, 0.0001247064, 0.0001227892, 0.0001047597, 
    0.0001011013, 6.257946e-05, 5.363954e-05, 5.402164e-05, 4.383698e-05,
  1.010828e-05, 2.714729e-05, 3.676465e-05, 1.806793e-05, 7.579599e-05, 
    0.0001296027, 0.0001306377, 0.0001186662, 0.0001401844, 0.0001654998, 
    0.0001649421, 0.0001530634, 9.258561e-05, 5.446827e-05, 4.843769e-05,
  3.231405e-06, 7.938656e-06, 2.414376e-05, 2.436611e-05, 0.0001100544, 
    0.0001526808, 0.0001507291, 0.0001400904, 0.0001438858, 0.0001611428, 
    0.0001869105, 0.0001614798, 0.0001753925, 0.0001281298, 7.592246e-05,
  3.227072e-06, 8.520581e-06, 2.793669e-05, 2.26843e-05, 8.735798e-05, 
    0.0001385513, 0.0001882284, 0.0001448079, 0.0002007678, 0.0001750771, 
    0.0001326285, 0.000116397, 9.20522e-05, 0.000134755, 8.73687e-05,
  2.645149e-06, 4.660556e-06, 7.33208e-06, 1.832644e-05, 5.647989e-05, 
    9.310436e-05, 0.0001335995, 0.0001782379, 0.0001770379, 0.0001877159, 
    0.0001524901, 9.718927e-05, 0.0001865664, 0.0001302719, 0.0001287997,
  6.605474e-08, 7.179269e-06, 1.980857e-06, 7.85325e-06, 5.188364e-05, 
    6.396853e-05, 0.0001013789, 0.0001402308, 0.0001831942, 0.0002035402, 
    0.0001765167, 0.0001774006, 0.0001378435, 0.0001174772, 0.0001280797,
  5.318788e-08, 2.699848e-07, 1.039129e-06, 4.744939e-07, 2.111735e-05, 
    6.735316e-05, 7.939769e-05, 9.305139e-05, 0.0001088467, 0.0001045747, 
    0.0001054087, 9.865452e-05, 9.204568e-05, 9.626066e-05, 6.803707e-05,
  2.384019e-10, 7.170735e-11, 1.75944e-07, 1.709397e-07, 7.243553e-07, 
    2.198245e-05, 6.082364e-05, 6.086634e-05, 5.280485e-05, 4.354193e-05, 
    4.906692e-05, 4.966391e-05, 4.95142e-05, 3.335242e-05, 2.856929e-05,
  4.91007e-11, 2.428794e-11, 3.356384e-08, 9.809378e-08, 3.491934e-07, 
    3.473855e-06, 2.759885e-05, 2.821487e-05, 3.099007e-05, 2.728185e-05, 
    2.399142e-05, 2.278865e-05, 1.930447e-05, 1.780862e-05, 1.609275e-05,
  6.938234e-11, 2.492256e-10, 7.651177e-10, 6.90966e-08, 2.943959e-08, 
    2.6613e-07, 7.186949e-06, 2.215497e-05, 2.638636e-05, 3.104464e-05, 
    2.204954e-05, 1.853908e-05, 1.735021e-05, 2.683856e-05, 2.575742e-05,
  2.333426e-05, 1.263628e-05, 4.546365e-06, 1.348237e-05, 3.124652e-05, 
    2.362432e-05, 2.466054e-05, 2.435746e-05, 3.795036e-05, 3.518941e-05, 
    3.365927e-05, 5.236604e-05, 6.403964e-05, 8.863067e-05, 9.392272e-05,
  9.382221e-06, 1.513338e-05, 2.695098e-06, 1.717026e-06, 5.427262e-05, 
    5.9074e-05, 3.283875e-05, 3.049882e-05, 4.067121e-05, 3.563081e-05, 
    4.122777e-05, 4.413626e-05, 5.389827e-05, 7.129239e-05, 8.450778e-05,
  1.223652e-06, 3.351096e-06, 1.671522e-05, 5.160363e-06, 4.398111e-05, 
    8.43345e-05, 6.044085e-05, 6.515706e-05, 3.818702e-05, 3.920243e-05, 
    4.479441e-05, 4.235663e-05, 5.771309e-05, 7.032557e-05, 7.67033e-05,
  5.52185e-07, 4.160393e-06, 3.029976e-05, 8.939389e-06, 4.862925e-05, 
    7.451747e-05, 0.0001313549, 0.0001374889, 7.79583e-05, 4.687565e-05, 
    3.760444e-05, 3.852934e-05, 4.054225e-05, 4.694963e-05, 5.348435e-05,
  6.712475e-08, 6.986657e-07, 1.054741e-05, 1.967564e-05, 3.465188e-05, 
    6.949193e-05, 0.0001209086, 0.0001620916, 0.0001242939, 8.628629e-05, 
    6.633793e-05, 4.178367e-05, 3.455345e-05, 3.675451e-05, 6.032664e-05,
  4.380289e-10, 1.275686e-07, 1.50185e-06, 7.546022e-06, 3.372948e-05, 
    6.532542e-05, 0.0001034869, 0.0001612278, 0.0001608602, 0.0001266822, 
    0.000110493, 8.292864e-05, 7.986865e-05, 8.079004e-05, 4.999694e-05,
  1.080737e-10, 3.875593e-10, 1.830917e-07, 6.703724e-07, 2.881154e-05, 
    7.591212e-05, 0.0001120697, 0.000175442, 0.000213395, 0.0001886826, 
    0.0001808769, 0.0001712913, 0.0001521689, 0.0001016204, 9.78508e-05,
  3.495488e-12, 1.997571e-11, 1.009733e-08, 9.510563e-08, 4.459741e-07, 
    5.644085e-05, 0.0001294382, 0.0001574355, 0.0002051707, 0.0001983151, 
    0.000197976, 0.0001993898, 0.0001952219, 0.0001629709, 0.0001452692,
  2.629429e-12, 9.110344e-13, 3.669176e-12, 3.527296e-12, 2.391578e-08, 
    3.382748e-06, 0.0001019559, 0.0001717297, 0.0002168187, 0.0001987559, 
    0.0002144023, 0.0002149922, 0.0001693971, 0.0001478027, 0.0001434961,
  8.91612e-13, 6.492526e-13, 9.892662e-11, 5.140169e-10, 5.216417e-10, 
    6.816603e-07, 3.800435e-05, 0.0001142865, 0.0002424477, 0.0002718192, 
    0.0001940767, 0.0001568067, 0.0001818594, 0.0001468064, 0.0001326084,
  4.899433e-08, 1.260722e-08, 5.964973e-09, 2.194651e-09, 6.394727e-07, 
    1.907301e-06, 3.6962e-06, 3.765881e-06, 5.389008e-06, 5.707124e-06, 
    6.90003e-06, 9.087585e-06, 1.173926e-05, 1.258699e-05, 1.36879e-05,
  5.41328e-09, 8.222359e-09, 1.172979e-07, 4.965493e-10, 3.238654e-06, 
    4.514772e-06, 3.43802e-06, 4.04103e-06, 6.520473e-06, 5.396093e-06, 
    6.258047e-06, 9.913449e-06, 1.236418e-05, 1.745062e-05, 2.481262e-05,
  4.529668e-09, 1.023703e-08, 5.410177e-09, 1.386252e-09, 2.301287e-06, 
    7.730891e-06, 4.058227e-06, 4.286479e-06, 6.565338e-06, 7.069471e-06, 
    5.582001e-06, 6.347331e-06, 1.049389e-05, 1.538038e-05, 1.974712e-05,
  4.311051e-09, 9.453872e-09, 1.574993e-08, 3.530362e-07, 3.118405e-06, 
    9.859956e-06, 6.438283e-06, 5.431747e-06, 6.744775e-06, 7.134561e-06, 
    6.014527e-06, 5.644601e-06, 9.423189e-06, 1.156678e-05, 1.278384e-05,
  6.983844e-09, 3.995601e-09, 5.386589e-09, 1.98624e-07, 1.644033e-06, 
    7.919302e-06, 1.089874e-05, 6.047575e-06, 5.83292e-06, 8.595128e-06, 
    9.384534e-06, 6.668593e-06, 7.57405e-06, 1.116203e-05, 1.584989e-05,
  4.311629e-09, 6.505124e-09, 3.683283e-09, 1.384038e-09, 1.237672e-06, 
    9.63707e-06, 1.249602e-05, 7.867178e-06, 6.061785e-06, 8.118265e-06, 
    1.133244e-05, 1.100408e-05, 1.04511e-05, 1.220786e-05, 1.965352e-05,
  4.922347e-10, 4.98902e-09, 6.225671e-09, 1.667592e-09, 4.460987e-07, 
    4.809705e-06, 1.314336e-05, 1.44193e-05, 6.703533e-06, 8.059817e-06, 
    1.247859e-05, 1.231674e-05, 1.100046e-05, 1.172777e-05, 1.506675e-05,
  2.183182e-10, 7.28241e-10, 3.773228e-09, 4.46863e-09, 2.270812e-09, 
    8.608293e-07, 1.434402e-05, 1.773462e-05, 1.445968e-05, 6.500681e-06, 
    7.536295e-06, 1.265556e-05, 1.287156e-05, 1.156864e-05, 1.484781e-05,
  3.028513e-17, 1.756143e-11, 1.842065e-09, 1.493707e-09, 2.688939e-10, 
    1.808184e-07, 6.165195e-06, 1.884173e-05, 2.172688e-05, 9.553268e-06, 
    8.920599e-06, 9.288991e-06, 1.245113e-05, 1.587498e-05, 1.631347e-05,
  1.451566e-22, 2.269832e-15, 4.27605e-11, 1.13094e-09, 1.361642e-09, 
    3.75994e-09, 2.124588e-06, 1.386183e-05, 2.710537e-05, 2.431893e-05, 
    1.432321e-05, 8.111694e-06, 1.006874e-05, 1.333234e-05, 1.600419e-05,
  1.361742e-07, 1.042288e-07, 7.208982e-08, 4.771295e-08, 8.732239e-07, 
    6.222697e-06, 1.719215e-05, 4.509209e-05, 6.926111e-05, 0.000101939, 
    0.0001110976, 4.844907e-05, 1.265514e-05, 2.881747e-07, 4.708474e-07,
  3.022408e-07, 8.229221e-08, 4.45483e-08, 3.928544e-08, 2.984782e-06, 
    1.286038e-05, 2.987806e-05, 4.25834e-05, 7.715329e-05, 0.0001062068, 
    7.264504e-05, 2.364938e-05, 3.30038e-06, 8.370653e-07, 1.07434e-06,
  9.434801e-07, 2.466504e-08, 3.201383e-08, 2.14599e-08, 3.996646e-06, 
    1.570434e-05, 2.771109e-05, 4.693085e-05, 9.344822e-05, 9.752417e-05, 
    4.675631e-05, 1.156156e-05, 1.013556e-06, 9.589113e-07, 1.479381e-06,
  2.750386e-08, 1.227404e-08, 2.40432e-08, 1.829093e-08, 2.290253e-06, 
    1.424319e-05, 2.504566e-05, 4.83183e-05, 0.0001050985, 0.0001139581, 
    2.345687e-05, 1.634248e-06, 1.13866e-06, 1.773708e-06, 2.985642e-06,
  2.919256e-09, 6.158083e-09, 1.24893e-08, 1.506384e-08, 5.057871e-07, 
    8.985717e-06, 1.999732e-05, 4.643964e-05, 0.0001023129, 9.017687e-05, 
    1.7752e-05, 1.824298e-06, 1.208348e-06, 1.269073e-06, 4.53266e-06,
  3.472909e-09, 5.26003e-09, 8.050794e-09, 1.076232e-08, 8.021861e-08, 
    5.619407e-06, 1.546111e-05, 4.264815e-05, 8.906791e-05, 8.879966e-05, 
    1.489671e-05, 5.247667e-07, 8.602339e-07, 2.762617e-06, 4.307095e-06,
  7.437581e-10, 1.786336e-09, 7.28462e-09, 1.045869e-08, 4.475719e-08, 
    1.953013e-06, 1.354795e-05, 3.614048e-05, 8.900761e-05, 8.239166e-05, 
    1.455245e-05, 7.992895e-07, 1.717081e-06, 3.187115e-06, 3.829261e-06,
  4.420874e-10, 1.475035e-09, 4.086623e-09, 7.117554e-09, 3.94442e-08, 
    3.990824e-07, 1.405302e-05, 3.371189e-05, 8.363128e-05, 7.925468e-05, 
    1.441141e-05, 1.143347e-06, 4.200514e-07, 2.970317e-06, 5.26339e-06,
  7.021801e-13, 3.703626e-11, 6.391088e-10, 4.182789e-09, 6.524043e-09, 
    2.622402e-08, 1.726595e-05, 3.219238e-05, 7.40169e-05, 7.36644e-05, 
    1.561181e-05, 1.354433e-06, 1.469088e-06, 4.622798e-06, 6.221205e-06,
  3.101129e-14, 2.056352e-11, 2.374473e-10, 6.66226e-10, 5.094912e-09, 
    1.508797e-08, 6.744491e-07, 2.658404e-05, 5.152558e-05, 6.288784e-05, 
    2.239806e-05, 4.17813e-06, 2.451242e-06, 4.66635e-06, 7.087093e-06,
  3.348329e-05, 4.405663e-05, 6.991749e-05, 8.56156e-05, 8.249181e-05, 
    7.39778e-05, 3.832178e-05, 3.199718e-05, 3.020882e-05, 7.334515e-05, 
    0.0002936159, 0.0005028815, 0.0005283501, 0.0003850793, 0.0002482506,
  6.036102e-05, 7.070503e-05, 7.248744e-05, 3.964649e-05, 7.21129e-05, 
    5.213427e-05, 4.909487e-05, 3.045341e-05, 2.779833e-05, 7.930979e-05, 
    0.0002998331, 0.0004583998, 0.0004266906, 0.0002975603, 0.0001918697,
  5.190478e-05, 4.360338e-05, 3.745838e-05, 2.518063e-05, 5.292328e-05, 
    3.751518e-05, 3.265906e-05, 2.865804e-05, 2.712814e-05, 0.0001729745, 
    0.0005413545, 0.0004805618, 0.0002739493, 0.0001826853, 0.0001183817,
  2.961945e-05, 2.617302e-05, 2.637809e-05, 1.759012e-05, 2.742709e-05, 
    3.659321e-05, 3.406292e-05, 2.396496e-05, 2.811269e-05, 0.0001666479, 
    0.00042815, 0.0003158124, 0.000265292, 0.0001005335, 9.377312e-05,
  1.13752e-05, 8.576503e-06, 3.810509e-06, 8.62752e-06, 1.076453e-05, 
    2.790754e-05, 2.130623e-05, 1.934418e-05, 3.405627e-05, 0.0003112988, 
    0.0002822307, 0.0001979516, 0.0001161981, 0.0001299358, 0.0001205624,
  3.99516e-06, 4.160799e-06, 4.933133e-06, 1.707117e-06, 9.907418e-07, 
    1.418768e-05, 1.250221e-05, 1.541359e-05, 4.99059e-05, 0.00020116, 
    0.0001660218, 0.0001414205, 0.0001802571, 0.000134767, 0.0001996187,
  1.746474e-06, 2.59928e-06, 3.525261e-06, 1.211728e-06, 1.462536e-06, 
    6.806496e-06, 1.071351e-05, 1.790562e-05, 4.643374e-05, 0.0001108382, 
    0.0001138782, 0.0001069129, 0.0001370257, 0.000152591, 0.0002251405,
  1.274114e-06, 1.630364e-06, 8.997449e-07, 8.868482e-07, 4.450556e-08, 
    6.915601e-06, 8.80465e-06, 1.176613e-05, 3.349415e-05, 7.838291e-05, 
    7.948519e-05, 0.0001052545, 0.0001316236, 0.0001643083, 0.0002180815,
  8.648308e-07, 1.682978e-06, 5.837703e-07, 3.748866e-07, 7.072897e-08, 
    1.278912e-07, 4.394898e-06, 6.414829e-06, 1.852589e-05, 4.936366e-05, 
    8.474564e-05, 0.0001059058, 0.0001695698, 0.0001953295, 0.0001468984,
  1.011151e-06, 1.797682e-06, 2.241025e-06, 1.387119e-06, 5.067567e-07, 
    6.408832e-07, 4.848555e-06, 7.070829e-06, 1.521033e-05, 4.076142e-05, 
    0.0001270389, 0.0002956686, 0.0002498227, 0.0001983822, 7.332607e-05,
  6.773914e-05, 9.77985e-05, 8.749474e-05, 0.000106872, 0.0001630649, 
    0.0001792685, 0.0001231152, 0.0001565863, 0.0001322418, 0.000181503, 
    0.0001612169, 0.0002440745, 0.0003000362, 0.0002965177, 0.0002531671,
  5.878481e-06, 1.838454e-05, 4.671175e-05, 5.958268e-05, 0.0001858047, 
    0.0002279261, 0.000247, 0.0001715021, 0.0001822553, 0.0001890508, 
    0.0001830725, 0.0002418208, 0.0001960266, 0.0001866604, 0.0001620876,
  3.731922e-06, 4.402489e-06, 1.31536e-05, 3.749648e-05, 0.0001446157, 
    0.0001822576, 0.0002556915, 0.0002819413, 0.0002133311, 0.0002813618, 
    0.0002354239, 0.0002045093, 0.0001886378, 0.0001397833, 0.0001002078,
  5.363935e-06, 5.40332e-06, 3.449999e-05, 2.138534e-05, 8.827491e-05, 
    0.0001580351, 0.0002191677, 0.0002815417, 0.0003031201, 0.0002570428, 
    0.00019901, 0.0001598214, 0.00015058, 0.0001134051, 0.0001014248,
  4.486183e-06, 6.356653e-06, 4.232212e-06, 2.834988e-05, 3.599383e-05, 
    9.926657e-05, 0.0001354124, 0.0001776409, 0.0001933159, 0.0001961767, 
    0.0001912998, 0.0001919767, 0.0001459128, 0.0001154979, 0.0001338918,
  4.116725e-06, 4.979969e-06, 7.731655e-06, 1.234193e-05, 1.51404e-05, 
    5.334124e-05, 6.823696e-05, 9.172304e-05, 0.000114897, 0.0001394824, 
    0.0001616934, 0.0001506973, 0.0001456515, 0.0001465824, 0.0001561275,
  1.538174e-06, 2.24047e-06, 2.930873e-06, 3.998482e-06, 1.437519e-05, 
    2.932636e-05, 4.622264e-05, 5.519401e-05, 6.485303e-05, 8.357444e-05, 
    0.0001110443, 0.0001098563, 9.878958e-05, 0.0001364216, 0.0002047926,
  2.029855e-07, 1.501847e-06, 5.611794e-07, 3.150506e-06, 7.121361e-07, 
    2.509225e-05, 3.403772e-05, 3.408259e-05, 4.54962e-05, 5.681875e-05, 
    7.158132e-05, 6.138553e-05, 8.667132e-05, 0.0002047296, 0.0002397146,
  3.901671e-07, 4.086629e-08, 1.684833e-07, 5.650702e-07, 1.035299e-06, 
    3.014621e-06, 3.013366e-05, 2.662066e-05, 3.939643e-05, 4.744326e-05, 
    4.456715e-05, 5.409083e-05, 0.0001459563, 0.0002003651, 0.0002687261,
  1.728718e-08, 1.033055e-07, 7.006419e-07, 9.499311e-07, 1.112474e-06, 
    1.248828e-06, 1.976081e-05, 2.290636e-05, 2.72876e-05, 2.39654e-05, 
    3.04577e-05, 8.847576e-05, 0.0001816634, 0.0002169341, 0.0002405502,
  3.563211e-05, 6.245034e-05, 4.864946e-05, 6.823809e-05, 7.661535e-05, 
    6.358767e-05, 3.277749e-05, 3.81992e-05, 7.339843e-05, 0.0001450134, 
    0.0002153251, 0.0003326342, 0.0002798662, 0.0002311488, 0.0002471008,
  2.646141e-06, 1.961134e-05, 3.736979e-05, 3.918634e-05, 9.195517e-05, 
    9.41987e-05, 7.246342e-05, 4.51531e-05, 3.992871e-05, 4.210385e-05, 
    8.154074e-05, 0.0001659578, 0.0002356565, 0.0002416595, 0.000219256,
  2.742919e-07, 4.686796e-07, 1.160431e-05, 2.194677e-05, 8.858871e-05, 
    0.0001071622, 9.914021e-05, 8.233114e-05, 6.01341e-05, 3.963972e-05, 
    3.745628e-05, 5.943868e-05, 8.511257e-05, 0.0001619734, 0.000167548,
  2.907728e-07, 2.716167e-07, 9.910149e-07, 1.151087e-05, 6.833067e-05, 
    0.000101581, 0.0001206121, 0.0001211954, 0.00010756, 7.531458e-05, 
    4.220934e-05, 2.645183e-05, 3.125122e-05, 4.495072e-05, 7.084377e-05,
  2.372532e-07, 2.04093e-07, 1.77529e-07, 1.894698e-06, 2.512123e-05, 
    7.729114e-05, 0.0001042653, 0.0001356229, 0.0001368573, 0.0001159931, 
    7.838069e-05, 5.544475e-05, 3.183491e-05, 2.658386e-05, 2.304179e-05,
  2.575875e-09, 1.387466e-08, 1.854544e-07, 5.233568e-07, 2.994993e-06, 
    3.777434e-05, 6.833814e-05, 0.000103033, 0.0001257231, 0.0001577221, 
    0.0001385808, 0.0001146608, 7.540967e-05, 5.912943e-05, 4.133866e-05,
  9.513382e-13, 1.047181e-11, 5.013995e-09, 1.992733e-10, 6.816113e-07, 
    9.893915e-06, 3.267993e-05, 5.913462e-05, 9.581535e-05, 0.0001272045, 
    0.0001634479, 0.0001549013, 0.000135711, 0.0001032485, 6.384875e-05,
  3.83308e-12, 9.562382e-14, 1.133107e-13, 2.329778e-13, 1.12915e-10, 
    1.292203e-06, 1.028325e-05, 2.851277e-05, 4.694446e-05, 6.715427e-05, 
    0.0001019905, 0.000115407, 0.0001289768, 0.0001184623, 0.0001029785,
  4.640963e-11, 2.848397e-11, 8.873602e-12, 6.150426e-12, 1.392812e-10, 
    2.58746e-10, 6.55531e-07, 8.166948e-06, 1.54379e-05, 2.354815e-05, 
    3.723723e-05, 6.8102e-05, 8.287235e-05, 9.174002e-05, 8.775473e-05,
  7.573198e-11, 2.222186e-10, 5.681039e-11, 6.349407e-11, 1.024342e-10, 
    5.019803e-10, 9.231988e-08, 1.239792e-07, 6.345507e-06, 1.041956e-05, 
    1.799437e-05, 2.439032e-05, 3.204724e-05, 4.479099e-05, 5.536716e-05,
  0.0001220758, 9.853116e-05, 3.758197e-05, 5.89035e-05, 9.645161e-05, 
    9.37459e-05, 4.827417e-05, 5.710493e-05, 9.216004e-05, 0.0001012747, 
    0.0001152976, 0.0001720655, 0.0002458717, 0.0002591505, 0.0001537973,
  8.413906e-05, 8.895963e-05, 5.82953e-05, 2.927123e-05, 0.0001447569, 
    0.0001460868, 0.0001004654, 5.869387e-05, 6.076326e-05, 5.413007e-05, 
    4.981197e-05, 5.221607e-05, 7.684641e-05, 0.0001077337, 0.0001536662,
  8.10413e-05, 7.381138e-05, 8.85103e-05, 2.073769e-05, 0.0001366899, 
    0.0002008408, 0.0001291849, 8.203663e-05, 6.232043e-05, 4.289486e-05, 
    2.677804e-05, 2.053228e-05, 2.341119e-05, 2.843481e-05, 3.637361e-05,
  4.142763e-05, 5.96221e-05, 2.889714e-05, 4.539996e-05, 0.0001124504, 
    0.0001650204, 0.0001682329, 0.0001233391, 0.0001050386, 8.792993e-05, 
    6.593095e-05, 4.215754e-05, 2.826797e-05, 1.610498e-05, 7.929176e-06,
  1.225422e-05, 2.28644e-05, 1.716212e-05, 1.286567e-05, 3.398911e-05, 
    0.0001080029, 0.0001315569, 0.0001241701, 0.0001019336, 9.689212e-05, 
    9.91976e-05, 7.155009e-05, 5.757638e-05, 4.351199e-05, 2.714931e-05,
  1.945509e-06, 2.232497e-06, 1.062446e-06, 1.226612e-06, 1.523245e-05, 
    6.389425e-05, 8.019162e-05, 8.43966e-05, 7.597537e-05, 6.95352e-05, 
    7.974146e-05, 7.759617e-05, 7.364589e-05, 6.631097e-05, 5.883822e-05,
  6.273644e-07, 1.831859e-06, 8.506268e-07, 5.194644e-08, 4.064427e-06, 
    3.524647e-05, 4.17901e-05, 4.26573e-05, 4.847061e-05, 4.979654e-05, 
    5.061471e-05, 4.740812e-05, 4.763438e-05, 5.342019e-05, 5.46927e-05,
  2.086651e-06, 1.099533e-06, 3.451403e-07, 2.691663e-07, 1.653223e-07, 
    7.867427e-06, 2.484628e-05, 3.177088e-05, 3.635739e-05, 3.88207e-05, 
    4.154862e-05, 3.778183e-05, 3.893306e-05, 4.294051e-05, 4.721929e-05,
  3.194698e-06, 2.506199e-06, 8.322265e-07, 5.418325e-07, 5.198332e-07, 
    5.022864e-07, 1.039062e-05, 2.031397e-05, 3.072923e-05, 3.823115e-05, 
    3.877373e-05, 4.418243e-05, 4.573325e-05, 4.333293e-05, 4.166783e-05,
  1.350026e-06, 1.19889e-06, 1.803802e-06, 1.737036e-06, 7.304405e-07, 
    6.803123e-07, 1.864695e-06, 6.968136e-06, 1.887669e-05, 2.654747e-05, 
    2.82975e-05, 3.471394e-05, 3.444761e-05, 3.172316e-05, 2.913199e-05,
  1.660557e-05, 6.90678e-06, 1.27485e-07, 5.204877e-06, 2.635121e-05, 
    3.020504e-05, 1.727682e-05, 1.365314e-05, 1.980944e-05, 1.374557e-05, 
    6.431923e-06, 1.035127e-05, 1.254922e-05, 1.367572e-05, 1.717202e-05,
  1.163196e-05, 1.160044e-05, 2.460448e-07, 1.505887e-07, 2.798894e-05, 
    3.983578e-05, 2.819674e-05, 2.196068e-05, 2.944306e-05, 2.442539e-05, 
    1.712267e-05, 1.747987e-05, 1.902176e-05, 9.898035e-06, 7.901143e-06,
  1.106069e-05, 1.667062e-05, 1.200917e-05, 2.597907e-06, 6.443086e-05, 
    0.0001036634, 6.827847e-05, 5.66073e-05, 5.868414e-05, 5.686345e-05, 
    4.419848e-05, 4.186483e-05, 4.294082e-05, 3.251459e-05, 2.045191e-05,
  2.193095e-05, 3.331133e-05, 5.021235e-05, 5.252431e-05, 0.0001307644, 
    0.000194219, 0.0001384886, 0.000106236, 9.225459e-05, 8.056482e-05, 
    6.96108e-05, 5.629075e-05, 4.025563e-05, 2.640215e-05, 2.254504e-05,
  3.384944e-05, 5.281893e-05, 4.206254e-05, 7.073311e-05, 0.0001315289, 
    0.0002648554, 0.0002312944, 0.0001473434, 0.0001218204, 8.640841e-05, 
    7.309749e-05, 5.953433e-05, 4.198082e-05, 2.651068e-05, 1.944577e-05,
  3.725151e-05, 5.077917e-05, 5.200035e-05, 8.232403e-05, 0.0001276702, 
    0.0002685687, 0.0002085555, 0.0001161767, 5.126237e-05, 3.015125e-05, 
    2.056229e-05, 2.675091e-05, 2.504095e-05, 2.8022e-05, 2.430456e-05,
  3.133782e-05, 3.913075e-05, 5.183154e-05, 0.0001289268, 0.0001923262, 
    0.0001667463, 0.0001139324, 8.215148e-05, 7.597116e-05, 4.636858e-05, 
    2.659935e-05, 2.426204e-05, 1.934168e-05, 2.148317e-05, 2.176935e-05,
  3.154659e-05, 4.133954e-05, 4.595292e-05, 0.0001564651, 0.0002210175, 
    0.0001097189, 7.148345e-05, 7.789719e-05, 9.901445e-05, 0.0001021598, 
    7.824918e-05, 3.910846e-05, 2.75951e-05, 2.00559e-05, 1.552765e-05,
  4.323088e-05, 5.154982e-05, 6.932866e-05, 0.000168617, 0.0002384319, 
    7.145595e-05, 4.837362e-05, 4.578237e-05, 4.437663e-05, 5.502692e-05, 
    6.253054e-05, 4.929294e-05, 3.411963e-05, 2.313277e-05, 1.779839e-05,
  3.457398e-05, 4.967198e-05, 8.131566e-05, 0.0001396539, 0.0001450714, 
    6.313642e-05, 2.43436e-05, 4.331991e-05, 4.279991e-05, 2.984716e-05, 
    2.699294e-05, 2.413837e-05, 2.358529e-05, 1.819088e-05, 1.593575e-05,
  3.83125e-07, 3.162683e-07, 2.365774e-07, 3.026393e-07, 5.41931e-06, 
    1.260249e-05, 1.166664e-05, 1.172358e-05, 1.682778e-05, 1.952441e-05, 
    2.19904e-05, 2.527476e-05, 2.810901e-05, 2.486406e-05, 2.443946e-05,
  1.757708e-08, 5.41045e-07, 1.354686e-07, 1.391568e-07, 4.144392e-06, 
    1.350451e-05, 1.436859e-05, 1.220479e-05, 1.466174e-05, 1.91515e-05, 
    1.832736e-05, 2.233792e-05, 2.852384e-05, 3.033486e-05, 3.124732e-05,
  3.950501e-09, 2.603962e-09, 4.427786e-09, 1.363882e-07, 2.014374e-06, 
    2.146144e-05, 2.397744e-05, 1.725299e-05, 1.431819e-05, 1.412305e-05, 
    1.090839e-05, 1.198826e-05, 1.5736e-05, 1.920575e-05, 2.275364e-05,
  1.282144e-09, 1.016286e-09, 5.608371e-07, 4.797956e-07, 4.639586e-06, 
    2.544426e-05, 3.05328e-05, 2.33485e-05, 1.945288e-05, 1.250284e-05, 
    8.557322e-06, 8.230612e-06, 6.955085e-06, 6.877966e-06, 6.243936e-06,
  3.19475e-09, 3.154465e-09, 1.579215e-06, 2.003489e-06, 1.358169e-06, 
    2.204711e-05, 3.362324e-05, 3.468072e-05, 2.964147e-05, 2.811047e-05, 
    2.346797e-05, 1.851658e-05, 1.14702e-05, 7.098564e-06, 1.000244e-06,
  2.142794e-09, 6.999179e-09, 2.264392e-08, 8.039498e-07, 4.74323e-06, 
    4.879507e-05, 4.946847e-05, 8.054783e-05, 5.774645e-05, 3.652818e-05, 
    2.584973e-05, 1.954945e-05, 2.149352e-05, 2.029624e-05, 1.619947e-05,
  7.673908e-10, 2.062099e-08, 3.115667e-08, 5.64622e-08, 8.940702e-06, 
    6.532852e-05, 0.0001567575, 0.0001096711, 5.642969e-05, 3.57715e-05, 
    1.402373e-05, 1.206169e-05, 1.037762e-05, 7.554634e-06, 9.835628e-06,
  8.589508e-11, 3.317514e-08, 5.931904e-08, 5.699816e-08, 8.964817e-06, 
    9.396981e-05, 0.0001540491, 0.0001017301, 7.186003e-05, 3.958453e-05, 
    3.650425e-05, 2.938571e-05, 1.279233e-05, 6.651479e-06, 7.598005e-06,
  1.857987e-10, 1.691729e-08, 7.169025e-09, 2.85914e-07, 2.709996e-05, 
    0.0001069765, 0.0001926618, 0.000117825, 5.550908e-05, 3.783661e-05, 
    3.400145e-05, 2.629132e-05, 2.443834e-05, 2.271786e-05, 1.679619e-05,
  2.116568e-11, 1.04569e-08, 1.149199e-06, 1.71636e-05, 5.960377e-05, 
    0.000148718, 0.0001443015, 0.0001614309, 8.312957e-05, 2.515104e-05, 
    1.086525e-05, 5.137362e-06, 9.515144e-06, 2.239635e-05, 2.794832e-05,
  3.74235e-11, 5.012459e-10, 1.080024e-09, 2.929044e-09, 1.018571e-07, 
    1.325565e-06, 2.54324e-06, 3.897743e-06, 1.13971e-05, 2.09328e-05, 
    3.525396e-05, 5.234868e-05, 6.434492e-05, 7.056808e-05, 7.755909e-05,
  1.263619e-09, 4.291052e-10, 5.297797e-10, 4.639523e-09, 2.008492e-08, 
    9.395759e-07, 1.355428e-06, 2.1602e-06, 7.116716e-06, 1.054881e-05, 
    2.133293e-05, 3.651378e-05, 4.806562e-05, 5.812548e-05, 6.590162e-05,
  2.782347e-10, 7.077817e-09, 9.757535e-09, 2.94711e-09, 5.943069e-08, 
    1.891242e-07, 9.167004e-07, 2.655776e-06, 7.420992e-06, 8.164756e-06, 
    9.47497e-06, 1.559017e-05, 2.636201e-05, 3.616995e-05, 4.355913e-05,
  9.800236e-10, 2.399779e-09, 2.524601e-09, 2.263677e-09, 8.617143e-09, 
    4.912744e-08, 6.366248e-08, 3.944691e-07, 5.574338e-06, 5.993705e-06, 
    4.911248e-06, 8.744327e-06, 1.441813e-05, 1.998795e-05, 2.153689e-05,
  8.035008e-11, 6.17806e-10, 1.825484e-09, 2.411131e-09, 3.515031e-09, 
    6.76324e-09, 9.13906e-09, 1.202892e-08, 1.757044e-06, 3.460339e-06, 
    4.786948e-06, 7.767585e-06, 1.217878e-05, 1.455455e-05, 1.577386e-05,
  5.47119e-11, 4.019924e-11, 2.631924e-10, 6.795037e-10, 1.249644e-09, 
    1.783148e-09, 2.570685e-09, 1.693642e-09, 2.768474e-08, 1.932797e-06, 
    3.861142e-06, 1.104133e-05, 1.025485e-05, 9.686971e-06, 9.098095e-06,
  3.049424e-11, 2.113497e-10, 3.511866e-10, 5.318112e-10, 4.060654e-10, 
    6.249574e-10, 9.648387e-10, 9.12255e-10, 7.174674e-07, 4.212276e-06, 
    6.734731e-06, 6.762358e-06, 7.343368e-06, 5.096552e-06, 5.273285e-06,
  4.949139e-10, 5.680848e-11, 1.739402e-10, 4.662847e-10, 2.560861e-10, 
    1.550771e-10, 5.306891e-10, 4.247977e-07, 3.50459e-06, 8.973387e-06, 
    9.166622e-06, 5.135197e-06, 3.116486e-06, 2.681399e-06, 1.934576e-06,
  5.716058e-10, 2.304731e-11, 2.892088e-10, 3.422378e-10, 5.217772e-11, 
    3.347888e-11, 2.319651e-10, 8.359222e-07, 8.189751e-06, 1.660906e-05, 
    1.226067e-05, 5.313842e-06, 1.394263e-06, 1.05788e-06, 4.516582e-07,
  3.235013e-10, 5.380687e-10, 2.653836e-09, 2.325293e-10, 5.730317e-11, 
    2.66256e-10, 3.255468e-08, 2.531852e-06, 1.908988e-05, 2.931045e-05, 
    1.762932e-05, 5.120964e-06, 1.515878e-06, 1.8201e-06, 6.461909e-06,
  7.635666e-10, 9.043018e-11, 4.683253e-11, 2.241766e-09, 6.230361e-09, 
    4.398066e-09, 9.686448e-08, 7.936106e-07, 1.627072e-06, 6.199886e-07, 
    1.041786e-06, 2.520001e-06, 3.527967e-06, 2.247542e-06, 2.228369e-06,
  4.080241e-12, 6.515497e-12, 3.166938e-11, 4.161153e-11, 9.781956e-11, 
    1.222159e-10, 7.798685e-08, 3.462888e-07, 2.15869e-06, 2.818043e-06, 
    2.145474e-06, 2.152691e-06, 2.699592e-06, 2.073025e-06, 2.814424e-06,
  8.286892e-25, 9.062031e-25, 2.815169e-25, 3.100252e-25, 5.350229e-12, 
    1.071857e-11, 7.029566e-10, 3.572283e-07, 2.296034e-06, 2.537384e-06, 
    2.664163e-06, 1.57749e-06, 2.158028e-06, 1.857479e-06, 2.442567e-06,
  2.299644e-25, 1.294431e-25, 1.060132e-25, 1.094897e-25, 1.082755e-25, 
    1.622024e-25, 5.602478e-11, 1.861167e-08, 1.64949e-06, 4.130895e-06, 
    3.064593e-06, 2.847665e-06, 1.961138e-06, 1.329367e-06, 1.116613e-06,
  1.416584e-25, 1.493452e-25, 1.086282e-25, 8.637575e-26, 1.284478e-25, 
    8.003071e-26, 1.339941e-25, 4.573165e-10, 8.434991e-07, 4.970887e-06, 
    3.435447e-06, 3.52438e-06, 2.205624e-06, 2.210147e-06, 2.2223e-06,
  1.613015e-25, 1.643474e-25, 1.63102e-25, 8.913493e-26, 1.006068e-25, 
    1.210265e-25, 1.407593e-25, 8.266578e-11, 1.05201e-08, 2.536012e-06, 
    3.600947e-06, 4.091349e-06, 3.934107e-06, 2.822469e-06, 4.133443e-06,
  1.360635e-25, 1.041575e-25, 1.160651e-25, 1.139738e-25, 1.166723e-25, 
    1.292389e-25, 1.211967e-14, 2.987703e-14, 5.893846e-10, 3.749842e-08, 
    2.412141e-06, 5.566395e-06, 4.799472e-06, 4.443722e-06, 5.009133e-06,
  4.672315e-26, 6.161107e-26, 6.148976e-26, 6.990611e-26, 1.266473e-25, 
    1.035946e-25, 1.287946e-25, 9.178198e-14, 3.728427e-14, 1.674524e-09, 
    7.56146e-07, 2.629328e-06, 7.486438e-06, 6.192809e-06, 5.429411e-06,
  4.706707e-26, 4.761207e-26, 5.123368e-26, 5.3627e-26, 7.129605e-17, 
    4.897669e-26, 5.642039e-26, 8.294049e-14, 1.645992e-13, 5.99566e-11, 
    2.483505e-09, 7.303355e-07, 5.277611e-06, 6.585292e-06, 7.110245e-06,
  1.361631e-17, 1.358989e-26, 3.861753e-27, 3.730208e-13, 7.502862e-12, 
    8.23219e-12, 2.826353e-13, 2.638783e-13, 5.201076e-13, 1.366379e-13, 
    1.50359e-11, 2.118506e-08, 1.6789e-06, 7.809133e-06, 5.221887e-06,
  2.262511e-10, 2.252681e-09, 2.38603e-08, 1.425361e-07, 8.9459e-07, 
    3.990639e-06, 4.374983e-06, 4.710298e-06, 9.525557e-06, 7.383115e-06, 
    7.598528e-06, 8.232812e-06, 7.983215e-06, 8.416226e-06, 6.471547e-06,
  5.272536e-12, 8.177042e-12, 4.783663e-10, 8.412582e-10, 2.945876e-09, 
    1.59527e-07, 3.064844e-07, 2.749463e-06, 3.452939e-06, 3.497784e-06, 
    3.117379e-06, 3.39544e-06, 4.606638e-06, 4.815067e-06, 3.386262e-06,
  1.364977e-14, 3.072542e-15, 4.302269e-14, 3.993683e-12, 2.435134e-10, 
    4.102292e-10, 2.552508e-10, 1.618207e-09, 5.018614e-08, 2.082438e-07, 
    1.332262e-06, 1.086179e-06, 2.954964e-06, 3.194208e-06, 2.328964e-06,
  3.878199e-12, 1.36248e-15, 3.294379e-22, 1.261402e-22, 9.2008e-23, 
    4.816199e-12, 5.608739e-12, 9.716584e-11, 1.885008e-09, 4.235786e-09, 
    1.701194e-08, 6.058859e-07, 1.079363e-06, 4.411638e-07, 1.758033e-06,
  2.008405e-10, 1.613659e-14, 2.072654e-22, 1.638096e-22, 1.146141e-22, 
    7.370095e-23, 1.109319e-22, 6.889192e-23, 4.385526e-18, 3.83183e-12, 
    3.421446e-10, 1.26071e-08, 9.019672e-08, 1.01417e-06, 5.957609e-07,
  3.033725e-10, 8.122019e-14, 3.299282e-17, 1.25619e-22, 8.242296e-23, 
    4.323276e-23, 3.561072e-23, 2.538958e-23, 5.331628e-23, 3.646417e-23, 
    4.83472e-17, 1.957405e-13, 1.373721e-09, 1.952735e-08, 3.102815e-09,
  3.376776e-11, 2.62962e-13, 1.090825e-22, 5.465514e-23, 4.097961e-23, 
    3.991855e-23, 1.176937e-23, 2.348787e-14, 5.404961e-24, 8.286062e-24, 
    1.109282e-23, 4.20786e-16, 5.366157e-14, 4.596967e-12, 4.601294e-09,
  1.628043e-10, 1.785059e-11, 5.000615e-17, 2.922983e-20, 2.694294e-23, 
    8.778853e-24, 3.679724e-24, 8.48144e-25, 2.679686e-25, 1.575208e-11, 
    1.33398e-11, 5.816893e-10, 5.401161e-11, 1.288253e-10, 1.537814e-10,
  1.700614e-09, 2.443971e-11, 5.333845e-12, 3.763919e-23, 1.406229e-23, 
    4.135529e-24, 1.736041e-24, 5.127713e-25, 8.394386e-14, 5.097953e-10, 
    3.275376e-09, 1.391097e-08, 2.868124e-08, 6.958916e-09, 1.791192e-08,
  3.635185e-12, 9.896632e-12, 1.065211e-16, 9.6806e-24, 1.09867e-23, 
    2.534146e-24, 3.658795e-25, 9.319316e-26, 2.635554e-11, 1.708794e-10, 
    5.59835e-12, 1.983811e-10, 3.831888e-08, 2.511104e-07, 2.004131e-07,
  4.335621e-06, 5.334516e-06, 5.13907e-06, 2.47702e-06, 4.603632e-06, 
    4.581654e-06, 5.116868e-06, 4.989478e-06, 5.633146e-06, 9.407523e-06, 
    5.22043e-06, 4.291069e-06, 5.866472e-06, 4.597554e-06, 5.720382e-06,
  5.610344e-06, 3.592522e-06, 2.742027e-06, 8.545952e-07, 9.873449e-07, 
    2.891531e-06, 1.66529e-06, 1.686586e-06, 5.037433e-06, 1.146054e-05, 
    9.436942e-06, 1.035464e-05, 9.085274e-06, 5.848044e-06, 4.183186e-06,
  4.145586e-06, 3.942276e-06, 1.944259e-06, 5.795119e-07, 5.706843e-07, 
    1.853919e-06, 2.744126e-06, 4.162323e-06, 5.788129e-06, 8.636699e-06, 
    1.157636e-05, 1.278249e-05, 1.076495e-05, 5.696266e-06, 8.760127e-06,
  5.22524e-06, 3.580611e-06, 1.172718e-06, 1.237213e-06, 1.79236e-07, 
    5.325323e-09, 1.429517e-06, 4.05993e-06, 7.063412e-06, 9.056856e-06, 
    7.81573e-06, 8.900777e-06, 4.712611e-06, 8.609186e-06, 7.129469e-06,
  4.486218e-06, 3.972766e-06, 5.764005e-07, 1.367517e-06, 5.507006e-07, 
    1.156862e-08, 2.318111e-07, 2.500461e-06, 4.363284e-06, 5.471878e-06, 
    1.039183e-05, 6.262863e-06, 2.704059e-06, 7.048095e-06, 8.994804e-06,
  6.993332e-06, 5.484019e-06, 1.157173e-06, 1.574126e-07, 7.32189e-09, 
    4.828846e-09, 3.778836e-09, 1.698647e-06, 3.039307e-06, 8.403117e-06, 
    1.065001e-05, 7.13477e-06, 3.916407e-06, 3.593739e-06, 6.125515e-06,
  5.86394e-06, 7.520824e-06, 2.611191e-06, 2.64278e-08, 2.001244e-09, 
    1.84032e-09, 5.534913e-09, 1.240807e-06, 3.672521e-06, 8.931435e-06, 
    1.22751e-05, 4.427814e-06, 2.921728e-06, 5.187489e-06, 4.868058e-06,
  5.15087e-06, 5.793859e-06, 2.336457e-06, 1.16366e-06, 7.555023e-09, 
    8.837266e-10, 4.762691e-09, 1.061998e-06, 4.100707e-06, 1.530745e-05, 
    1.3466e-05, 4.857628e-06, 4.173909e-06, 3.392453e-06, 5.893285e-06,
  1.076514e-05, 7.162809e-06, 6.589233e-07, 1.316852e-06, 4.460489e-07, 
    7.007097e-09, 1.3478e-08, 2.121457e-06, 8.976172e-06, 1.900563e-05, 
    1.271188e-05, 5.641479e-06, 4.91632e-06, 7.89697e-06, 9.457264e-06,
  8.039012e-06, 8.493168e-06, 5.815466e-06, 1.418782e-06, 3.297645e-07, 
    2.702864e-08, 8.040077e-09, 4.333256e-06, 1.516049e-05, 2.283322e-05, 
    1.239354e-05, 3.124337e-06, 5.633113e-06, 8.306665e-06, 9.519436e-06,
  1.324455e-05, 1.18504e-05, 8.128233e-06, 1.52903e-05, 9.579503e-05, 
    7.517156e-05, 4.911681e-05, 5.844796e-05, 6.918309e-05, 4.889059e-05, 
    3.382325e-05, 8.285917e-05, 0.0001279805, 0.00020948, 0.0001958905,
  1.321131e-05, 3.005086e-06, 5.167377e-06, 9.347606e-06, 8.868423e-05, 
    7.318717e-05, 5.424425e-05, 3.493514e-05, 4.984836e-05, 3.594099e-05, 
    3.453749e-05, 6.431022e-05, 0.0002178785, 0.0001638339, 0.000165347,
  8.807838e-06, 8.746712e-06, 2.551495e-06, 5.928606e-06, 7.24989e-05, 
    5.939884e-05, 6.751737e-05, 5.069417e-05, 3.458743e-05, 2.734674e-05, 
    4.152705e-05, 0.0001262711, 0.0002395971, 0.000153566, 0.0001178579,
  1.118794e-05, 9.721344e-06, 3.53488e-06, 4.183694e-06, 6.398753e-06, 
    6.088591e-05, 5.704337e-05, 3.829191e-05, 2.002232e-05, 1.798043e-05, 
    6.994598e-05, 0.0001977215, 0.0001206296, 9.824399e-05, 6.767914e-05,
  1.184918e-05, 1.122005e-05, 3.326511e-06, 4.056183e-06, 3.14265e-06, 
    3.722632e-06, 4.500271e-05, 2.452253e-05, 9.93701e-06, 3.019557e-05, 
    0.0001258899, 0.0001716144, 9.539705e-05, 0.0001072302, 3.247353e-05,
  5.340393e-06, 6.875144e-06, 8.862381e-06, 3.966186e-06, 3.785951e-06, 
    3.722759e-06, 1.118056e-06, 1.29489e-05, 1.64381e-05, 5.872529e-05, 
    0.000161375, 0.0001570783, 6.985628e-05, 0.0001242237, 5.16758e-05,
  4.995206e-06, 8.545195e-06, 1.031767e-05, 7.391817e-06, 3.467585e-06, 
    4.10758e-06, 1.031889e-06, 2.756208e-06, 2.433272e-05, 9.273733e-05, 
    0.0001227656, 9.47535e-05, 5.570599e-05, 5.411588e-05, 7.500554e-05,
  8.049842e-06, 9.721495e-06, 9.53515e-06, 8.275522e-06, 4.726116e-06, 
    3.308513e-06, 9.701702e-07, 2.900909e-06, 2.896061e-05, 7.609562e-05, 
    7.244837e-05, 4.493576e-05, 2.928121e-05, 3.345558e-05, 6.880389e-05,
  1.975589e-05, 1.593165e-05, 9.621803e-06, 1.25883e-05, 1.055852e-05, 
    2.058198e-06, 5.426136e-07, 2.431377e-06, 2.069898e-05, 4.371539e-05, 
    5.246605e-05, 3.354272e-05, 3.997845e-05, 4.557433e-05, 3.329653e-05,
  1.932709e-05, 2.456355e-05, 1.679599e-05, 9.967988e-06, 3.983677e-06, 
    2.019984e-06, 1.576216e-06, 3.566514e-06, 1.235533e-05, 3.272618e-05, 
    4.350053e-05, 3.76645e-05, 4.943044e-05, 4.220468e-05, 3.266888e-05 ;

 sftlf =
  0.1986115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.9611561, 0.1583273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7949425, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.7552791, 0.2484612, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 0.9872221, 0.4156101, 0.04560489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 0.8345782, 0.2958934, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.7792858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 0.9990003, 0.3505592, 0.06537855, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 0.8140894, 0.2409153, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 0.9453563, 0.02902743, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  1.522432, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  122.465, 2.830728, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  113.0215, 29.31339, 0.004701966, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  140.0874, 33.71546, 1.141547, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  141.9684, 87.21121, 14.52402, 0.1304746, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  165.7051, 185.2302, 111.1391, 5.227489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  172.6293, 232.1111, 238.8028, 89.74486, 0.6524738, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  149.5705, 217.5222, 183.4477, 142.7244, 6.651272, 0.2006134, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  253.9191, 270.7406, 160.8987, 135.4378, 83.93595, 3.422685, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  248.2018, 381.5977, 396.3867, 296.0411, 147.8827, 85.51294, 0.2661929, 0, 
    0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
