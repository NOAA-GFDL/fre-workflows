netcdf \00010101.atmos_daily.tile6.pv350K {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pv350K(time, grid_yt, grid_xt) ;
		pv350K:_FillValue = -1.e+10f ;
		pv350K:missing_value = -1.e+10f ;
		pv350K:units = "(K m**2) / (kg s)" ;
		pv350K:long_name = "350-K potential vorticity; needs x350 scaling" ;
		pv350K:cell_methods = "time: mean" ;
		pv350K:time_avg_info = "average_T1,average_T2,average_DT" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:11 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile6.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile6.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pv350K =
  -1.192704e-08, -1.222038e-08, -1.078178e-08, -9.503952e-09, -8.829477e-09, 
    -8.485541e-09, -8.530437e-09, -8.713566e-09, -9.092493e-09, 
    -9.520386e-09, -1.009853e-08, -1.086563e-08, -1.206397e-08, 
    -1.345365e-08, -1.499199e-08,
  -1.174462e-08, -1.219739e-08, -1.247998e-08, -1.118978e-08, -1.037073e-08, 
    -9.610524e-09, -9.376217e-09, -9.448387e-09, -9.839317e-09, 
    -1.043297e-08, -1.136466e-08, -1.220629e-08, -1.332611e-08, 
    -1.437819e-08, -1.599197e-08,
  -1.229698e-08, -1.200954e-08, -1.23332e-08, -1.265972e-08, -1.18147e-08, 
    -1.116237e-08, -1.057192e-08, -1.030033e-08, -1.046377e-08, 
    -1.097515e-08, -1.172085e-08, -1.269523e-08, -1.396637e-08, 
    -1.517626e-08, -1.643866e-08,
  -1.401007e-08, -1.29521e-08, -1.24328e-08, -1.273431e-08, -1.253714e-08, 
    -1.22151e-08, -1.175604e-08, -1.160744e-08, -1.147456e-08, -1.184564e-08, 
    -1.249285e-08, -1.332388e-08, -1.438905e-08, -1.574113e-08, -1.683406e-08,
  -1.595797e-08, -1.5145e-08, -1.354593e-08, -1.323775e-08, -1.341494e-08, 
    -1.262324e-08, -1.24976e-08, -1.219801e-08, -1.251226e-08, -1.262002e-08, 
    -1.310445e-08, -1.364056e-08, -1.429177e-08, -1.517749e-08, -1.638214e-08,
  -1.907113e-08, -1.763759e-08, -1.582922e-08, -1.429721e-08, -1.411816e-08, 
    -1.410577e-08, -1.295866e-08, -1.268698e-08, -1.258077e-08, 
    -1.324416e-08, -1.338398e-08, -1.405036e-08, -1.477228e-08, 
    -1.558022e-08, -1.654772e-08,
  -2.293096e-08, -2.083426e-08, -1.881268e-08, -1.652935e-08, -1.489401e-08, 
    -1.470345e-08, -1.453059e-08, -1.339385e-08, -1.282335e-08, 
    -1.306837e-08, -1.390151e-08, -1.430934e-08, -1.519975e-08, 
    -1.597719e-08, -1.658424e-08,
  -2.633989e-08, -2.50031e-08, -2.262027e-08, -1.986227e-08, -1.747393e-08, 
    -1.559918e-08, -1.518487e-08, -1.489009e-08, -1.388096e-08, 
    -1.312007e-08, -1.338868e-08, -1.440946e-08, -1.485548e-08, 
    -1.545989e-08, -1.584127e-08,
  -2.857653e-08, -2.803074e-08, -2.68078e-08, -2.40934e-08, -2.08355e-08, 
    -1.825718e-08, -1.618561e-08, -1.550399e-08, -1.496244e-08, 
    -1.398832e-08, -1.338497e-08, -1.342505e-08, -1.441275e-08, 
    -1.473316e-08, -1.503034e-08,
  -2.85782e-08, -2.99697e-08, -2.95416e-08, -2.837212e-08, -2.504207e-08, 
    -2.168875e-08, -1.924404e-08, -1.714704e-08, -1.574132e-08, 
    -1.518949e-08, -1.416444e-08, -1.371535e-08, -1.347217e-08, 
    -1.452983e-08, -1.458085e-08,
  -1.06172e-08, -9.427266e-09, -8.791789e-09, -8.036113e-09, -7.511957e-09, 
    -6.963967e-09, -6.562472e-09, -6.315294e-09, -6.238531e-09, 
    -6.256825e-09, -6.13949e-09, -6.340084e-09, -6.621415e-09, -7.290641e-09, 
    -8.037012e-09,
  -1.166864e-08, -1.053073e-08, -9.932638e-09, -9.522641e-09, -9.065614e-09, 
    -8.612483e-09, -8.131812e-09, -7.652068e-09, -7.364786e-09, 
    -7.059134e-09, -7.025638e-09, -7.205597e-09, -7.807333e-09, 
    -8.814868e-09, -1.008048e-08,
  -1.343823e-08, -1.157975e-08, -1.050418e-08, -1.011505e-08, -9.911037e-09, 
    -9.674742e-09, -9.427628e-09, -9.09862e-09, -8.756867e-09, -8.518104e-09, 
    -8.302586e-09, -8.582127e-09, -9.285978e-09, -1.039497e-08, -1.13955e-08,
  -1.690183e-08, -1.36093e-08, -1.206393e-08, -1.07597e-08, -1.031994e-08, 
    -1.023542e-08, -1.028987e-08, -1.026112e-08, -1.014042e-08, 
    -9.977416e-09, -1.002192e-08, -1.043463e-08, -1.116315e-08, 
    -1.196338e-08, -1.241638e-08,
  -1.981755e-08, -1.757602e-08, -1.483313e-08, -1.290197e-08, -1.138531e-08, 
    -1.076847e-08, -1.055975e-08, -1.069028e-08, -1.083019e-08, -1.1076e-08, 
    -1.154559e-08, -1.212183e-08, -1.276519e-08, -1.316765e-08, -1.406799e-08,
  -2.011654e-08, -2.041042e-08, -1.850769e-08, -1.668425e-08, -1.441193e-08, 
    -1.294603e-08, -1.199723e-08, -1.177946e-08, -1.184864e-08, 
    -1.224471e-08, -1.269109e-08, -1.336614e-08, -1.396324e-08, 
    -1.492219e-08, -1.612337e-08,
  -2.040056e-08, -2.031884e-08, -1.970767e-08, -1.921168e-08, -1.775493e-08, 
    -1.634503e-08, -1.510133e-08, -1.422233e-08, -1.390691e-08, 
    -1.401944e-08, -1.442388e-08, -1.505518e-08, -1.593785e-08, 
    -1.696977e-08, -1.812901e-08,
  -2.083943e-08, -2.02062e-08, -1.960082e-08, -1.936006e-08, -1.905165e-08, 
    -1.825672e-08, -1.748483e-08, -1.672796e-08, -1.623268e-08, 
    -1.617418e-08, -1.658618e-08, -1.722408e-08, -1.818522e-08, 
    -1.911309e-08, -1.981338e-08,
  -2.190034e-08, -2.062102e-08, -1.988252e-08, -1.918619e-08, -1.901055e-08, 
    -1.898391e-08, -1.863283e-08, -1.84513e-08, -1.825777e-08, -1.838682e-08, 
    -1.874367e-08, -1.929481e-08, -1.981947e-08, -2.013298e-08, -1.979171e-08,
  -2.306816e-08, -2.143764e-08, -2.062637e-08, -1.967098e-08, -1.886619e-08, 
    -1.870233e-08, -1.87042e-08, -1.862796e-08, -1.861009e-08, -1.877743e-08, 
    -1.898657e-08, -1.923678e-08, -1.937948e-08, -1.911418e-08, -1.905345e-08,
  -3.411441e-09, -3.125722e-09, -3.129671e-09, -3.040129e-09, -2.879462e-09, 
    -2.674092e-09, -2.57309e-09, -2.598999e-09, -2.770844e-09, -3.018332e-09, 
    -3.519609e-09, -4.4782e-09, -5.993643e-09, -7.510624e-09, -8.837516e-09,
  -3.992332e-09, -3.498113e-09, -3.365766e-09, -3.29358e-09, -3.250978e-09, 
    -3.167625e-09, -3.083386e-09, -3.108269e-09, -3.282304e-09, 
    -3.448232e-09, -3.847743e-09, -4.724678e-09, -6.051505e-09, -7.44131e-09, 
    -8.776542e-09,
  -4.968137e-09, -4.25484e-09, -3.901691e-09, -3.718467e-09, -3.669846e-09, 
    -3.665161e-09, -3.682569e-09, -3.761618e-09, -3.943029e-09, 
    -4.204094e-09, -4.613075e-09, -5.352859e-09, -6.589484e-09, 
    -7.863768e-09, -9.142504e-09,
  -6.21223e-09, -5.409722e-09, -4.872172e-09, -4.470158e-09, -4.295225e-09, 
    -4.290294e-09, -4.318729e-09, -4.386281e-09, -4.546877e-09, 
    -4.876553e-09, -5.317681e-09, -5.896548e-09, -6.899467e-09, 
    -8.187867e-09, -9.634874e-09,
  -7.709414e-09, -6.855882e-09, -6.269997e-09, -5.692605e-09, -5.226255e-09, 
    -4.924634e-09, -4.918011e-09, -5.047002e-09, -5.129726e-09, 
    -5.365237e-09, -5.809498e-09, -6.289675e-09, -7.23226e-09, -8.541537e-09, 
    -9.716452e-09,
  -9.463699e-09, -8.407107e-09, -7.869867e-09, -7.322008e-09, -6.808079e-09, 
    -6.471098e-09, -6.300485e-09, -6.326217e-09, -6.479e-09, -6.687496e-09, 
    -6.977414e-09, -7.327726e-09, -7.955054e-09, -8.955894e-09, -9.844773e-09,
  -1.144547e-08, -1.005168e-08, -9.310984e-09, -8.92372e-09, -8.621325e-09, 
    -8.335647e-09, -8.114172e-09, -8.054319e-09, -8.100368e-09, 
    -8.175457e-09, -8.306345e-09, -8.540355e-09, -8.98833e-09, -9.955399e-09, 
    -1.073459e-08,
  -1.422966e-08, -1.244271e-08, -1.131065e-08, -1.036994e-08, -9.97633e-09, 
    -9.836241e-09, -9.947718e-09, -1.006555e-08, -1.030299e-08, 
    -1.047799e-08, -1.05966e-08, -1.078086e-08, -1.123743e-08, -1.189862e-08, 
    -1.252399e-08,
  -1.725169e-08, -1.550777e-08, -1.42898e-08, -1.310212e-08, -1.237681e-08, 
    -1.165826e-08, -1.130186e-08, -1.124985e-08, -1.142979e-08, 
    -1.161822e-08, -1.196763e-08, -1.226569e-08, -1.265251e-08, 
    -1.304185e-08, -1.368733e-08,
  -1.914508e-08, -1.848023e-08, -1.73584e-08, -1.630266e-08, -1.555745e-08, 
    -1.506661e-08, -1.466856e-08, -1.389333e-08, -1.355563e-08, 
    -1.331444e-08, -1.337233e-08, -1.347724e-08, -1.360646e-08, 
    -1.370524e-08, -1.412789e-08,
  -1.762029e-09, -1.731263e-09, -2.059218e-09, -2.652036e-09, -3.68292e-09, 
    -4.919435e-09, -6.452634e-09, -8.556083e-09, -1.140541e-08, -1.49254e-08, 
    -1.816217e-08, -2.164633e-08, -2.506645e-08, -2.92162e-08, -3.109058e-08,
  -2.040443e-09, -2.068578e-09, -2.27896e-09, -2.537666e-09, -3.253474e-09, 
    -4.43633e-09, -5.930152e-09, -7.714725e-09, -9.970561e-09, -1.303732e-08, 
    -1.631366e-08, -1.948055e-08, -2.286835e-08, -2.73946e-08, -2.996683e-08,
  -2.386308e-09, -2.362954e-09, -2.459924e-09, -2.615772e-09, -3.189096e-09, 
    -4.065179e-09, -5.443365e-09, -7.172128e-09, -9.01188e-09, -1.147012e-08, 
    -1.436894e-08, -1.755143e-08, -2.0616e-08, -2.487758e-08, -2.869789e-08,
  -2.649033e-09, -2.535894e-09, -2.716556e-09, -2.757319e-09, -3.132222e-09, 
    -3.830802e-09, -5.11553e-09, -6.590752e-09, -8.234133e-09, -1.033132e-08, 
    -1.273138e-08, -1.569425e-08, -1.880864e-08, -2.228924e-08, -2.648147e-08,
  -3.343209e-09, -3.00519e-09, -2.903656e-09, -2.989099e-09, -3.327127e-09, 
    -3.812657e-09, -4.749152e-09, -6.011089e-09, -7.615172e-09, 
    -9.332133e-09, -1.157338e-08, -1.396833e-08, -1.680062e-08, 
    -1.984996e-08, -2.361987e-08,
  -3.933368e-09, -3.640724e-09, -3.491832e-09, -3.393566e-09, -3.671406e-09, 
    -4.159374e-09, -4.781222e-09, -5.70212e-09, -7.132125e-09, -8.692379e-09, 
    -1.063288e-08, -1.294878e-08, -1.493062e-08, -1.750728e-08, -2.082979e-08,
  -5.868358e-09, -4.692578e-09, -4.292112e-09, -4.323897e-09, -4.384469e-09, 
    -4.421479e-09, -4.787623e-09, -5.374594e-09, -6.574418e-09, 
    -8.003215e-09, -9.757746e-09, -1.231041e-08, -1.416457e-08, 
    -1.565687e-08, -1.8604e-08,
  -8.532611e-09, -6.947412e-09, -6.000302e-09, -5.389403e-09, -5.154917e-09, 
    -5.193566e-09, -5.191173e-09, -5.569178e-09, -6.410681e-09, 
    -7.711744e-09, -9.158647e-09, -1.177227e-08, -1.35507e-08, -1.471435e-08, 
    -1.68234e-08,
  -1.187395e-08, -9.779247e-09, -8.546335e-09, -7.260387e-09, -6.502844e-09, 
    -6.16237e-09, -6.124998e-09, -6.383372e-09, -6.974008e-09, -8.068184e-09, 
    -8.953033e-09, -1.091255e-08, -1.277395e-08, -1.380159e-08, -1.601254e-08,
  -1.612431e-08, -1.374318e-08, -1.201522e-08, -1.029966e-08, -9.086954e-09, 
    -8.054866e-09, -7.447444e-09, -7.246781e-09, -7.645681e-09, 
    -8.326732e-09, -8.872936e-09, -1.041894e-08, -1.17667e-08, -1.263343e-08, 
    -1.435114e-08,
  -1.538845e-08, -1.580991e-08, -1.636083e-08, -1.696874e-08, -1.746025e-08, 
    -1.77647e-08, -1.76819e-08, -1.734305e-08, -1.611364e-08, -1.482699e-08, 
    -1.351997e-08, -1.183864e-08, -1.03089e-08, -8.869428e-09, -8.045259e-09,
  -1.630689e-08, -1.67976e-08, -1.741575e-08, -1.803645e-08, -1.883113e-08, 
    -1.942323e-08, -1.968656e-08, -1.930423e-08, -1.866733e-08, 
    -1.767561e-08, -1.615515e-08, -1.468739e-08, -1.286163e-08, 
    -1.122906e-08, -9.789134e-09,
  -1.789953e-08, -1.841107e-08, -1.893844e-08, -1.945896e-08, -2.032272e-08, 
    -2.1151e-08, -2.164538e-08, -2.181176e-08, -2.134882e-08, -2.069673e-08, 
    -1.970695e-08, -1.806649e-08, -1.627226e-08, -1.42753e-08, -1.233867e-08,
  -1.812221e-08, -1.918615e-08, -2.015098e-08, -2.062164e-08, -2.124882e-08, 
    -2.204917e-08, -2.271948e-08, -2.281286e-08, -2.299231e-08, 
    -2.284327e-08, -2.215366e-08, -2.122445e-08, -1.928074e-08, 
    -1.712535e-08, -1.503906e-08,
  -1.629757e-08, -1.855731e-08, -2.018527e-08, -2.114061e-08, -2.202042e-08, 
    -2.302569e-08, -2.357001e-08, -2.364945e-08, -2.396862e-08, 
    -2.423604e-08, -2.432083e-08, -2.370741e-08, -2.233475e-08, 
    -2.028104e-08, -1.74992e-08,
  -1.358176e-08, -1.61342e-08, -1.886704e-08, -2.011455e-08, -2.144421e-08, 
    -2.268864e-08, -2.382408e-08, -2.41284e-08, -2.473201e-08, -2.54857e-08, 
    -2.571564e-08, -2.629952e-08, -2.567209e-08, -2.382894e-08, -2.146232e-08,
  -1.19377e-08, -1.457274e-08, -1.675844e-08, -1.880808e-08, -2.063425e-08, 
    -2.228762e-08, -2.364727e-08, -2.453288e-08, -2.512385e-08, 
    -2.621881e-08, -2.700082e-08, -2.71132e-08, -2.793974e-08, -2.748222e-08, 
    -2.473823e-08,
  -1.069804e-08, -1.219546e-08, -1.349364e-08, -1.616585e-08, -1.829855e-08, 
    -2.067154e-08, -2.284348e-08, -2.417177e-08, -2.491433e-08, -2.57384e-08, 
    -2.713423e-08, -2.812216e-08, -2.786947e-08, -2.866751e-08, -2.82094e-08,
  -9.498668e-09, -1.001148e-08, -1.15581e-08, -1.357415e-08, -1.5092e-08, 
    -1.717712e-08, -2.005632e-08, -2.285682e-08, -2.497483e-08, 
    -2.608629e-08, -2.658361e-08, -2.756249e-08, -2.836167e-08, 
    -2.775235e-08, -2.798151e-08,
  -8.259651e-09, -8.624921e-09, -9.257329e-09, -1.019749e-08, -1.158492e-08, 
    -1.293004e-08, -1.517068e-08, -1.814845e-08, -2.115737e-08, -2.36447e-08, 
    -2.590019e-08, -2.710287e-08, -2.786359e-08, -2.769756e-08, -2.700545e-08,
  -5.910881e-09, -6.874974e-09, -8.184775e-09, -9.718576e-09, -1.157792e-08, 
    -1.364983e-08, -1.569803e-08, -1.752374e-08, -1.928827e-08, 
    -2.084659e-08, -2.227695e-08, -2.355136e-08, -2.460117e-08, 
    -2.519044e-08, -2.553486e-08,
  -5.526355e-09, -6.140489e-09, -7.363846e-09, -8.692117e-09, -1.030178e-08, 
    -1.228579e-08, -1.436993e-08, -1.638582e-08, -1.832211e-08, 
    -2.010847e-08, -2.174656e-08, -2.336536e-08, -2.465432e-08, 
    -2.557189e-08, -2.626765e-08,
  -5.630947e-09, -5.756022e-09, -6.614513e-09, -7.762788e-09, -9.138334e-09, 
    -1.084197e-08, -1.286134e-08, -1.498642e-08, -1.72238e-08, -1.926944e-08, 
    -2.108773e-08, -2.263144e-08, -2.396928e-08, -2.500655e-08, -2.58074e-08,
  -6.206409e-09, -5.671383e-09, -6.192841e-09, -6.958913e-09, -8.053823e-09, 
    -9.47566e-09, -1.118453e-08, -1.311893e-08, -1.536379e-08, -1.790981e-08, 
    -2.01112e-08, -2.177713e-08, -2.327222e-08, -2.462783e-08, -2.564707e-08,
  -7.862877e-09, -6.369727e-09, -6.078985e-09, -6.492262e-09, -7.260598e-09, 
    -8.277712e-09, -9.662755e-09, -1.137237e-08, -1.328086e-08, 
    -1.570355e-08, -1.841448e-08, -2.074238e-08, -2.252334e-08, 
    -2.390951e-08, -2.508087e-08,
  -1.03058e-08, -8.478361e-09, -7.055758e-09, -6.604814e-09, -6.859544e-09, 
    -7.42558e-09, -8.425697e-09, -9.797949e-09, -1.148895e-08, -1.361377e-08, 
    -1.606459e-08, -1.883807e-08, -2.103125e-08, -2.29756e-08, -2.438441e-08,
  -1.266764e-08, -1.090852e-08, -9.17337e-09, -7.964116e-09, -7.27941e-09, 
    -6.939454e-09, -7.489765e-09, -8.57258e-09, -9.91735e-09, -1.154606e-08, 
    -1.370919e-08, -1.633513e-08, -1.913276e-08, -2.124452e-08, -2.324828e-08,
  -1.520685e-08, -1.310576e-08, -1.123284e-08, -9.881664e-09, -8.83764e-09, 
    -7.898582e-09, -7.197513e-09, -7.798065e-09, -8.801266e-09, -1.00156e-08, 
    -1.165364e-08, -1.378624e-08, -1.631884e-08, -1.915379e-08, -2.138138e-08,
  -1.604813e-08, -1.432178e-08, -1.338136e-08, -1.226122e-08, -1.08494e-08, 
    -9.933113e-09, -8.801612e-09, -7.991853e-09, -7.958515e-09, 
    -8.833974e-09, -1.00458e-08, -1.173972e-08, -1.384642e-08, -1.624158e-08, 
    -1.903953e-08,
  -1.586917e-08, -1.562268e-08, -1.562025e-08, -1.461287e-08, -1.342643e-08, 
    -1.239181e-08, -1.115248e-08, -1.008595e-08, -9.21003e-09, -8.775581e-09, 
    -8.934709e-09, -9.938989e-09, -1.173915e-08, -1.386959e-08, -1.601775e-08,
  -2.125405e-08, -2.201581e-08, -2.305325e-08, -2.387941e-08, -2.398873e-08, 
    -2.441378e-08, -2.436259e-08, -2.426985e-08, -2.398786e-08, 
    -2.364883e-08, -2.332512e-08, -2.279401e-08, -2.227772e-08, 
    -2.164599e-08, -2.083116e-08,
  -2.052131e-08, -2.170074e-08, -2.29541e-08, -2.38731e-08, -2.426392e-08, 
    -2.487151e-08, -2.482154e-08, -2.460353e-08, -2.438525e-08, 
    -2.442071e-08, -2.423573e-08, -2.383766e-08, -2.339016e-08, 
    -2.294119e-08, -2.224276e-08,
  -1.99721e-08, -2.109388e-08, -2.258813e-08, -2.361953e-08, -2.421395e-08, 
    -2.514919e-08, -2.525458e-08, -2.529708e-08, -2.506975e-08, 
    -2.492509e-08, -2.47731e-08, -2.470459e-08, -2.4111e-08, -2.363774e-08, 
    -2.309309e-08,
  -1.910312e-08, -2.008653e-08, -2.168529e-08, -2.297002e-08, -2.382189e-08, 
    -2.483583e-08, -2.538649e-08, -2.578775e-08, -2.569002e-08, 
    -2.575536e-08, -2.548711e-08, -2.534673e-08, -2.52604e-08, -2.503058e-08, 
    -2.428511e-08,
  -1.792791e-08, -1.89724e-08, -2.038581e-08, -2.188716e-08, -2.300777e-08, 
    -2.422362e-08, -2.498283e-08, -2.594507e-08, -2.644183e-08, 
    -2.641772e-08, -2.657275e-08, -2.64042e-08, -2.594467e-08, -2.57295e-08, 
    -2.547834e-08,
  -1.643632e-08, -1.779284e-08, -1.917875e-08, -2.047813e-08, -2.171815e-08, 
    -2.321367e-08, -2.429674e-08, -2.522541e-08, -2.626244e-08, 
    -2.706846e-08, -2.735766e-08, -2.731302e-08, -2.721976e-08, 
    -2.713213e-08, -2.650276e-08,
  -1.500466e-08, -1.626146e-08, -1.782865e-08, -1.917511e-08, -2.033138e-08, 
    -2.161508e-08, -2.305317e-08, -2.449627e-08, -2.543669e-08, 
    -2.649387e-08, -2.750396e-08, -2.807827e-08, -2.832353e-08, 
    -2.824552e-08, -2.845889e-08,
  -1.323443e-08, -1.496346e-08, -1.634123e-08, -1.778494e-08, -1.898736e-08, 
    -2.006695e-08, -2.129158e-08, -2.273272e-08, -2.445329e-08, 
    -2.562428e-08, -2.676101e-08, -2.744549e-08, -2.832422e-08, 
    -2.854418e-08, -2.857882e-08,
  -1.152457e-08, -1.319746e-08, -1.467173e-08, -1.613578e-08, -1.747108e-08, 
    -1.862811e-08, -1.975161e-08, -2.096807e-08, -2.23979e-08, -2.399257e-08, 
    -2.565294e-08, -2.670903e-08, -2.748789e-08, -2.828207e-08, -2.840695e-08,
  -1.005564e-08, -1.14683e-08, -1.292208e-08, -1.431237e-08, -1.57574e-08, 
    -1.701523e-08, -1.813718e-08, -1.929881e-08, -2.032858e-08, -2.17253e-08, 
    -2.311195e-08, -2.480875e-08, -2.604751e-08, -2.711335e-08, -2.801051e-08,
  -2.36433e-08, -2.413471e-08, -2.440121e-08, -2.482839e-08, -2.460125e-08, 
    -2.376545e-08, -2.259055e-08, -2.090108e-08, -1.88495e-08, -1.652346e-08, 
    -1.406119e-08, -1.157767e-08, -9.37022e-09, -7.412757e-09, -5.735268e-09,
  -2.383196e-08, -2.420688e-08, -2.479146e-08, -2.531872e-08, -2.561213e-08, 
    -2.538248e-08, -2.5046e-08, -2.404386e-08, -2.233932e-08, -2.018891e-08, 
    -1.779815e-08, -1.516407e-08, -1.248794e-08, -1.005086e-08, -7.932456e-09,
  -2.396964e-08, -2.417262e-08, -2.438844e-08, -2.505121e-08, -2.536274e-08, 
    -2.511455e-08, -2.480911e-08, -2.457956e-08, -2.40714e-08, -2.294949e-08, 
    -2.109904e-08, -1.876948e-08, -1.613014e-08, -1.336505e-08, -1.095746e-08,
  -2.321137e-08, -2.390688e-08, -2.429014e-08, -2.466696e-08, -2.504772e-08, 
    -2.521168e-08, -2.504476e-08, -2.493208e-08, -2.43851e-08, -2.380733e-08, 
    -2.287042e-08, -2.12905e-08, -1.935628e-08, -1.677732e-08, -1.412073e-08,
  -2.360709e-08, -2.318015e-08, -2.374904e-08, -2.448489e-08, -2.489677e-08, 
    -2.496444e-08, -2.496066e-08, -2.497194e-08, -2.502209e-08, 
    -2.449053e-08, -2.417639e-08, -2.323001e-08, -2.182475e-08, 
    -1.976101e-08, -1.747505e-08,
  -2.428794e-08, -2.353602e-08, -2.333517e-08, -2.375065e-08, -2.436524e-08, 
    -2.486227e-08, -2.497505e-08, -2.474157e-08, -2.475972e-08, -2.46505e-08, 
    -2.44377e-08, -2.43281e-08, -2.369145e-08, -2.235662e-08, -2.031411e-08,
  -2.336935e-08, -2.391631e-08, -2.363083e-08, -2.364319e-08, -2.378765e-08, 
    -2.420286e-08, -2.438625e-08, -2.471518e-08, -2.456169e-08, -2.4271e-08, 
    -2.389312e-08, -2.426715e-08, -2.426543e-08, -2.396221e-08, -2.278649e-08,
  -2.165479e-08, -2.312044e-08, -2.394345e-08, -2.360762e-08, -2.342818e-08, 
    -2.358217e-08, -2.388877e-08, -2.390577e-08, -2.428265e-08, 
    -2.415234e-08, -2.326624e-08, -2.332458e-08, -2.345011e-08, 
    -2.402283e-08, -2.406305e-08,
  -1.95445e-08, -2.070234e-08, -2.291617e-08, -2.389344e-08, -2.357014e-08, 
    -2.316796e-08, -2.32996e-08, -2.341809e-08, -2.362418e-08, -2.391083e-08, 
    -2.354267e-08, -2.297002e-08, -2.275709e-08, -2.320088e-08, -2.400849e-08,
  -1.795495e-08, -1.907209e-08, -2.051074e-08, -2.253396e-08, -2.336111e-08, 
    -2.327272e-08, -2.298191e-08, -2.286721e-08, -2.286004e-08, 
    -2.325171e-08, -2.36198e-08, -2.348609e-08, -2.299005e-08, -2.268275e-08, 
    -2.324195e-08,
  -1.678318e-08, -1.457191e-08, -1.309399e-08, -1.1155e-08, -9.439884e-09, 
    -7.938444e-09, -6.665623e-09, -5.625411e-09, -4.807923e-09, 
    -4.132841e-09, -3.628048e-09, -3.412718e-09, -3.334999e-09, 
    -3.272989e-09, -3.265792e-09,
  -1.985528e-08, -1.781026e-08, -1.611487e-08, -1.415482e-08, -1.217816e-08, 
    -1.027445e-08, -8.603579e-09, -7.24857e-09, -6.171102e-09, -5.270968e-09, 
    -4.523266e-09, -3.966418e-09, -3.703136e-09, -3.620579e-09, -3.587007e-09,
  -2.245746e-08, -2.065374e-08, -1.910089e-08, -1.721815e-08, -1.527936e-08, 
    -1.318877e-08, -1.126187e-08, -9.41334e-09, -7.962655e-09, -6.814109e-09, 
    -5.925481e-09, -5.1366e-09, -4.496225e-09, -4.111898e-09, -3.917937e-09,
  -2.478976e-08, -2.350752e-08, -2.197144e-08, -1.998933e-08, -1.821387e-08, 
    -1.612384e-08, -1.416582e-08, -1.209484e-08, -1.022027e-08, 
    -8.613945e-09, -7.349096e-09, -6.428334e-09, -5.673337e-09, 
    -5.043817e-09, -4.620825e-09,
  -2.600642e-08, -2.548954e-08, -2.450891e-08, -2.303883e-08, -2.111583e-08, 
    -1.903319e-08, -1.700876e-08, -1.504456e-08, -1.303911e-08, 
    -1.116079e-08, -9.470926e-09, -8.04932e-09, -7.043218e-09, -6.221093e-09, 
    -5.576587e-09,
  -2.655033e-08, -2.689627e-08, -2.657912e-08, -2.546914e-08, -2.40831e-08, 
    -2.21313e-08, -1.98723e-08, -1.776758e-08, -1.57611e-08, -1.384867e-08, 
    -1.198416e-08, -1.035356e-08, -8.903508e-09, -7.879913e-09, -7.028111e-09,
  -2.621957e-08, -2.684454e-08, -2.770029e-08, -2.773122e-08, -2.715733e-08, 
    -2.556879e-08, -2.336503e-08, -2.081967e-08, -1.842688e-08, -1.64876e-08, 
    -1.453203e-08, -1.27467e-08, -1.106895e-08, -9.692417e-09, -8.69442e-09,
  -2.557749e-08, -2.610187e-08, -2.671521e-08, -2.731145e-08, -2.800897e-08, 
    -2.795248e-08, -2.687141e-08, -2.456715e-08, -2.181817e-08, 
    -1.915007e-08, -1.718806e-08, -1.53039e-08, -1.349397e-08, -1.182976e-08, 
    -1.049674e-08,
  -2.527175e-08, -2.557741e-08, -2.628032e-08, -2.643157e-08, -2.678057e-08, 
    -2.755533e-08, -2.758568e-08, -2.70128e-08, -2.573758e-08, -2.273218e-08, 
    -1.992634e-08, -1.770326e-08, -1.598671e-08, -1.420111e-08, -1.256729e-08,
  -2.378353e-08, -2.560729e-08, -2.653398e-08, -2.701143e-08, -2.668205e-08, 
    -2.66912e-08, -2.699632e-08, -2.695311e-08, -2.664694e-08, -2.593609e-08, 
    -2.362171e-08, -2.063242e-08, -1.840128e-08, -1.650058e-08, -1.496964e-08,
  -4.641712e-09, -4.391553e-09, -4.462442e-09, -4.529372e-09, -4.785461e-09, 
    -5.157831e-09, -5.770804e-09, -6.41961e-09, -7.018341e-09, -7.658583e-09, 
    -8.436003e-09, -9.309726e-09, -1.043672e-08, -1.208292e-08, -1.430261e-08,
  -5.293654e-09, -4.812336e-09, -4.781124e-09, -4.798244e-09, -5.084333e-09, 
    -5.48873e-09, -6.040496e-09, -6.609856e-09, -7.21348e-09, -7.904117e-09, 
    -8.65149e-09, -9.855153e-09, -1.146214e-08, -1.36849e-08, -1.595871e-08,
  -6.24521e-09, -5.464065e-09, -5.303506e-09, -5.181074e-09, -5.401869e-09, 
    -5.751369e-09, -6.281623e-09, -6.818073e-09, -7.420265e-09, 
    -8.076209e-09, -8.929563e-09, -1.037795e-08, -1.247353e-08, 
    -1.487108e-08, -1.70509e-08,
  -7.494461e-09, -6.369042e-09, -6.012954e-09, -5.653831e-09, -5.689123e-09, 
    -5.967873e-09, -6.481172e-09, -7.056745e-09, -7.642981e-09, 
    -8.285631e-09, -9.294691e-09, -1.095686e-08, -1.292759e-08, 
    -1.509216e-08, -1.718263e-08,
  -9.734129e-09, -8.055423e-09, -7.329943e-09, -6.586293e-09, -6.370858e-09, 
    -6.407997e-09, -6.695393e-09, -7.147017e-09, -7.740162e-09, 
    -8.535452e-09, -9.63672e-09, -1.12967e-08, -1.334697e-08, -1.520737e-08, 
    -1.701806e-08,
  -1.293301e-08, -1.074771e-08, -9.447401e-09, -8.167898e-09, -7.413058e-09, 
    -7.011923e-09, -7.076161e-09, -7.431479e-09, -7.964669e-09, 
    -8.552879e-09, -9.504841e-09, -1.116635e-08, -1.303494e-08, -1.48398e-08, 
    -1.659928e-08,
  -1.693851e-08, -1.491154e-08, -1.320939e-08, -1.13132e-08, -9.65891e-09, 
    -8.646788e-09, -8.150826e-09, -8.049422e-09, -8.314556e-09, 
    -8.831814e-09, -9.622028e-09, -1.085626e-08, -1.261247e-08, 
    -1.441116e-08, -1.653964e-08,
  -2.005784e-08, -1.852229e-08, -1.723306e-08, -1.556979e-08, -1.359041e-08, 
    -1.154363e-08, -9.828409e-09, -8.861466e-09, -8.822742e-09, 
    -9.053826e-09, -9.471524e-09, -1.039674e-08, -1.196159e-08, 
    -1.382907e-08, -1.583378e-08,
  -2.310632e-08, -2.187082e-08, -2.056231e-08, -1.90973e-08, -1.773354e-08, 
    -1.595512e-08, -1.384459e-08, -1.181146e-08, -1.031359e-08, 
    -9.648224e-09, -9.936229e-09, -1.037569e-08, -1.11621e-08, -1.279366e-08, 
    -1.484112e-08,
  -2.560308e-08, -2.492471e-08, -2.401776e-08, -2.249508e-08, -2.086657e-08, 
    -1.926204e-08, -1.762746e-08, -1.574821e-08, -1.342e-08, -1.14075e-08, 
    -1.059438e-08, -1.024472e-08, -1.103268e-08, -1.194164e-08, -1.372012e-08,
  -1.054362e-08, -1.206209e-08, -1.328879e-08, -1.485785e-08, -1.591096e-08, 
    -1.667553e-08, -1.711322e-08, -1.749828e-08, -1.834476e-08, 
    -1.945808e-08, -2.022848e-08, -2.098635e-08, -2.155123e-08, 
    -2.167209e-08, -2.14533e-08,
  -1.07124e-08, -1.232964e-08, -1.371605e-08, -1.519544e-08, -1.632298e-08, 
    -1.717459e-08, -1.80125e-08, -1.93787e-08, -2.087328e-08, -2.106515e-08, 
    -2.135218e-08, -2.130697e-08, -2.128454e-08, -2.124823e-08, -2.102475e-08,
  -1.084383e-08, -1.237324e-08, -1.381272e-08, -1.537062e-08, -1.651099e-08, 
    -1.766487e-08, -1.919265e-08, -2.090916e-08, -2.139323e-08, 
    -2.127903e-08, -2.167274e-08, -2.174456e-08, -2.191019e-08, 
    -2.173609e-08, -2.169859e-08,
  -1.090769e-08, -1.251388e-08, -1.408872e-08, -1.560141e-08, -1.683277e-08, 
    -1.844244e-08, -2.012265e-08, -2.117683e-08, -2.10843e-08, -2.174668e-08, 
    -2.295197e-08, -2.400488e-08, -2.458055e-08, -2.442601e-08, -2.391985e-08,
  -1.098745e-08, -1.266327e-08, -1.432586e-08, -1.580003e-08, -1.733449e-08, 
    -1.920525e-08, -2.080202e-08, -2.138217e-08, -2.235104e-08, 
    -2.478544e-08, -2.701612e-08, -2.827448e-08, -2.825251e-08, 
    -2.771133e-08, -2.676265e-08,
  -1.116046e-08, -1.295213e-08, -1.45738e-08, -1.604296e-08, -1.77371e-08, 
    -1.966186e-08, -2.094702e-08, -2.228304e-08, -2.517846e-08, 
    -2.800497e-08, -2.983152e-08, -3.022964e-08, -2.952352e-08, 
    -2.894489e-08, -2.859804e-08,
  -1.130933e-08, -1.312548e-08, -1.466142e-08, -1.613056e-08, -1.79582e-08, 
    -1.980701e-08, -2.1276e-08, -2.340419e-08, -2.637e-08, -2.903728e-08, 
    -3.072724e-08, -3.08812e-08, -2.985206e-08, -2.995489e-08, -2.905314e-08,
  -1.158275e-08, -1.338524e-08, -1.470687e-08, -1.613277e-08, -1.784161e-08, 
    -1.956925e-08, -2.110134e-08, -2.322117e-08, -2.600856e-08, 
    -2.876464e-08, -2.988651e-08, -3.083376e-08, -3.119472e-08, 
    -3.028405e-08, -2.960996e-08,
  -1.179315e-08, -1.345598e-08, -1.463939e-08, -1.59625e-08, -1.751815e-08, 
    -1.903486e-08, -2.045329e-08, -2.222467e-08, -2.504514e-08, 
    -2.716631e-08, -2.860649e-08, -3.031611e-08, -3.067276e-08, 
    -3.051981e-08, -2.999533e-08,
  -1.206434e-08, -1.345795e-08, -1.442309e-08, -1.553333e-08, -1.686082e-08, 
    -1.832989e-08, -1.953987e-08, -2.12092e-08, -2.368891e-08, -2.517244e-08, 
    -2.681049e-08, -2.951322e-08, -3.067626e-08, -3.103506e-08, -3.06686e-08,
  -7.620556e-09, -8.064251e-09, -8.563592e-09, -9.370901e-09, -1.04966e-08, 
    -1.171024e-08, -1.28596e-08, -1.397101e-08, -1.500477e-08, -1.59599e-08, 
    -1.693065e-08, -1.800021e-08, -1.921449e-08, -2.054295e-08, -2.198215e-08,
  -8.779453e-09, -9.21381e-09, -9.910542e-09, -1.089949e-08, -1.19364e-08, 
    -1.302272e-08, -1.410907e-08, -1.512644e-08, -1.60128e-08, -1.692034e-08, 
    -1.783139e-08, -1.893206e-08, -2.022785e-08, -2.169064e-08, -2.315829e-08,
  -9.874461e-09, -1.036105e-08, -1.134195e-08, -1.239722e-08, -1.338358e-08, 
    -1.448428e-08, -1.539076e-08, -1.61698e-08, -1.692028e-08, -1.778193e-08, 
    -1.876554e-08, -1.998958e-08, -2.130528e-08, -2.266502e-08, -2.405592e-08,
  -1.099583e-08, -1.168172e-08, -1.287001e-08, -1.375919e-08, -1.476093e-08, 
    -1.572611e-08, -1.647872e-08, -1.712569e-08, -1.783826e-08, 
    -1.872082e-08, -1.969899e-08, -2.083439e-08, -2.205381e-08, 
    -2.342056e-08, -2.476037e-08,
  -1.211898e-08, -1.304222e-08, -1.402456e-08, -1.482064e-08, -1.576001e-08, 
    -1.662142e-08, -1.719891e-08, -1.788789e-08, -1.870551e-08, 
    -1.959649e-08, -2.062066e-08, -2.174642e-08, -2.2866e-08, -2.398202e-08, 
    -2.508472e-08,
  -1.316165e-08, -1.407776e-08, -1.485949e-08, -1.568088e-08, -1.663321e-08, 
    -1.733547e-08, -1.793355e-08, -1.872997e-08, -1.952067e-08, 
    -2.038949e-08, -2.138266e-08, -2.233173e-08, -2.320826e-08, 
    -2.426911e-08, -2.529328e-08,
  -1.389268e-08, -1.476879e-08, -1.556554e-08, -1.64802e-08, -1.736552e-08, 
    -1.800524e-08, -1.863879e-08, -1.936649e-08, -2.0178e-08, -2.116209e-08, 
    -2.202156e-08, -2.282318e-08, -2.38317e-08, -2.472298e-08, -2.537516e-08,
  -1.432002e-08, -1.526536e-08, -1.615273e-08, -1.706394e-08, -1.810029e-08, 
    -1.883436e-08, -1.959439e-08, -2.060317e-08, -2.140555e-08, 
    -2.208762e-08, -2.273642e-08, -2.351566e-08, -2.403368e-08, 
    -2.464379e-08, -2.52925e-08,
  -1.466842e-08, -1.568729e-08, -1.665752e-08, -1.770276e-08, -1.878351e-08, 
    -1.953733e-08, -2.040291e-08, -2.148217e-08, -2.240733e-08, 
    -2.348607e-08, -2.403986e-08, -2.446367e-08, -2.497991e-08, 
    -2.534988e-08, -2.564234e-08,
  -1.487393e-08, -1.598383e-08, -1.704641e-08, -1.817656e-08, -1.940287e-08, 
    -2.025595e-08, -2.140798e-08, -2.306968e-08, -2.410726e-08, -2.47509e-08, 
    -2.502903e-08, -2.568181e-08, -2.581988e-08, -2.598225e-08, -2.600139e-08,
  -6.242421e-09, -7.414824e-09, -8.56182e-09, -9.777956e-09, -1.109134e-08, 
    -1.24109e-08, -1.373671e-08, -1.504783e-08, -1.642941e-08, -1.77657e-08, 
    -1.916933e-08, -2.05071e-08, -2.163883e-08, -2.278164e-08, -2.382405e-08,
  -6.66686e-09, -7.838272e-09, -8.977048e-09, -1.019428e-08, -1.142194e-08, 
    -1.26501e-08, -1.388332e-08, -1.511981e-08, -1.64407e-08, -1.77924e-08, 
    -1.919736e-08, -2.047571e-08, -2.167342e-08, -2.286102e-08, -2.399393e-08,
  -7.084831e-09, -8.226896e-09, -9.451611e-09, -1.066558e-08, -1.187754e-08, 
    -1.301046e-08, -1.409239e-08, -1.522185e-08, -1.648826e-08, 
    -1.780594e-08, -1.914487e-08, -2.040111e-08, -2.167485e-08, -2.2936e-08, 
    -2.409671e-08,
  -7.477856e-09, -8.675997e-09, -9.949011e-09, -1.118142e-08, -1.234086e-08, 
    -1.339674e-08, -1.434312e-08, -1.539095e-08, -1.657886e-08, 
    -1.781386e-08, -1.910283e-08, -2.038284e-08, -2.173001e-08, -2.30212e-08, 
    -2.426245e-08,
  -8.119255e-09, -9.317278e-09, -1.05967e-08, -1.177864e-08, -1.283386e-08, 
    -1.375565e-08, -1.465688e-08, -1.566637e-08, -1.67648e-08, -1.791898e-08, 
    -1.915999e-08, -2.046236e-08, -2.181412e-08, -2.314269e-08, -2.456341e-08,
  -9.0388e-09, -1.01331e-08, -1.131136e-08, -1.231136e-08, -1.323505e-08, 
    -1.411461e-08, -1.499084e-08, -1.595502e-08, -1.700923e-08, 
    -1.810519e-08, -1.93225e-08, -2.059153e-08, -2.195593e-08, -2.333655e-08, 
    -2.496526e-08,
  -9.932985e-09, -1.093284e-08, -1.191673e-08, -1.27704e-08, -1.364299e-08, 
    -1.448176e-08, -1.532907e-08, -1.631014e-08, -1.732888e-08, 
    -1.841928e-08, -1.958666e-08, -2.080319e-08, -2.213129e-08, 
    -2.351393e-08, -2.537113e-08,
  -1.06289e-08, -1.158611e-08, -1.245622e-08, -1.325728e-08, -1.408486e-08, 
    -1.487834e-08, -1.573714e-08, -1.671109e-08, -1.772487e-08, 
    -1.881868e-08, -1.997044e-08, -2.105082e-08, -2.241364e-08, 
    -2.382741e-08, -2.575075e-08,
  -1.11911e-08, -1.217528e-08, -1.299748e-08, -1.378211e-08, -1.461016e-08, 
    -1.538083e-08, -1.623627e-08, -1.723549e-08, -1.827202e-08, 
    -1.937497e-08, -2.041119e-08, -2.148646e-08, -2.279246e-08, 
    -2.431117e-08, -2.641501e-08,
  -1.174806e-08, -1.275183e-08, -1.356821e-08, -1.439391e-08, -1.516209e-08, 
    -1.591911e-08, -1.68574e-08, -1.788255e-08, -1.889884e-08, -1.997091e-08, 
    -2.096312e-08, -2.199538e-08, -2.336425e-08, -2.495862e-08, -2.686589e-08,
  -1.814757e-08, -1.827032e-08, -1.834017e-08, -1.85751e-08, -1.871921e-08, 
    -1.896304e-08, -1.900168e-08, -1.907104e-08, -1.904703e-08, 
    -1.897008e-08, -1.875015e-08, -1.855041e-08, -1.838691e-08, 
    -1.834584e-08, -1.855332e-08,
  -1.889181e-08, -1.897058e-08, -1.893809e-08, -1.897836e-08, -1.891714e-08, 
    -1.899457e-08, -1.902833e-08, -1.914654e-08, -1.919317e-08, -1.92131e-08, 
    -1.911167e-08, -1.905024e-08, -1.898088e-08, -1.916999e-08, -1.952033e-08,
  -1.965268e-08, -1.952312e-08, -1.965535e-08, -1.961152e-08, -1.944215e-08, 
    -1.940912e-08, -1.942172e-08, -1.954719e-08, -1.957518e-08, 
    -1.958054e-08, -1.959335e-08, -1.965747e-08, -1.97454e-08, -2.001557e-08, 
    -2.038473e-08,
  -2.032926e-08, -2.019486e-08, -2.025042e-08, -2.021346e-08, -2.022204e-08, 
    -2.010627e-08, -2.012449e-08, -2.00905e-08, -2.01264e-08, -2.010106e-08, 
    -2.02385e-08, -2.033863e-08, -2.059464e-08, -2.093789e-08, -2.132398e-08,
  -2.061627e-08, -2.07171e-08, -2.082872e-08, -2.085434e-08, -2.093344e-08, 
    -2.090145e-08, -2.086774e-08, -2.080217e-08, -2.086308e-08, 
    -2.093747e-08, -2.107219e-08, -2.116775e-08, -2.156501e-08, 
    -2.199038e-08, -2.246629e-08,
  -2.041603e-08, -2.097008e-08, -2.119559e-08, -2.128742e-08, -2.135091e-08, 
    -2.147037e-08, -2.147939e-08, -2.156335e-08, -2.155955e-08, 
    -2.168213e-08, -2.18524e-08, -2.210453e-08, -2.256349e-08, -2.307111e-08, 
    -2.351653e-08,
  -2.023025e-08, -2.110436e-08, -2.158235e-08, -2.184532e-08, -2.196475e-08, 
    -2.202314e-08, -2.209114e-08, -2.21703e-08, -2.230726e-08, -2.244295e-08, 
    -2.269364e-08, -2.298072e-08, -2.346345e-08, -2.392694e-08, -2.439874e-08,
  -1.997061e-08, -2.0984e-08, -2.164664e-08, -2.209145e-08, -2.226992e-08, 
    -2.236024e-08, -2.255532e-08, -2.27614e-08, -2.289404e-08, -2.306613e-08, 
    -2.342502e-08, -2.383565e-08, -2.433514e-08, -2.482971e-08, -2.544861e-08,
  -1.970758e-08, -2.093809e-08, -2.16856e-08, -2.223253e-08, -2.262118e-08, 
    -2.289252e-08, -2.31557e-08, -2.338317e-08, -2.356583e-08, -2.385317e-08, 
    -2.425749e-08, -2.464423e-08, -2.510601e-08, -2.570201e-08, -2.63347e-08,
  -1.93421e-08, -2.06972e-08, -2.151112e-08, -2.216467e-08, -2.287559e-08, 
    -2.338124e-08, -2.376432e-08, -2.411941e-08, -2.443138e-08, 
    -2.475844e-08, -2.499447e-08, -2.529464e-08, -2.571634e-08, 
    -2.631769e-08, -2.680266e-08,
  -1.649202e-08, -1.657517e-08, -1.654389e-08, -1.659768e-08, -1.655938e-08, 
    -1.657073e-08, -1.641897e-08, -1.620687e-08, -1.591043e-08, 
    -1.578054e-08, -1.579695e-08, -1.595167e-08, -1.599894e-08, 
    -1.597153e-08, -1.612014e-08,
  -1.668184e-08, -1.660551e-08, -1.660358e-08, -1.6557e-08, -1.663381e-08, 
    -1.666677e-08, -1.66942e-08, -1.652961e-08, -1.624454e-08, -1.582006e-08, 
    -1.564556e-08, -1.567587e-08, -1.573488e-08, -1.574403e-08, -1.568743e-08,
  -1.686202e-08, -1.673308e-08, -1.665618e-08, -1.655182e-08, -1.657275e-08, 
    -1.666637e-08, -1.681829e-08, -1.682105e-08, -1.634481e-08, 
    -1.607048e-08, -1.577935e-08, -1.56322e-08, -1.566113e-08, -1.566857e-08, 
    -1.572853e-08,
  -1.688248e-08, -1.684749e-08, -1.682843e-08, -1.666002e-08, -1.658334e-08, 
    -1.65656e-08, -1.677327e-08, -1.688606e-08, -1.669861e-08, -1.639965e-08, 
    -1.620741e-08, -1.593431e-08, -1.586115e-08, -1.578666e-08, -1.587758e-08,
  -1.704328e-08, -1.69222e-08, -1.706002e-08, -1.699389e-08, -1.683224e-08, 
    -1.669409e-08, -1.691182e-08, -1.706188e-08, -1.7195e-08, -1.684698e-08, 
    -1.677934e-08, -1.636179e-08, -1.625352e-08, -1.616976e-08, -1.617173e-08,
  -1.766212e-08, -1.731379e-08, -1.73519e-08, -1.7491e-08, -1.745601e-08, 
    -1.737801e-08, -1.749183e-08, -1.768449e-08, -1.785471e-08, 
    -1.756943e-08, -1.751882e-08, -1.710414e-08, -1.691142e-08, 
    -1.672403e-08, -1.671363e-08,
  -1.846693e-08, -1.786838e-08, -1.760837e-08, -1.76281e-08, -1.776439e-08, 
    -1.788264e-08, -1.798498e-08, -1.825102e-08, -1.835407e-08, 
    -1.815837e-08, -1.812226e-08, -1.782566e-08, -1.758206e-08, 
    -1.751048e-08, -1.736963e-08,
  -1.929099e-08, -1.86726e-08, -1.816768e-08, -1.788713e-08, -1.784806e-08, 
    -1.791233e-08, -1.806901e-08, -1.83069e-08, -1.852304e-08, -1.853249e-08, 
    -1.860897e-08, -1.860514e-08, -1.836927e-08, -1.834959e-08, -1.804302e-08,
  -2.012791e-08, -1.953057e-08, -1.899572e-08, -1.850969e-08, -1.813952e-08, 
    -1.79681e-08, -1.808935e-08, -1.814855e-08, -1.833764e-08, -1.845744e-08, 
    -1.875468e-08, -1.912347e-08, -1.924024e-08, -1.946024e-08, -1.915506e-08,
  -2.091902e-08, -2.024868e-08, -1.976412e-08, -1.930161e-08, -1.878661e-08, 
    -1.845392e-08, -1.833092e-08, -1.832545e-08, -1.84908e-08, -1.854323e-08, 
    -1.885203e-08, -1.928327e-08, -1.980294e-08, -2.048986e-08, -2.073626e-08,
  -1.635716e-08, -1.590462e-08, -1.570659e-08, -1.563406e-08, -1.513268e-08, 
    -1.438426e-08, -1.405997e-08, -1.359765e-08, -1.327616e-08, 
    -1.346431e-08, -1.335568e-08, -1.332754e-08, -1.329893e-08, 
    -1.346473e-08, -1.365502e-08,
  -1.663607e-08, -1.608769e-08, -1.563888e-08, -1.539012e-08, -1.504702e-08, 
    -1.461432e-08, -1.407206e-08, -1.384864e-08, -1.350665e-08, 
    -1.360231e-08, -1.378796e-08, -1.382732e-08, -1.378225e-08, 
    -1.388666e-08, -1.402407e-08,
  -1.70583e-08, -1.642752e-08, -1.583695e-08, -1.553381e-08, -1.513288e-08, 
    -1.487778e-08, -1.426458e-08, -1.420358e-08, -1.375585e-08, 
    -1.384368e-08, -1.394114e-08, -1.411435e-08, -1.404566e-08, 
    -1.415996e-08, -1.428544e-08,
  -1.75947e-08, -1.664331e-08, -1.604868e-08, -1.54788e-08, -1.503736e-08, 
    -1.482649e-08, -1.450669e-08, -1.460973e-08, -1.394997e-08, 
    -1.402541e-08, -1.393964e-08, -1.425304e-08, -1.421779e-08, 
    -1.431262e-08, -1.435231e-08,
  -1.786944e-08, -1.670963e-08, -1.604662e-08, -1.542003e-08, -1.507616e-08, 
    -1.484072e-08, -1.465429e-08, -1.482308e-08, -1.433676e-08, 
    -1.417607e-08, -1.413696e-08, -1.433256e-08, -1.422459e-08, 
    -1.441982e-08, -1.46088e-08,
  -1.816329e-08, -1.692286e-08, -1.62702e-08, -1.537136e-08, -1.519815e-08, 
    -1.504973e-08, -1.501624e-08, -1.508192e-08, -1.467869e-08, 
    -1.434154e-08, -1.404337e-08, -1.416987e-08, -1.424233e-08, 
    -1.463711e-08, -1.482517e-08,
  -1.820997e-08, -1.714938e-08, -1.67556e-08, -1.551806e-08, -1.544939e-08, 
    -1.537098e-08, -1.536978e-08, -1.558483e-08, -1.501042e-08, 
    -1.462518e-08, -1.413864e-08, -1.427005e-08, -1.435531e-08, 
    -1.486991e-08, -1.503051e-08,
  -1.805062e-08, -1.714785e-08, -1.706549e-08, -1.617772e-08, -1.584827e-08, 
    -1.602153e-08, -1.595703e-08, -1.617722e-08, -1.555392e-08, 
    -1.511179e-08, -1.465722e-08, -1.44377e-08, -1.445948e-08, -1.503575e-08, 
    -1.531036e-08,
  -1.783018e-08, -1.686089e-08, -1.676163e-08, -1.632299e-08, -1.603924e-08, 
    -1.615519e-08, -1.610186e-08, -1.615367e-08, -1.591879e-08, 
    -1.568972e-08, -1.55234e-08, -1.490944e-08, -1.479956e-08, -1.498861e-08, 
    -1.539584e-08,
  -1.796946e-08, -1.709065e-08, -1.676089e-08, -1.638463e-08, -1.602305e-08, 
    -1.625128e-08, -1.6201e-08, -1.630409e-08, -1.605723e-08, -1.613537e-08, 
    -1.60994e-08, -1.565939e-08, -1.54363e-08, -1.524563e-08, -1.540014e-08,
  -1.38698e-08, -1.332158e-08, -1.266769e-08, -1.266558e-08, -1.288422e-08, 
    -1.315929e-08, -1.317726e-08, -1.289144e-08, -1.296558e-08, 
    -1.294613e-08, -1.315291e-08, -1.352943e-08, -1.380574e-08, 
    -1.417117e-08, -1.444985e-08,
  -1.44035e-08, -1.399913e-08, -1.325463e-08, -1.280867e-08, -1.290033e-08, 
    -1.331015e-08, -1.363075e-08, -1.351104e-08, -1.353826e-08, -1.35758e-08, 
    -1.371474e-08, -1.400283e-08, -1.426685e-08, -1.459662e-08, -1.484687e-08,
  -1.519871e-08, -1.42818e-08, -1.375001e-08, -1.320789e-08, -1.299625e-08, 
    -1.328406e-08, -1.373552e-08, -1.386011e-08, -1.381295e-08, 
    -1.386546e-08, -1.391414e-08, -1.40884e-08, -1.451977e-08, -1.482879e-08, 
    -1.515005e-08,
  -1.588741e-08, -1.472177e-08, -1.436469e-08, -1.353794e-08, -1.33557e-08, 
    -1.325726e-08, -1.368319e-08, -1.409046e-08, -1.4119e-08, -1.418059e-08, 
    -1.404622e-08, -1.421532e-08, -1.455924e-08, -1.498132e-08, -1.529766e-08,
  -1.626429e-08, -1.510168e-08, -1.43596e-08, -1.344006e-08, -1.344327e-08, 
    -1.31534e-08, -1.35822e-08, -1.42342e-08, -1.426687e-08, -1.424362e-08, 
    -1.42515e-08, -1.441394e-08, -1.469388e-08, -1.503894e-08, -1.530594e-08,
  -1.659221e-08, -1.524589e-08, -1.433797e-08, -1.337615e-08, -1.34141e-08, 
    -1.327987e-08, -1.388856e-08, -1.428181e-08, -1.431254e-08, 
    -1.439026e-08, -1.454137e-08, -1.463351e-08, -1.481074e-08, 
    -1.498037e-08, -1.528542e-08,
  -1.630482e-08, -1.52027e-08, -1.439606e-08, -1.342652e-08, -1.353524e-08, 
    -1.365416e-08, -1.4052e-08, -1.425984e-08, -1.429636e-08, -1.449878e-08, 
    -1.46441e-08, -1.473992e-08, -1.486486e-08, -1.505825e-08, -1.535567e-08,
  -1.611755e-08, -1.514739e-08, -1.459613e-08, -1.366213e-08, -1.356215e-08, 
    -1.368313e-08, -1.397436e-08, -1.418077e-08, -1.429432e-08, 
    -1.476541e-08, -1.470943e-08, -1.481733e-08, -1.497865e-08, 
    -1.509951e-08, -1.54251e-08,
  -1.610915e-08, -1.509568e-08, -1.459189e-08, -1.371656e-08, -1.365603e-08, 
    -1.387731e-08, -1.377352e-08, -1.409798e-08, -1.431961e-08, 
    -1.478915e-08, -1.481709e-08, -1.501539e-08, -1.501432e-08, 
    -1.521491e-08, -1.551652e-08,
  -1.637876e-08, -1.512686e-08, -1.477476e-08, -1.405082e-08, -1.40192e-08, 
    -1.36415e-08, -1.360823e-08, -1.398399e-08, -1.427869e-08, -1.493259e-08, 
    -1.502217e-08, -1.517029e-08, -1.521211e-08, -1.534089e-08, -1.560178e-08,
  -1.338283e-08, -1.317317e-08, -1.315196e-08, -1.345588e-08, -1.395644e-08, 
    -1.428971e-08, -1.435398e-08, -1.455125e-08, -1.449824e-08, 
    -1.427194e-08, -1.391639e-08, -1.363075e-08, -1.375469e-08, 
    -1.401175e-08, -1.445176e-08,
  -1.3562e-08, -1.352271e-08, -1.331483e-08, -1.339335e-08, -1.385965e-08, 
    -1.419989e-08, -1.422656e-08, -1.451504e-08, -1.463303e-08, 
    -1.469275e-08, -1.449727e-08, -1.433887e-08, -1.439058e-08, 
    -1.461475e-08, -1.492483e-08,
  -1.367739e-08, -1.355621e-08, -1.362431e-08, -1.359825e-08, -1.395117e-08, 
    -1.436801e-08, -1.441945e-08, -1.441988e-08, -1.462592e-08, 
    -1.474342e-08, -1.47797e-08, -1.486837e-08, -1.501268e-08, -1.532104e-08, 
    -1.579371e-08,
  -1.414056e-08, -1.347324e-08, -1.378632e-08, -1.381426e-08, -1.391557e-08, 
    -1.440882e-08, -1.46657e-08, -1.46008e-08, -1.478095e-08, -1.472537e-08, 
    -1.499533e-08, -1.515394e-08, -1.555465e-08, -1.607185e-08, -1.674617e-08,
  -1.526315e-08, -1.369582e-08, -1.357023e-08, -1.39571e-08, -1.408489e-08, 
    -1.443424e-08, -1.472433e-08, -1.47653e-08, -1.483457e-08, -1.487759e-08, 
    -1.505243e-08, -1.530782e-08, -1.578198e-08, -1.641836e-08, -1.730184e-08,
  -1.642562e-08, -1.426017e-08, -1.341315e-08, -1.395108e-08, -1.433104e-08, 
    -1.424907e-08, -1.464656e-08, -1.495978e-08, -1.502503e-08, 
    -1.504583e-08, -1.507795e-08, -1.537469e-08, -1.576806e-08, 
    -1.658358e-08, -1.755506e-08,
  -1.707527e-08, -1.49009e-08, -1.342189e-08, -1.365271e-08, -1.434123e-08, 
    -1.43037e-08, -1.466827e-08, -1.505326e-08, -1.51455e-08, -1.515934e-08, 
    -1.520438e-08, -1.533275e-08, -1.576088e-08, -1.66127e-08, -1.782412e-08,
  -1.749948e-08, -1.548304e-08, -1.363902e-08, -1.33931e-08, -1.421494e-08, 
    -1.436558e-08, -1.46636e-08, -1.500514e-08, -1.522756e-08, -1.531266e-08, 
    -1.532842e-08, -1.53003e-08, -1.570985e-08, -1.650366e-08, -1.770725e-08,
  -1.763046e-08, -1.587899e-08, -1.392101e-08, -1.314899e-08, -1.404704e-08, 
    -1.454762e-08, -1.463935e-08, -1.493602e-08, -1.525163e-08, 
    -1.550127e-08, -1.545495e-08, -1.541503e-08, -1.576542e-08, 
    -1.628056e-08, -1.736941e-08,
  -1.762186e-08, -1.606137e-08, -1.421614e-08, -1.307924e-08, -1.398478e-08, 
    -1.45423e-08, -1.465227e-08, -1.486373e-08, -1.525438e-08, -1.564346e-08, 
    -1.568081e-08, -1.563045e-08, -1.575954e-08, -1.614248e-08, -1.69424e-08,
  -1.480718e-08, -1.643543e-08, -1.674541e-08, -1.609906e-08, -1.488239e-08, 
    -1.402216e-08, -1.291065e-08, -1.235381e-08, -1.205758e-08, 
    -1.201442e-08, -1.255818e-08, -1.331749e-08, -1.377972e-08, 
    -1.391869e-08, -1.352178e-08,
  -1.482521e-08, -1.596155e-08, -1.648187e-08, -1.638961e-08, -1.53183e-08, 
    -1.458524e-08, -1.370116e-08, -1.304083e-08, -1.289396e-08, 
    -1.309105e-08, -1.343295e-08, -1.380344e-08, -1.424608e-08, 
    -1.430275e-08, -1.396743e-08,
  -1.463215e-08, -1.546488e-08, -1.647624e-08, -1.699828e-08, -1.635773e-08, 
    -1.531854e-08, -1.473748e-08, -1.410661e-08, -1.393421e-08, 
    -1.399401e-08, -1.394932e-08, -1.445652e-08, -1.489937e-08, 
    -1.476499e-08, -1.458193e-08,
  -1.450114e-08, -1.500949e-08, -1.631455e-08, -1.69543e-08, -1.688147e-08, 
    -1.591255e-08, -1.536682e-08, -1.491249e-08, -1.474955e-08, 
    -1.467245e-08, -1.463204e-08, -1.520735e-08, -1.542976e-08, 
    -1.524791e-08, -1.548785e-08,
  -1.454339e-08, -1.488983e-08, -1.614242e-08, -1.673438e-08, -1.704775e-08, 
    -1.643494e-08, -1.575035e-08, -1.531237e-08, -1.527185e-08, -1.51102e-08, 
    -1.534828e-08, -1.591747e-08, -1.607913e-08, -1.613513e-08, -1.657274e-08,
  -1.483062e-08, -1.492705e-08, -1.601659e-08, -1.672571e-08, -1.713227e-08, 
    -1.6952e-08, -1.621895e-08, -1.586167e-08, -1.585962e-08, -1.569603e-08, 
    -1.612409e-08, -1.664023e-08, -1.677202e-08, -1.719307e-08, -1.794155e-08,
  -1.516317e-08, -1.514024e-08, -1.592017e-08, -1.67806e-08, -1.711753e-08, 
    -1.713958e-08, -1.654306e-08, -1.615382e-08, -1.610014e-08, -1.6012e-08, 
    -1.647129e-08, -1.712347e-08, -1.75364e-08, -1.860895e-08, -2.022467e-08,
  -1.547336e-08, -1.544286e-08, -1.582552e-08, -1.679726e-08, -1.705549e-08, 
    -1.724613e-08, -1.686795e-08, -1.655697e-08, -1.637598e-08, 
    -1.627419e-08, -1.684076e-08, -1.774715e-08, -1.873155e-08, 
    -2.017519e-08, -2.248758e-08,
  -1.595786e-08, -1.573639e-08, -1.570675e-08, -1.668474e-08, -1.695448e-08, 
    -1.723953e-08, -1.725683e-08, -1.706818e-08, -1.683611e-08, 
    -1.683963e-08, -1.742036e-08, -1.862482e-08, -1.998285e-08, 
    -2.165393e-08, -2.426678e-08,
  -1.634526e-08, -1.599252e-08, -1.563416e-08, -1.661198e-08, -1.701571e-08, 
    -1.72865e-08, -1.747916e-08, -1.743763e-08, -1.728601e-08, -1.745559e-08, 
    -1.814119e-08, -1.931515e-08, -2.090948e-08, -2.276564e-08, -2.490301e-08,
  -1.554873e-08, -1.150116e-08, -8.229439e-09, -6.919358e-09, -6.376885e-09, 
    -6.219238e-09, -6.165227e-09, -5.976634e-09, -6.366718e-09, 
    -6.681592e-09, -6.78525e-09, -6.922562e-09, -7.290534e-09, -8.111078e-09, 
    -9.12118e-09,
  -1.62145e-08, -1.215977e-08, -8.297333e-09, -7.38688e-09, -6.599653e-09, 
    -6.365035e-09, -6.181308e-09, -6.081439e-09, -6.504017e-09, 
    -6.831962e-09, -6.9724e-09, -7.194501e-09, -7.84408e-09, -9.048042e-09, 
    -1.026562e-08,
  -1.650027e-08, -1.21191e-08, -8.576211e-09, -7.920272e-09, -7.134547e-09, 
    -6.823541e-09, -6.679334e-09, -6.526328e-09, -6.82329e-09, -7.113822e-09, 
    -7.412661e-09, -7.853939e-09, -8.828894e-09, -1.017743e-08, -1.156939e-08,
  -1.65577e-08, -1.230746e-08, -8.854602e-09, -8.083051e-09, -7.582544e-09, 
    -7.57267e-09, -7.555951e-09, -7.276077e-09, -7.374787e-09, -7.690025e-09, 
    -8.228816e-09, -8.919961e-09, -1.021917e-08, -1.144362e-08, -1.304001e-08,
  -1.632297e-08, -1.240029e-08, -9.245722e-09, -8.382356e-09, -7.993687e-09, 
    -8.427854e-09, -8.271176e-09, -8.051973e-09, -8.029506e-09, 
    -8.546325e-09, -9.301045e-09, -1.02388e-08, -1.122743e-08, -1.247074e-08, 
    -1.450665e-08,
  -1.59852e-08, -1.248226e-08, -9.561425e-09, -8.574966e-09, -8.395915e-09, 
    -9.207821e-09, -8.891879e-09, -8.604708e-09, -8.632422e-09, 
    -9.322755e-09, -1.023141e-08, -1.105079e-08, -1.202727e-08, 
    -1.372148e-08, -1.668922e-08,
  -1.55848e-08, -1.247549e-08, -9.896038e-09, -8.815603e-09, -8.917665e-09, 
    -9.833227e-09, -9.271729e-09, -8.967116e-09, -9.203024e-09, 
    -1.006558e-08, -1.098655e-08, -1.175284e-08, -1.321103e-08, 
    -1.551371e-08, -1.938318e-08,
  -1.474719e-08, -1.266566e-08, -1.023871e-08, -9.218655e-09, -9.438335e-09, 
    -1.027935e-08, -9.403072e-09, -9.236011e-09, -9.828357e-09, 
    -1.070842e-08, -1.160055e-08, -1.267764e-08, -1.455732e-08, 
    -1.734803e-08, -2.228176e-08,
  -1.417791e-08, -1.297168e-08, -1.049962e-08, -9.680694e-09, -9.986619e-09, 
    -1.0354e-08, -9.510424e-09, -9.635365e-09, -1.04507e-08, -1.129585e-08, 
    -1.244739e-08, -1.389426e-08, -1.608743e-08, -1.968648e-08, -2.485562e-08,
  -1.436048e-08, -1.313829e-08, -1.090017e-08, -1.041422e-08, -1.046368e-08, 
    -1.010003e-08, -9.707069e-09, -1.008924e-08, -1.104098e-08, 
    -1.200789e-08, -1.335231e-08, -1.496574e-08, -1.757156e-08, 
    -2.226844e-08, -2.61544e-08,
  -8.717831e-09, -6.515014e-09, -6.59975e-09, -7.096892e-09, -7.866474e-09, 
    -8.663271e-09, -9.403822e-09, -1.043581e-08, -1.15485e-08, -1.305678e-08, 
    -1.483975e-08, -1.654923e-08, -1.792406e-08, -1.880675e-08, -1.945033e-08,
  -9.248497e-09, -6.673209e-09, -6.466064e-09, -7.083538e-09, -7.973603e-09, 
    -8.820138e-09, -9.756877e-09, -1.095754e-08, -1.230322e-08, 
    -1.403506e-08, -1.578512e-08, -1.74944e-08, -1.899195e-08, -2.024717e-08, 
    -2.122736e-08,
  -9.797392e-09, -6.91717e-09, -6.37186e-09, -7.019192e-09, -8.004853e-09, 
    -8.990027e-09, -1.006599e-08, -1.1563e-08, -1.316674e-08, -1.493599e-08, 
    -1.653178e-08, -1.855493e-08, -2.034444e-08, -2.166208e-08, -2.279096e-08,
  -1.051741e-08, -7.171721e-09, -6.286613e-09, -6.829986e-09, -7.966207e-09, 
    -9.185097e-09, -1.049101e-08, -1.218405e-08, -1.387778e-08, 
    -1.563613e-08, -1.76776e-08, -1.994823e-08, -2.157775e-08, -2.30988e-08, 
    -2.453052e-08,
  -1.134025e-08, -7.425625e-09, -6.26972e-09, -6.719898e-09, -7.997787e-09, 
    -9.323658e-09, -1.079126e-08, -1.275132e-08, -1.454984e-08, 
    -1.671386e-08, -1.887166e-08, -2.103948e-08, -2.284786e-08, -2.47351e-08, 
    -2.60492e-08,
  -1.222979e-08, -7.598982e-09, -6.284473e-09, -6.58012e-09, -7.929766e-09, 
    -9.479184e-09, -1.125736e-08, -1.33168e-08, -1.530353e-08, -1.760947e-08, 
    -1.9722e-08, -2.199498e-08, -2.406494e-08, -2.577939e-08, -2.709618e-08,
  -1.256827e-08, -7.863099e-09, -6.328837e-09, -6.455183e-09, -7.827621e-09, 
    -9.584179e-09, -1.145052e-08, -1.368767e-08, -1.599726e-08, 
    -1.840718e-08, -2.060509e-08, -2.299607e-08, -2.50147e-08, -2.670489e-08, 
    -2.787196e-08,
  -1.268169e-08, -8.13055e-09, -6.386847e-09, -6.340602e-09, -7.674067e-09, 
    -9.628742e-09, -1.162298e-08, -1.408267e-08, -1.664534e-08, 
    -1.909351e-08, -2.140391e-08, -2.391705e-08, -2.573121e-08, 
    -2.742283e-08, -2.830046e-08,
  -1.227311e-08, -8.344796e-09, -6.53067e-09, -6.299728e-09, -7.542234e-09, 
    -9.607619e-09, -1.17461e-08, -1.437544e-08, -1.709146e-08, -1.97646e-08, 
    -2.23793e-08, -2.476278e-08, -2.639997e-08, -2.786729e-08, -2.863058e-08,
  -1.166849e-08, -8.440385e-09, -6.675192e-09, -6.299193e-09, -7.414418e-09, 
    -9.546829e-09, -1.186301e-08, -1.461226e-08, -1.749742e-08, 
    -2.045255e-08, -2.312323e-08, -2.533248e-08, -2.683613e-08, 
    -2.799979e-08, -2.883263e-08,
  -1.554934e-08, -1.75866e-08, -1.971879e-08, -2.13285e-08, -2.265864e-08, 
    -2.437482e-08, -2.543249e-08, -2.557348e-08, -2.594244e-08, 
    -2.618452e-08, -2.620334e-08, -2.621553e-08, -2.617744e-08, 
    -2.628682e-08, -2.667525e-08,
  -1.620129e-08, -1.792294e-08, -2.006346e-08, -2.189108e-08, -2.325695e-08, 
    -2.507043e-08, -2.645402e-08, -2.674805e-08, -2.695899e-08, 
    -2.697818e-08, -2.696276e-08, -2.725556e-08, -2.718225e-08, -2.66147e-08, 
    -2.656546e-08,
  -1.65754e-08, -1.787131e-08, -2.019478e-08, -2.238972e-08, -2.38539e-08, 
    -2.577591e-08, -2.738446e-08, -2.76798e-08, -2.772077e-08, -2.758475e-08, 
    -2.751325e-08, -2.761091e-08, -2.717778e-08, -2.625688e-08, -2.582065e-08,
  -1.645325e-08, -1.764819e-08, -2.00843e-08, -2.277625e-08, -2.436332e-08, 
    -2.635712e-08, -2.79327e-08, -2.843156e-08, -2.836782e-08, -2.786432e-08, 
    -2.746757e-08, -2.696757e-08, -2.639548e-08, -2.555112e-08, -2.484938e-08,
  -1.61445e-08, -1.732888e-08, -1.969576e-08, -2.276878e-08, -2.457038e-08, 
    -2.65566e-08, -2.833786e-08, -2.89906e-08, -2.885857e-08, -2.77879e-08, 
    -2.712961e-08, -2.615048e-08, -2.532518e-08, -2.404676e-08, -2.339637e-08,
  -1.558459e-08, -1.691567e-08, -1.921257e-08, -2.258164e-08, -2.477682e-08, 
    -2.660725e-08, -2.844733e-08, -2.909802e-08, -2.877535e-08, 
    -2.742467e-08, -2.652379e-08, -2.518976e-08, -2.42947e-08, -2.298009e-08, 
    -2.182449e-08,
  -1.489431e-08, -1.640676e-08, -1.865698e-08, -2.218584e-08, -2.47399e-08, 
    -2.646193e-08, -2.850004e-08, -2.910111e-08, -2.845013e-08, 
    -2.697213e-08, -2.576265e-08, -2.421699e-08, -2.315772e-08, 
    -2.196948e-08, -2.071003e-08,
  -1.408016e-08, -1.588157e-08, -1.806422e-08, -2.154994e-08, -2.441971e-08, 
    -2.637305e-08, -2.852313e-08, -2.88358e-08, -2.789249e-08, -2.639659e-08, 
    -2.49479e-08, -2.335756e-08, -2.218407e-08, -2.093431e-08, -1.954219e-08,
  -1.339624e-08, -1.525884e-08, -1.737452e-08, -2.084857e-08, -2.395306e-08, 
    -2.621768e-08, -2.846986e-08, -2.860478e-08, -2.745321e-08, 
    -2.595763e-08, -2.438788e-08, -2.274706e-08, -2.157555e-08, 
    -2.046437e-08, -1.902895e-08,
  -1.302566e-08, -1.472193e-08, -1.674023e-08, -1.994237e-08, -2.334272e-08, 
    -2.601839e-08, -2.821886e-08, -2.814035e-08, -2.701491e-08, 
    -2.548272e-08, -2.395574e-08, -2.22842e-08, -2.114519e-08, -2.015468e-08, 
    -1.886854e-08,
  -2.88555e-08, -2.980375e-08, -2.701468e-08, -2.476792e-08, -2.249608e-08, 
    -1.993411e-08, -1.803175e-08, -1.765949e-08, -1.753385e-08, 
    -1.784719e-08, -1.851764e-08, -1.937322e-08, -2.056727e-08, 
    -2.137673e-08, -2.173478e-08,
  -2.903566e-08, -3.032176e-08, -2.773073e-08, -2.561096e-08, -2.311566e-08, 
    -1.994571e-08, -1.792321e-08, -1.680389e-08, -1.626618e-08, 
    -1.642756e-08, -1.728854e-08, -1.805616e-08, -1.943482e-08, 
    -2.094951e-08, -2.212799e-08,
  -2.781554e-08, -2.988112e-08, -2.783174e-08, -2.529264e-08, -2.304152e-08, 
    -1.971041e-08, -1.774641e-08, -1.635794e-08, -1.554534e-08, 
    -1.541022e-08, -1.595026e-08, -1.655309e-08, -1.761659e-08, 
    -1.905656e-08, -2.061683e-08,
  -2.727526e-08, -2.902765e-08, -2.790899e-08, -2.522202e-08, -2.290774e-08, 
    -1.976346e-08, -1.759402e-08, -1.587459e-08, -1.50019e-08, -1.479092e-08, 
    -1.509294e-08, -1.548821e-08, -1.6182e-08, -1.717933e-08, -1.844592e-08,
  -2.636945e-08, -2.656736e-08, -2.630084e-08, -2.450658e-08, -2.284727e-08, 
    -1.991188e-08, -1.782721e-08, -1.586753e-08, -1.478991e-08, 
    -1.450256e-08, -1.453797e-08, -1.458426e-08, -1.481541e-08, 
    -1.531262e-08, -1.588075e-08,
  -2.603467e-08, -2.541715e-08, -2.526876e-08, -2.368813e-08, -2.244219e-08, 
    -2.000002e-08, -1.820004e-08, -1.66041e-08, -1.574261e-08, -1.535754e-08, 
    -1.488555e-08, -1.481095e-08, -1.460067e-08, -1.473745e-08, -1.502464e-08,
  -2.487679e-08, -2.485292e-08, -2.410228e-08, -2.329601e-08, -2.211258e-08, 
    -2.01048e-08, -1.868805e-08, -1.773287e-08, -1.738779e-08, -1.732896e-08, 
    -1.665884e-08, -1.617518e-08, -1.557947e-08, -1.512569e-08, -1.503182e-08,
  -2.409159e-08, -2.418071e-08, -2.319235e-08, -2.315197e-08, -2.196564e-08, 
    -2.027735e-08, -1.90074e-08, -1.855677e-08, -1.87543e-08, -1.890638e-08, 
    -1.859427e-08, -1.806496e-08, -1.781925e-08, -1.731251e-08, -1.702355e-08,
  -2.318454e-08, -2.350036e-08, -2.273541e-08, -2.316215e-08, -2.194916e-08, 
    -2.037215e-08, -1.93791e-08, -1.921127e-08, -1.975534e-08, -2.010156e-08, 
    -1.996503e-08, -1.989197e-08, -1.977793e-08, -1.96854e-08, -1.942117e-08,
  -2.266632e-08, -2.311377e-08, -2.25323e-08, -2.352892e-08, -2.234786e-08, 
    -2.102157e-08, -2.05392e-08, -2.102348e-08, -2.147297e-08, -2.179319e-08, 
    -2.175335e-08, -2.190118e-08, -2.179324e-08, -2.17738e-08, -2.149921e-08,
  -2.063033e-08, -1.987134e-08, -2.083787e-08, -2.243192e-08, -2.347257e-08, 
    -2.450974e-08, -2.446457e-08, -2.426835e-08, -2.360152e-08, 
    -2.296761e-08, -2.208304e-08, -2.128706e-08, -2.029851e-08, -1.95849e-08, 
    -1.907423e-08,
  -2.104782e-08, -2.012768e-08, -2.087594e-08, -2.235291e-08, -2.343976e-08, 
    -2.465398e-08, -2.50462e-08, -2.52973e-08, -2.493364e-08, -2.469575e-08, 
    -2.412173e-08, -2.347396e-08, -2.245275e-08, -2.138139e-08, -2.047965e-08,
  -2.116618e-08, -2.049175e-08, -2.054152e-08, -2.163161e-08, -2.234474e-08, 
    -2.319544e-08, -2.372036e-08, -2.402825e-08, -2.437149e-08, 
    -2.486708e-08, -2.501858e-08, -2.483401e-08, -2.420587e-08, 
    -2.328482e-08, -2.238008e-08,
  -2.105327e-08, -2.020439e-08, -1.996478e-08, -2.058142e-08, -2.109413e-08, 
    -2.184754e-08, -2.259303e-08, -2.312604e-08, -2.323238e-08, 
    -2.387791e-08, -2.431619e-08, -2.466698e-08, -2.465533e-08, 
    -2.427886e-08, -2.371307e-08,
  -2.119848e-08, -1.990811e-08, -1.943575e-08, -1.995505e-08, -2.072403e-08, 
    -2.165475e-08, -2.267099e-08, -2.365144e-08, -2.38439e-08, -2.420587e-08, 
    -2.459733e-08, -2.507324e-08, -2.545455e-08, -2.49637e-08, -2.472465e-08,
  -2.145907e-08, -1.971811e-08, -1.904781e-08, -2.008353e-08, -2.105767e-08, 
    -2.240208e-08, -2.360402e-08, -2.452283e-08, -2.472671e-08, 
    -2.498629e-08, -2.576356e-08, -2.608572e-08, -2.686521e-08, 
    -2.650504e-08, -2.58429e-08,
  -2.144866e-08, -1.977505e-08, -1.91207e-08, -2.066752e-08, -2.216111e-08, 
    -2.367914e-08, -2.463977e-08, -2.4864e-08, -2.516778e-08, -2.538249e-08, 
    -2.622648e-08, -2.664175e-08, -2.775437e-08, -2.792613e-08, -2.743036e-08,
  -2.149197e-08, -2.021761e-08, -1.937405e-08, -2.135853e-08, -2.323076e-08, 
    -2.497395e-08, -2.564152e-08, -2.562561e-08, -2.557614e-08, -2.60019e-08, 
    -2.667454e-08, -2.680493e-08, -2.773012e-08, -2.838851e-08, -2.828224e-08,
  -2.190002e-08, -2.068713e-08, -1.994892e-08, -2.215522e-08, -2.448296e-08, 
    -2.643974e-08, -2.635331e-08, -2.624544e-08, -2.596288e-08, 
    -2.589854e-08, -2.656104e-08, -2.686474e-08, -2.716386e-08, 
    -2.813687e-08, -2.837588e-08,
  -2.243415e-08, -2.133861e-08, -2.06479e-08, -2.263731e-08, -2.580392e-08, 
    -2.725589e-08, -2.656289e-08, -2.63236e-08, -2.59571e-08, -2.56194e-08, 
    -2.599817e-08, -2.649148e-08, -2.65454e-08, -2.735548e-08, -2.806176e-08,
  -2.729741e-08, -2.910227e-08, -2.929399e-08, -2.964386e-08, -2.855759e-08, 
    -2.799009e-08, -2.757132e-08, -2.772951e-08, -2.747223e-08, 
    -2.725433e-08, -2.71005e-08, -2.647718e-08, -2.528012e-08, -2.405381e-08, 
    -2.297246e-08,
  -2.61622e-08, -2.725217e-08, -2.817939e-08, -2.865776e-08, -2.889039e-08, 
    -2.844102e-08, -2.757777e-08, -2.780565e-08, -2.751469e-08, 
    -2.704596e-08, -2.70643e-08, -2.696032e-08, -2.627884e-08, -2.544509e-08, 
    -2.46484e-08,
  -2.607267e-08, -2.692787e-08, -2.775812e-08, -2.843785e-08, -2.921195e-08, 
    -2.948906e-08, -2.826493e-08, -2.774078e-08, -2.759044e-08, 
    -2.699953e-08, -2.623979e-08, -2.604818e-08, -2.582958e-08, 
    -2.533604e-08, -2.519633e-08,
  -2.602933e-08, -2.676715e-08, -2.710581e-08, -2.759885e-08, -2.867952e-08, 
    -2.979786e-08, -2.972575e-08, -2.881576e-08, -2.808378e-08, 
    -2.733472e-08, -2.646276e-08, -2.572585e-08, -2.548195e-08, 
    -2.498202e-08, -2.506664e-08,
  -2.58541e-08, -2.667415e-08, -2.661822e-08, -2.696395e-08, -2.796424e-08, 
    -2.915318e-08, -2.984118e-08, -2.964225e-08, -2.888991e-08, 
    -2.809282e-08, -2.664439e-08, -2.571462e-08, -2.520721e-08, 
    -2.472513e-08, -2.434584e-08,
  -2.592424e-08, -2.67013e-08, -2.655032e-08, -2.671263e-08, -2.739837e-08, 
    -2.866661e-08, -2.974062e-08, -3.017659e-08, -2.960473e-08, 
    -2.857662e-08, -2.748686e-08, -2.582401e-08, -2.521842e-08, 
    -2.459574e-08, -2.391071e-08,
  -2.576076e-08, -2.681615e-08, -2.649727e-08, -2.642328e-08, -2.711689e-08, 
    -2.829212e-08, -2.94709e-08, -3.014301e-08, -3.019537e-08, -2.900521e-08, 
    -2.781668e-08, -2.627839e-08, -2.531666e-08, -2.470394e-08, -2.370752e-08,
  -2.558469e-08, -2.677951e-08, -2.668994e-08, -2.639604e-08, -2.686611e-08, 
    -2.802673e-08, -2.95481e-08, -3.019223e-08, -3.037289e-08, -2.956313e-08, 
    -2.818736e-08, -2.640988e-08, -2.546033e-08, -2.475563e-08, -2.356577e-08,
  -2.519929e-08, -2.664455e-08, -2.695913e-08, -2.655453e-08, -2.673587e-08, 
    -2.7704e-08, -2.931918e-08, -3.009364e-08, -3.042129e-08, -2.9822e-08, 
    -2.854187e-08, -2.669739e-08, -2.538745e-08, -2.482726e-08, -2.351649e-08,
  -2.498448e-08, -2.638515e-08, -2.703057e-08, -2.678558e-08, -2.665964e-08, 
    -2.751163e-08, -2.907821e-08, -3.004147e-08, -3.037465e-08, 
    -3.006895e-08, -2.885088e-08, -2.709767e-08, -2.568674e-08, 
    -2.497306e-08, -2.380367e-08,
  -2.677282e-08, -2.577014e-08, -2.467577e-08, -2.335395e-08, -2.189403e-08, 
    -2.057269e-08, -1.938542e-08, -1.83864e-08, -1.780905e-08, -1.750518e-08, 
    -1.751718e-08, -1.762705e-08, -1.823883e-08, -1.824021e-08, -1.833909e-08,
  -2.75778e-08, -2.687223e-08, -2.613764e-08, -2.476075e-08, -2.350296e-08, 
    -2.212169e-08, -2.066949e-08, -1.891622e-08, -1.763464e-08, 
    -1.691625e-08, -1.655222e-08, -1.647755e-08, -1.658997e-08, 
    -1.719424e-08, -1.792372e-08,
  -2.838079e-08, -2.77968e-08, -2.743219e-08, -2.606794e-08, -2.491427e-08, 
    -2.369381e-08, -2.269726e-08, -2.106437e-08, -1.874508e-08, 
    -1.703629e-08, -1.597701e-08, -1.574537e-08, -1.580507e-08, 
    -1.586975e-08, -1.643775e-08,
  -2.912335e-08, -2.892656e-08, -2.851624e-08, -2.754471e-08, -2.603562e-08, 
    -2.470374e-08, -2.375151e-08, -2.319317e-08, -2.143756e-08, 
    -1.885829e-08, -1.651566e-08, -1.534837e-08, -1.518706e-08, 
    -1.537423e-08, -1.60402e-08,
  -2.891938e-08, -2.920299e-08, -2.924181e-08, -2.875876e-08, -2.773661e-08, 
    -2.606087e-08, -2.462432e-08, -2.379737e-08, -2.303746e-08, 
    -2.127689e-08, -1.855462e-08, -1.622558e-08, -1.486552e-08, 
    -1.457272e-08, -1.476534e-08,
  -2.908411e-08, -2.945218e-08, -2.966567e-08, -2.929256e-08, -2.88891e-08, 
    -2.770376e-08, -2.613062e-08, -2.478961e-08, -2.400492e-08, -2.29895e-08, 
    -2.09949e-08, -1.814198e-08, -1.584704e-08, -1.451722e-08, -1.457734e-08,
  -2.88032e-08, -2.922317e-08, -2.965105e-08, -2.980642e-08, -2.953098e-08, 
    -2.889841e-08, -2.769789e-08, -2.627567e-08, -2.478936e-08, 
    -2.396948e-08, -2.291213e-08, -2.059785e-08, -1.759556e-08, 
    -1.506004e-08, -1.435607e-08,
  -2.879095e-08, -2.911807e-08, -2.949879e-08, -2.946042e-08, -2.968773e-08, 
    -2.938862e-08, -2.885536e-08, -2.811114e-08, -2.66917e-08, -2.477764e-08, 
    -2.398176e-08, -2.288346e-08, -2.042707e-08, -1.704995e-08, -1.471541e-08,
  -2.841205e-08, -2.884402e-08, -2.966343e-08, -2.96514e-08, -2.963821e-08, 
    -2.964043e-08, -2.910958e-08, -2.897296e-08, -2.86309e-08, -2.690171e-08, 
    -2.498822e-08, -2.402631e-08, -2.267146e-08, -1.982235e-08, -1.652806e-08,
  -2.811836e-08, -2.80325e-08, -2.907596e-08, -2.981309e-08, -2.974099e-08, 
    -2.974716e-08, -2.963657e-08, -2.929889e-08, -2.948483e-08, 
    -2.887383e-08, -2.698063e-08, -2.542404e-08, -2.40095e-08, -2.203584e-08, 
    -1.891219e-08,
  -1.535982e-08, -1.500209e-08, -1.482396e-08, -1.484907e-08, -1.506055e-08, 
    -1.533111e-08, -1.58404e-08, -1.655606e-08, -1.728039e-08, -1.784037e-08, 
    -1.860202e-08, -1.932893e-08, -1.971887e-08, -1.9897e-08, -2.003354e-08,
  -1.647653e-08, -1.596495e-08, -1.587383e-08, -1.569235e-08, -1.554958e-08, 
    -1.568341e-08, -1.615268e-08, -1.70077e-08, -1.796181e-08, -1.864017e-08, 
    -1.9477e-08, -2.042373e-08, -2.103622e-08, -2.116947e-08, -2.11502e-08,
  -1.752207e-08, -1.690476e-08, -1.675547e-08, -1.645343e-08, -1.6291e-08, 
    -1.62844e-08, -1.661201e-08, -1.742729e-08, -1.858364e-08, -1.947306e-08, 
    -2.032791e-08, -2.141332e-08, -2.236167e-08, -2.269127e-08, -2.233059e-08,
  -1.868867e-08, -1.799025e-08, -1.763423e-08, -1.725933e-08, -1.694449e-08, 
    -1.692925e-08, -1.705077e-08, -1.753611e-08, -1.846741e-08, 
    -1.964258e-08, -2.089473e-08, -2.229777e-08, -2.34652e-08, -2.417941e-08, 
    -2.393415e-08,
  -1.996164e-08, -1.931533e-08, -1.8777e-08, -1.825394e-08, -1.787237e-08, 
    -1.800269e-08, -1.820066e-08, -1.85278e-08, -1.912427e-08, -2.015052e-08, 
    -2.165059e-08, -2.304474e-08, -2.388093e-08, -2.477027e-08, -2.468271e-08,
  -2.126499e-08, -2.068661e-08, -2.015864e-08, -1.961315e-08, -1.908761e-08, 
    -1.877735e-08, -1.884096e-08, -1.909628e-08, -1.936663e-08, 
    -1.975284e-08, -2.080369e-08, -2.21478e-08, -2.394128e-08, -2.462686e-08, 
    -2.497113e-08,
  -2.328786e-08, -2.260554e-08, -2.191122e-08, -2.116458e-08, -2.035623e-08, 
    -1.968813e-08, -1.905052e-08, -1.884228e-08, -1.900644e-08, -1.91316e-08, 
    -1.947013e-08, -1.96631e-08, -2.073442e-08, -2.184639e-08, -2.369252e-08,
  -2.658875e-08, -2.609046e-08, -2.498511e-08, -2.385468e-08, -2.24468e-08, 
    -2.112964e-08, -1.994813e-08, -1.885844e-08, -1.813168e-08, 
    -1.812108e-08, -1.850413e-08, -1.876025e-08, -1.944712e-08, 
    -1.992694e-08, -2.105318e-08,
  -3.137547e-08, -3.153763e-08, -3.059346e-08, -2.955646e-08, -2.794766e-08, 
    -2.612969e-08, -2.43408e-08, -2.238607e-08, -2.091388e-08, -1.96313e-08, 
    -1.923773e-08, -1.894276e-08, -1.919454e-08, -1.982064e-08, -1.950546e-08,
  -3.408171e-08, -3.418025e-08, -3.456674e-08, -3.397706e-08, -3.270216e-08, 
    -3.02969e-08, -2.851197e-08, -2.64734e-08, -2.459877e-08, -2.290842e-08, 
    -2.161275e-08, -2.072421e-08, -1.959105e-08, -1.971612e-08, -2.024873e-08,
  -1.881339e-08, -1.988043e-08, -1.986745e-08, -2.054335e-08, -2.135421e-08, 
    -2.433251e-08, -2.582749e-08, -2.720174e-08, -2.812751e-08, 
    -2.712133e-08, -2.533414e-08, -2.249585e-08, -1.939575e-08, 
    -1.651618e-08, -1.523877e-08,
  -1.892347e-08, -1.991201e-08, -1.987014e-08, -2.063657e-08, -2.137678e-08, 
    -2.340466e-08, -2.483322e-08, -2.703166e-08, -2.849107e-08, 
    -2.784797e-08, -2.659387e-08, -2.412569e-08, -2.117785e-08, 
    -1.803672e-08, -1.55397e-08,
  -1.910857e-08, -1.983656e-08, -1.970972e-08, -2.048626e-08, -2.117727e-08, 
    -2.305246e-08, -2.44635e-08, -2.711622e-08, -2.775051e-08, -2.741185e-08, 
    -2.604332e-08, -2.431042e-08, -2.190813e-08, -1.949957e-08, -1.671578e-08,
  -1.898059e-08, -1.953277e-08, -1.971903e-08, -2.058957e-08, -2.133415e-08, 
    -2.295488e-08, -2.458721e-08, -2.74487e-08, -2.707008e-08, -2.572854e-08, 
    -2.510187e-08, -2.388285e-08, -2.204293e-08, -1.99584e-08, -1.79352e-08,
  -1.906446e-08, -1.927434e-08, -1.939342e-08, -2.042102e-08, -2.137678e-08, 
    -2.307326e-08, -2.522708e-08, -2.775571e-08, -2.649516e-08, 
    -2.528556e-08, -2.433213e-08, -2.274304e-08, -2.096421e-08, 
    -1.961096e-08, -1.82903e-08,
  -1.899231e-08, -1.895287e-08, -1.964904e-08, -2.090098e-08, -2.189555e-08, 
    -2.384367e-08, -2.659432e-08, -2.592853e-08, -2.486678e-08, 
    -2.367109e-08, -2.272119e-08, -2.127322e-08, -1.979273e-08, -1.90079e-08, 
    -1.789393e-08,
  -1.906453e-08, -1.897445e-08, -1.994914e-08, -2.110453e-08, -2.217074e-08, 
    -2.462553e-08, -2.549218e-08, -2.421532e-08, -2.403043e-08, 
    -2.253049e-08, -2.141378e-08, -2.007489e-08, -1.913736e-08, 
    -1.848682e-08, -1.783125e-08,
  -1.918755e-08, -1.921641e-08, -2.029118e-08, -2.117268e-08, -2.186644e-08, 
    -2.25311e-08, -2.206233e-08, -2.386807e-08, -2.316904e-08, -2.220449e-08, 
    -2.130942e-08, -2.036501e-08, -1.942982e-08, -1.860986e-08, -1.774042e-08,
  -1.945397e-08, -1.962938e-08, -2.051258e-08, -2.143463e-08, -2.262573e-08, 
    -2.513568e-08, -2.698101e-08, -2.540609e-08, -2.39891e-08, -2.20828e-08, 
    -2.10071e-08, -2.003058e-08, -1.925123e-08, -1.838735e-08, -1.753262e-08,
  -2.039539e-08, -2.120629e-08, -2.253718e-08, -2.401365e-08, -2.679213e-08, 
    -2.982242e-08, -2.753844e-08, -2.649835e-08, -2.3966e-08, -2.150511e-08, 
    -2.002967e-08, -1.941454e-08, -1.896856e-08, -1.832147e-08, -1.744129e-08,
  -2.193268e-08, -2.445424e-08, -2.626719e-08, -2.573696e-08, -2.293273e-08, 
    -2.311019e-08, -2.525004e-08, -2.556217e-08, -2.398546e-08, 
    -2.265875e-08, -2.162251e-08, -2.170242e-08, -2.169417e-08, -2.17971e-08, 
    -2.190638e-08,
  -2.110223e-08, -2.3418e-08, -2.518554e-08, -2.466646e-08, -2.205574e-08, 
    -2.234159e-08, -2.484194e-08, -2.617257e-08, -2.453433e-08, 
    -2.306751e-08, -2.186578e-08, -2.184059e-08, -2.160174e-08, -2.14222e-08, 
    -2.148897e-08,
  -2.019558e-08, -2.228236e-08, -2.403482e-08, -2.397684e-08, -2.155531e-08, 
    -2.145846e-08, -2.38997e-08, -2.645585e-08, -2.465907e-08, -2.288988e-08, 
    -2.190115e-08, -2.1827e-08, -2.154495e-08, -2.129651e-08, -2.13106e-08,
  -1.93104e-08, -2.117727e-08, -2.284934e-08, -2.321763e-08, -2.152462e-08, 
    -2.117665e-08, -2.350824e-08, -2.640444e-08, -2.431171e-08, 
    -2.281735e-08, -2.201046e-08, -2.187404e-08, -2.153846e-08, 
    -2.124175e-08, -2.128465e-08,
  -1.831786e-08, -2.017565e-08, -2.173844e-08, -2.242615e-08, -2.150774e-08, 
    -2.119932e-08, -2.380565e-08, -2.628694e-08, -2.338554e-08, 
    -2.273343e-08, -2.199526e-08, -2.198485e-08, -2.165507e-08, 
    -2.132101e-08, -2.133901e-08,
  -1.709653e-08, -1.923846e-08, -2.076016e-08, -2.176063e-08, -2.14755e-08, 
    -2.110972e-08, -2.448296e-08, -2.569931e-08, -2.29224e-08, -2.265933e-08, 
    -2.20903e-08, -2.21959e-08, -2.19457e-08, -2.161009e-08, -2.154011e-08,
  -1.589858e-08, -1.836129e-08, -1.996582e-08, -2.119334e-08, -2.147232e-08, 
    -2.110779e-08, -2.463119e-08, -2.460501e-08, -2.222668e-08, 
    -2.273328e-08, -2.221557e-08, -2.244119e-08, -2.231321e-08, 
    -2.207418e-08, -2.19717e-08,
  -1.496172e-08, -1.751934e-08, -1.931708e-08, -2.077133e-08, -2.14934e-08, 
    -2.175754e-08, -2.430332e-08, -2.392978e-08, -2.142231e-08, 
    -2.283286e-08, -2.253413e-08, -2.28402e-08, -2.284665e-08, -2.267081e-08, 
    -2.267107e-08,
  -1.446073e-08, -1.678898e-08, -1.880417e-08, -2.044582e-08, -2.148098e-08, 
    -2.254571e-08, -2.418013e-08, -2.282207e-08, -2.094827e-08, 
    -2.255062e-08, -2.296104e-08, -2.330553e-08, -2.346442e-08, 
    -2.346928e-08, -2.355774e-08,
  -1.429675e-08, -1.621854e-08, -1.838062e-08, -2.03116e-08, -2.173878e-08, 
    -2.319142e-08, -2.366839e-08, -2.230202e-08, -2.054336e-08, 
    -2.207275e-08, -2.319854e-08, -2.363801e-08, -2.403564e-08, 
    -2.434243e-08, -2.468659e-08,
  -2.639294e-08, -2.635421e-08, -2.469051e-08, -2.401122e-08, -2.292942e-08, 
    -2.171037e-08, -1.986868e-08, -1.784621e-08, -1.613481e-08, 
    -1.484181e-08, -1.39674e-08, -1.317361e-08, -1.246834e-08, -1.201512e-08, 
    -1.187403e-08,
  -2.63284e-08, -2.515757e-08, -2.397822e-08, -2.366157e-08, -2.281466e-08, 
    -2.191745e-08, -2.007123e-08, -1.820934e-08, -1.658675e-08, -1.52193e-08, 
    -1.434576e-08, -1.35569e-08, -1.286747e-08, -1.227018e-08, -1.188604e-08,
  -2.578764e-08, -2.489357e-08, -2.405311e-08, -2.345924e-08, -2.30783e-08, 
    -2.215909e-08, -2.043594e-08, -1.847985e-08, -1.682959e-08, 
    -1.559624e-08, -1.476472e-08, -1.398678e-08, -1.329299e-08, 
    -1.263421e-08, -1.212694e-08,
  -2.552759e-08, -2.48274e-08, -2.451454e-08, -2.363167e-08, -2.305134e-08, 
    -2.249018e-08, -2.090463e-08, -1.912512e-08, -1.747472e-08, 
    -1.616845e-08, -1.512856e-08, -1.427026e-08, -1.371037e-08, -1.30706e-08, 
    -1.23677e-08,
  -2.531352e-08, -2.492525e-08, -2.504441e-08, -2.416185e-08, -2.322909e-08, 
    -2.258241e-08, -2.134343e-08, -1.966053e-08, -1.806399e-08, 
    -1.663702e-08, -1.547881e-08, -1.437081e-08, -1.383713e-08, 
    -1.337616e-08, -1.270291e-08,
  -2.520091e-08, -2.521014e-08, -2.541746e-08, -2.44423e-08, -2.345484e-08, 
    -2.280014e-08, -2.185983e-08, -2.035454e-08, -1.876445e-08, -1.7236e-08, 
    -1.592766e-08, -1.473066e-08, -1.393989e-08, -1.348524e-08, -1.29082e-08,
  -2.540764e-08, -2.582352e-08, -2.586916e-08, -2.468546e-08, -2.366613e-08, 
    -2.280245e-08, -2.214331e-08, -2.081653e-08, -1.944636e-08, 
    -1.782532e-08, -1.643776e-08, -1.515867e-08, -1.421311e-08, 
    -1.350136e-08, -1.298649e-08,
  -2.546524e-08, -2.602698e-08, -2.639524e-08, -2.50872e-08, -2.407174e-08, 
    -2.298581e-08, -2.251116e-08, -2.123835e-08, -2.009092e-08, 
    -1.847464e-08, -1.707311e-08, -1.575737e-08, -1.46641e-08, -1.374661e-08, 
    -1.310567e-08,
  -2.531207e-08, -2.606966e-08, -2.664582e-08, -2.55092e-08, -2.449528e-08, 
    -2.323789e-08, -2.272113e-08, -2.164566e-08, -2.067007e-08, 
    -1.917634e-08, -1.776011e-08, -1.641376e-08, -1.51677e-08, -1.414491e-08, 
    -1.325248e-08,
  -2.488599e-08, -2.578622e-08, -2.665113e-08, -2.586825e-08, -2.498449e-08, 
    -2.374546e-08, -2.301201e-08, -2.210924e-08, -2.115841e-08, 
    -1.995582e-08, -1.85759e-08, -1.718515e-08, -1.574886e-08, -1.460047e-08, 
    -1.354229e-08,
  -1.984719e-08, -2.127145e-08, -2.0013e-08, -1.963327e-08, -1.671718e-08, 
    -1.426354e-08, -1.358045e-08, -1.396575e-08, -1.292737e-08, 
    -1.198286e-08, -1.16291e-08, -1.159491e-08, -1.191437e-08, -1.2553e-08, 
    -1.333935e-08,
  -1.99205e-08, -2.024875e-08, -1.921015e-08, -1.847555e-08, -1.556303e-08, 
    -1.365531e-08, -1.404971e-08, -1.383632e-08, -1.275464e-08, 
    -1.210618e-08, -1.186543e-08, -1.190434e-08, -1.240833e-08, 
    -1.316898e-08, -1.421328e-08,
  -1.917887e-08, -1.927498e-08, -1.844875e-08, -1.728076e-08, -1.473884e-08, 
    -1.368759e-08, -1.432798e-08, -1.342707e-08, -1.274126e-08, 
    -1.219902e-08, -1.200682e-08, -1.213135e-08, -1.277798e-08, 
    -1.369933e-08, -1.503279e-08,
  -1.862753e-08, -1.860733e-08, -1.775403e-08, -1.641146e-08, -1.410189e-08, 
    -1.39388e-08, -1.431377e-08, -1.305582e-08, -1.238705e-08, -1.195144e-08, 
    -1.199448e-08, -1.234845e-08, -1.321141e-08, -1.441928e-08, -1.585087e-08,
  -1.833848e-08, -1.81058e-08, -1.702646e-08, -1.537658e-08, -1.371964e-08, 
    -1.42026e-08, -1.395074e-08, -1.276258e-08, -1.217739e-08, -1.191788e-08, 
    -1.202505e-08, -1.25866e-08, -1.372559e-08, -1.51925e-08, -1.645769e-08,
  -1.803891e-08, -1.740616e-08, -1.586331e-08, -1.437113e-08, -1.370622e-08, 
    -1.415649e-08, -1.35019e-08, -1.250117e-08, -1.20108e-08, -1.193102e-08, 
    -1.205435e-08, -1.291404e-08, -1.441534e-08, -1.580401e-08, -1.702413e-08,
  -1.747021e-08, -1.641479e-08, -1.492834e-08, -1.383324e-08, -1.395539e-08, 
    -1.404018e-08, -1.307473e-08, -1.221659e-08, -1.194918e-08, 
    -1.196535e-08, -1.22377e-08, -1.341049e-08, -1.503698e-08, -1.641614e-08, 
    -1.779861e-08,
  -1.679783e-08, -1.559053e-08, -1.452995e-08, -1.390459e-08, -1.406928e-08, 
    -1.388264e-08, -1.258929e-08, -1.192582e-08, -1.201621e-08, 
    -1.207008e-08, -1.253322e-08, -1.401724e-08, -1.563551e-08, 
    -1.729572e-08, -1.895077e-08,
  -1.645812e-08, -1.538003e-08, -1.445009e-08, -1.429513e-08, -1.399004e-08, 
    -1.335593e-08, -1.211641e-08, -1.189271e-08, -1.217058e-08, 
    -1.221175e-08, -1.289627e-08, -1.467365e-08, -1.648492e-08, 
    -1.843182e-08, -2.00361e-08,
  -1.662139e-08, -1.560789e-08, -1.467788e-08, -1.425067e-08, -1.359824e-08, 
    -1.267915e-08, -1.178478e-08, -1.197043e-08, -1.218372e-08, 
    -1.243385e-08, -1.337684e-08, -1.53176e-08, -1.715627e-08, -1.897849e-08, 
    -2.047557e-08,
  -1.458835e-08, -1.495528e-08, -1.606243e-08, -1.838595e-08, -2.037392e-08, 
    -1.973994e-08, -1.756383e-08, -1.697452e-08, -1.788808e-08, 
    -1.864668e-08, -1.886745e-08, -1.911121e-08, -1.942671e-08, 
    -1.920823e-08, -1.853454e-08,
  -1.497843e-08, -1.522646e-08, -1.646034e-08, -1.91359e-08, -2.056262e-08, 
    -1.949961e-08, -1.681815e-08, -1.713752e-08, -1.846854e-08, 
    -1.947319e-08, -1.995398e-08, -2.042876e-08, -2.05218e-08, -2.020282e-08, 
    -1.913337e-08,
  -1.529765e-08, -1.547867e-08, -1.694359e-08, -1.990691e-08, -2.073488e-08, 
    -1.873776e-08, -1.660174e-08, -1.783148e-08, -1.924359e-08, 
    -2.048871e-08, -2.118744e-08, -2.186064e-08, -2.174384e-08, -2.1047e-08, 
    -1.989805e-08,
  -1.545367e-08, -1.578153e-08, -1.761883e-08, -2.082414e-08, -2.069205e-08, 
    -1.774364e-08, -1.662967e-08, -1.853249e-08, -2.010524e-08, 
    -2.134586e-08, -2.220656e-08, -2.277674e-08, -2.247577e-08, -2.1671e-08, 
    -2.065807e-08,
  -1.56953e-08, -1.616801e-08, -1.853082e-08, -2.167018e-08, -2.033372e-08, 
    -1.690263e-08, -1.717543e-08, -1.962553e-08, -2.112006e-08, -2.23268e-08, 
    -2.294817e-08, -2.325073e-08, -2.284105e-08, -2.227098e-08, -2.168592e-08,
  -1.601301e-08, -1.679908e-08, -1.984377e-08, -2.221178e-08, -1.944816e-08, 
    -1.665739e-08, -1.827177e-08, -2.070303e-08, -2.195019e-08, 
    -2.276322e-08, -2.354383e-08, -2.368281e-08, -2.35595e-08, -2.318983e-08, 
    -2.295936e-08,
  -1.651915e-08, -1.771784e-08, -2.113766e-08, -2.218749e-08, -1.83889e-08, 
    -1.696889e-08, -1.940997e-08, -2.169237e-08, -2.270323e-08, 
    -2.350707e-08, -2.449665e-08, -2.471299e-08, -2.469278e-08, 
    -2.450197e-08, -2.433521e-08,
  -1.730526e-08, -1.902783e-08, -2.235654e-08, -2.168788e-08, -1.760501e-08, 
    -1.75361e-08, -2.059428e-08, -2.260398e-08, -2.362202e-08, -2.484395e-08, 
    -2.570303e-08, -2.57837e-08, -2.565189e-08, -2.561232e-08, -2.546924e-08,
  -1.83974e-08, -2.035588e-08, -2.29454e-08, -2.066319e-08, -1.743428e-08, 
    -1.854108e-08, -2.15698e-08, -2.350558e-08, -2.500533e-08, -2.614773e-08, 
    -2.673447e-08, -2.684865e-08, -2.694304e-08, -2.706334e-08, -2.692038e-08,
  -1.947437e-08, -2.159087e-08, -2.287345e-08, -1.967502e-08, -1.778031e-08, 
    -1.938096e-08, -2.256549e-08, -2.482451e-08, -2.6508e-08, -2.752313e-08, 
    -2.796141e-08, -2.781256e-08, -2.771128e-08, -2.763919e-08, -2.757566e-08,
  -1.7805e-08, -1.760964e-08, -1.769284e-08, -1.878051e-08, -1.94428e-08, 
    -1.9999e-08, -2.123435e-08, -2.202911e-08, -2.232914e-08, -2.231635e-08, 
    -2.161791e-08, -2.023502e-08, -1.830414e-08, -1.664782e-08, -1.516666e-08,
  -1.809164e-08, -1.792601e-08, -1.811499e-08, -1.945089e-08, -2.012369e-08, 
    -2.107671e-08, -2.284762e-08, -2.371629e-08, -2.4309e-08, -2.407675e-08, 
    -2.386191e-08, -2.259029e-08, -2.089743e-08, -1.902224e-08, -1.697976e-08,
  -1.830994e-08, -1.80759e-08, -1.839963e-08, -1.98214e-08, -2.071817e-08, 
    -2.212959e-08, -2.384771e-08, -2.474983e-08, -2.549677e-08, 
    -2.555417e-08, -2.517078e-08, -2.431715e-08, -2.31061e-08, -2.135218e-08, 
    -1.954818e-08,
  -1.84762e-08, -1.82169e-08, -1.866027e-08, -2.018336e-08, -2.137711e-08, 
    -2.310562e-08, -2.483068e-08, -2.563153e-08, -2.659367e-08, 
    -2.692043e-08, -2.680315e-08, -2.579297e-08, -2.487088e-08, -2.34657e-08, 
    -2.175424e-08,
  -1.864139e-08, -1.837585e-08, -1.886385e-08, -2.041368e-08, -2.193035e-08, 
    -2.399565e-08, -2.562372e-08, -2.638366e-08, -2.720458e-08, 
    -2.804387e-08, -2.833086e-08, -2.779688e-08, -2.666382e-08, 
    -2.557237e-08, -2.386856e-08,
  -1.885495e-08, -1.853967e-08, -1.898257e-08, -2.057851e-08, -2.244266e-08, 
    -2.487594e-08, -2.628444e-08, -2.676123e-08, -2.742685e-08, 
    -2.858499e-08, -2.918715e-08, -2.914341e-08, -2.834021e-08, 
    -2.741037e-08, -2.580961e-08,
  -1.908251e-08, -1.872021e-08, -1.902377e-08, -2.067294e-08, -2.288701e-08, 
    -2.565338e-08, -2.675138e-08, -2.695041e-08, -2.781618e-08, 
    -2.894074e-08, -2.966553e-08, -2.967291e-08, -2.937215e-08, 
    -2.873625e-08, -2.783445e-08,
  -1.931034e-08, -1.887052e-08, -1.901351e-08, -2.068029e-08, -2.32759e-08, 
    -2.638398e-08, -2.725426e-08, -2.730563e-08, -2.819951e-08, 
    -2.894093e-08, -2.971156e-08, -2.988482e-08, -2.982571e-08, 
    -2.958662e-08, -2.917535e-08,
  -1.952956e-08, -1.902142e-08, -1.898766e-08, -2.060118e-08, -2.359183e-08, 
    -2.699721e-08, -2.770274e-08, -2.786021e-08, -2.845164e-08, 
    -2.890402e-08, -2.930721e-08, -2.971389e-08, -2.970367e-08, 
    -2.974564e-08, -2.965843e-08,
  -1.976633e-08, -1.91186e-08, -1.892015e-08, -2.049207e-08, -2.380064e-08, 
    -2.75518e-08, -2.819873e-08, -2.824987e-08, -2.853736e-08, -2.850008e-08, 
    -2.879123e-08, -2.922549e-08, -2.946315e-08, -2.95454e-08, -2.962142e-08,
  -2.504292e-08, -2.701645e-08, -2.709341e-08, -2.648145e-08, -2.54115e-08, 
    -2.360345e-08, -2.122049e-08, -1.878713e-08, -1.66621e-08, -1.470736e-08, 
    -1.299885e-08, -1.189764e-08, -1.117372e-08, -1.051569e-08, -1.016894e-08,
  -2.567417e-08, -2.782155e-08, -2.877457e-08, -2.872828e-08, -2.776069e-08, 
    -2.606482e-08, -2.384699e-08, -2.113575e-08, -1.861122e-08, 
    -1.650034e-08, -1.438196e-08, -1.274283e-08, -1.175139e-08, 
    -1.086247e-08, -1.030626e-08,
  -2.582409e-08, -2.797434e-08, -2.924081e-08, -2.973989e-08, -2.912502e-08, 
    -2.749841e-08, -2.543071e-08, -2.304303e-08, -2.016334e-08, 
    -1.770559e-08, -1.54655e-08, -1.37274e-08, -1.239422e-08, -1.123031e-08, 
    -1.049592e-08,
  -2.613578e-08, -2.832796e-08, -2.974404e-08, -3.03058e-08, -3.026363e-08, 
    -2.964298e-08, -2.776852e-08, -2.525837e-08, -2.273127e-08, 
    -1.958446e-08, -1.684507e-08, -1.489521e-08, -1.320068e-08, 
    -1.171832e-08, -1.06034e-08,
  -2.62218e-08, -2.847618e-08, -2.98562e-08, -3.028956e-08, -2.996702e-08, 
    -2.980449e-08, -2.931053e-08, -2.688781e-08, -2.439347e-08, 
    -2.153713e-08, -1.857996e-08, -1.625119e-08, -1.428988e-08, 
    -1.241368e-08, -1.10382e-08,
  -2.611287e-08, -2.87298e-08, -3.018142e-08, -3.10339e-08, -3.042015e-08, 
    -3.00276e-08, -3.030232e-08, -2.911004e-08, -2.658138e-08, -2.326682e-08, 
    -2.053125e-08, -1.791523e-08, -1.573167e-08, -1.338038e-08, -1.160895e-08,
  -2.589164e-08, -2.887788e-08, -3.06675e-08, -3.136823e-08, -3.102122e-08, 
    -3.032641e-08, -3.059234e-08, -3.022756e-08, -2.865671e-08, -2.54104e-08, 
    -2.211777e-08, -1.967997e-08, -1.732842e-08, -1.497905e-08, -1.254917e-08,
  -2.562752e-08, -2.891685e-08, -3.111372e-08, -3.190711e-08, -3.156486e-08, 
    -3.073746e-08, -3.074719e-08, -3.070446e-08, -2.941058e-08, 
    -2.773555e-08, -2.40305e-08, -2.136985e-08, -1.901404e-08, -1.658171e-08, 
    -1.413184e-08,
  -2.520199e-08, -2.875859e-08, -3.144681e-08, -3.242832e-08, -3.193311e-08, 
    -3.098147e-08, -3.099078e-08, -3.098737e-08, -3.006553e-08, 
    -2.868548e-08, -2.623283e-08, -2.307355e-08, -2.078824e-08, 
    -1.833337e-08, -1.575436e-08,
  -2.467109e-08, -2.846159e-08, -3.155467e-08, -3.2849e-08, -3.220234e-08, 
    -3.127234e-08, -3.103069e-08, -3.092175e-08, -3.032369e-08, 
    -2.943553e-08, -2.750162e-08, -2.499152e-08, -2.235489e-08, 
    -2.009708e-08, -1.76017e-08,
  -1.17299e-08, -1.072487e-08, -1.017712e-08, -9.308734e-09, -8.563977e-09, 
    -7.908763e-09, -7.4997e-09, -7.231357e-09, -6.984572e-09, -6.813709e-09, 
    -6.736022e-09, -6.685136e-09, -6.626364e-09, -6.480435e-09, -6.383353e-09,
  -1.278105e-08, -1.189079e-08, -1.104297e-08, -1.0015e-08, -9.062176e-09, 
    -8.205028e-09, -7.712623e-09, -7.352032e-09, -7.069264e-09, 
    -6.821187e-09, -6.616486e-09, -6.514352e-09, -6.375862e-09, 
    -6.297269e-09, -6.239481e-09,
  -1.350839e-08, -1.254555e-08, -1.154259e-08, -1.056084e-08, -9.566228e-09, 
    -8.66204e-09, -8.013561e-09, -7.664159e-09, -7.404932e-09, -7.150757e-09, 
    -6.872108e-09, -6.704693e-09, -6.522135e-09, -6.405846e-09, -6.282403e-09,
  -1.429358e-08, -1.32264e-08, -1.218865e-08, -1.117434e-08, -1.025943e-08, 
    -9.309096e-09, -8.619456e-09, -8.202639e-09, -7.942014e-09, 
    -7.653875e-09, -7.250652e-09, -6.92259e-09, -6.64316e-09, -6.507304e-09, 
    -6.420944e-09,
  -1.507184e-08, -1.401281e-08, -1.295917e-08, -1.187623e-08, -1.102336e-08, 
    -1.014171e-08, -9.429298e-09, -9.035521e-09, -8.722376e-09, 
    -8.486817e-09, -8.110925e-09, -7.657931e-09, -7.240098e-09, 
    -6.831395e-09, -6.641021e-09,
  -1.563396e-08, -1.46625e-08, -1.378644e-08, -1.276912e-08, -1.192688e-08, 
    -1.109026e-08, -1.027281e-08, -9.709575e-09, -9.422382e-09, 
    -9.191225e-09, -8.910337e-09, -8.472774e-09, -8.068856e-09, 
    -7.574345e-09, -7.112872e-09,
  -1.639802e-08, -1.54146e-08, -1.458213e-08, -1.383403e-08, -1.30054e-08, 
    -1.229983e-08, -1.150816e-08, -1.083333e-08, -1.03808e-08, -1.01076e-08, 
    -9.857634e-09, -9.387837e-09, -8.954237e-09, -8.515015e-09, -8.023867e-09,
  -1.723497e-08, -1.632078e-08, -1.545016e-08, -1.483466e-08, -1.415199e-08, 
    -1.351666e-08, -1.277069e-08, -1.221607e-08, -1.172075e-08, 
    -1.136273e-08, -1.107121e-08, -1.066951e-08, -1.0069e-08, -9.527965e-09, 
    -9.015963e-09,
  -1.795155e-08, -1.717468e-08, -1.638574e-08, -1.592039e-08, -1.535751e-08, 
    -1.481271e-08, -1.403442e-08, -1.346885e-08, -1.308881e-08, 
    -1.279517e-08, -1.26148e-08, -1.231766e-08, -1.181196e-08, -1.111572e-08, 
    -1.033822e-08,
  -1.878336e-08, -1.791656e-08, -1.724371e-08, -1.689943e-08, -1.65268e-08, 
    -1.617629e-08, -1.555619e-08, -1.497554e-08, -1.453859e-08, 
    -1.422944e-08, -1.408725e-08, -1.395738e-08, -1.365556e-08, 
    -1.313596e-08, -1.235506e-08,
  -8.731539e-09, -7.913601e-09, -7.319813e-09, -6.757075e-09, -6.276457e-09, 
    -5.667408e-09, -5.041246e-09, -4.412559e-09, -3.846238e-09, 
    -3.355524e-09, -2.97e-09, -2.700299e-09, -2.519288e-09, -2.422326e-09, 
    -2.434478e-09,
  -9.508511e-09, -8.56088e-09, -7.923575e-09, -7.346798e-09, -6.886582e-09, 
    -6.335907e-09, -5.766056e-09, -5.155392e-09, -4.541237e-09, 
    -3.951188e-09, -3.472542e-09, -3.086265e-09, -2.793082e-09, 
    -2.597616e-09, -2.485104e-09,
  -1.038536e-08, -9.333041e-09, -8.69343e-09, -8.012263e-09, -7.470752e-09, 
    -6.886751e-09, -6.308609e-09, -5.772183e-09, -5.240705e-09, 
    -4.657902e-09, -4.14282e-09, -3.754257e-09, -3.449914e-09, -3.232693e-09, 
    -3.06546e-09,
  -1.18938e-08, -1.055094e-08, -9.74326e-09, -9.023228e-09, -8.416923e-09, 
    -7.843985e-09, -7.194029e-09, -6.50973e-09, -5.929175e-09, -5.37388e-09, 
    -4.74975e-09, -4.23104e-09, -3.877819e-09, -3.648461e-09, -3.467175e-09,
  -1.368301e-08, -1.232441e-08, -1.119145e-08, -1.029768e-08, -9.507574e-09, 
    -8.829478e-09, -8.182885e-09, -7.558572e-09, -6.950956e-09, 
    -6.422334e-09, -5.894531e-09, -5.315639e-09, -4.825949e-09, 
    -4.546081e-09, -4.269426e-09,
  -1.574444e-08, -1.458604e-08, -1.335445e-08, -1.208721e-08, -1.105748e-08, 
    -1.00734e-08, -9.330241e-09, -8.625412e-09, -7.971908e-09, -7.294924e-09, 
    -6.726467e-09, -6.150501e-09, -5.5716e-09, -5.109349e-09, -4.871572e-09,
  -1.775071e-08, -1.671656e-08, -1.568408e-08, -1.424773e-08, -1.285575e-08, 
    -1.156255e-08, -1.050549e-08, -9.647896e-09, -8.855024e-09, 
    -8.088878e-09, -7.399316e-09, -6.763095e-09, -6.136723e-09, 
    -5.599411e-09, -5.137387e-09,
  -1.993912e-08, -1.911752e-08, -1.823838e-08, -1.687399e-08, -1.52946e-08, 
    -1.356123e-08, -1.216814e-08, -1.09341e-08, -9.904879e-09, -9.020441e-09, 
    -8.226836e-09, -7.57083e-09, -7.00134e-09, -6.479096e-09, -5.971664e-09,
  -2.206571e-08, -2.147252e-08, -2.075022e-08, -1.960071e-08, -1.826923e-08, 
    -1.64601e-08, -1.471044e-08, -1.308324e-08, -1.174069e-08, -1.059441e-08, 
    -9.727357e-09, -8.97049e-09, -8.213628e-09, -7.51188e-09, -7.00647e-09,
  -2.442266e-08, -2.401841e-08, -2.338153e-08, -2.233662e-08, -2.124019e-08, 
    -1.996552e-08, -1.829678e-08, -1.649453e-08, -1.478922e-08, 
    -1.337597e-08, -1.214747e-08, -1.122816e-08, -1.06137e-08, -1.001807e-08, 
    -9.383801e-09,
  -4.891043e-09, -4.850969e-09, -5.084062e-09, -5.402361e-09, -5.781848e-09, 
    -6.057919e-09, -6.262386e-09, -6.370643e-09, -6.412649e-09, 
    -6.433392e-09, -6.466518e-09, -6.575767e-09, -6.746005e-09, 
    -6.901239e-09, -7.041694e-09,
  -5.152723e-09, -5.43067e-09, -5.864594e-09, -6.234099e-09, -6.648497e-09, 
    -7.008221e-09, -7.342439e-09, -7.572943e-09, -7.734487e-09, 
    -7.843473e-09, -7.96698e-09, -8.136928e-09, -8.387057e-09, -8.622201e-09, 
    -8.837877e-09,
  -5.476425e-09, -5.952155e-09, -6.514772e-09, -7.016614e-09, -7.517998e-09, 
    -8.082602e-09, -8.596336e-09, -9.0586e-09, -9.420631e-09, -9.761659e-09, 
    -1.008231e-08, -1.044503e-08, -1.080167e-08, -1.118237e-08, -1.149333e-08,
  -5.779313e-09, -6.364604e-09, -7.141578e-09, -7.833915e-09, -8.509107e-09, 
    -9.238589e-09, -9.885462e-09, -1.049042e-08, -1.102015e-08, 
    -1.149569e-08, -1.18828e-08, -1.221092e-08, -1.250284e-08, -1.274639e-08, 
    -1.296034e-08,
  -6.365323e-09, -6.773436e-09, -7.546408e-09, -8.448337e-09, -9.331187e-09, 
    -1.02389e-08, -1.108453e-08, -1.190938e-08, -1.263091e-08, -1.331406e-08, 
    -1.394959e-08, -1.450611e-08, -1.502172e-08, -1.5484e-08, -1.590338e-08,
  -7.286709e-09, -7.598076e-09, -8.638787e-09, -9.584078e-09, -1.048861e-08, 
    -1.143635e-08, -1.228707e-08, -1.309746e-08, -1.382129e-08, 
    -1.452038e-08, -1.518668e-08, -1.582834e-08, -1.649079e-08, 
    -1.713136e-08, -1.7823e-08,
  -9.157067e-09, -9.578335e-09, -1.068869e-08, -1.135807e-08, -1.22001e-08, 
    -1.288493e-08, -1.352094e-08, -1.402103e-08, -1.453013e-08, 
    -1.498034e-08, -1.5455e-08, -1.586995e-08, -1.639822e-08, -1.691849e-08, 
    -1.746628e-08,
  -1.146459e-08, -1.20742e-08, -1.291088e-08, -1.334368e-08, -1.389824e-08, 
    -1.433565e-08, -1.474071e-08, -1.524278e-08, -1.583585e-08, 
    -1.635482e-08, -1.680857e-08, -1.721567e-08, -1.762059e-08, -1.79998e-08, 
    -1.8317e-08,
  -1.37995e-08, -1.430054e-08, -1.496836e-08, -1.526332e-08, -1.575039e-08, 
    -1.614072e-08, -1.661745e-08, -1.718508e-08, -1.776498e-08, 
    -1.821237e-08, -1.850999e-08, -1.878228e-08, -1.903634e-08, 
    -1.933405e-08, -1.958042e-08,
  -1.629547e-08, -1.673163e-08, -1.711477e-08, -1.734512e-08, -1.775097e-08, 
    -1.830337e-08, -1.883975e-08, -1.947704e-08, -1.992162e-08, 
    -2.022498e-08, -2.035391e-08, -2.041925e-08, -2.046765e-08, -2.04928e-08, 
    -2.053712e-08,
  -9.989904e-09, -1.005422e-08, -1.017247e-08, -1.015824e-08, -1.009857e-08, 
    -1.006597e-08, -9.936497e-09, -9.740054e-09, -9.447071e-09, 
    -9.051718e-09, -8.627677e-09, -8.226079e-09, -7.840709e-09, -7.48718e-09, 
    -7.157804e-09,
  -1.09833e-08, -1.118002e-08, -1.132487e-08, -1.144797e-08, -1.148781e-08, 
    -1.156533e-08, -1.152263e-08, -1.141098e-08, -1.117959e-08, 
    -1.072823e-08, -1.018167e-08, -9.537324e-09, -8.963355e-09, 
    -8.434483e-09, -7.995447e-09,
  -1.227187e-08, -1.2418e-08, -1.264557e-08, -1.285885e-08, -1.316162e-08, 
    -1.342562e-08, -1.362915e-08, -1.363336e-08, -1.355258e-08, 
    -1.329309e-08, -1.287705e-08, -1.230069e-08, -1.145031e-08, -1.05533e-08, 
    -9.639092e-09,
  -1.340504e-08, -1.359213e-08, -1.416184e-08, -1.446403e-08, -1.483239e-08, 
    -1.498709e-08, -1.514702e-08, -1.512122e-08, -1.502842e-08, 
    -1.480892e-08, -1.450441e-08, -1.408367e-08, -1.359395e-08, 
    -1.300456e-08, -1.229423e-08,
  -1.479219e-08, -1.553438e-08, -1.61347e-08, -1.6238e-08, -1.639104e-08, 
    -1.645779e-08, -1.659803e-08, -1.645743e-08, -1.631644e-08, 
    -1.598794e-08, -1.561983e-08, -1.515326e-08, -1.475564e-08, 
    -1.438795e-08, -1.401527e-08,
  -1.714207e-08, -1.739992e-08, -1.747335e-08, -1.739641e-08, -1.753589e-08, 
    -1.741555e-08, -1.741474e-08, -1.715421e-08, -1.695051e-08, -1.64755e-08, 
    -1.59748e-08, -1.533522e-08, -1.479571e-08, -1.431729e-08, -1.404429e-08,
  -1.758138e-08, -1.783046e-08, -1.762211e-08, -1.721373e-08, -1.702012e-08, 
    -1.66682e-08, -1.64474e-08, -1.602507e-08, -1.567297e-08, -1.520203e-08, 
    -1.474441e-08, -1.42753e-08, -1.386976e-08, -1.350777e-08, -1.322486e-08,
  -1.801525e-08, -1.785749e-08, -1.715312e-08, -1.691519e-08, -1.662206e-08, 
    -1.643669e-08, -1.625051e-08, -1.586964e-08, -1.55896e-08, -1.517366e-08, 
    -1.476223e-08, -1.436012e-08, -1.398891e-08, -1.362858e-08, -1.3336e-08,
  -1.784162e-08, -1.735233e-08, -1.700983e-08, -1.709122e-08, -1.71278e-08, 
    -1.694879e-08, -1.642976e-08, -1.60698e-08, -1.560754e-08, -1.532521e-08, 
    -1.504536e-08, -1.48022e-08, -1.454164e-08, -1.424173e-08, -1.390204e-08,
  -1.722523e-08, -1.736609e-08, -1.758563e-08, -1.774247e-08, -1.74525e-08, 
    -1.68219e-08, -1.623267e-08, -1.571616e-08, -1.534737e-08, -1.513098e-08, 
    -1.495001e-08, -1.483067e-08, -1.472383e-08, -1.456254e-08, -1.433424e-08,
  -1.093009e-08, -1.072217e-08, -1.085114e-08, -1.060122e-08, -1.046068e-08, 
    -1.007176e-08, -9.6462e-09, -9.10835e-09, -8.716084e-09, -8.389654e-09, 
    -8.050755e-09, -7.733695e-09, -7.363781e-09, -7.095909e-09, -6.86404e-09,
  -1.174026e-08, -1.16923e-08, -1.187915e-08, -1.172104e-08, -1.158498e-08, 
    -1.128564e-08, -1.087233e-08, -1.032898e-08, -9.696773e-09, 
    -9.217762e-09, -8.776605e-09, -8.405739e-09, -8.120272e-09, 
    -7.897753e-09, -7.742598e-09,
  -1.219475e-08, -1.235278e-08, -1.254609e-08, -1.250266e-08, -1.253558e-08, 
    -1.225184e-08, -1.198882e-08, -1.151159e-08, -1.09679e-08, -1.032046e-08, 
    -9.798068e-09, -9.201099e-09, -8.749925e-09, -8.374444e-09, -8.210109e-09,
  -1.193489e-08, -1.22954e-08, -1.241378e-08, -1.221074e-08, -1.199561e-08, 
    -1.150163e-08, -1.123623e-08, -1.125057e-08, -1.117323e-08, 
    -1.099478e-08, -1.064066e-08, -1.019606e-08, -9.824621e-09, 
    -9.350513e-09, -8.860163e-09,
  -1.249635e-08, -1.296628e-08, -1.300505e-08, -1.286748e-08, -1.263056e-08, 
    -1.196844e-08, -1.114039e-08, -1.05018e-08, -1.007023e-08, -9.832394e-09, 
    -9.971547e-09, -1.005181e-08, -1.013211e-08, -9.989099e-09, -9.694992e-09,
  -1.328322e-08, -1.347233e-08, -1.361739e-08, -1.355476e-08, -1.349073e-08, 
    -1.287568e-08, -1.192423e-08, -1.101541e-08, -1.031352e-08, 
    -9.777391e-09, -9.487497e-09, -9.280559e-09, -9.234711e-09, 
    -9.367532e-09, -9.565227e-09,
  -1.359993e-08, -1.370714e-08, -1.400657e-08, -1.407552e-08, -1.403403e-08, 
    -1.367123e-08, -1.296355e-08, -1.220226e-08, -1.141973e-08, 
    -1.074608e-08, -1.025981e-08, -9.866671e-09, -9.560557e-09, 
    -9.217438e-09, -9.097053e-09,
  -1.371246e-08, -1.405733e-08, -1.415768e-08, -1.406835e-08, -1.39586e-08, 
    -1.356154e-08, -1.28636e-08, -1.240731e-08, -1.209223e-08, -1.188244e-08, 
    -1.168566e-08, -1.133613e-08, -1.085288e-08, -1.029574e-08, -9.751479e-09,
  -1.388561e-08, -1.424609e-08, -1.427164e-08, -1.414487e-08, -1.401843e-08, 
    -1.389901e-08, -1.348135e-08, -1.304768e-08, -1.266518e-08, 
    -1.234984e-08, -1.221806e-08, -1.223283e-08, -1.214593e-08, 
    -1.178151e-08, -1.124632e-08,
  -1.410418e-08, -1.438897e-08, -1.410746e-08, -1.393006e-08, -1.418773e-08, 
    -1.43301e-08, -1.416889e-08, -1.415348e-08, -1.393544e-08, -1.364333e-08, 
    -1.324184e-08, -1.284259e-08, -1.255259e-08, -1.241504e-08, -1.22649e-08,
  -1.126327e-08, -1.154466e-08, -1.159935e-08, -1.149937e-08, -1.137927e-08, 
    -1.131235e-08, -1.127274e-08, -1.139343e-08, -1.170654e-08, 
    -1.211203e-08, -1.251199e-08, -1.292838e-08, -1.327951e-08, 
    -1.354555e-08, -1.382716e-08,
  -1.08354e-08, -1.116787e-08, -1.144004e-08, -1.141357e-08, -1.131544e-08, 
    -1.11887e-08, -1.110193e-08, -1.108793e-08, -1.121729e-08, -1.14559e-08, 
    -1.181121e-08, -1.226534e-08, -1.277363e-08, -1.328085e-08, -1.380936e-08,
  -1.074262e-08, -1.109346e-08, -1.142495e-08, -1.165695e-08, -1.173977e-08, 
    -1.166026e-08, -1.154608e-08, -1.144351e-08, -1.138955e-08, 
    -1.143026e-08, -1.153963e-08, -1.173625e-08, -1.210359e-08, 
    -1.254808e-08, -1.302821e-08,
  -1.083262e-08, -1.102025e-08, -1.130623e-08, -1.143874e-08, -1.1648e-08, 
    -1.179431e-08, -1.184407e-08, -1.176692e-08, -1.176573e-08, 
    -1.181719e-08, -1.186563e-08, -1.186929e-08, -1.196349e-08, 
    -1.211142e-08, -1.235597e-08,
  -1.125954e-08, -1.130242e-08, -1.135387e-08, -1.124765e-08, -1.132259e-08, 
    -1.153761e-08, -1.188156e-08, -1.207856e-08, -1.216641e-08, 
    -1.227641e-08, -1.250428e-08, -1.257984e-08, -1.259972e-08, 
    -1.263247e-08, -1.270127e-08,
  -1.173545e-08, -1.176025e-08, -1.157535e-08, -1.127136e-08, -1.106341e-08, 
    -1.106781e-08, -1.134091e-08, -1.165558e-08, -1.193257e-08, 
    -1.215059e-08, -1.24089e-08, -1.274569e-08, -1.295333e-08, -1.310477e-08, 
    -1.317009e-08,
  -1.230087e-08, -1.218072e-08, -1.171447e-08, -1.123866e-08, -1.087703e-08, 
    -1.06637e-08, -1.078241e-08, -1.10086e-08, -1.132694e-08, -1.167728e-08, 
    -1.1918e-08, -1.219442e-08, -1.255099e-08, -1.284069e-08, -1.303017e-08,
  -1.292538e-08, -1.275938e-08, -1.211855e-08, -1.143021e-08, -1.073706e-08, 
    -1.015001e-08, -1.010867e-08, -1.02155e-08, -1.036926e-08, -1.066579e-08, 
    -1.090701e-08, -1.112612e-08, -1.139821e-08, -1.178592e-08, -1.214725e-08,
  -1.361753e-08, -1.364624e-08, -1.316549e-08, -1.231771e-08, -1.134767e-08, 
    -1.030774e-08, -9.819781e-09, -9.571297e-09, -9.509634e-09, 
    -9.551742e-09, -9.649295e-09, -9.693744e-09, -9.779589e-09, 
    -9.891542e-09, -1.013819e-08,
  -1.432391e-08, -1.468053e-08, -1.407748e-08, -1.315488e-08, -1.178119e-08, 
    -1.081744e-08, -1.031405e-08, -9.933738e-09, -9.783993e-09, -9.6562e-09, 
    -9.605357e-09, -9.526817e-09, -9.489034e-09, -9.396661e-09, -9.355e-09,
  -1.485893e-08, -1.525141e-08, -1.542751e-08, -1.563709e-08, -1.555802e-08, 
    -1.541107e-08, -1.513685e-08, -1.469687e-08, -1.431721e-08, 
    -1.390445e-08, -1.369612e-08, -1.325057e-08, -1.283925e-08, 
    -1.207117e-08, -1.127592e-08,
  -1.423651e-08, -1.44475e-08, -1.441699e-08, -1.475205e-08, -1.492602e-08, 
    -1.49835e-08, -1.487323e-08, -1.461835e-08, -1.43028e-08, -1.38709e-08, 
    -1.351509e-08, -1.304782e-08, -1.252397e-08, -1.183236e-08, -1.095572e-08,
  -1.338778e-08, -1.343716e-08, -1.339667e-08, -1.346179e-08, -1.35597e-08, 
    -1.369904e-08, -1.375509e-08, -1.372929e-08, -1.355603e-08, 
    -1.330255e-08, -1.296091e-08, -1.254419e-08, -1.202447e-08, 
    -1.137832e-08, -1.068837e-08,
  -1.276353e-08, -1.269376e-08, -1.240899e-08, -1.253225e-08, -1.260488e-08, 
    -1.283012e-08, -1.302552e-08, -1.312477e-08, -1.310229e-08, 
    -1.294015e-08, -1.258582e-08, -1.220697e-08, -1.175229e-08, 
    -1.132341e-08, -1.081025e-08,
  -1.225124e-08, -1.220281e-08, -1.19425e-08, -1.183908e-08, -1.174713e-08, 
    -1.171624e-08, -1.174991e-08, -1.186627e-08, -1.189833e-08, 
    -1.185776e-08, -1.166528e-08, -1.139842e-08, -1.102663e-08, 
    -1.057001e-08, -9.928382e-09,
  -1.134254e-08, -1.162015e-08, -1.146407e-08, -1.139548e-08, -1.121932e-08, 
    -1.108052e-08, -1.09042e-08, -1.081254e-08, -1.068517e-08, -1.059512e-08, 
    -1.042222e-08, -1.021142e-08, -9.877087e-09, -9.487811e-09, -9.044086e-09,
  -1.032551e-08, -1.062203e-08, -1.072372e-08, -1.071181e-08, -1.069609e-08, 
    -1.061393e-08, -1.049909e-08, -1.035998e-08, -1.023451e-08, 
    -1.006656e-08, -9.906921e-09, -9.668432e-09, -9.417137e-09, -9.06679e-09, 
    -8.686679e-09,
  -9.808098e-09, -9.871707e-09, -9.895372e-09, -9.881832e-09, -9.870361e-09, 
    -9.810941e-09, -9.728368e-09, -9.603001e-09, -9.506325e-09, 
    -9.404205e-09, -9.306535e-09, -9.18906e-09, -9.031452e-09, -8.790073e-09, 
    -8.493659e-09,
  -9.745307e-09, -9.606571e-09, -9.539432e-09, -9.443037e-09, -9.391705e-09, 
    -9.326862e-09, -9.291296e-09, -9.216678e-09, -9.145834e-09, 
    -9.061025e-09, -8.966883e-09, -8.871702e-09, -8.768863e-09, 
    -8.596732e-09, -8.359439e-09,
  -9.555209e-09, -9.420947e-09, -9.331385e-09, -9.225991e-09, -9.153439e-09, 
    -9.081322e-09, -9.026617e-09, -8.982005e-09, -8.94926e-09, -8.913086e-09, 
    -8.871116e-09, -8.811765e-09, -8.729158e-09, -8.628333e-09, -8.475759e-09,
  -1.087998e-08, -1.044194e-08, -9.954808e-09, -9.389514e-09, -8.853246e-09, 
    -8.227588e-09, -7.625545e-09, -7.016621e-09, -6.403099e-09, 
    -5.784986e-09, -5.127764e-09, -4.528688e-09, -4.076531e-09, 
    -3.900746e-09, -4.065755e-09,
  -9.814205e-09, -9.77098e-09, -9.437926e-09, -9.078247e-09, -8.550915e-09, 
    -8.032105e-09, -7.449704e-09, -6.934485e-09, -6.339155e-09, 
    -5.727642e-09, -5.027185e-09, -4.431954e-09, -4.045693e-09, 
    -3.926331e-09, -4.254389e-09,
  -8.555419e-09, -8.623056e-09, -8.551557e-09, -8.311051e-09, -8.010739e-09, 
    -7.652181e-09, -7.206054e-09, -6.694456e-09, -6.087283e-09, 
    -5.433274e-09, -4.773774e-09, -4.278902e-09, -4.010717e-09, 
    -3.991882e-09, -4.453464e-09,
  -7.881319e-09, -7.889755e-09, -7.953136e-09, -7.939597e-09, -7.77644e-09, 
    -7.49904e-09, -7.115783e-09, -6.610354e-09, -6.030219e-09, -5.424625e-09, 
    -4.85572e-09, -4.388982e-09, -4.159337e-09, -4.13456e-09, -4.698147e-09,
  -7.17721e-09, -7.033037e-09, -6.982409e-09, -6.94165e-09, -6.89451e-09, 
    -6.770019e-09, -6.545524e-09, -6.198122e-09, -5.725157e-09, 
    -5.219279e-09, -4.698251e-09, -4.304522e-09, -4.101112e-09, 
    -4.174416e-09, -4.820334e-09,
  -6.598305e-09, -6.450848e-09, -6.403785e-09, -6.283197e-09, -6.241171e-09, 
    -6.140464e-09, -5.952189e-09, -5.643957e-09, -5.233139e-09, 
    -4.808657e-09, -4.409247e-09, -4.113317e-09, -3.987926e-09, 
    -4.182319e-09, -4.893567e-09,
  -6.351705e-09, -5.989297e-09, -5.842835e-09, -5.646581e-09, -5.580947e-09, 
    -5.432775e-09, -5.289726e-09, -5.001215e-09, -4.683681e-09, 
    -4.384805e-09, -4.128978e-09, -3.952493e-09, -3.963105e-09, -4.25013e-09, 
    -4.926792e-09,
  -6.397742e-09, -5.96782e-09, -5.664495e-09, -5.358555e-09, -5.167078e-09, 
    -4.986735e-09, -4.84413e-09, -4.627042e-09, -4.372996e-09, -4.117175e-09, 
    -3.923328e-09, -3.823614e-09, -3.951051e-09, -4.305193e-09, -4.92714e-09,
  -6.779826e-09, -6.282252e-09, -5.934754e-09, -5.537085e-09, -5.264124e-09, 
    -4.995615e-09, -4.762421e-09, -4.515028e-09, -4.259625e-09, 
    -4.021002e-09, -3.851123e-09, -3.812499e-09, -3.975354e-09, 
    -4.304025e-09, -4.890755e-09,
  -7.834741e-09, -7.256449e-09, -6.820466e-09, -6.312994e-09, -5.86715e-09, 
    -5.439092e-09, -5.065429e-09, -4.748458e-09, -4.449225e-09, 
    -4.180969e-09, -3.989265e-09, -3.950235e-09, -4.071445e-09, 
    -4.352521e-09, -4.852315e-09,
  -5.576622e-09, -5.457142e-09, -5.391288e-09, -5.362957e-09, -5.304817e-09, 
    -5.346894e-09, -5.423182e-09, -5.536597e-09, -5.540336e-09, 
    -5.492958e-09, -5.443196e-09, -5.725405e-09, -6.859803e-09, 
    -9.011782e-09, -1.25672e-08,
  -6.035004e-09, -5.699507e-09, -5.454091e-09, -5.308844e-09, -5.283787e-09, 
    -5.266498e-09, -5.432358e-09, -5.4975e-09, -5.355156e-09, -5.27643e-09, 
    -5.216083e-09, -5.494163e-09, -6.599956e-09, -8.546557e-09, -1.174706e-08,
  -6.007479e-09, -5.839862e-09, -5.593148e-09, -5.412269e-09, -5.318945e-09, 
    -5.249884e-09, -5.347828e-09, -5.415075e-09, -5.152866e-09, 
    -4.999284e-09, -4.960549e-09, -5.264276e-09, -6.366483e-09, 
    -8.203198e-09, -1.115761e-08,
  -5.885105e-09, -5.990927e-09, -5.685072e-09, -5.49959e-09, -5.318116e-09, 
    -5.236716e-09, -5.248759e-09, -5.221994e-09, -4.942892e-09, 
    -4.738522e-09, -4.700058e-09, -5.098442e-09, -6.170851e-09, 
    -7.845733e-09, -1.06527e-08,
  -5.446399e-09, -5.793708e-09, -5.696167e-09, -5.478697e-09, -5.252597e-09, 
    -5.15496e-09, -5.121619e-09, -5.035967e-09, -4.694471e-09, -4.464323e-09, 
    -4.419077e-09, -4.926037e-09, -5.997558e-09, -7.57082e-09, -1.033953e-08,
  -4.911669e-09, -5.347252e-09, -5.25375e-09, -5.273789e-09, -5.07581e-09, 
    -4.938572e-09, -4.870649e-09, -4.782096e-09, -4.431446e-09, 
    -4.201824e-09, -4.179951e-09, -4.732902e-09, -5.857764e-09, 
    -7.465015e-09, -1.017989e-08,
  -4.274566e-09, -4.695413e-09, -4.759801e-09, -4.840478e-09, -4.729511e-09, 
    -4.640018e-09, -4.590944e-09, -4.469961e-09, -4.164012e-09, 
    -3.998004e-09, -3.993585e-09, -4.612207e-09, -5.781272e-09, 
    -7.503319e-09, -1.031439e-08,
  -3.786664e-09, -4.112068e-09, -4.320597e-09, -4.388792e-09, -4.361208e-09, 
    -4.301679e-09, -4.278182e-09, -4.151238e-09, -3.932334e-09, 
    -3.851945e-09, -3.898279e-09, -4.548943e-09, -5.817551e-09, 
    -7.740083e-09, -1.056832e-08,
  -3.454927e-09, -3.651196e-09, -3.855409e-09, -3.990607e-09, -4.002793e-09, 
    -4.02108e-09, -4.000166e-09, -3.927421e-09, -3.850803e-09, -3.908214e-09, 
    -3.965891e-09, -4.633514e-09, -5.988678e-09, -8.247044e-09, -1.111907e-08,
  -3.455248e-09, -3.52632e-09, -3.672157e-09, -3.838301e-09, -3.868961e-09, 
    -3.880824e-09, -3.850452e-09, -3.82825e-09, -3.895865e-09, -4.093543e-09, 
    -4.257354e-09, -5.033144e-09, -6.480351e-09, -8.891181e-09, -1.146982e-08,
  -4.951852e-09, -5.200692e-09, -5.477396e-09, -5.88462e-09, -6.711247e-09, 
    -7.830036e-09, -9.010892e-09, -1.014372e-08, -1.156457e-08, 
    -1.281003e-08, -1.458265e-08, -1.615425e-08, -1.820795e-08, 
    -2.066766e-08, -2.365888e-08,
  -4.771167e-09, -5.057703e-09, -5.240616e-09, -5.481601e-09, -6.044614e-09, 
    -6.982194e-09, -8.150311e-09, -9.336816e-09, -1.082361e-08, 
    -1.220788e-08, -1.377138e-08, -1.563609e-08, -1.764095e-08, 
    -2.018637e-08, -2.346337e-08,
  -4.71e-09, -4.892335e-09, -5.084289e-09, -5.189062e-09, -5.530119e-09, 
    -6.320635e-09, -7.361084e-09, -8.524547e-09, -9.99644e-09, -1.15334e-08, 
    -1.315559e-08, -1.497713e-08, -1.693133e-08, -1.96624e-08, -2.319092e-08,
  -4.914039e-09, -4.858553e-09, -4.94419e-09, -5.001935e-09, -5.14617e-09, 
    -5.733973e-09, -6.675442e-09, -7.730105e-09, -9.21113e-09, -1.075031e-08, 
    -1.241114e-08, -1.438333e-08, -1.641521e-08, -1.904664e-08, -2.279971e-08,
  -5.294409e-09, -5.031318e-09, -4.98036e-09, -4.926837e-09, -4.966371e-09, 
    -5.334456e-09, -6.068271e-09, -6.968001e-09, -8.412957e-09, 
    -9.998659e-09, -1.164035e-08, -1.381767e-08, -1.590087e-08, 
    -1.848771e-08, -2.227719e-08,
  -5.594163e-09, -5.255433e-09, -5.082412e-09, -4.955733e-09, -4.904605e-09, 
    -5.08905e-09, -5.642545e-09, -6.360715e-09, -7.648103e-09, -9.241856e-09, 
    -1.089119e-08, -1.31652e-08, -1.552168e-08, -1.803204e-08, -2.188914e-08,
  -5.83116e-09, -5.561934e-09, -5.170141e-09, -5.166454e-09, -4.922287e-09, 
    -5.010568e-09, -5.307155e-09, -5.863947e-09, -6.997478e-09, 
    -8.576932e-09, -1.020453e-08, -1.251874e-08, -1.513487e-08, 
    -1.778702e-08, -2.145771e-08,
  -6.000757e-09, -5.805937e-09, -5.287485e-09, -5.218192e-09, -4.992192e-09, 
    -5.064611e-09, -5.187938e-09, -5.510632e-09, -6.454276e-09, 
    -7.985894e-09, -9.527525e-09, -1.184734e-08, -1.476495e-08, 
    -1.750592e-08, -2.121633e-08,
  -5.909035e-09, -5.826264e-09, -5.408721e-09, -5.1794e-09, -5.057949e-09, 
    -5.165498e-09, -5.130472e-09, -5.356246e-09, -6.050263e-09, 
    -7.465337e-09, -8.948454e-09, -1.118451e-08, -1.428837e-08, 
    -1.736609e-08, -2.094793e-08,
  -5.821903e-09, -5.755417e-09, -5.466967e-09, -5.188495e-09, -5.109034e-09, 
    -5.108796e-09, -5.073763e-09, -5.251095e-09, -5.797952e-09, 
    -7.068528e-09, -8.492665e-09, -1.057998e-08, -1.378166e-08, 
    -1.714511e-08, -2.080728e-08,
  -1.063678e-08, -1.145042e-08, -1.246011e-08, -1.328881e-08, -1.319015e-08, 
    -1.282758e-08, -1.212256e-08, -1.245138e-08, -1.2698e-08, -1.259983e-08, 
    -1.194661e-08, -9.682008e-09, -1.087494e-08, -1.326141e-08, -1.537846e-08,
  -9.963687e-09, -1.111401e-08, -1.228958e-08, -1.353793e-08, -1.401641e-08, 
    -1.340567e-08, -1.262205e-08, -1.279308e-08, -1.359902e-08, 
    -1.467893e-08, -1.319702e-08, -1.107452e-08, -1.210791e-08, 
    -1.334694e-08, -1.482032e-08,
  -9.509773e-09, -1.04118e-08, -1.186441e-08, -1.327802e-08, -1.406036e-08, 
    -1.349486e-08, -1.310779e-08, -1.343589e-08, -1.446792e-08, 
    -1.641191e-08, -1.407481e-08, -1.252217e-08, -1.364162e-08, 
    -1.436196e-08, -1.480604e-08,
  -8.869803e-09, -9.95052e-09, -1.132597e-08, -1.258929e-08, -1.34453e-08, 
    -1.321725e-08, -1.337777e-08, -1.360756e-08, -1.514525e-08, 
    -1.768598e-08, -1.545982e-08, -1.520322e-08, -1.640238e-08, 
    -1.505452e-08, -1.492063e-08,
  -8.291167e-09, -9.456288e-09, -1.088821e-08, -1.210039e-08, -1.269742e-08, 
    -1.258741e-08, -1.286835e-08, -1.328332e-08, -1.473865e-08, 
    -1.808742e-08, -1.646601e-08, -1.645814e-08, -1.716952e-08, 
    -1.563598e-08, -1.500668e-08,
  -7.770829e-09, -9.109968e-09, -1.056739e-08, -1.178713e-08, -1.221907e-08, 
    -1.199582e-08, -1.248275e-08, -1.308132e-08, -1.473783e-08, -1.78192e-08, 
    -1.632488e-08, -1.652486e-08, -1.672862e-08, -1.518048e-08, -1.601865e-08,
  -7.262897e-09, -8.714596e-09, -1.034714e-08, -1.134116e-08, -1.168559e-08, 
    -1.165399e-08, -1.246164e-08, -1.305482e-08, -1.483468e-08, 
    -1.721311e-08, -1.579592e-08, -1.558132e-08, -1.565068e-08, 
    -1.552016e-08, -1.83382e-08,
  -6.839703e-09, -8.301011e-09, -9.896426e-09, -1.08364e-08, -1.132953e-08, 
    -1.160875e-08, -1.24124e-08, -1.317052e-08, -1.483138e-08, -1.59349e-08, 
    -1.492081e-08, -1.551375e-08, -1.636745e-08, -1.776678e-08, -2.065199e-08,
  -6.496102e-09, -7.835537e-09, -9.390178e-09, -1.047657e-08, -1.088815e-08, 
    -1.1328e-08, -1.219244e-08, -1.296994e-08, -1.428517e-08, -1.467205e-08, 
    -1.457532e-08, -1.633432e-08, -1.759513e-08, -1.950681e-08, -2.444997e-08,
  -6.219915e-09, -7.469101e-09, -8.960766e-09, -1.009063e-08, -1.041768e-08, 
    -1.082449e-08, -1.171334e-08, -1.264573e-08, -1.375444e-08, 
    -1.391167e-08, -1.498884e-08, -1.695163e-08, -1.896334e-08, 
    -2.351243e-08, -2.909328e-08,
  -1.109614e-08, -1.121235e-08, -1.135979e-08, -1.16065e-08, -1.199319e-08, 
    -1.250089e-08, -1.31343e-08, -1.401649e-08, -1.479568e-08, -1.540724e-08, 
    -1.608355e-08, -1.65068e-08, -1.679729e-08, -1.69385e-08, -1.696145e-08,
  -1.186711e-08, -1.175187e-08, -1.18363e-08, -1.178948e-08, -1.19581e-08, 
    -1.237135e-08, -1.282924e-08, -1.344631e-08, -1.415976e-08, 
    -1.478053e-08, -1.534441e-08, -1.582564e-08, -1.626358e-08, 
    -1.655224e-08, -1.663758e-08,
  -1.231894e-08, -1.223684e-08, -1.231707e-08, -1.230339e-08, -1.249729e-08, 
    -1.251138e-08, -1.270129e-08, -1.299404e-08, -1.359221e-08, 
    -1.409985e-08, -1.472686e-08, -1.515588e-08, -1.554232e-08, 
    -1.590683e-08, -1.617773e-08,
  -1.353178e-08, -1.326611e-08, -1.322418e-08, -1.316023e-08, -1.297744e-08, 
    -1.234135e-08, -1.2312e-08, -1.266253e-08, -1.304628e-08, -1.343545e-08, 
    -1.406472e-08, -1.450025e-08, -1.490292e-08, -1.528705e-08, -1.568111e-08,
  -1.383477e-08, -1.359384e-08, -1.337594e-08, -1.30598e-08, -1.249794e-08, 
    -1.182064e-08, -1.203867e-08, -1.224899e-08, -1.260133e-08, 
    -1.280389e-08, -1.331677e-08, -1.383025e-08, -1.421904e-08, 
    -1.468345e-08, -1.510205e-08,
  -1.335132e-08, -1.328301e-08, -1.292155e-08, -1.243317e-08, -1.191984e-08, 
    -1.181207e-08, -1.202467e-08, -1.228422e-08, -1.243382e-08, 
    -1.266404e-08, -1.311155e-08, -1.353348e-08, -1.391951e-08, 
    -1.432384e-08, -1.467218e-08,
  -1.303809e-08, -1.306479e-08, -1.270024e-08, -1.167222e-08, -1.151506e-08, 
    -1.143848e-08, -1.209598e-08, -1.246571e-08, -1.242767e-08, 
    -1.245137e-08, -1.273236e-08, -1.303897e-08, -1.335066e-08, 
    -1.393079e-08, -1.436704e-08,
  -1.30714e-08, -1.309968e-08, -1.258322e-08, -1.178297e-08, -1.159456e-08, 
    -1.167268e-08, -1.208216e-08, -1.207371e-08, -1.206727e-08, 
    -1.215663e-08, -1.244774e-08, -1.274182e-08, -1.327916e-08, 
    -1.384106e-08, -1.438004e-08,
  -1.335928e-08, -1.34795e-08, -1.29565e-08, -1.250588e-08, -1.224651e-08, 
    -1.220843e-08, -1.211181e-08, -1.205718e-08, -1.224306e-08, 
    -1.240564e-08, -1.271645e-08, -1.295269e-08, -1.343776e-08, 
    -1.392023e-08, -1.446353e-08,
  -1.377165e-08, -1.412083e-08, -1.386806e-08, -1.375406e-08, -1.358167e-08, 
    -1.336271e-08, -1.315154e-08, -1.307264e-08, -1.30815e-08, -1.308575e-08, 
    -1.335801e-08, -1.348009e-08, -1.392371e-08, -1.449617e-08, -1.527607e-08,
  -1.469812e-08, -1.597189e-08, -1.607926e-08, -1.5773e-08, -1.536649e-08, 
    -1.520626e-08, -1.531683e-08, -1.638635e-08, -1.808803e-08, 
    -1.930337e-08, -2.050304e-08, -2.18795e-08, -2.467937e-08, -2.745387e-08, 
    -2.788346e-08,
  -1.357601e-08, -1.459302e-08, -1.536769e-08, -1.612471e-08, -1.608e-08, 
    -1.558801e-08, -1.546412e-08, -1.642719e-08, -1.761631e-08, 
    -1.864768e-08, -1.969638e-08, -2.106521e-08, -2.289346e-08, 
    -2.540103e-08, -2.628125e-08,
  -1.308561e-08, -1.375339e-08, -1.458192e-08, -1.50432e-08, -1.571334e-08, 
    -1.605791e-08, -1.563939e-08, -1.616507e-08, -1.707185e-08, 
    -1.795581e-08, -1.887143e-08, -2.007588e-08, -2.156362e-08, 
    -2.364596e-08, -2.497468e-08,
  -1.327038e-08, -1.354659e-08, -1.389339e-08, -1.437702e-08, -1.501525e-08, 
    -1.541641e-08, -1.556246e-08, -1.652728e-08, -1.725084e-08, 
    -1.811121e-08, -1.861866e-08, -1.953624e-08, -2.049053e-08, 
    -2.199264e-08, -2.368741e-08,
  -1.441558e-08, -1.424502e-08, -1.442588e-08, -1.474147e-08, -1.517817e-08, 
    -1.555632e-08, -1.596444e-08, -1.683075e-08, -1.717595e-08, 
    -1.798161e-08, -1.84616e-08, -1.924378e-08, -1.983688e-08, -2.065861e-08, 
    -2.187491e-08,
  -1.449996e-08, -1.456056e-08, -1.484043e-08, -1.483603e-08, -1.517158e-08, 
    -1.560786e-08, -1.613188e-08, -1.682028e-08, -1.729063e-08, -1.81178e-08, 
    -1.833322e-08, -1.881869e-08, -1.915449e-08, -1.961202e-08, -2.050005e-08,
  -1.369801e-08, -1.414571e-08, -1.453839e-08, -1.475011e-08, -1.508825e-08, 
    -1.547953e-08, -1.600839e-08, -1.650172e-08, -1.702658e-08, 
    -1.744222e-08, -1.762556e-08, -1.805723e-08, -1.830236e-08, 
    -1.862328e-08, -1.911767e-08,
  -1.347644e-08, -1.366596e-08, -1.39442e-08, -1.427521e-08, -1.462549e-08, 
    -1.494212e-08, -1.528559e-08, -1.565222e-08, -1.605007e-08, 
    -1.631002e-08, -1.671021e-08, -1.716217e-08, -1.737389e-08, 
    -1.771287e-08, -1.800482e-08,
  -1.410361e-08, -1.383345e-08, -1.388822e-08, -1.390433e-08, -1.426222e-08, 
    -1.449665e-08, -1.485662e-08, -1.503196e-08, -1.521787e-08, 
    -1.542251e-08, -1.572292e-08, -1.599425e-08, -1.648758e-08, 
    -1.682603e-08, -1.713256e-08,
  -1.5567e-08, -1.498336e-08, -1.481709e-08, -1.46037e-08, -1.460199e-08, 
    -1.453937e-08, -1.462106e-08, -1.478595e-08, -1.491544e-08, 
    -1.503749e-08, -1.522721e-08, -1.556758e-08, -1.590754e-08, 
    -1.618428e-08, -1.64916e-08,
  -1.222351e-08, -1.206581e-08, -1.235824e-08, -1.294611e-08, -1.388727e-08, 
    -1.546436e-08, -1.823088e-08, -2.180898e-08, -2.379551e-08, -2.63502e-08, 
    -3.060885e-08, -3.085088e-08, -2.762771e-08, -2.479403e-08, -2.035085e-08,
  -1.305389e-08, -1.256335e-08, -1.282844e-08, -1.319197e-08, -1.408823e-08, 
    -1.556789e-08, -1.843038e-08, -2.179456e-08, -2.339353e-08, 
    -2.621964e-08, -2.997241e-08, -3.003176e-08, -2.832915e-08, 
    -2.601216e-08, -2.242664e-08,
  -1.477093e-08, -1.380382e-08, -1.362377e-08, -1.364522e-08, -1.44034e-08, 
    -1.564238e-08, -1.836223e-08, -2.115782e-08, -2.261623e-08, 
    -2.531947e-08, -2.895532e-08, -2.952427e-08, -2.918246e-08, 
    -2.681591e-08, -2.364132e-08,
  -1.721426e-08, -1.592232e-08, -1.531572e-08, -1.512536e-08, -1.539904e-08, 
    -1.654877e-08, -1.860876e-08, -2.081694e-08, -2.166708e-08, 
    -2.438237e-08, -2.807819e-08, -2.895002e-08, -2.921879e-08, 
    -2.735588e-08, -2.479515e-08,
  -1.923304e-08, -1.839912e-08, -1.74089e-08, -1.704329e-08, -1.705471e-08, 
    -1.754434e-08, -1.882482e-08, -2.006703e-08, -2.079687e-08, 
    -2.349706e-08, -2.681657e-08, -2.737298e-08, -2.817157e-08, 
    -2.726619e-08, -2.556256e-08,
  -1.903444e-08, -1.939926e-08, -1.912773e-08, -1.888177e-08, -1.878789e-08, 
    -1.913295e-08, -1.952203e-08, -2.009911e-08, -2.085206e-08, 
    -2.334177e-08, -2.545954e-08, -2.642644e-08, -2.783475e-08, 
    -2.763282e-08, -2.587383e-08,
  -1.794051e-08, -1.893095e-08, -1.921433e-08, -1.968739e-08, -1.995575e-08, 
    -2.018437e-08, -1.997547e-08, -2.010091e-08, -2.086434e-08, 
    -2.205118e-08, -2.361394e-08, -2.500428e-08, -2.678967e-08, 
    -2.656185e-08, -2.505666e-08,
  -1.75732e-08, -1.762989e-08, -1.805167e-08, -1.885968e-08, -1.980727e-08, 
    -2.033487e-08, -2.03346e-08, -2.029403e-08, -2.052681e-08, -2.097459e-08, 
    -2.206445e-08, -2.369441e-08, -2.588173e-08, -2.560572e-08, -2.452865e-08,
  -1.799716e-08, -1.754156e-08, -1.738977e-08, -1.721195e-08, -1.796924e-08, 
    -1.86923e-08, -1.932129e-08, -1.944602e-08, -1.970089e-08, -1.999856e-08, 
    -2.111533e-08, -2.320326e-08, -2.437616e-08, -2.403935e-08, -2.337328e-08,
  -1.8538e-08, -1.801989e-08, -1.757292e-08, -1.759972e-08, -1.728516e-08, 
    -1.771853e-08, -1.82319e-08, -1.915942e-08, -1.940159e-08, -2.032775e-08, 
    -2.117388e-08, -2.24194e-08, -2.272125e-08, -2.267555e-08, -2.256947e-08,
  -1.46495e-08, -1.493549e-08, -1.610483e-08, -1.745737e-08, -1.915625e-08, 
    -2.080856e-08, -2.207843e-08, -2.340764e-08, -2.569465e-08, 
    -2.639515e-08, -2.302698e-08, -1.960218e-08, -1.678008e-08, 
    -1.152317e-08, -6.615164e-09,
  -1.502192e-08, -1.502331e-08, -1.610564e-08, -1.69536e-08, -1.898396e-08, 
    -2.044001e-08, -2.274487e-08, -2.471273e-08, -2.840527e-08, 
    -2.849242e-08, -2.339493e-08, -2.091348e-08, -1.891096e-08, 
    -1.428671e-08, -8.546556e-09,
  -1.529608e-08, -1.488943e-08, -1.542266e-08, -1.63584e-08, -1.88485e-08, 
    -2.123298e-08, -2.416095e-08, -2.695944e-08, -2.898166e-08, 
    -2.846766e-08, -2.346437e-08, -2.158171e-08, -1.98604e-08, -1.592223e-08, 
    -1.002324e-08,
  -1.690303e-08, -1.666326e-08, -1.742904e-08, -1.867338e-08, -2.115343e-08, 
    -2.375573e-08, -2.558705e-08, -2.808366e-08, -2.873117e-08, 
    -2.843523e-08, -2.466202e-08, -2.238758e-08, -2.070211e-08, 
    -1.779803e-08, -1.183139e-08,
  -2.147702e-08, -2.111102e-08, -2.182061e-08, -2.281187e-08, -2.437091e-08, 
    -2.557358e-08, -2.646293e-08, -2.866331e-08, -2.903882e-08, -2.86402e-08, 
    -2.573334e-08, -2.304921e-08, -2.15253e-08, -1.89587e-08, -1.32117e-08,
  -2.681924e-08, -2.563855e-08, -2.570143e-08, -2.596659e-08, -2.63063e-08, 
    -2.696094e-08, -2.799023e-08, -2.964654e-08, -3.003302e-08, 
    -2.923406e-08, -2.723449e-08, -2.42228e-08, -2.227265e-08, -1.999004e-08, 
    -1.439642e-08,
  -2.834911e-08, -2.84397e-08, -2.820073e-08, -2.79104e-08, -2.798059e-08, 
    -2.826964e-08, -2.876699e-08, -2.998129e-08, -3.018248e-08, 
    -2.956755e-08, -2.808122e-08, -2.462922e-08, -2.278786e-08, 
    -2.062191e-08, -1.525291e-08,
  -2.621659e-08, -2.7271e-08, -2.812095e-08, -2.839511e-08, -2.891956e-08, 
    -2.925432e-08, -2.994559e-08, -3.038629e-08, -3.047122e-08, 
    -2.907846e-08, -2.696748e-08, -2.452153e-08, -2.318773e-08, 
    -2.077688e-08, -1.588888e-08,
  -2.249295e-08, -2.420777e-08, -2.503562e-08, -2.598859e-08, -2.678362e-08, 
    -2.72486e-08, -2.77668e-08, -2.73896e-08, -2.673033e-08, -2.534679e-08, 
    -2.446237e-08, -2.330821e-08, -2.232684e-08, -2.089511e-08, -1.608745e-08,
  -2.068061e-08, -2.11782e-08, -2.17278e-08, -2.219315e-08, -2.272259e-08, 
    -2.305312e-08, -2.316487e-08, -2.333093e-08, -2.336019e-08, 
    -2.316895e-08, -2.242004e-08, -2.19544e-08, -2.17792e-08, -2.036555e-08, 
    -1.614293e-08,
  -1.778653e-08, -1.767655e-08, -1.821461e-08, -1.994596e-08, -2.157159e-08, 
    -2.465481e-08, -2.613322e-08, -2.678703e-08, -2.384599e-08, 
    -2.107825e-08, -1.640074e-08, -9.931238e-09, -4.204264e-09, 
    -2.491607e-09, -2.172545e-09,
  -1.77367e-08, -1.80036e-08, -1.907133e-08, -2.038965e-08, -2.262435e-08, 
    -2.579382e-08, -2.775469e-08, -2.76603e-08, -2.585583e-08, -2.310454e-08, 
    -1.953883e-08, -1.4243e-08, -6.550342e-09, -2.934289e-09, -2.351241e-09,
  -1.60329e-08, -1.737578e-08, -1.850764e-08, -2.015621e-08, -2.31314e-08, 
    -2.575796e-08, -2.701681e-08, -2.614319e-08, -2.54812e-08, -2.300363e-08, 
    -2.039921e-08, -1.635794e-08, -8.675609e-09, -3.667625e-09, -2.612208e-09,
  -1.674225e-08, -1.746895e-08, -1.872377e-08, -1.982357e-08, -2.258885e-08, 
    -2.416533e-08, -2.559532e-08, -2.546958e-08, -2.616303e-08, 
    -2.396368e-08, -2.173237e-08, -1.834314e-08, -1.084496e-08, 
    -4.686667e-09, -2.952851e-09,
  -1.854099e-08, -1.827371e-08, -1.863681e-08, -1.940866e-08, -2.121296e-08, 
    -2.254118e-08, -2.435073e-08, -2.462244e-08, -2.445998e-08, 
    -2.367278e-08, -2.171426e-08, -1.930292e-08, -1.254281e-08, 
    -5.903669e-09, -3.330109e-09,
  -1.957739e-08, -1.921804e-08, -1.904614e-08, -1.947075e-08, -2.120823e-08, 
    -2.323519e-08, -2.50788e-08, -2.452929e-08, -2.419431e-08, -2.420194e-08, 
    -2.206698e-08, -1.983489e-08, -1.419945e-08, -7.02531e-09, -3.751389e-09,
  -2.277869e-08, -2.157122e-08, -2.201898e-08, -2.215963e-08, -2.38589e-08, 
    -2.434408e-08, -2.471639e-08, -2.343995e-08, -2.368636e-08, 
    -2.248517e-08, -2.155267e-08, -2.029459e-08, -1.50196e-08, -8.113536e-09, 
    -4.167623e-09,
  -2.487365e-08, -2.4931e-08, -2.546111e-08, -2.534262e-08, -2.58007e-08, 
    -2.506488e-08, -2.489998e-08, -2.40003e-08, -2.393921e-08, -2.258381e-08, 
    -2.09378e-08, -1.996362e-08, -1.563051e-08, -8.669378e-09, -4.639518e-09,
  -2.26404e-08, -2.276696e-08, -2.267706e-08, -2.295392e-08, -2.322772e-08, 
    -2.28374e-08, -2.257919e-08, -2.225159e-08, -2.112195e-08, -2.014036e-08, 
    -2.006297e-08, -1.963786e-08, -1.53983e-08, -9.166037e-09, -4.931139e-09,
  -1.979103e-08, -1.973335e-08, -1.946889e-08, -1.92798e-08, -1.911439e-08, 
    -1.901155e-08, -1.898915e-08, -1.923498e-08, -1.934441e-08, 
    -1.972673e-08, -1.969335e-08, -1.906049e-08, -1.526491e-08, 
    -8.984691e-09, -5.175404e-09,
  -1.684958e-08, -1.581024e-08, -1.594753e-08, -1.636554e-08, -1.628194e-08, 
    -1.639099e-08, -1.344815e-08, -1.113845e-08, -8.905308e-09, 
    -6.991519e-09, -5.646765e-09, -5.470205e-09, -5.489587e-09, 
    -5.078642e-09, -4.724071e-09,
  -1.843861e-08, -1.808419e-08, -1.991787e-08, -2.066322e-08, -2.257327e-08, 
    -2.259483e-08, -2.018395e-08, -1.551186e-08, -1.104025e-08, 
    -8.437997e-09, -6.226316e-09, -5.595311e-09, -5.575842e-09, 
    -5.039241e-09, -4.682793e-09,
  -2.089428e-08, -2.165049e-08, -2.375965e-08, -2.535647e-08, -2.830197e-08, 
    -2.641278e-08, -2.252884e-08, -1.889254e-08, -1.451182e-08, 
    -9.901837e-09, -7.579342e-09, -6.081724e-09, -5.880906e-09, 
    -5.315929e-09, -5.203552e-09,
  -2.160533e-08, -2.272543e-08, -2.509003e-08, -2.701978e-08, -2.874275e-08, 
    -2.641803e-08, -2.258979e-08, -1.985672e-08, -1.66596e-08, -1.21043e-08, 
    -8.624088e-09, -6.621795e-09, -6.035076e-09, -5.653305e-09, -5.788574e-09,
  -2.339312e-08, -2.447715e-08, -2.652524e-08, -2.792131e-08, -2.839178e-08, 
    -2.594672e-08, -2.229591e-08, -2.075621e-08, -1.794992e-08, 
    -1.397064e-08, -1.019155e-08, -7.408437e-09, -6.256521e-09, 
    -5.811453e-09, -5.724829e-09,
  -2.567339e-08, -2.662359e-08, -2.923925e-08, -2.913533e-08, -2.851335e-08, 
    -2.469961e-08, -2.394434e-08, -2.083335e-08, -1.832619e-08, 
    -1.444181e-08, -1.114058e-08, -8.258351e-09, -6.316106e-09, 
    -5.666098e-09, -5.441044e-09,
  -2.859815e-08, -2.828156e-08, -2.837966e-08, -2.61379e-08, -2.485054e-08, 
    -2.36147e-08, -2.148475e-08, -1.905654e-08, -1.73564e-08, -1.48091e-08, 
    -1.179903e-08, -8.927998e-09, -6.538225e-09, -6.01566e-09, -5.658805e-09,
  -2.356373e-08, -2.383203e-08, -2.396753e-08, -2.246423e-08, -2.181216e-08, 
    -2.083157e-08, -1.937801e-08, -1.852882e-08, -1.659433e-08, 
    -1.441954e-08, -1.200389e-08, -9.17661e-09, -6.458221e-09, -5.898097e-09, 
    -5.618615e-09,
  -2.211214e-08, -2.165977e-08, -2.145677e-08, -2.02324e-08, -1.935725e-08, 
    -1.866609e-08, -1.797641e-08, -1.708484e-08, -1.535242e-08, 
    -1.403677e-08, -1.178758e-08, -9.510192e-09, -6.605089e-09, 
    -5.784706e-09, -5.464608e-09,
  -2.179595e-08, -2.1424e-08, -2.097882e-08, -1.969562e-08, -1.857137e-08, 
    -1.760673e-08, -1.693716e-08, -1.600746e-08, -1.480654e-08, 
    -1.345259e-08, -1.145244e-08, -9.287306e-09, -6.534354e-09, 
    -5.618685e-09, -5.402613e-09,
  -9.448514e-09, -8.619776e-09, -8.288982e-09, -7.990609e-09, -7.595867e-09, 
    -5.997486e-09, -5.353696e-09, -5.171773e-09, -6.196936e-09, 
    -7.755992e-09, -1.032891e-08, -1.15876e-08, -1.255717e-08, -1.345366e-08, 
    -1.362473e-08,
  -1.304064e-08, -1.20128e-08, -1.10059e-08, -9.843455e-09, -9.20034e-09, 
    -8.281557e-09, -7.220599e-09, -6.760018e-09, -6.893692e-09, 
    -7.411137e-09, -8.436177e-09, -1.012577e-08, -1.143485e-08, 
    -1.222113e-08, -1.248323e-08,
  -1.467326e-08, -1.539542e-08, -1.493047e-08, -1.373517e-08, -1.228125e-08, 
    -1.03177e-08, -9.009611e-09, -7.820933e-09, -7.565266e-09, -8.09067e-09, 
    -8.389892e-09, -9.61273e-09, -1.069336e-08, -1.150012e-08, -1.152711e-08,
  -1.199608e-08, -1.275181e-08, -1.38928e-08, -1.474527e-08, -1.384916e-08, 
    -1.216848e-08, -1.035752e-08, -9.041632e-09, -7.903226e-09, 
    -7.950146e-09, -8.049017e-09, -8.357165e-09, -9.361438e-09, 
    -1.050763e-08, -1.060959e-08,
  -9.440468e-09, -9.413693e-09, -9.438937e-09, -1.001476e-08, -1.165662e-08, 
    -1.203148e-08, -1.145691e-08, -9.996987e-09, -8.740627e-09, 
    -7.889487e-09, -7.692047e-09, -7.361378e-09, -7.966598e-09, 
    -9.213601e-09, -9.800845e-09,
  -1.038993e-08, -8.560408e-09, -8.088264e-09, -7.955113e-09, -8.354619e-09, 
    -8.842052e-09, -8.934002e-09, -8.584642e-09, -8.169953e-09, 
    -7.638311e-09, -7.177733e-09, -6.697741e-09, -6.841446e-09, 
    -7.673641e-09, -8.408867e-09,
  -1.124316e-08, -8.167985e-09, -6.98237e-09, -6.177303e-09, -6.313987e-09, 
    -6.724018e-09, -6.933484e-09, -7.093607e-09, -6.983008e-09, 
    -7.021881e-09, -6.570436e-09, -6.149968e-09, -5.906885e-09, 
    -6.475296e-09, -7.08027e-09,
  -1.268088e-08, -8.952556e-09, -6.697298e-09, -5.722843e-09, -5.296508e-09, 
    -5.480734e-09, -5.503769e-09, -5.591979e-09, -5.801669e-09, 
    -6.006854e-09, -5.630951e-09, -5.237393e-09, -5.215462e-09, 
    -5.502015e-09, -5.920743e-09,
  -1.332145e-08, -1.025938e-08, -6.73624e-09, -5.46402e-09, -4.838443e-09, 
    -4.8485e-09, -4.724547e-09, -4.785716e-09, -4.844688e-09, -4.904067e-09, 
    -4.803319e-09, -4.785597e-09, -4.755075e-09, -4.921497e-09, -5.127795e-09,
  -1.374002e-08, -1.152958e-08, -7.242708e-09, -5.33882e-09, -4.468855e-09, 
    -4.374127e-09, -4.189915e-09, -4.294959e-09, -4.196727e-09, 
    -4.070253e-09, -4.013352e-09, -4.171489e-09, -4.403796e-09, 
    -4.543762e-09, -4.709622e-09,
  -7.983232e-09, -7.985206e-09, -7.501385e-09, -7.578576e-09, -7.38288e-09, 
    -6.907724e-09, -6.152502e-09, -6.538894e-09, -6.557085e-09, 
    -5.760961e-09, -4.788819e-09, -3.940024e-09, -3.748183e-09, -3.52566e-09, 
    -3.255474e-09,
  -8.015195e-09, -8.369605e-09, -7.747154e-09, -7.55164e-09, -7.26719e-09, 
    -6.881995e-09, -6.440787e-09, -6.757666e-09, -6.958801e-09, 
    -6.530892e-09, -5.718214e-09, -4.654968e-09, -4.24324e-09, -4.095816e-09, 
    -3.869265e-09,
  -7.555325e-09, -8.383966e-09, -8.297364e-09, -7.869795e-09, -7.669395e-09, 
    -7.274364e-09, -7.039576e-09, -7.240927e-09, -7.386591e-09, 
    -7.121419e-09, -6.668953e-09, -5.593988e-09, -4.914551e-09, 
    -4.632121e-09, -4.367179e-09,
  -7.365905e-09, -8.064253e-09, -8.672634e-09, -8.435722e-09, -8.055391e-09, 
    -7.78679e-09, -7.643609e-09, -7.544465e-09, -7.615229e-09, -7.606373e-09, 
    -7.411046e-09, -6.867743e-09, -6.135013e-09, -5.423352e-09, -5.004752e-09,
  -7.421266e-09, -7.933583e-09, -8.47867e-09, -8.97324e-09, -8.865345e-09, 
    -8.487471e-09, -8.189435e-09, -7.925738e-09, -7.941165e-09, 
    -7.942596e-09, -8.053928e-09, -8.041009e-09, -7.572026e-09, 
    -6.776836e-09, -6.043876e-09,
  -7.658953e-09, -8.160772e-09, -8.394647e-09, -8.773666e-09, -9.069669e-09, 
    -9.073912e-09, -8.881701e-09, -8.612671e-09, -8.687135e-09, 
    -8.823245e-09, -9.050853e-09, -9.232651e-09, -9.072235e-09, 
    -8.468225e-09, -7.6865e-09,
  -7.964144e-09, -8.482611e-09, -8.792185e-09, -9.230356e-09, -9.707778e-09, 
    -1.003906e-08, -1.015993e-08, -1.01538e-08, -1.027915e-08, -1.033228e-08, 
    -1.044303e-08, -1.04232e-08, -1.030883e-08, -9.9049e-09, -9.091793e-09,
  -8.164776e-09, -8.968267e-09, -9.476872e-09, -9.813259e-09, -1.033932e-08, 
    -1.075134e-08, -1.098685e-08, -1.109728e-08, -1.113183e-08, 
    -1.117763e-08, -1.132119e-08, -1.126697e-08, -1.102458e-08, 
    -1.066355e-08, -1.003535e-08,
  -8.361035e-09, -9.430769e-09, -1.028295e-08, -1.085138e-08, -1.108815e-08, 
    -1.143884e-08, -1.152354e-08, -1.160127e-08, -1.166359e-08, 
    -1.166546e-08, -1.172383e-08, -1.151515e-08, -1.128409e-08, -1.10823e-08, 
    -1.084789e-08,
  -7.918677e-09, -9.072582e-09, -1.023304e-08, -1.102164e-08, -1.150886e-08, 
    -1.190236e-08, -1.208782e-08, -1.215993e-08, -1.222011e-08, 
    -1.218698e-08, -1.222217e-08, -1.203761e-08, -1.178987e-08, 
    -1.144091e-08, -1.120303e-08,
  -3.912704e-09, -3.442663e-09, -3.018934e-09, -2.608518e-09, -2.310844e-09, 
    -2.210862e-09, -2.20798e-09, -2.153409e-09, -1.96576e-09, -1.830916e-09, 
    -1.713519e-09, -1.774572e-09, -1.795553e-09, -1.801275e-09, -1.821816e-09,
  -4.263367e-09, -3.766348e-09, -3.365664e-09, -2.89887e-09, -2.495227e-09, 
    -2.254578e-09, -2.195093e-09, -2.153872e-09, -1.980033e-09, 
    -1.842545e-09, -1.690856e-09, -1.69081e-09, -1.68586e-09, -1.720092e-09, 
    -1.846432e-09,
  -4.608909e-09, -4.04601e-09, -3.664772e-09, -3.285472e-09, -2.787768e-09, 
    -2.430754e-09, -2.2521e-09, -2.205222e-09, -2.054815e-09, -1.867791e-09, 
    -1.723955e-09, -1.652391e-09, -1.648201e-09, -1.700448e-09, -1.996115e-09,
  -4.990315e-09, -4.435389e-09, -3.965516e-09, -3.59919e-09, -3.129867e-09, 
    -2.676814e-09, -2.410916e-09, -2.276877e-09, -2.184177e-09, 
    -2.017121e-09, -1.878053e-09, -1.791966e-09, -1.811218e-09, 
    -1.969153e-09, -2.314057e-09,
  -5.255461e-09, -4.761147e-09, -4.352251e-09, -3.90273e-09, -3.447536e-09, 
    -2.946944e-09, -2.58481e-09, -2.377696e-09, -2.301887e-09, -2.233578e-09, 
    -2.13908e-09, -2.07456e-09, -2.097405e-09, -2.289252e-09, -2.585357e-09,
  -5.718289e-09, -5.117835e-09, -4.742448e-09, -4.276355e-09, -3.753516e-09, 
    -3.22522e-09, -2.84987e-09, -2.585014e-09, -2.386511e-09, -2.273978e-09, 
    -2.191684e-09, -2.171666e-09, -2.235991e-09, -2.420783e-09, -2.6064e-09,
  -6.494055e-09, -5.615588e-09, -5.22078e-09, -4.807098e-09, -4.312138e-09, 
    -3.717214e-09, -3.263556e-09, -2.876182e-09, -2.60135e-09, -2.388131e-09, 
    -2.292611e-09, -2.24556e-09, -2.317832e-09, -2.511267e-09, -2.626896e-09,
  -7.675355e-09, -6.15979e-09, -5.558935e-09, -5.179865e-09, -4.809724e-09, 
    -4.321179e-09, -3.823976e-09, -3.386689e-09, -3.032515e-09, 
    -2.763294e-09, -2.599009e-09, -2.546047e-09, -2.619646e-09, -2.70349e-09, 
    -2.448335e-09,
  -9.002133e-09, -7.175633e-09, -5.964733e-09, -5.312053e-09, -4.888088e-09, 
    -4.488225e-09, -4.102152e-09, -3.704101e-09, -3.326939e-09, 
    -3.014177e-09, -2.836639e-09, -2.794927e-09, -2.864831e-09, 
    -2.670394e-09, -2.286044e-09,
  -1.03152e-08, -8.558557e-09, -6.959584e-09, -5.86408e-09, -5.203959e-09, 
    -4.805286e-09, -4.392688e-09, -3.993263e-09, -3.670419e-09, -3.44094e-09, 
    -3.338001e-09, -3.287061e-09, -3.101363e-09, -2.779702e-09, -2.49712e-09,
  -1.572523e-09, -1.468656e-09, -1.401124e-09, -1.352507e-09, -1.287093e-09, 
    -1.199003e-09, -1.123283e-09, -1.051401e-09, -9.913018e-10, 
    -9.578973e-10, -9.310355e-10, -9.420107e-10, -9.552594e-10, 
    -9.654046e-10, -9.683259e-10,
  -1.637149e-09, -1.505571e-09, -1.425766e-09, -1.374132e-09, -1.317446e-09, 
    -1.258614e-09, -1.208836e-09, -1.142106e-09, -1.081483e-09, 
    -1.037308e-09, -1.002947e-09, -9.898405e-10, -9.878161e-10, 
    -9.691704e-10, -9.521409e-10,
  -1.742343e-09, -1.593843e-09, -1.496189e-09, -1.417482e-09, -1.374547e-09, 
    -1.333919e-09, -1.304829e-09, -1.266406e-09, -1.240352e-09, 
    -1.207335e-09, -1.177076e-09, -1.133631e-09, -1.080428e-09, 
    -1.023164e-09, -1.0186e-09,
  -2.024143e-09, -1.840087e-09, -1.660983e-09, -1.547135e-09, -1.489925e-09, 
    -1.4533e-09, -1.428898e-09, -1.41968e-09, -1.424842e-09, -1.428675e-09, 
    -1.427039e-09, -1.418639e-09, -1.415872e-09, -1.445536e-09, -1.522301e-09,
  -2.416641e-09, -2.207227e-09, -1.944032e-09, -1.77639e-09, -1.71552e-09, 
    -1.690763e-09, -1.666094e-09, -1.661523e-09, -1.675105e-09, 
    -1.722418e-09, -1.761762e-09, -1.812977e-09, -1.902954e-09, 
    -2.046409e-09, -2.246007e-09,
  -2.742218e-09, -2.5821e-09, -2.274838e-09, -2.096428e-09, -2.040359e-09, 
    -2.033969e-09, -2.010073e-09, -1.982635e-09, -2.005256e-09, 
    -2.063028e-09, -2.163402e-09, -2.292768e-09, -2.492934e-09, -2.7219e-09, 
    -2.953901e-09,
  -2.984851e-09, -2.931834e-09, -2.719575e-09, -2.496211e-09, -2.436422e-09, 
    -2.47184e-09, -2.539934e-09, -2.585872e-09, -2.659147e-09, -2.793326e-09, 
    -2.968773e-09, -3.204777e-09, -3.458107e-09, -3.754974e-09, -4.068063e-09,
  -3.192523e-09, -3.184299e-09, -3.132569e-09, -3.060721e-09, -2.996016e-09, 
    -2.983635e-09, -3.066881e-09, -3.167899e-09, -3.315596e-09, 
    -3.532284e-09, -3.824786e-09, -4.211093e-09, -4.683743e-09, -5.12248e-09, 
    -5.437629e-09,
  -3.337377e-09, -3.284969e-09, -3.216502e-09, -3.206619e-09, -3.265555e-09, 
    -3.435507e-09, -3.728988e-09, -4.207049e-09, -4.772042e-09, 
    -5.335098e-09, -5.784563e-09, -6.147164e-09, -6.460831e-09, -6.83445e-09, 
    -7.231151e-09,
  -3.490032e-09, -3.477603e-09, -3.67461e-09, -4.013732e-09, -4.486083e-09, 
    -4.990242e-09, -5.570897e-09, -6.180579e-09, -6.773222e-09, 
    -7.254553e-09, -7.653617e-09, -8.055173e-09, -8.537802e-09, 
    -9.178055e-09, -9.85837e-09,
  -3.352732e-09, -2.440052e-09, -2.080958e-09, -1.556305e-09, -1.438337e-09, 
    -1.293451e-09, -1.100491e-09, -1.059638e-09, -1.205758e-09, 
    -1.332498e-09, -1.400472e-09, -1.412493e-09, -1.397385e-09, 
    -1.423605e-09, -1.471347e-09,
  -4.535796e-09, -3.227086e-09, -2.82115e-09, -2.237335e-09, -1.826475e-09, 
    -1.608082e-09, -1.399332e-09, -1.149107e-09, -1.058068e-09, 
    -1.158858e-09, -1.277525e-09, -1.340095e-09, -1.345082e-09, -1.31986e-09, 
    -1.328281e-09,
  -6.394998e-09, -4.67654e-09, -3.901067e-09, -3.251652e-09, -2.698177e-09, 
    -2.172561e-09, -1.929652e-09, -1.690581e-09, -1.38971e-09, -1.18995e-09, 
    -1.209567e-09, -1.319396e-09, -1.432149e-09, -1.451058e-09, -1.456873e-09,
  -8.823675e-09, -6.677257e-09, -5.357839e-09, -4.399379e-09, -3.763099e-09, 
    -3.180193e-09, -2.565524e-09, -2.205244e-09, -2.067717e-09, 
    -1.788281e-09, -1.561864e-09, -1.455201e-09, -1.505762e-09, 
    -1.543557e-09, -1.61948e-09,
  -1.212461e-08, -9.804716e-09, -7.838987e-09, -6.179691e-09, -4.979692e-09, 
    -4.280834e-09, -3.724406e-09, -3.023248e-09, -2.524439e-09, 
    -2.351356e-09, -2.202275e-09, -1.958566e-09, -1.823337e-09, 
    -1.832706e-09, -1.835251e-09,
  -1.409709e-08, -1.374143e-08, -1.171088e-08, -9.330313e-09, -7.286533e-09, 
    -5.711034e-09, -4.774332e-09, -4.172238e-09, -3.509461e-09, 
    -2.909753e-09, -2.659328e-09, -2.52653e-09, -2.271756e-09, -1.998023e-09, 
    -1.911757e-09,
  -1.407227e-08, -1.537909e-08, -1.595582e-08, -1.431649e-08, -1.185299e-08, 
    -9.30742e-09, -7.258131e-09, -5.758273e-09, -4.927323e-09, -4.185536e-09, 
    -3.439091e-09, -3.048596e-09, -2.88792e-09, -2.82781e-09, -2.651863e-09,
  -1.443523e-08, -1.475482e-08, -1.61101e-08, -1.744471e-08, -1.737724e-08, 
    -1.535584e-08, -1.265247e-08, -1.011917e-08, -8.065638e-09, 
    -6.524135e-09, -5.516512e-09, -4.551862e-09, -3.855663e-09, 
    -3.640865e-09, -3.531418e-09,
  -1.704191e-08, -1.639837e-08, -1.684991e-08, -1.782271e-08, -1.927252e-08, 
    -2.035147e-08, -1.997804e-08, -1.80042e-08, -1.542967e-08, -1.307046e-08, 
    -1.093153e-08, -9.265191e-09, -7.699581e-09, -6.337182e-09, -5.484063e-09,
  -1.834614e-08, -1.739482e-08, -1.680552e-08, -1.659558e-08, -1.721611e-08, 
    -1.815822e-08, -1.916254e-08, -1.981323e-08, -1.938612e-08, 
    -1.799145e-08, -1.598459e-08, -1.425228e-08, -1.270158e-08, -1.13631e-08, 
    -9.902152e-09,
  -3.811062e-09, -2.874116e-09, -2.604551e-09, -2.70944e-09, -3.035568e-09, 
    -3.378068e-09, -3.574715e-09, -3.684631e-09, -3.731688e-09, 
    -3.683027e-09, -3.54859e-09, -3.407838e-09, -3.303937e-09, -3.244401e-09, 
    -3.163841e-09,
  -4.959993e-09, -3.70268e-09, -2.924021e-09, -2.455572e-09, -2.567413e-09, 
    -2.889054e-09, -3.26234e-09, -3.470079e-09, -3.585681e-09, -3.630336e-09, 
    -3.569609e-09, -3.483859e-09, -3.358163e-09, -3.308867e-09, -3.293227e-09,
  -6.349731e-09, -4.924165e-09, -4.014146e-09, -3.029183e-09, -2.511457e-09, 
    -2.510737e-09, -2.763473e-09, -3.053519e-09, -3.262496e-09, 
    -3.379061e-09, -3.430251e-09, -3.422443e-09, -3.380277e-09, -3.29478e-09, 
    -3.28278e-09,
  -7.852664e-09, -6.244461e-09, -5.249984e-09, -4.068929e-09, -3.197353e-09, 
    -2.581031e-09, -2.551007e-09, -2.710872e-09, -2.960038e-09, 
    -3.103339e-09, -3.190734e-09, -3.200822e-09, -3.231605e-09, 
    -3.238647e-09, -3.231188e-09,
  -9.991044e-09, -7.78101e-09, -6.673815e-09, -5.338312e-09, -4.199398e-09, 
    -3.350545e-09, -2.672111e-09, -2.509301e-09, -2.660683e-09, -2.87728e-09, 
    -2.991443e-09, -3.056908e-09, -3.057485e-09, -3.084054e-09, -3.150582e-09,
  -1.23981e-08, -9.859995e-09, -8.237017e-09, -6.987772e-09, -5.667404e-09, 
    -4.470079e-09, -3.554969e-09, -2.860507e-09, -2.509329e-09, -2.58985e-09, 
    -2.77753e-09, -2.914036e-09, -2.961914e-09, -2.995541e-09, -3.062868e-09,
  -1.464269e-08, -1.236084e-08, -1.028316e-08, -8.583789e-09, -7.322155e-09, 
    -6.060166e-09, -4.881762e-09, -3.843295e-09, -3.166846e-09, 
    -2.708789e-09, -2.557641e-09, -2.680365e-09, -2.783219e-09, 
    -2.835232e-09, -2.870674e-09,
  -1.626225e-08, -1.474722e-08, -1.272852e-08, -1.072104e-08, -9.10389e-09, 
    -7.66045e-09, -6.500582e-09, -5.38404e-09, -4.29577e-09, -3.596519e-09, 
    -3.067408e-09, -2.774998e-09, -2.765742e-09, -2.819927e-09, -2.897821e-09,
  -1.704909e-08, -1.649688e-08, -1.516474e-08, -1.310841e-08, -1.129901e-08, 
    -9.591194e-09, -8.115657e-09, -6.916304e-09, -5.99536e-09, -4.929589e-09, 
    -4.19311e-09, -3.611087e-09, -3.219247e-09, -3.052544e-09, -3.059641e-09,
  -1.7854e-08, -1.723526e-08, -1.687489e-08, -1.553044e-08, -1.370506e-08, 
    -1.18481e-08, -1.024284e-08, -8.671998e-09, -7.471157e-09, -6.629507e-09, 
    -5.752231e-09, -4.931763e-09, -4.341735e-09, -3.955518e-09, -3.74793e-09,
  -3.536382e-09, -2.721479e-09, -2.211973e-09, -1.80193e-09, -1.46586e-09, 
    -1.07986e-09, -8.806096e-10, -7.577272e-10, -7.722983e-10, -7.64895e-10, 
    -6.826344e-10, -6.025641e-10, -6.416614e-10, -6.4985e-10, -6.499162e-10,
  -4.465001e-09, -3.302168e-09, -2.691071e-09, -2.154436e-09, -1.844089e-09, 
    -1.511784e-09, -1.163507e-09, -8.48318e-10, -5.82159e-10, -4.774863e-10, 
    -4.138621e-10, -4.339137e-10, -4.588521e-10, -5.547058e-10, -6.787678e-10,
  -5.393389e-09, -4.000834e-09, -3.155656e-09, -2.473008e-09, -2.090325e-09, 
    -1.830187e-09, -1.61909e-09, -1.342672e-09, -1.03581e-09, -7.547375e-10, 
    -5.762272e-10, -5.231803e-10, -5.408824e-10, -6.611651e-10, -7.987174e-10,
  -6.334924e-09, -4.95241e-09, -3.821941e-09, -3.03313e-09, -2.412445e-09, 
    -2.052387e-09, -1.849051e-09, -1.702027e-09, -1.544357e-09, 
    -1.355504e-09, -1.153452e-09, -9.619435e-10, -9.638833e-10, 
    -9.517575e-10, -1.049796e-09,
  -7.24262e-09, -5.978607e-09, -4.612318e-09, -3.614575e-09, -2.937038e-09, 
    -2.375945e-09, -2.059273e-09, -1.870502e-09, -1.778715e-09, 
    -1.665179e-09, -1.570215e-09, -1.449453e-09, -1.403815e-09, -1.34549e-09, 
    -1.433674e-09,
  -8.171997e-09, -6.980679e-09, -5.762649e-09, -4.286635e-09, -3.52849e-09, 
    -2.881547e-09, -2.373402e-09, -2.072871e-09, -1.912562e-09, 
    -1.862013e-09, -1.829842e-09, -1.827206e-09, -1.767887e-09, 
    -1.763138e-09, -1.763131e-09,
  -8.80048e-09, -7.705303e-09, -6.854151e-09, -5.359619e-09, -4.136086e-09, 
    -3.508432e-09, -2.918025e-09, -2.437828e-09, -2.135722e-09, 
    -1.953789e-09, -1.866801e-09, -1.841164e-09, -1.836009e-09, -1.84113e-09, 
    -1.820842e-09,
  -9.615051e-09, -8.357891e-09, -7.611986e-09, -6.587913e-09, -5.077143e-09, 
    -4.089085e-09, -3.537527e-09, -2.967032e-09, -2.497217e-09, 
    -2.217639e-09, -2.001014e-09, -1.921274e-09, -1.895374e-09, 
    -1.905165e-09, -1.894303e-09,
  -1.039065e-08, -9.162447e-09, -8.226593e-09, -7.467048e-09, -6.362187e-09, 
    -4.987137e-09, -4.214134e-09, -3.656762e-09, -3.112377e-09, -2.66253e-09, 
    -2.38047e-09, -2.193516e-09, -2.112762e-09, -2.072198e-09, -2.103217e-09,
  -1.116357e-08, -9.878813e-09, -8.894148e-09, -8.06472e-09, -7.340192e-09, 
    -6.171194e-09, -5.071083e-09, -4.394628e-09, -3.880761e-09, 
    -3.404187e-09, -2.999012e-09, -2.751218e-09, -2.571046e-09, 
    -2.515488e-09, -2.596298e-09,
  -1.052776e-09, -9.2175e-10, -8.938573e-10, -9.603834e-10, -1.144611e-09, 
    -1.357988e-09, -1.595294e-09, -1.856538e-09, -2.185339e-09, 
    -2.469856e-09, -2.798157e-09, -3.0828e-09, -3.382896e-09, -3.660082e-09, 
    -4.065216e-09,
  -1.260165e-09, -1.119055e-09, -1.107924e-09, -1.119114e-09, -1.279676e-09, 
    -1.47286e-09, -1.735498e-09, -2.013092e-09, -2.299735e-09, -2.571421e-09, 
    -2.898283e-09, -3.199285e-09, -3.524528e-09, -3.835995e-09, -4.277843e-09,
  -1.486296e-09, -1.255853e-09, -1.250711e-09, -1.293327e-09, -1.40317e-09, 
    -1.59479e-09, -1.837627e-09, -2.119447e-09, -2.404497e-09, -2.687866e-09, 
    -3.010598e-09, -3.304847e-09, -3.647906e-09, -4.010391e-09, -4.476888e-09,
  -1.748271e-09, -1.454691e-09, -1.408605e-09, -1.448657e-09, -1.546813e-09, 
    -1.741713e-09, -1.971814e-09, -2.233484e-09, -2.520037e-09, 
    -2.803102e-09, -3.09931e-09, -3.417726e-09, -3.81582e-09, -4.211611e-09, 
    -4.713802e-09,
  -2.001137e-09, -1.682082e-09, -1.604437e-09, -1.618089e-09, -1.695688e-09, 
    -1.869038e-09, -2.112144e-09, -2.359772e-09, -2.616988e-09, 
    -2.915606e-09, -3.208326e-09, -3.56037e-09, -3.99399e-09, -4.439465e-09, 
    -4.994771e-09,
  -2.318764e-09, -1.880514e-09, -1.78011e-09, -1.770468e-09, -1.832115e-09, 
    -1.983328e-09, -2.229297e-09, -2.482983e-09, -2.734601e-09, 
    -3.028787e-09, -3.302607e-09, -3.679934e-09, -4.152201e-09, 
    -4.655465e-09, -5.336198e-09,
  -2.579658e-09, -2.15991e-09, -1.971639e-09, -1.934208e-09, -1.97504e-09, 
    -2.117229e-09, -2.333885e-09, -2.597888e-09, -2.845359e-09, 
    -3.125986e-09, -3.443594e-09, -3.80388e-09, -4.31198e-09, -4.905235e-09, 
    -5.68591e-09,
  -2.842811e-09, -2.403548e-09, -2.204922e-09, -2.084983e-09, -2.112087e-09, 
    -2.217489e-09, -2.423583e-09, -2.698745e-09, -2.963521e-09, 
    -3.241777e-09, -3.557678e-09, -3.920095e-09, -4.516246e-09, -5.20935e-09, 
    -6.033173e-09,
  -3.117237e-09, -2.617172e-09, -2.398369e-09, -2.298957e-09, -2.277913e-09, 
    -2.30713e-09, -2.471858e-09, -2.729019e-09, -3.050264e-09, -3.303536e-09, 
    -3.619152e-09, -4.066806e-09, -4.725785e-09, -5.502818e-09, -6.352105e-09,
  -3.484478e-09, -2.841565e-09, -2.557518e-09, -2.453932e-09, -2.444691e-09, 
    -2.480869e-09, -2.59728e-09, -2.839118e-09, -3.146626e-09, -3.423194e-09, 
    -3.745229e-09, -4.263986e-09, -4.944481e-09, -5.754236e-09, -6.645523e-09,
  -3.22008e-09, -3.247591e-09, -3.202727e-09, -3.079678e-09, -3.074819e-09, 
    -3.007962e-09, -3.093696e-09, -3.168815e-09, -3.274748e-09, 
    -3.360458e-09, -3.5067e-09, -3.769711e-09, -4.488108e-09, -5.394646e-09, 
    -6.501728e-09,
  -3.234041e-09, -3.22236e-09, -3.17458e-09, -3.061505e-09, -2.984091e-09, 
    -2.955558e-09, -3.110934e-09, -3.236355e-09, -3.395034e-09, 
    -3.420489e-09, -3.591949e-09, -3.924051e-09, -4.801455e-09, 
    -5.793593e-09, -6.941239e-09,
  -3.353459e-09, -3.293642e-09, -3.212101e-09, -3.080539e-09, -2.984334e-09, 
    -3.004303e-09, -3.208734e-09, -3.343122e-09, -3.486661e-09, 
    -3.486609e-09, -3.689732e-09, -4.211262e-09, -5.260241e-09, 
    -6.274834e-09, -7.504598e-09,
  -3.429297e-09, -3.373606e-09, -3.258225e-09, -3.099537e-09, -2.999853e-09, 
    -3.069222e-09, -3.309458e-09, -3.453528e-09, -3.525944e-09, 
    -3.509635e-09, -3.795841e-09, -4.584954e-09, -5.72019e-09, -6.729955e-09, 
    -8.129169e-09,
  -3.47809e-09, -3.429591e-09, -3.298489e-09, -3.129157e-09, -3.031687e-09, 
    -3.154053e-09, -3.366205e-09, -3.529682e-09, -3.600487e-09, 
    -3.607681e-09, -4.056049e-09, -5.026114e-09, -6.159158e-09, 
    -7.133942e-09, -8.82983e-09,
  -3.590343e-09, -3.515997e-09, -3.396595e-09, -3.193102e-09, -3.111804e-09, 
    -3.2419e-09, -3.470557e-09, -3.636404e-09, -3.648917e-09, -3.758092e-09, 
    -4.438876e-09, -5.497228e-09, -6.635571e-09, -7.757348e-09, -9.731143e-09,
  -3.66988e-09, -3.614417e-09, -3.52274e-09, -3.311296e-09, -3.234006e-09, 
    -3.394573e-09, -3.613069e-09, -3.676587e-09, -3.746324e-09, 
    -4.020584e-09, -4.846472e-09, -6.002962e-09, -7.137228e-09, 
    -8.512639e-09, -1.076082e-08,
  -3.744297e-09, -3.724055e-09, -3.669588e-09, -3.473444e-09, -3.387237e-09, 
    -3.530145e-09, -3.700817e-09, -3.76513e-09, -3.920777e-09, -4.360068e-09, 
    -5.308938e-09, -6.535468e-09, -7.76879e-09, -9.552907e-09, -1.179508e-08,
  -3.825691e-09, -3.843259e-09, -3.833754e-09, -3.61284e-09, -3.523364e-09, 
    -3.711938e-09, -3.877225e-09, -3.889236e-09, -4.085494e-09, -4.77839e-09, 
    -5.841963e-09, -7.114872e-09, -8.604315e-09, -1.064063e-08, -1.265409e-08,
  -3.886266e-09, -3.950422e-09, -3.987609e-09, -3.730687e-09, -3.658767e-09, 
    -3.843385e-09, -3.99902e-09, -4.031736e-09, -4.439685e-09, -5.30473e-09, 
    -6.441092e-09, -7.814313e-09, -9.504805e-09, -1.160814e-08, -1.343751e-08,
  -3.001123e-09, -2.634239e-09, -2.616027e-09, -2.910176e-09, -3.102912e-09, 
    -3.250554e-09, -3.582531e-09, -4.040185e-09, -4.760354e-09, 
    -5.578044e-09, -6.287546e-09, -6.940597e-09, -7.994214e-09, 
    -9.302838e-09, -1.096559e-08,
  -3.136247e-09, -2.792837e-09, -2.63916e-09, -2.849938e-09, -3.058755e-09, 
    -3.21893e-09, -3.590916e-09, -4.141538e-09, -4.92035e-09, -5.706107e-09, 
    -6.356883e-09, -7.017538e-09, -8.03079e-09, -9.289818e-09, -1.096859e-08,
  -3.212334e-09, -2.951908e-09, -2.716285e-09, -2.845655e-09, -3.045181e-09, 
    -3.215677e-09, -3.633248e-09, -4.279687e-09, -5.06642e-09, -5.819582e-09, 
    -6.434802e-09, -7.078425e-09, -8.033903e-09, -9.327295e-09, -1.110013e-08,
  -3.273347e-09, -3.10997e-09, -2.836993e-09, -2.909637e-09, -3.038482e-09, 
    -3.26064e-09, -3.683917e-09, -4.42487e-09, -5.215247e-09, -5.927888e-09, 
    -6.542302e-09, -7.200566e-09, -8.107731e-09, -9.383878e-09, -1.121353e-08,
  -3.254889e-09, -3.233388e-09, -2.958325e-09, -2.963744e-09, -3.116176e-09, 
    -3.351013e-09, -3.786051e-09, -4.554154e-09, -5.346222e-09, 
    -6.029163e-09, -6.688188e-09, -7.317572e-09, -8.270366e-09, 
    -9.577549e-09, -1.135455e-08,
  -3.268557e-09, -3.31369e-09, -3.104004e-09, -3.081529e-09, -3.235101e-09, 
    -3.450527e-09, -3.921942e-09, -4.704846e-09, -5.479098e-09, -6.16882e-09, 
    -6.839971e-09, -7.386626e-09, -8.422214e-09, -9.776204e-09, -1.155984e-08,
  -3.293064e-09, -3.346808e-09, -3.259777e-09, -3.237623e-09, -3.441498e-09, 
    -3.690795e-09, -4.176322e-09, -4.828263e-09, -5.585016e-09, 
    -6.346825e-09, -6.914251e-09, -7.438441e-09, -8.647832e-09, 
    -1.009746e-08, -1.184608e-08,
  -3.36611e-09, -3.462271e-09, -3.462335e-09, -3.474737e-09, -3.739372e-09, 
    -3.986612e-09, -4.402876e-09, -4.969029e-09, -5.788446e-09, 
    -6.523176e-09, -6.985318e-09, -7.565926e-09, -8.950396e-09, 
    -1.044593e-08, -1.224531e-08,
  -3.447231e-09, -3.584062e-09, -3.650925e-09, -3.757612e-09, -4.079087e-09, 
    -4.268498e-09, -4.626653e-09, -5.154586e-09, -5.953573e-09, 
    -6.617717e-09, -7.047854e-09, -7.798167e-09, -9.345649e-09, 
    -1.082298e-08, -1.264008e-08,
  -3.574608e-09, -3.75657e-09, -3.924706e-09, -4.149943e-09, -4.412209e-09, 
    -4.535412e-09, -4.830203e-09, -5.34688e-09, -6.102705e-09, -6.700225e-09, 
    -7.193522e-09, -8.224827e-09, -9.76617e-09, -1.121633e-08, -1.300876e-08,
  -3.981751e-09, -4.023365e-09, -3.889042e-09, -3.528121e-09, -3.125857e-09, 
    -2.757889e-09, -2.615625e-09, -2.681134e-09, -2.784694e-09, 
    -3.160728e-09, -4.126757e-09, -5.32203e-09, -7.010264e-09, -9.720301e-09, 
    -1.346419e-08,
  -3.831026e-09, -4.061526e-09, -4.018555e-09, -3.737133e-09, -3.370991e-09, 
    -3.00118e-09, -2.814499e-09, -2.858255e-09, -2.954877e-09, -3.296743e-09, 
    -4.14918e-09, -5.353141e-09, -7.170024e-09, -9.875842e-09, -1.373047e-08,
  -3.794837e-09, -4.03749e-09, -4.082921e-09, -3.908655e-09, -3.574018e-09, 
    -3.226342e-09, -3.046636e-09, -3.079981e-09, -3.148887e-09, -3.46999e-09, 
    -4.219406e-09, -5.393745e-09, -7.2512e-09, -9.948158e-09, -1.385068e-08,
  -3.699723e-09, -4.005486e-09, -4.116476e-09, -4.043443e-09, -3.753779e-09, 
    -3.44048e-09, -3.280201e-09, -3.26599e-09, -3.312578e-09, -3.646829e-09, 
    -4.328407e-09, -5.429982e-09, -7.330139e-09, -1.0001e-08, -1.389422e-08,
  -3.371488e-09, -3.989758e-09, -4.110488e-09, -4.127941e-09, -3.89935e-09, 
    -3.617489e-09, -3.482608e-09, -3.443501e-09, -3.520253e-09, 
    -3.786777e-09, -4.418761e-09, -5.468789e-09, -7.366455e-09, 
    -1.000057e-08, -1.386664e-08,
  -3.016208e-09, -3.859895e-09, -4.156382e-09, -4.183607e-09, -4.026514e-09, 
    -3.773789e-09, -3.66332e-09, -3.621999e-09, -3.68479e-09, -3.921148e-09, 
    -4.551029e-09, -5.52667e-09, -7.406386e-09, -9.997237e-09, -1.38257e-08,
  -2.9703e-09, -3.598467e-09, -4.147564e-09, -4.266671e-09, -4.133756e-09, 
    -3.887595e-09, -3.838017e-09, -3.82618e-09, -3.868659e-09, -4.091387e-09, 
    -4.683168e-09, -5.61537e-09, -7.489202e-09, -1.000085e-08, -1.369774e-08,
  -3.041898e-09, -3.268964e-09, -4.079141e-09, -4.370527e-09, -4.219995e-09, 
    -3.997863e-09, -4.005174e-09, -4.012992e-09, -4.065408e-09, 
    -4.283007e-09, -4.829727e-09, -5.744311e-09, -7.565576e-09, 
    -1.000901e-08, -1.374069e-08,
  -3.145241e-09, -3.078252e-09, -3.933617e-09, -4.47197e-09, -4.325711e-09, 
    -4.115623e-09, -4.148541e-09, -4.19409e-09, -4.265329e-09, -4.456192e-09, 
    -4.975851e-09, -5.886971e-09, -7.633051e-09, -1.000624e-08, -1.368282e-08,
  -3.180404e-09, -3.00283e-09, -3.823129e-09, -4.544681e-09, -4.434728e-09, 
    -4.251645e-09, -4.302148e-09, -4.372189e-09, -4.467101e-09, 
    -4.640209e-09, -5.135643e-09, -6.007383e-09, -7.679144e-09, 
    -9.992381e-09, -1.360629e-08,
  -2.656837e-09, -2.565134e-09, -2.580114e-09, -2.680766e-09, -2.975062e-09, 
    -3.53267e-09, -4.539662e-09, -5.935004e-09, -7.653523e-09, -9.837504e-09, 
    -1.220375e-08, -1.501445e-08, -1.827961e-08, -2.155292e-08, -2.426171e-08,
  -2.578637e-09, -2.504771e-09, -2.539471e-09, -2.604968e-09, -2.853427e-09, 
    -3.394884e-09, -4.392868e-09, -5.740215e-09, -7.46879e-09, -9.76101e-09, 
    -1.229187e-08, -1.545328e-08, -1.876388e-08, -2.192641e-08, -2.453014e-08,
  -2.53781e-09, -2.451144e-09, -2.477807e-09, -2.525026e-09, -2.74886e-09, 
    -3.286816e-09, -4.271237e-09, -5.633265e-09, -7.380119e-09, 
    -9.673008e-09, -1.241103e-08, -1.581628e-08, -1.920419e-08, 
    -2.229488e-08, -2.483144e-08,
  -2.611177e-09, -2.382539e-09, -2.405323e-09, -2.445014e-09, -2.67673e-09, 
    -3.176361e-09, -4.152307e-09, -5.502474e-09, -7.23294e-09, -9.566955e-09, 
    -1.247255e-08, -1.601191e-08, -1.947296e-08, -2.266126e-08, -2.537143e-08,
  -2.758923e-09, -2.402057e-09, -2.318528e-09, -2.351349e-09, -2.594182e-09, 
    -3.077262e-09, -4.033964e-09, -5.418158e-09, -7.118436e-09, 
    -9.478789e-09, -1.244075e-08, -1.602953e-08, -1.968483e-08, 
    -2.323343e-08, -2.632062e-08,
  -2.855382e-09, -2.540603e-09, -2.24561e-09, -2.288902e-09, -2.480696e-09, 
    -2.954214e-09, -3.921303e-09, -5.315082e-09, -7.041623e-09, 
    -9.362053e-09, -1.229683e-08, -1.60053e-08, -2.005883e-08, -2.401884e-08, 
    -2.717413e-08,
  -2.862481e-09, -2.729674e-09, -2.252376e-09, -2.229217e-09, -2.362915e-09, 
    -2.848471e-09, -3.805411e-09, -5.264162e-09, -6.950532e-09, 
    -9.195485e-09, -1.204418e-08, -1.596278e-08, -2.040193e-08, 
    -2.456103e-08, -2.780096e-08,
  -2.862718e-09, -2.909699e-09, -2.344637e-09, -2.178373e-09, -2.287739e-09, 
    -2.72144e-09, -3.69583e-09, -5.173408e-09, -6.866998e-09, -8.933701e-09, 
    -1.173548e-08, -1.587787e-08, -2.056112e-08, -2.498389e-08, -2.854303e-08,
  -3.025711e-09, -3.000213e-09, -2.502308e-09, -2.17105e-09, -2.226347e-09, 
    -2.61366e-09, -3.555706e-09, -5.006923e-09, -6.558605e-09, -8.583781e-09, 
    -1.134707e-08, -1.567616e-08, -2.052277e-08, -2.525971e-08, -2.898858e-08,
  -3.168013e-09, -2.970816e-09, -2.65628e-09, -2.193968e-09, -2.174342e-09, 
    -2.531894e-09, -3.384203e-09, -4.718279e-09, -6.220825e-09, 
    -8.191492e-09, -1.090688e-08, -1.537123e-08, -2.042152e-08, 
    -2.543712e-08, -2.899761e-08,
  -4.477906e-09, -5.581443e-09, -6.451149e-09, -7.131979e-09, -7.917849e-09, 
    -9.405699e-09, -1.153825e-08, -1.389528e-08, -1.599352e-08, 
    -1.723285e-08, -1.767775e-08, -1.824959e-08, -1.820088e-08, 
    -1.810274e-08, -1.752966e-08,
  -4.855728e-09, -5.998895e-09, -6.847271e-09, -7.57586e-09, -8.550471e-09, 
    -1.019342e-08, -1.255497e-08, -1.4863e-08, -1.661637e-08, -1.740049e-08, 
    -1.781084e-08, -1.80791e-08, -1.768285e-08, -1.778436e-08, -1.848805e-08,
  -5.296297e-09, -6.43999e-09, -7.258928e-09, -8.114507e-09, -9.174123e-09, 
    -1.107378e-08, -1.357933e-08, -1.587552e-08, -1.722168e-08, 
    -1.779336e-08, -1.797683e-08, -1.772483e-08, -1.765612e-08, 
    -1.836472e-08, -2.257433e-08,
  -5.672898e-09, -6.806953e-09, -7.635038e-09, -8.604958e-09, -9.773943e-09, 
    -1.215944e-08, -1.468601e-08, -1.666397e-08, -1.76126e-08, -1.78843e-08, 
    -1.785068e-08, -1.739056e-08, -1.81633e-08, -2.21731e-08, -2.84517e-08,
  -5.941873e-09, -7.082811e-09, -7.957307e-09, -9.061005e-09, -1.059992e-08, 
    -1.336268e-08, -1.556087e-08, -1.715305e-08, -1.77889e-08, -1.803525e-08, 
    -1.744213e-08, -1.788983e-08, -2.230124e-08, -2.829481e-08, -3.156928e-08,
  -6.232325e-09, -7.250937e-09, -8.334584e-09, -9.50382e-09, -1.190368e-08, 
    -1.45518e-08, -1.632252e-08, -1.745247e-08, -1.795005e-08, -1.773192e-08, 
    -1.801034e-08, -2.204341e-08, -2.808436e-08, -3.161473e-08, -2.981043e-08,
  -6.540033e-09, -7.431853e-09, -8.685661e-09, -1.030126e-08, -1.311662e-08, 
    -1.545202e-08, -1.663508e-08, -1.768708e-08, -1.772034e-08, 
    -1.826825e-08, -2.130471e-08, -2.749436e-08, -3.14491e-08, -3.01234e-08, 
    -2.961855e-08,
  -6.754923e-09, -7.526021e-09, -9.113005e-09, -1.120088e-08, -1.420151e-08, 
    -1.59232e-08, -1.699732e-08, -1.748743e-08, -1.816328e-08, -2.090434e-08, 
    -2.736304e-08, -3.112508e-08, -3.067402e-08, -3.026021e-08, -3.009196e-08,
  -6.745025e-09, -7.805419e-09, -9.482043e-09, -1.208122e-08, -1.506874e-08, 
    -1.61855e-08, -1.694213e-08, -1.778255e-08, -2.043114e-08, -2.635468e-08, 
    -3.003383e-08, -3.090201e-08, -3.018645e-08, -3.066168e-08, -2.997119e-08,
  -6.765246e-09, -7.956042e-09, -9.765524e-09, -1.309229e-08, -1.520276e-08, 
    -1.618917e-08, -1.707407e-08, -1.965805e-08, -2.474759e-08, 
    -2.879411e-08, -3.027097e-08, -3.005849e-08, -3.050827e-08, 
    -2.995814e-08, -2.953371e-08,
  -2.856541e-09, -2.97649e-09, -4.483464e-09, -6.045551e-09, -7.009208e-09, 
    -7.377806e-09, -8.251724e-09, -9.998464e-09, -1.205198e-08, 
    -1.457405e-08, -1.670475e-08, -1.894454e-08, -2.028183e-08, 
    -2.154117e-08, -2.242215e-08,
  -3.252153e-09, -3.251576e-09, -4.675418e-09, -5.96821e-09, -7.202769e-09, 
    -7.922988e-09, -8.86453e-09, -1.064645e-08, -1.272963e-08, -1.560797e-08, 
    -1.780011e-08, -1.95069e-08, -2.048672e-08, -2.187577e-08, -2.228778e-08,
  -3.524878e-09, -3.948624e-09, -5.000973e-09, -5.871782e-09, -7.420147e-09, 
    -8.603894e-09, -9.685799e-09, -1.142708e-08, -1.369041e-08, 
    -1.680747e-08, -1.853793e-08, -1.994709e-08, -2.080238e-08, 
    -2.179049e-08, -2.171821e-08,
  -4.354133e-09, -4.919311e-09, -5.088442e-09, -6.007825e-09, -7.927524e-09, 
    -9.780363e-09, -1.074964e-08, -1.258439e-08, -1.492497e-08, 
    -1.778679e-08, -1.924401e-08, -2.045318e-08, -2.070269e-08, 
    -2.134985e-08, -2.1017e-08,
  -4.883829e-09, -5.144946e-09, -5.692503e-09, -6.526288e-09, -8.908002e-09, 
    -1.102072e-08, -1.204156e-08, -1.38268e-08, -1.619403e-08, -1.874994e-08, 
    -2.004459e-08, -2.043747e-08, -2.045242e-08, -2.106276e-08, -2.092919e-08,
  -5.261363e-09, -5.671894e-09, -6.685597e-09, -7.690937e-09, -1.019026e-08, 
    -1.241233e-08, -1.323656e-08, -1.522288e-08, -1.773397e-08, 
    -1.971724e-08, -2.029296e-08, -2.036781e-08, -2.020354e-08, 
    -2.090847e-08, -2.135095e-08,
  -6.170248e-09, -7.084028e-09, -8.037411e-09, -9.161036e-09, -1.188517e-08, 
    -1.360517e-08, -1.476161e-08, -1.70655e-08, -1.922223e-08, -1.974252e-08, 
    -1.995475e-08, -1.976574e-08, -2.078827e-08, -2.268881e-08, -2.30043e-08,
  -7.838952e-09, -8.463029e-09, -9.384172e-09, -1.110176e-08, -1.351421e-08, 
    -1.509685e-08, -1.636728e-08, -1.823449e-08, -1.880805e-08, 
    -1.906852e-08, -1.966578e-08, -2.181057e-08, -2.333873e-08, 
    -2.428485e-08, -2.45405e-08,
  -9.294333e-09, -9.912516e-09, -1.111134e-08, -1.311451e-08, -1.54385e-08, 
    -1.663511e-08, -1.781643e-08, -1.852857e-08, -1.900287e-08, 
    -2.023758e-08, -2.27249e-08, -2.404459e-08, -2.522171e-08, -2.567796e-08, 
    -2.459932e-08,
  -1.062613e-08, -1.162136e-08, -1.324793e-08, -1.589206e-08, -1.73116e-08, 
    -1.80263e-08, -1.864334e-08, -1.928463e-08, -2.056395e-08, -2.31566e-08, 
    -2.485985e-08, -2.622282e-08, -2.632963e-08, -2.50124e-08, -2.316312e-08,
  -7.319038e-09, -8.571595e-09, -1.031632e-08, -1.101711e-08, -1.209561e-08, 
    -1.378477e-08, -1.396253e-08, -1.56832e-08, -1.733241e-08, -1.44502e-08, 
    -1.427366e-08, -1.58875e-08, -1.74419e-08, -1.798308e-08, -1.693677e-08,
  -6.620373e-09, -7.995887e-09, -1.017594e-08, -1.143015e-08, -1.21843e-08, 
    -1.348232e-08, -1.370259e-08, -1.494052e-08, -1.611596e-08, 
    -1.484648e-08, -1.564011e-08, -1.602743e-08, -1.717213e-08, 
    -1.764233e-08, -1.666157e-08,
  -5.380745e-09, -6.133268e-09, -8.762912e-09, -1.075445e-08, -1.256801e-08, 
    -1.298104e-08, -1.269502e-08, -1.493243e-08, -1.67456e-08, -1.541438e-08, 
    -1.60609e-08, -1.578136e-08, -1.670743e-08, -1.731325e-08, -1.680272e-08,
  -3.892973e-09, -4.403393e-09, -6.725425e-09, -9.916894e-09, -1.248399e-08, 
    -1.175491e-08, -1.19337e-08, -1.449986e-08, -1.663676e-08, -1.553812e-08, 
    -1.607483e-08, -1.571606e-08, -1.652562e-08, -1.683847e-08, -1.770229e-08,
  -3.652503e-09, -5.12121e-09, -8.281509e-09, -1.035288e-08, -1.154641e-08, 
    -1.0644e-08, -1.161354e-08, -1.439738e-08, -1.679535e-08, -1.544671e-08, 
    -1.571357e-08, -1.58407e-08, -1.619348e-08, -1.703668e-08, -1.797913e-08,
  -5.138452e-09, -7.479454e-09, -1.015681e-08, -1.048125e-08, -1.059354e-08, 
    -9.733515e-09, -1.182594e-08, -1.535915e-08, -1.611643e-08, 
    -1.571482e-08, -1.584524e-08, -1.65753e-08, -1.723747e-08, -1.744649e-08, 
    -1.859915e-08,
  -6.783662e-09, -8.33287e-09, -9.518772e-09, -1.009326e-08, -9.713836e-09, 
    -9.531895e-09, -1.294882e-08, -1.627204e-08, -1.618324e-08, 
    -1.633928e-08, -1.701069e-08, -1.845994e-08, -1.835119e-08, 
    -1.850501e-08, -1.889082e-08,
  -7.09826e-09, -7.735664e-09, -8.773789e-09, -9.366286e-09, -9.334068e-09, 
    -1.084433e-08, -1.503006e-08, -1.657479e-08, -1.723643e-08, 
    -1.787067e-08, -1.909972e-08, -1.953426e-08, -1.898731e-08, 
    -1.850074e-08, -1.82898e-08,
  -7.007549e-09, -7.699755e-09, -8.689683e-09, -9.210217e-09, -1.071806e-08, 
    -1.377698e-08, -1.649383e-08, -1.687132e-08, -1.856696e-08, 
    -1.937488e-08, -1.994315e-08, -1.950326e-08, -1.86365e-08, -1.832189e-08, 
    -1.84363e-08,
  -7.022049e-09, -7.791933e-09, -9.47656e-09, -1.100281e-08, -1.32016e-08, 
    -1.60109e-08, -1.719667e-08, -1.791209e-08, -1.960021e-08, -2.019972e-08, 
    -1.999512e-08, -1.918723e-08, -1.889914e-08, -1.891773e-08, -1.914298e-08,
  -8.764173e-09, -9.105264e-09, -9.327669e-09, -9.862588e-09, -1.056803e-08, 
    -1.160412e-08, -1.306852e-08, -1.502969e-08, -1.673068e-08, 
    -1.858498e-08, -2.077354e-08, -2.212705e-08, -2.310037e-08, 
    -2.394929e-08, -2.393602e-08,
  -9.355545e-09, -9.753975e-09, -1.009216e-08, -1.075451e-08, -1.145025e-08, 
    -1.249853e-08, -1.398154e-08, -1.575734e-08, -1.746828e-08, 
    -1.934866e-08, -2.105737e-08, -2.264978e-08, -2.369309e-08, 
    -2.393926e-08, -2.350734e-08,
  -9.953944e-09, -1.03084e-08, -1.101122e-08, -1.155642e-08, -1.237657e-08, 
    -1.343053e-08, -1.482271e-08, -1.634852e-08, -1.783467e-08, -1.96977e-08, 
    -2.109546e-08, -2.249336e-08, -2.383224e-08, -2.332808e-08, -2.25686e-08,
  -1.083964e-08, -1.10716e-08, -1.189984e-08, -1.260456e-08, -1.319491e-08, 
    -1.409386e-08, -1.540423e-08, -1.70974e-08, -1.811668e-08, -1.944568e-08, 
    -2.072907e-08, -2.218328e-08, -2.360719e-08, -2.276522e-08, -2.149057e-08,
  -1.131231e-08, -1.159573e-08, -1.232356e-08, -1.294947e-08, -1.405967e-08, 
    -1.484129e-08, -1.613924e-08, -1.775705e-08, -1.839039e-08, 
    -1.907363e-08, -1.997032e-08, -2.170522e-08, -2.287985e-08, 
    -2.133705e-08, -2.060154e-08,
  -1.117179e-08, -1.212159e-08, -1.278048e-08, -1.346747e-08, -1.537834e-08, 
    -1.539835e-08, -1.624915e-08, -1.759541e-08, -1.845728e-08, -1.8807e-08, 
    -1.975762e-08, -2.157562e-08, -2.204803e-08, -1.970156e-08, -2.020601e-08,
  -1.163386e-08, -1.285284e-08, -1.323719e-08, -1.426362e-08, -1.572979e-08, 
    -1.561072e-08, -1.628384e-08, -1.762359e-08, -1.851258e-08, -1.85634e-08, 
    -1.930382e-08, -2.126876e-08, -2.058162e-08, -1.837027e-08, -1.979682e-08,
  -1.235725e-08, -1.326577e-08, -1.429589e-08, -1.502272e-08, -1.558136e-08, 
    -1.509602e-08, -1.577359e-08, -1.735812e-08, -1.813183e-08, 
    -1.825789e-08, -1.885739e-08, -2.041912e-08, -1.865834e-08, 
    -1.808448e-08, -1.966113e-08,
  -1.289835e-08, -1.406305e-08, -1.512424e-08, -1.46459e-08, -1.48086e-08, 
    -1.48554e-08, -1.601239e-08, -1.692626e-08, -1.745672e-08, -1.728243e-08, 
    -1.874182e-08, -1.933535e-08, -1.72795e-08, -1.814311e-08, -1.975855e-08,
  -1.388736e-08, -1.454514e-08, -1.447072e-08, -1.361674e-08, -1.392335e-08, 
    -1.509996e-08, -1.641446e-08, -1.613415e-08, -1.727003e-08, 
    -1.700382e-08, -1.879114e-08, -1.749615e-08, -1.706679e-08, 
    -1.816989e-08, -1.946506e-08,
  -1.574421e-08, -1.752429e-08, -1.836712e-08, -1.903138e-08, -1.934684e-08, 
    -1.994784e-08, -2.077287e-08, -2.161778e-08, -2.235194e-08, 
    -2.243669e-08, -2.264277e-08, -2.279871e-08, -2.275597e-08, 
    -2.290583e-08, -2.292141e-08,
  -1.563838e-08, -1.714828e-08, -1.766763e-08, -1.813218e-08, -1.848124e-08, 
    -1.931441e-08, -2.035528e-08, -2.137833e-08, -2.185744e-08, 
    -2.214481e-08, -2.256597e-08, -2.271395e-08, -2.308899e-08, -2.32603e-08, 
    -2.354059e-08,
  -1.542648e-08, -1.666185e-08, -1.706086e-08, -1.754651e-08, -1.803211e-08, 
    -1.899274e-08, -2.026507e-08, -2.122673e-08, -2.155788e-08, 
    -2.206212e-08, -2.232404e-08, -2.237747e-08, -2.274064e-08, 
    -2.293241e-08, -2.331603e-08,
  -1.503107e-08, -1.616609e-08, -1.675452e-08, -1.732162e-08, -1.769615e-08, 
    -1.880683e-08, -2.006411e-08, -2.108787e-08, -2.148552e-08, 
    -2.228358e-08, -2.268236e-08, -2.271796e-08, -2.311847e-08, 
    -2.296031e-08, -2.334813e-08,
  -1.461513e-08, -1.571613e-08, -1.647372e-08, -1.709452e-08, -1.737989e-08, 
    -1.849712e-08, -1.968615e-08, -2.087408e-08, -2.141841e-08, 
    -2.254504e-08, -2.305598e-08, -2.304703e-08, -2.320666e-08, 
    -2.269897e-08, -2.315116e-08,
  -1.42508e-08, -1.529883e-08, -1.617575e-08, -1.68114e-08, -1.696583e-08, 
    -1.808229e-08, -1.936824e-08, -2.08858e-08, -2.108012e-08, -2.253154e-08, 
    -2.292796e-08, -2.286336e-08, -2.253947e-08, -2.233293e-08, -2.265174e-08,
  -1.384424e-08, -1.485504e-08, -1.586849e-08, -1.657402e-08, -1.665844e-08, 
    -1.777686e-08, -1.938531e-08, -2.065273e-08, -2.101786e-08, 
    -2.243882e-08, -2.278981e-08, -2.283529e-08, -2.220114e-08, 
    -2.201533e-08, -2.237514e-08,
  -1.343086e-08, -1.43976e-08, -1.552711e-08, -1.632823e-08, -1.629344e-08, 
    -1.748312e-08, -1.920067e-08, -2.055702e-08, -2.107928e-08, 
    -2.226816e-08, -2.235693e-08, -2.274948e-08, -2.204561e-08, -2.19071e-08, 
    -2.225791e-08,
  -1.302268e-08, -1.397789e-08, -1.520145e-08, -1.606366e-08, -1.598411e-08, 
    -1.708943e-08, -1.889549e-08, -2.024859e-08, -2.121605e-08, 
    -2.200618e-08, -2.217404e-08, -2.231367e-08, -2.195548e-08, 
    -2.144903e-08, -2.193267e-08,
  -1.253328e-08, -1.364063e-08, -1.487514e-08, -1.573748e-08, -1.574711e-08, 
    -1.671837e-08, -1.854036e-08, -1.993557e-08, -2.092296e-08, 
    -2.164695e-08, -2.188786e-08, -2.233325e-08, -2.1688e-08, -2.101105e-08, 
    -2.197125e-08,
  -2.096581e-08, -2.409992e-08, -2.567575e-08, -2.66449e-08, -2.64094e-08, 
    -2.582421e-08, -2.469927e-08, -2.307243e-08, -2.176447e-08, -2.07461e-08, 
    -2.013565e-08, -1.989015e-08, -1.969312e-08, -1.973467e-08, -2.0047e-08,
  -2.449575e-08, -2.661633e-08, -2.683124e-08, -2.662635e-08, -2.584484e-08, 
    -2.539579e-08, -2.445451e-08, -2.348772e-08, -2.256482e-08, 
    -2.181981e-08, -2.113556e-08, -2.045601e-08, -1.990726e-08, 
    -1.966003e-08, -1.961163e-08,
  -2.775885e-08, -2.861411e-08, -2.822634e-08, -2.801963e-08, -2.757952e-08, 
    -2.717081e-08, -2.636249e-08, -2.568837e-08, -2.513204e-08, 
    -2.490899e-08, -2.474536e-08, -2.436974e-08, -2.387208e-08, 
    -2.344597e-08, -2.30117e-08,
  -2.719902e-08, -2.762066e-08, -2.737292e-08, -2.756278e-08, -2.739829e-08, 
    -2.715626e-08, -2.693324e-08, -2.669261e-08, -2.650206e-08, 
    -2.638395e-08, -2.629837e-08, -2.621034e-08, -2.619547e-08, 
    -2.615319e-08, -2.599407e-08,
  -2.597379e-08, -2.652582e-08, -2.643903e-08, -2.639287e-08, -2.624435e-08, 
    -2.612919e-08, -2.628165e-08, -2.650075e-08, -2.678973e-08, 
    -2.704138e-08, -2.725725e-08, -2.746687e-08, -2.776076e-08, 
    -2.800637e-08, -2.804873e-08,
  -2.500917e-08, -2.541489e-08, -2.518031e-08, -2.520712e-08, -2.517371e-08, 
    -2.553379e-08, -2.589361e-08, -2.611426e-08, -2.612815e-08, 
    -2.610957e-08, -2.5979e-08, -2.610409e-08, -2.627629e-08, -2.652494e-08, 
    -2.635489e-08,
  -2.477237e-08, -2.467791e-08, -2.433528e-08, -2.420754e-08, -2.413363e-08, 
    -2.435198e-08, -2.439103e-08, -2.412451e-08, -2.39585e-08, -2.392205e-08, 
    -2.387822e-08, -2.40321e-08, -2.437292e-08, -2.481048e-08, -2.489058e-08,
  -2.483536e-08, -2.470705e-08, -2.415135e-08, -2.395967e-08, -2.407584e-08, 
    -2.418408e-08, -2.377936e-08, -2.352819e-08, -2.339467e-08, 
    -2.338635e-08, -2.32485e-08, -2.324074e-08, -2.350039e-08, -2.402415e-08, 
    -2.42106e-08,
  -2.466685e-08, -2.468005e-08, -2.384563e-08, -2.363713e-08, -2.359675e-08, 
    -2.320186e-08, -2.280466e-08, -2.297066e-08, -2.30181e-08, -2.290181e-08, 
    -2.270258e-08, -2.263601e-08, -2.283876e-08, -2.319459e-08, -2.355587e-08,
  -2.461966e-08, -2.475196e-08, -2.385742e-08, -2.374325e-08, -2.338917e-08, 
    -2.28306e-08, -2.277719e-08, -2.305649e-08, -2.310803e-08, -2.261048e-08, 
    -2.208999e-08, -2.204327e-08, -2.201047e-08, -2.237804e-08, -2.290225e-08,
  -7.083378e-09, -6.836431e-09, -6.652606e-09, -6.440648e-09, -6.28528e-09, 
    -6.129651e-09, -6.04276e-09, -6.058066e-09, -6.218929e-09, -6.420426e-09, 
    -6.689985e-09, -6.965013e-09, -7.353635e-09, -7.857784e-09, -8.689401e-09,
  -7.605901e-09, -7.422096e-09, -7.467424e-09, -7.407265e-09, -7.435115e-09, 
    -7.440288e-09, -7.508182e-09, -7.622076e-09, -7.755719e-09, 
    -7.944835e-09, -8.207505e-09, -8.488489e-09, -8.864644e-09, -9.46604e-09, 
    -1.036775e-08,
  -9.379559e-09, -8.825955e-09, -8.66225e-09, -8.451776e-09, -8.410344e-09, 
    -8.400807e-09, -8.512302e-09, -8.622683e-09, -8.776034e-09, 
    -8.991221e-09, -9.282387e-09, -9.667008e-09, -1.02105e-08, -1.085235e-08, 
    -1.150106e-08,
  -1.265809e-08, -1.147185e-08, -1.101709e-08, -1.049214e-08, -1.029995e-08, 
    -1.010616e-08, -1.0068e-08, -1.009576e-08, -1.020899e-08, -1.0395e-08, 
    -1.067931e-08, -1.103625e-08, -1.141778e-08, -1.189846e-08, -1.247872e-08,
  -1.760098e-08, -1.608819e-08, -1.50739e-08, -1.414333e-08, -1.35034e-08, 
    -1.300701e-08, -1.268137e-08, -1.245862e-08, -1.233927e-08, -1.23194e-08, 
    -1.236603e-08, -1.248828e-08, -1.279237e-08, -1.315578e-08, -1.366181e-08,
  -2.007943e-08, -1.929298e-08, -1.861935e-08, -1.792601e-08, -1.718686e-08, 
    -1.653035e-08, -1.591427e-08, -1.542436e-08, -1.503451e-08, 
    -1.476723e-08, -1.470992e-08, -1.476194e-08, -1.491424e-08, 
    -1.527991e-08, -1.582919e-08,
  -2.019036e-08, -1.961833e-08, -1.946182e-08, -1.899597e-08, -1.85557e-08, 
    -1.808223e-08, -1.761992e-08, -1.719255e-08, -1.68388e-08, -1.66548e-08, 
    -1.662983e-08, -1.672264e-08, -1.697624e-08, -1.725676e-08, -1.76036e-08,
  -2.200757e-08, -2.142314e-08, -2.108897e-08, -2.061477e-08, -2.022154e-08, 
    -1.974119e-08, -1.938388e-08, -1.908365e-08, -1.887871e-08, 
    -1.879308e-08, -1.880309e-08, -1.886589e-08, -1.898581e-08, 
    -1.921149e-08, -1.960266e-08,
  -2.34999e-08, -2.309391e-08, -2.264267e-08, -2.220493e-08, -2.187074e-08, 
    -2.147974e-08, -2.111045e-08, -2.081273e-08, -2.064071e-08, -2.05512e-08, 
    -2.058168e-08, -2.06956e-08, -2.090492e-08, -2.120466e-08, -2.159112e-08,
  -2.383299e-08, -2.351224e-08, -2.318098e-08, -2.295215e-08, -2.283465e-08, 
    -2.264584e-08, -2.244995e-08, -2.228501e-08, -2.222372e-08, 
    -2.224277e-08, -2.231129e-08, -2.243717e-08, -2.257159e-08, 
    -2.279427e-08, -2.29243e-08,
  -2.715842e-09, -2.403088e-09, -2.337306e-09, -2.167848e-09, -1.972766e-09, 
    -2.028677e-09, -2.25157e-09, -2.558574e-09, -3.582521e-09, -4.396985e-09, 
    -4.764253e-09, -6.128095e-09, -7.599812e-09, -8.700307e-09, -9.4908e-09,
  -3.354965e-09, -3.240397e-09, -3.382223e-09, -3.242187e-09, -3.175214e-09, 
    -3.150125e-09, -3.091942e-09, -3.265651e-09, -3.955233e-09, 
    -4.767842e-09, -5.30562e-09, -6.343814e-09, -7.409589e-09, -8.579754e-09, 
    -9.597606e-09,
  -3.452309e-09, -3.460709e-09, -3.485665e-09, -3.50894e-09, -3.68948e-09, 
    -3.792662e-09, -3.818488e-09, -4.009231e-09, -4.655191e-09, 
    -5.504492e-09, -5.963381e-09, -6.399576e-09, -7.289862e-09, 
    -8.596444e-09, -9.823538e-09,
  -4.374427e-09, -4.170075e-09, -3.858414e-09, -3.727e-09, -3.836717e-09, 
    -4.111001e-09, -4.474053e-09, -4.942713e-09, -5.458004e-09, 
    -6.198904e-09, -6.670627e-09, -6.829551e-09, -7.431368e-09, 
    -8.465629e-09, -9.912442e-09,
  -5.747421e-09, -5.689314e-09, -5.309368e-09, -4.984378e-09, -4.974584e-09, 
    -5.141217e-09, -5.54496e-09, -6.010878e-09, -6.438312e-09, -6.880839e-09, 
    -6.967838e-09, -7.008954e-09, -7.538823e-09, -8.516643e-09, -1.038923e-08,
  -6.620592e-09, -6.642543e-09, -6.525986e-09, -6.391538e-09, -6.565129e-09, 
    -6.749096e-09, -6.924035e-09, -7.117865e-09, -7.285765e-09, 
    -7.370144e-09, -7.374123e-09, -7.60921e-09, -8.190773e-09, -9.360664e-09, 
    -1.112815e-08,
  -8.10426e-09, -7.702713e-09, -7.552308e-09, -7.401359e-09, -7.559267e-09, 
    -7.668938e-09, -7.787052e-09, -7.808953e-09, -7.910102e-09, 
    -8.128617e-09, -8.386597e-09, -8.63165e-09, -9.280258e-09, -1.035312e-08, 
    -1.185188e-08,
  -1.000161e-08, -9.371882e-09, -8.869923e-09, -8.628064e-09, -8.609942e-09, 
    -8.582918e-09, -8.597523e-09, -8.763932e-09, -9.026999e-09, 
    -9.300466e-09, -9.453167e-09, -9.665909e-09, -1.037735e-08, 
    -1.133024e-08, -1.273839e-08,
  -1.165658e-08, -1.097906e-08, -1.0475e-08, -9.976594e-09, -9.780646e-09, 
    -9.681893e-09, -9.758587e-09, -9.878061e-09, -1.008924e-08, 
    -1.027487e-08, -1.059653e-08, -1.118346e-08, -1.170189e-08, 
    -1.264237e-08, -1.377783e-08,
  -1.383413e-08, -1.295447e-08, -1.238426e-08, -1.179902e-08, -1.156392e-08, 
    -1.136047e-08, -1.132434e-08, -1.132344e-08, -1.151891e-08, 
    -1.187449e-08, -1.236666e-08, -1.287583e-08, -1.336807e-08, 
    -1.425687e-08, -1.502768e-08,
  -2.073927e-09, -2.057127e-09, -2.278756e-09, -2.836018e-09, -3.520335e-09, 
    -4.150553e-09, -4.986858e-09, -6.379116e-09, -7.889879e-09, 
    -9.321188e-09, -1.113214e-08, -1.311331e-08, -1.466703e-08, 
    -1.592129e-08, -1.622502e-08,
  -2.116119e-09, -2.200664e-09, -2.401597e-09, -2.848607e-09, -3.487323e-09, 
    -4.140043e-09, -4.902776e-09, -6.148873e-09, -7.684657e-09, 
    -9.207589e-09, -1.09099e-08, -1.290197e-08, -1.453924e-08, -1.572479e-08, 
    -1.627645e-08,
  -2.347512e-09, -2.649915e-09, -2.905587e-09, -3.154712e-09, -3.659051e-09, 
    -4.33479e-09, -4.81322e-09, -5.940596e-09, -7.371827e-09, -9.032431e-09, 
    -1.070993e-08, -1.270341e-08, -1.427073e-08, -1.537816e-08, -1.600253e-08,
  -2.847944e-09, -3.088822e-09, -3.362967e-09, -3.552361e-09, -3.993363e-09, 
    -4.465691e-09, -4.984531e-09, -5.770958e-09, -7.12772e-09, -8.84832e-09, 
    -1.054269e-08, -1.242243e-08, -1.403989e-08, -1.506941e-08, -1.58103e-08,
  -3.231865e-09, -3.422188e-09, -3.656206e-09, -3.956175e-09, -4.401847e-09, 
    -4.732694e-09, -5.05479e-09, -5.59352e-09, -6.929931e-09, -8.683516e-09, 
    -1.03401e-08, -1.223316e-08, -1.383956e-08, -1.473809e-08, -1.537951e-08,
  -3.777574e-09, -3.895384e-09, -4.002659e-09, -4.273682e-09, -4.73583e-09, 
    -4.821556e-09, -5.083387e-09, -5.534425e-09, -6.954621e-09, 
    -8.475644e-09, -1.01626e-08, -1.195308e-08, -1.362313e-08, -1.451721e-08, 
    -1.506566e-08,
  -5.030003e-09, -4.754728e-09, -4.569679e-09, -4.559896e-09, -4.617383e-09, 
    -4.703419e-09, -5.154491e-09, -5.773825e-09, -7.00109e-09, -8.327636e-09, 
    -9.968049e-09, -1.181636e-08, -1.344461e-08, -1.422566e-08, -1.464496e-08,
  -5.170161e-09, -5.009364e-09, -4.85284e-09, -4.57697e-09, -4.458546e-09, 
    -4.715801e-09, -5.404976e-09, -6.11053e-09, -7.081246e-09, -8.310971e-09, 
    -9.848199e-09, -1.153575e-08, -1.324382e-08, -1.397034e-08, -1.4407e-08,
  -4.563799e-09, -4.623697e-09, -4.54463e-09, -4.412091e-09, -4.603216e-09, 
    -5.172771e-09, -5.849474e-09, -6.400266e-09, -7.293317e-09, 
    -8.535439e-09, -9.892136e-09, -1.148498e-08, -1.297445e-08, 
    -1.365415e-08, -1.404694e-08,
  -4.516316e-09, -4.422759e-09, -4.279654e-09, -4.435874e-09, -5.015965e-09, 
    -5.740397e-09, -6.243277e-09, -6.783627e-09, -7.76385e-09, -9.05625e-09, 
    -1.021118e-08, -1.14466e-08, -1.268574e-08, -1.342454e-08, -1.396015e-08,
  -1.137885e-08, -1.230762e-08, -1.271078e-08, -1.273169e-08, -1.252691e-08, 
    -1.242173e-08, -1.209857e-08, -1.14067e-08, -1.006501e-08, -8.619786e-09, 
    -7.456703e-09, -6.113178e-09, -4.944055e-09, -3.831208e-09, -2.937277e-09,
  -1.173704e-08, -1.267595e-08, -1.318308e-08, -1.345231e-08, -1.355428e-08, 
    -1.346436e-08, -1.322771e-08, -1.270717e-08, -1.153996e-08, 
    -1.012249e-08, -8.944671e-09, -7.577637e-09, -6.327365e-09, 
    -5.003496e-09, -3.856041e-09,
  -1.156644e-08, -1.257835e-08, -1.325348e-08, -1.346805e-08, -1.383468e-08, 
    -1.385253e-08, -1.370393e-08, -1.334865e-08, -1.247752e-08, 
    -1.112785e-08, -1.012454e-08, -8.749765e-09, -7.435941e-09, 
    -6.150372e-09, -4.891246e-09,
  -1.148258e-08, -1.257487e-08, -1.34296e-08, -1.381944e-08, -1.431274e-08, 
    -1.45065e-08, -1.448104e-08, -1.421547e-08, -1.338499e-08, -1.224049e-08, 
    -1.122958e-08, -1.006034e-08, -8.740019e-09, -7.483623e-09, -6.09612e-09,
  -1.101521e-08, -1.207722e-08, -1.328812e-08, -1.39225e-08, -1.458791e-08, 
    -1.496771e-08, -1.496742e-08, -1.490738e-08, -1.420038e-08, 
    -1.319792e-08, -1.220385e-08, -1.106056e-08, -9.784704e-09, 
    -8.630374e-09, -7.348647e-09,
  -1.005108e-08, -1.135569e-08, -1.296903e-08, -1.392621e-08, -1.479537e-08, 
    -1.529468e-08, -1.550711e-08, -1.555811e-08, -1.501731e-08, 
    -1.408805e-08, -1.319383e-08, -1.213734e-08, -1.097512e-08, 
    -9.787673e-09, -8.612515e-09,
  -8.988485e-09, -1.068836e-08, -1.264014e-08, -1.371053e-08, -1.476466e-08, 
    -1.541694e-08, -1.601478e-08, -1.630479e-08, -1.586609e-08, 
    -1.497559e-08, -1.411696e-08, -1.317726e-08, -1.210752e-08, 
    -1.084439e-08, -9.72908e-09,
  -7.963881e-09, -9.89089e-09, -1.190798e-08, -1.346864e-08, -1.46201e-08, 
    -1.555004e-08, -1.628082e-08, -1.681983e-08, -1.654055e-08, 
    -1.571624e-08, -1.496946e-08, -1.4237e-08, -1.32732e-08, -1.205144e-08, 
    -1.09008e-08,
  -7.363033e-09, -9.022578e-09, -1.117408e-08, -1.28843e-08, -1.427882e-08, 
    -1.563288e-08, -1.655176e-08, -1.71881e-08, -1.728476e-08, -1.630814e-08, 
    -1.561504e-08, -1.505287e-08, -1.427877e-08, -1.310901e-08, -1.203176e-08,
  -7.111556e-09, -8.410216e-09, -1.036166e-08, -1.250503e-08, -1.407301e-08, 
    -1.543182e-08, -1.668018e-08, -1.749114e-08, -1.776607e-08, 
    -1.687509e-08, -1.623462e-08, -1.586232e-08, -1.532701e-08, 
    -1.413727e-08, -1.31465e-08,
  -2.415805e-09, -1.562248e-09, -1.111623e-09, -8.389187e-10, -7.472081e-10, 
    -7.262199e-10, -7.377896e-10, -7.888172e-10, -8.568328e-10, 
    -9.140924e-10, -9.305299e-10, -8.96167e-10, -8.485954e-10, -8.076146e-10, 
    -7.810817e-10,
  -3.394308e-09, -2.138171e-09, -1.461082e-09, -1.049114e-09, -8.210194e-10, 
    -7.930771e-10, -7.807673e-10, -8.220455e-10, -8.682303e-10, 
    -9.199342e-10, -9.25671e-10, -8.87712e-10, -8.318702e-10, -7.842447e-10, 
    -7.619513e-10,
  -4.222511e-09, -2.645565e-09, -1.755748e-09, -1.306849e-09, -9.585238e-10, 
    -8.67759e-10, -8.388548e-10, -8.573004e-10, -8.910028e-10, -9.403437e-10, 
    -9.353484e-10, -8.93104e-10, -8.285528e-10, -7.8072e-10, -7.73639e-10,
  -5.113638e-09, -3.511522e-09, -2.221265e-09, -1.609113e-09, -1.197073e-09, 
    -9.871556e-10, -9.285304e-10, -9.166077e-10, -9.287845e-10, 
    -9.629876e-10, -9.476551e-10, -8.940335e-10, -8.240605e-10, 
    -7.844455e-10, -7.926932e-10,
  -5.899541e-09, -4.413888e-09, -2.831593e-09, -1.968788e-09, -1.493554e-09, 
    -1.152845e-09, -1.032959e-09, -1.000357e-09, -9.862965e-10, 
    -9.898911e-10, -9.531719e-10, -8.868711e-10, -8.120524e-10, 
    -7.793643e-10, -8.122311e-10,
  -6.867602e-09, -5.33427e-09, -3.707256e-09, -2.461926e-09, -1.86192e-09, 
    -1.38739e-09, -1.148913e-09, -1.074056e-09, -1.039884e-09, -1.011397e-09, 
    -9.587301e-10, -8.772987e-10, -8.001561e-10, -7.807002e-10, -8.502263e-10,
  -7.649698e-09, -6.373979e-09, -4.665596e-09, -3.199762e-09, -2.326809e-09, 
    -1.704993e-09, -1.326538e-09, -1.14651e-09, -1.093331e-09, -1.038834e-09, 
    -9.637739e-10, -8.801544e-10, -8.096579e-10, -8.121191e-10, -9.070621e-10,
  -8.664315e-09, -7.535442e-09, -5.762054e-09, -4.11818e-09, -2.936175e-09, 
    -2.120729e-09, -1.594069e-09, -1.275388e-09, -1.144235e-09, 
    -1.074419e-09, -9.76035e-10, -8.983636e-10, -8.395796e-10, -8.617547e-10, 
    -9.723488e-10,
  -9.708251e-09, -8.659018e-09, -7.009143e-09, -5.182943e-09, -3.745888e-09, 
    -2.663949e-09, -1.965177e-09, -1.492671e-09, -1.216565e-09, 
    -1.109994e-09, -1.012082e-09, -9.275841e-10, -8.911188e-10, 
    -9.233969e-10, -1.05348e-09,
  -1.067634e-08, -9.604483e-09, -8.413057e-09, -6.352421e-09, -4.696539e-09, 
    -3.385704e-09, -2.507573e-09, -1.842666e-09, -1.410293e-09, 
    -1.185609e-09, -1.062905e-09, -9.845236e-10, -9.619044e-10, 
    -1.005772e-09, -1.137122e-09,
  -1.366121e-09, -1.400582e-09, -1.335423e-09, -1.259287e-09, -1.225201e-09, 
    -1.250703e-09, -1.287769e-09, -1.300169e-09, -1.346071e-09, 
    -1.550419e-09, -2.116747e-09, -3.162727e-09, -4.682324e-09, 
    -6.393495e-09, -8.085958e-09,
  -1.388827e-09, -1.405539e-09, -1.342938e-09, -1.280249e-09, -1.249406e-09, 
    -1.259142e-09, -1.291611e-09, -1.312797e-09, -1.396749e-09, 
    -1.712351e-09, -2.43171e-09, -3.662742e-09, -5.322918e-09, -7.113046e-09, 
    -8.868457e-09,
  -1.447101e-09, -1.439009e-09, -1.363884e-09, -1.296219e-09, -1.251079e-09, 
    -1.263202e-09, -1.296477e-09, -1.336711e-09, -1.464699e-09, 
    -1.870976e-09, -2.733602e-09, -4.178301e-09, -5.95935e-09, -7.831276e-09, 
    -9.621316e-09,
  -1.522474e-09, -1.48671e-09, -1.389742e-09, -1.302371e-09, -1.254476e-09, 
    -1.260839e-09, -1.297003e-09, -1.355105e-09, -1.522195e-09, 
    -2.021656e-09, -3.026476e-09, -4.645011e-09, -6.530827e-09, 
    -8.466165e-09, -1.036046e-08,
  -1.581079e-09, -1.520346e-09, -1.401158e-09, -1.303439e-09, -1.250327e-09, 
    -1.259166e-09, -1.307626e-09, -1.372273e-09, -1.576771e-09, 
    -2.172336e-09, -3.336437e-09, -5.102219e-09, -7.091508e-09, 
    -9.098352e-09, -1.118952e-08,
  -1.617909e-09, -1.536918e-09, -1.395212e-09, -1.301276e-09, -1.245498e-09, 
    -1.263999e-09, -1.316938e-09, -1.392673e-09, -1.64045e-09, -2.318788e-09, 
    -3.643865e-09, -5.557262e-09, -7.667518e-09, -9.808438e-09, -1.206259e-08,
  -1.627867e-09, -1.52684e-09, -1.370561e-09, -1.296008e-09, -1.237647e-09, 
    -1.266847e-09, -1.332801e-09, -1.415962e-09, -1.699594e-09, 
    -2.462898e-09, -3.952505e-09, -6.021105e-09, -8.268609e-09, 
    -1.052783e-08, -1.28792e-08,
  -1.624914e-09, -1.492417e-09, -1.345609e-09, -1.287752e-09, -1.237817e-09, 
    -1.279151e-09, -1.344495e-09, -1.431829e-09, -1.753243e-09, 
    -2.594554e-09, -4.25911e-09, -6.493452e-09, -8.845531e-09, -1.121705e-08, 
    -1.360786e-08,
  -1.60107e-09, -1.447756e-09, -1.31422e-09, -1.275245e-09, -1.239547e-09, 
    -1.291662e-09, -1.354794e-09, -1.450217e-09, -1.791531e-09, 
    -2.722846e-09, -4.558931e-09, -6.942962e-09, -9.395632e-09, 
    -1.181307e-08, -1.425857e-08,
  -1.565699e-09, -1.413742e-09, -1.283048e-09, -1.252544e-09, -1.239689e-09, 
    -1.300183e-09, -1.361408e-09, -1.458037e-09, -1.816369e-09, 
    -2.849908e-09, -4.85683e-09, -7.354093e-09, -9.897821e-09, -1.229983e-08, 
    -1.490565e-08,
  -1.589556e-09, -1.765471e-09, -2.145618e-09, -2.74969e-09, -3.919756e-09, 
    -5.749314e-09, -7.631482e-09, -9.340407e-09, -1.134743e-08, 
    -1.419734e-08, -1.689191e-08, -1.887884e-08, -2.048559e-08, 
    -2.169558e-08, -2.263513e-08,
  -1.666608e-09, -1.877611e-09, -2.32513e-09, -3.112833e-09, -4.683754e-09, 
    -6.692717e-09, -8.749407e-09, -1.093536e-08, -1.349598e-08, 
    -1.618438e-08, -1.820876e-08, -1.990445e-08, -2.123402e-08, 
    -2.179381e-08, -2.105871e-08,
  -1.730501e-09, -1.979171e-09, -2.517231e-09, -3.521112e-09, -5.409983e-09, 
    -7.677249e-09, -1.013944e-08, -1.265761e-08, -1.527454e-08, 
    -1.749961e-08, -1.930212e-08, -2.083865e-08, -2.132269e-08, 
    -2.078871e-08, -2.05243e-08,
  -1.803907e-09, -2.065738e-09, -2.695147e-09, -3.951337e-09, -6.130748e-09, 
    -8.629369e-09, -1.130612e-08, -1.382843e-08, -1.634671e-08, 
    -1.834753e-08, -2.015521e-08, -2.069321e-08, -2.03598e-08, -2.044402e-08, 
    -2.068959e-08,
  -1.856228e-09, -2.129102e-09, -2.869988e-09, -4.37293e-09, -6.792477e-09, 
    -9.390146e-09, -1.21566e-08, -1.480096e-08, -1.725751e-08, -1.915011e-08, 
    -1.985186e-08, -1.994314e-08, -2.044087e-08, -2.132072e-08, -2.302057e-08,
  -1.88973e-09, -2.197452e-09, -3.057094e-09, -4.756075e-09, -7.34091e-09, 
    -1.000259e-08, -1.291867e-08, -1.569804e-08, -1.780894e-08, 
    -1.877214e-08, -1.946769e-08, -2.042843e-08, -2.182524e-08, 
    -2.374645e-08, -2.496328e-08,
  -1.916091e-09, -2.26387e-09, -3.249923e-09, -5.097953e-09, -7.765732e-09, 
    -1.051072e-08, -1.364812e-08, -1.621506e-08, -1.759279e-08, -1.86792e-08, 
    -2.014814e-08, -2.19116e-08, -2.394103e-08, -2.527228e-08, -2.634833e-08,
  -1.924495e-09, -2.332867e-09, -3.394709e-09, -5.326132e-09, -8.087641e-09, 
    -1.094097e-08, -1.414517e-08, -1.620431e-08, -1.748347e-08, 
    -1.934327e-08, -2.15228e-08, -2.360033e-08, -2.529154e-08, -2.669487e-08, 
    -2.764056e-08,
  -1.936862e-09, -2.364201e-09, -3.514317e-09, -5.504627e-09, -8.288359e-09, 
    -1.122461e-08, -1.427895e-08, -1.606007e-08, -1.789082e-08, 
    -2.051627e-08, -2.288448e-08, -2.495776e-08, -2.650274e-08, 
    -2.786829e-08, -2.842037e-08,
  -1.923712e-09, -2.395617e-09, -3.577742e-09, -5.619027e-09, -8.364273e-09, 
    -1.136709e-08, -1.423841e-08, -1.612482e-08, -1.866905e-08, -2.15684e-08, 
    -2.40384e-08, -2.592069e-08, -2.752524e-08, -2.864827e-08, -2.89057e-08,
  -4.530814e-09, -6.5511e-09, -9.052319e-09, -1.073145e-08, -1.166483e-08, 
    -1.252014e-08, -1.325582e-08, -1.416427e-08, -1.564548e-08, 
    -1.702917e-08, -1.855164e-08, -2.109166e-08, -2.242141e-08, 
    -2.279881e-08, -2.28581e-08,
  -5.581065e-09, -7.691953e-09, -1.035363e-08, -1.127813e-08, -1.202118e-08, 
    -1.294144e-08, -1.39452e-08, -1.536673e-08, -1.682935e-08, -1.846116e-08, 
    -2.090486e-08, -2.255975e-08, -2.313452e-08, -2.314229e-08, -2.223647e-08,
  -6.682607e-09, -8.878583e-09, -1.114553e-08, -1.145681e-08, -1.256809e-08, 
    -1.372165e-08, -1.501841e-08, -1.662941e-08, -1.826327e-08, 
    -2.057485e-08, -2.236831e-08, -2.325263e-08, -2.312984e-08, 
    -2.236136e-08, -2.029884e-08,
  -7.684245e-09, -9.763394e-09, -1.130943e-08, -1.165044e-08, -1.320042e-08, 
    -1.451898e-08, -1.593038e-08, -1.793884e-08, -1.99866e-08, -2.19335e-08, 
    -2.32446e-08, -2.315321e-08, -2.238949e-08, -2.072233e-08, -1.744705e-08,
  -8.394386e-09, -1.011475e-08, -1.110934e-08, -1.215383e-08, -1.404478e-08, 
    -1.545004e-08, -1.740493e-08, -1.969559e-08, -2.147446e-08, 
    -2.311343e-08, -2.295292e-08, -2.227836e-08, -2.083639e-08, 
    -1.843721e-08, -1.785966e-08,
  -8.84491e-09, -1.030154e-08, -1.121184e-08, -1.294267e-08, -1.498764e-08, 
    -1.670367e-08, -1.90929e-08, -2.114586e-08, -2.257042e-08, -2.255843e-08, 
    -2.207806e-08, -2.090026e-08, -1.943156e-08, -1.926665e-08, -2.114708e-08,
  -9.136315e-09, -1.033154e-08, -1.168928e-08, -1.391703e-08, -1.618989e-08, 
    -1.818482e-08, -2.07629e-08, -2.211939e-08, -2.216175e-08, -2.183194e-08, 
    -2.098718e-08, -2.036503e-08, -2.048443e-08, -2.239646e-08, -2.486831e-08,
  -9.272823e-09, -1.04756e-08, -1.238644e-08, -1.505926e-08, -1.746193e-08, 
    -1.980927e-08, -2.178857e-08, -2.175568e-08, -2.148329e-08, 
    -2.095788e-08, -2.109949e-08, -2.143945e-08, -2.332522e-08, 
    -2.552611e-08, -2.625385e-08,
  -9.384999e-09, -1.079424e-08, -1.329954e-08, -1.641377e-08, -1.885603e-08, 
    -2.100717e-08, -2.180376e-08, -2.113354e-08, -2.082402e-08, 
    -2.165314e-08, -2.24243e-08, -2.381623e-08, -2.608484e-08, -2.717506e-08, 
    -2.666138e-08,
  -9.480789e-09, -1.129619e-08, -1.441588e-08, -1.766059e-08, -1.996719e-08, 
    -2.16217e-08, -2.107115e-08, -2.060493e-08, -2.173944e-08, -2.335973e-08, 
    -2.420932e-08, -2.631889e-08, -2.77702e-08, -2.777197e-08, -2.70436e-08,
  -1.128367e-08, -1.269589e-08, -1.374526e-08, -1.486638e-08, -1.592902e-08, 
    -1.747784e-08, -1.938781e-08, -2.2652e-08, -2.247422e-08, -2.44655e-08, 
    -2.358766e-08, -2.089472e-08, -1.933367e-08, -1.832634e-08, -1.794976e-08,
  -1.10308e-08, -1.239976e-08, -1.344684e-08, -1.45436e-08, -1.562848e-08, 
    -1.720416e-08, -1.989142e-08, -2.219226e-08, -2.10928e-08, -2.325058e-08, 
    -2.678454e-08, -1.985825e-08, -1.887764e-08, -1.829678e-08, -1.79582e-08,
  -1.095714e-08, -1.218845e-08, -1.316756e-08, -1.419341e-08, -1.525667e-08, 
    -1.711461e-08, -1.979921e-08, -2.064823e-08, -2.058797e-08, 
    -2.229896e-08, -2.626435e-08, -1.900415e-08, -1.870065e-08, 
    -1.831574e-08, -1.814551e-08,
  -1.099137e-08, -1.2124e-08, -1.305411e-08, -1.401886e-08, -1.512873e-08, 
    -1.704182e-08, -1.982315e-08, -2.044488e-08, -2.095038e-08, 
    -2.072592e-08, -2.374865e-08, -1.865767e-08, -1.876326e-08, 
    -1.860648e-08, -1.800922e-08,
  -1.113802e-08, -1.219155e-08, -1.306218e-08, -1.399521e-08, -1.509204e-08, 
    -1.701857e-08, -2.018067e-08, -2.067748e-08, -2.08922e-08, -1.946123e-08, 
    -2.168929e-08, -1.894408e-08, -1.885872e-08, -1.901929e-08, -1.761355e-08,
  -1.13098e-08, -1.230258e-08, -1.314043e-08, -1.403374e-08, -1.518219e-08, 
    -1.710127e-08, -2.103118e-08, -2.055388e-08, -1.94475e-08, -1.888028e-08, 
    -2.045451e-08, -1.953681e-08, -1.938336e-08, -1.894699e-08, -1.673996e-08,
  -1.160022e-08, -1.247229e-08, -1.325095e-08, -1.416356e-08, -1.529165e-08, 
    -1.755742e-08, -2.180937e-08, -1.960042e-08, -1.818215e-08, 
    -1.903797e-08, -2.018982e-08, -1.98542e-08, -1.966079e-08, -1.854897e-08, 
    -1.606942e-08,
  -1.180665e-08, -1.262923e-08, -1.345133e-08, -1.431305e-08, -1.554591e-08, 
    -1.814213e-08, -2.128813e-08, -1.842106e-08, -1.816765e-08, 
    -1.963438e-08, -2.08506e-08, -2.026347e-08, -1.975859e-08, -1.748535e-08, 
    -1.588904e-08,
  -1.199036e-08, -1.277984e-08, -1.36386e-08, -1.450609e-08, -1.598252e-08, 
    -1.866509e-08, -2.030062e-08, -1.818014e-08, -1.882603e-08, 
    -2.060847e-08, -2.121214e-08, -2.038075e-08, -1.91263e-08, -1.659544e-08, 
    -1.606806e-08,
  -1.214476e-08, -1.294041e-08, -1.386485e-08, -1.475417e-08, -1.659149e-08, 
    -1.882068e-08, -1.936571e-08, -1.870207e-08, -1.987739e-08, -2.15897e-08, 
    -2.136495e-08, -2.015126e-08, -1.815517e-08, -1.631274e-08, -1.64213e-08,
  -2.163369e-08, -2.377598e-08, -2.49959e-08, -2.556615e-08, -2.702028e-08, 
    -2.632258e-08, -2.386605e-08, -1.899629e-08, -1.704183e-08, 
    -1.608173e-08, -1.446308e-08, -1.29358e-08, -1.201882e-08, -1.131439e-08, 
    -1.103667e-08,
  -2.130684e-08, -2.315237e-08, -2.444644e-08, -2.530217e-08, -2.714718e-08, 
    -3.089878e-08, -2.330667e-08, -2.083424e-08, -1.769826e-08, 
    -1.686712e-08, -1.388889e-08, -1.206013e-08, -1.115318e-08, 
    -1.046163e-08, -9.780043e-09,
  -2.084828e-08, -2.25246e-08, -2.361226e-08, -2.458737e-08, -2.585052e-08, 
    -2.994096e-08, -1.975932e-08, -2.057204e-08, -1.961023e-08, 
    -1.850572e-08, -1.43079e-08, -1.168304e-08, -1.069554e-08, -9.929058e-09, 
    -8.996075e-09,
  -1.975093e-08, -2.190352e-08, -2.290703e-08, -2.401651e-08, -2.498853e-08, 
    -2.772054e-08, -2.111456e-08, -1.862336e-08, -1.906679e-08, 
    -1.983892e-08, -1.468224e-08, -1.159617e-08, -1.096588e-08, 
    -9.911329e-09, -8.899412e-09,
  -1.834944e-08, -2.089963e-08, -2.235093e-08, -2.3094e-08, -2.448492e-08, 
    -2.56368e-08, -2.150335e-08, -1.90017e-08, -1.941153e-08, -1.974404e-08, 
    -1.430065e-08, -1.19837e-08, -1.143206e-08, -1.042464e-08, -9.548602e-09,
  -1.707801e-08, -1.968215e-08, -2.162147e-08, -2.236768e-08, -2.372506e-08, 
    -2.508457e-08, -2.12619e-08, -2.082465e-08, -2.056246e-08, -1.937611e-08, 
    -1.439332e-08, -1.245668e-08, -1.164988e-08, -1.07321e-08, -1.012453e-08,
  -1.603535e-08, -1.869727e-08, -2.059135e-08, -2.164432e-08, -2.302745e-08, 
    -2.401798e-08, -2.168986e-08, -2.198162e-08, -2.095704e-08, 
    -1.786793e-08, -1.366418e-08, -1.24939e-08, -1.1903e-08, -1.116887e-08, 
    -1.070132e-08,
  -1.540445e-08, -1.797312e-08, -1.981923e-08, -2.080751e-08, -2.235252e-08, 
    -2.359726e-08, -2.27705e-08, -2.248647e-08, -2.06727e-08, -1.621834e-08, 
    -1.391127e-08, -1.305839e-08, -1.238199e-08, -1.166499e-08, -1.160486e-08,
  -1.506099e-08, -1.746314e-08, -1.912105e-08, -2.017365e-08, -2.198998e-08, 
    -2.333988e-08, -2.396569e-08, -2.237545e-08, -1.996537e-08, 
    -1.524124e-08, -1.425386e-08, -1.311712e-08, -1.262207e-08, 
    -1.208604e-08, -1.236226e-08,
  -1.488275e-08, -1.712496e-08, -1.86167e-08, -1.966399e-08, -2.17738e-08, 
    -2.36961e-08, -2.46348e-08, -2.172747e-08, -1.899199e-08, -1.492461e-08, 
    -1.435237e-08, -1.339483e-08, -1.315365e-08, -1.299517e-08, -1.348457e-08,
  -1.698062e-08, -1.651457e-08, -1.5341e-08, -1.420847e-08, -1.278547e-08, 
    -1.177166e-08, -1.179852e-08, -1.184575e-08, -1.193596e-08, -1.20813e-08, 
    -1.205365e-08, -1.219389e-08, -1.215086e-08, -1.207133e-08, -1.16565e-08,
  -1.762013e-08, -1.733395e-08, -1.632336e-08, -1.518668e-08, -1.378201e-08, 
    -1.166342e-08, -1.109674e-08, -1.097743e-08, -1.09184e-08, -1.100227e-08, 
    -1.10186e-08, -1.115383e-08, -1.127939e-08, -1.143817e-08, -1.14607e-08,
  -1.867355e-08, -1.81388e-08, -1.758275e-08, -1.645342e-08, -1.471832e-08, 
    -1.225189e-08, -1.103437e-08, -1.069371e-08, -1.073328e-08, -1.0541e-08, 
    -1.059614e-08, -1.069063e-08, -1.07468e-08, -1.077748e-08, -1.081133e-08,
  -2.003206e-08, -1.919127e-08, -1.858975e-08, -1.751391e-08, -1.605392e-08, 
    -1.310955e-08, -1.112339e-08, -1.045614e-08, -1.042912e-08, 
    -1.003116e-08, -9.992973e-09, -9.968442e-09, -1.009681e-08, 
    -1.011353e-08, -1.029757e-08,
  -2.095371e-08, -2.081087e-08, -1.959339e-08, -1.849742e-08, -1.74404e-08, 
    -1.444871e-08, -1.122548e-08, -1.039246e-08, -1.006376e-08, 
    -9.727905e-09, -9.555437e-09, -9.521994e-09, -9.729777e-09, 
    -9.790097e-09, -1.01028e-08,
  -2.155826e-08, -2.201299e-08, -2.122945e-08, -1.954794e-08, -1.842092e-08, 
    -1.584846e-08, -1.161781e-08, -1.052739e-08, -1.010975e-08, 
    -9.732208e-09, -9.516291e-09, -9.586818e-09, -9.761306e-09, 
    -1.006802e-08, -1.07144e-08,
  -2.144804e-08, -2.198833e-08, -2.278193e-08, -2.100737e-08, -1.945183e-08, 
    -1.736618e-08, -1.245919e-08, -1.084917e-08, -1.036686e-08, 
    -9.930339e-09, -9.683899e-09, -9.857501e-09, -1.023505e-08, -1.10173e-08, 
    -1.195574e-08,
  -2.083901e-08, -2.120638e-08, -2.342325e-08, -2.28943e-08, -2.055466e-08, 
    -1.893247e-08, -1.348229e-08, -1.108998e-08, -1.056198e-08, 
    -1.029416e-08, -1.021409e-08, -1.070138e-08, -1.137985e-08, 
    -1.222226e-08, -1.300222e-08,
  -1.953217e-08, -2.015856e-08, -2.295064e-08, -2.412125e-08, -2.201803e-08, 
    -2.019773e-08, -1.472145e-08, -1.127991e-08, -1.085396e-08, 
    -1.090504e-08, -1.095219e-08, -1.160655e-08, -1.228412e-08, 
    -1.302472e-08, -1.365923e-08,
  -1.842177e-08, -1.914899e-08, -2.183559e-08, -2.430611e-08, -2.333825e-08, 
    -2.152363e-08, -1.603171e-08, -1.158233e-08, -1.129591e-08, -1.14978e-08, 
    -1.164938e-08, -1.238605e-08, -1.305529e-08, -1.367162e-08, -1.442271e-08,
  -7.898112e-09, -7.972062e-09, -8.163177e-09, -8.371259e-09, -8.584786e-09, 
    -8.861148e-09, -9.200548e-09, -9.412774e-09, -9.604314e-09, 
    -9.661743e-09, -9.649367e-09, -9.647567e-09, -9.745615e-09, 
    -9.966578e-09, -1.027723e-08,
  -8.665211e-09, -8.738564e-09, -9.007601e-09, -9.311855e-09, -9.491306e-09, 
    -9.642101e-09, -9.866679e-09, -9.908056e-09, -9.880655e-09, 
    -9.798351e-09, -9.89461e-09, -1.014795e-08, -1.044593e-08, -1.09159e-08, 
    -1.149048e-08,
  -9.251227e-09, -9.328217e-09, -9.624394e-09, -9.894574e-09, -9.960615e-09, 
    -9.931838e-09, -9.916267e-09, -9.875356e-09, -9.95133e-09, -1.012919e-08, 
    -1.045069e-08, -1.089113e-08, -1.150217e-08, -1.23187e-08, -1.3292e-08,
  -9.572672e-09, -9.631884e-09, -9.868919e-09, -9.925066e-09, -9.923175e-09, 
    -9.74981e-09, -9.820942e-09, -1.001297e-08, -1.034382e-08, -1.064051e-08, 
    -1.112362e-08, -1.185859e-08, -1.283203e-08, -1.389816e-08, -1.490538e-08,
  -9.862748e-09, -9.721409e-09, -9.661166e-09, -9.562565e-09, -9.570579e-09, 
    -9.50091e-09, -9.793486e-09, -1.018001e-08, -1.061235e-08, -1.117492e-08, 
    -1.200578e-08, -1.29258e-08, -1.415645e-08, -1.527352e-08, -1.64118e-08,
  -9.834356e-09, -9.588125e-09, -9.414981e-09, -9.311627e-09, -9.462403e-09, 
    -9.53719e-09, -1.005079e-08, -1.065734e-08, -1.133229e-08, -1.219886e-08, 
    -1.306372e-08, -1.402956e-08, -1.512105e-08, -1.622485e-08, -1.732237e-08,
  -9.850409e-09, -9.581302e-09, -9.309753e-09, -9.292936e-09, -9.468344e-09, 
    -9.883714e-09, -1.053999e-08, -1.132253e-08, -1.210076e-08, 
    -1.306719e-08, -1.379156e-08, -1.475767e-08, -1.603438e-08, 
    -1.730147e-08, -1.808261e-08,
  -1.002469e-08, -9.686963e-09, -9.52347e-09, -9.468677e-09, -9.761423e-09, 
    -1.042096e-08, -1.121181e-08, -1.202775e-08, -1.298884e-08, 
    -1.388851e-08, -1.488975e-08, -1.617514e-08, -1.724211e-08, 
    -1.785637e-08, -1.81853e-08,
  -1.048073e-08, -9.893815e-09, -9.741672e-09, -9.763741e-09, -1.014076e-08, 
    -1.08675e-08, -1.156689e-08, -1.26399e-08, -1.366606e-08, -1.492925e-08, 
    -1.619835e-08, -1.69873e-08, -1.734126e-08, -1.7637e-08, -1.840095e-08,
  -1.104659e-08, -1.027675e-08, -1.005441e-08, -1.004471e-08, -1.042439e-08, 
    -1.103468e-08, -1.199769e-08, -1.334757e-08, -1.490275e-08, 
    -1.654355e-08, -1.730575e-08, -1.777918e-08, -1.797093e-08, 
    -1.866468e-08, -1.917783e-08,
  -7.735879e-09, -7.616535e-09, -7.562541e-09, -7.509777e-09, -7.461802e-09, 
    -7.457103e-09, -7.476568e-09, -7.456399e-09, -7.447196e-09, 
    -7.419454e-09, -7.323003e-09, -7.191559e-09, -7.049051e-09, 
    -6.916391e-09, -6.824293e-09,
  -9.530738e-09, -9.820646e-09, -1.001922e-08, -1.013618e-08, -1.018762e-08, 
    -1.018091e-08, -1.0125e-08, -9.884377e-09, -9.829071e-09, -9.629061e-09, 
    -9.47315e-09, -9.189164e-09, -8.950061e-09, -8.661971e-09, -8.426818e-09,
  -1.004559e-08, -1.031804e-08, -1.067106e-08, -1.090348e-08, -1.100885e-08, 
    -1.088822e-08, -1.057064e-08, -1.026402e-08, -1.008121e-08, 
    -9.750001e-09, -9.600748e-09, -9.215059e-09, -8.943257e-09, 
    -8.554638e-09, -8.266835e-09,
  -1.005951e-08, -1.025329e-08, -1.052294e-08, -1.075361e-08, -1.096087e-08, 
    -1.110576e-08, -1.079129e-08, -1.054642e-08, -1.041006e-08, 
    -1.002513e-08, -9.909344e-09, -9.51432e-09, -9.111049e-09, -8.591901e-09, 
    -8.273364e-09,
  -1.063205e-08, -1.088026e-08, -1.113166e-08, -1.141447e-08, -1.183655e-08, 
    -1.198331e-08, -1.191697e-08, -1.185662e-08, -1.173524e-08, 
    -1.141035e-08, -1.120185e-08, -1.07095e-08, -1.010222e-08, -9.506369e-09, 
    -9.042837e-09,
  -1.101958e-08, -1.142768e-08, -1.196745e-08, -1.251055e-08, -1.287327e-08, 
    -1.303763e-08, -1.303414e-08, -1.328242e-08, -1.302673e-08, -1.26594e-08, 
    -1.210397e-08, -1.154735e-08, -1.060314e-08, -9.959701e-09, -9.196011e-09,
  -1.132999e-08, -1.22188e-08, -1.309698e-08, -1.392888e-08, -1.426414e-08, 
    -1.44896e-08, -1.437082e-08, -1.422259e-08, -1.371642e-08, -1.343044e-08, 
    -1.264379e-08, -1.206725e-08, -1.123936e-08, -1.029952e-08, -9.300122e-09,
  -1.221724e-08, -1.288895e-08, -1.392753e-08, -1.483302e-08, -1.515428e-08, 
    -1.549476e-08, -1.539081e-08, -1.505974e-08, -1.401652e-08, 
    -1.342069e-08, -1.260634e-08, -1.247012e-08, -1.151529e-08, 
    -1.045722e-08, -9.342455e-09,
  -1.238971e-08, -1.317386e-08, -1.430623e-08, -1.553857e-08, -1.589666e-08, 
    -1.62242e-08, -1.593371e-08, -1.559205e-08, -1.446865e-08, -1.368834e-08, 
    -1.275865e-08, -1.220173e-08, -1.133101e-08, -1.061042e-08, -9.437343e-09,
  -1.203126e-08, -1.32404e-08, -1.445996e-08, -1.581926e-08, -1.642152e-08, 
    -1.68358e-08, -1.624272e-08, -1.616958e-08, -1.510126e-08, -1.417274e-08, 
    -1.295913e-08, -1.210406e-08, -1.14273e-08, -1.061194e-08, -9.525264e-09,
  -1.049269e-09, -9.310964e-10, -9.335243e-10, -9.817681e-10, -1.020793e-09, 
    -1.035315e-09, -1.035365e-09, -1.031483e-09, -1.049323e-09, 
    -1.071114e-09, -1.105186e-09, -1.249548e-09, -1.482481e-09, 
    -1.859232e-09, -2.436477e-09,
  -1.279645e-09, -1.041671e-09, -9.035984e-10, -8.802884e-10, -9.27559e-10, 
    -9.739692e-10, -1.010273e-09, -1.055401e-09, -1.104519e-09, 
    -1.136654e-09, -1.247675e-09, -1.406873e-09, -1.704343e-09, 
    -2.183756e-09, -2.883849e-09,
  -1.966086e-09, -1.523197e-09, -1.238306e-09, -1.051559e-09, -9.91441e-10, 
    -1.017768e-09, -1.068268e-09, -1.122878e-09, -1.201774e-09, 
    -1.297343e-09, -1.453908e-09, -1.668528e-09, -2.012806e-09, 
    -2.567266e-09, -3.317291e-09,
  -2.902518e-09, -2.207395e-09, -1.888708e-09, -1.537356e-09, -1.302665e-09, 
    -1.201304e-09, -1.238229e-09, -1.30402e-09, -1.399131e-09, -1.533815e-09, 
    -1.710539e-09, -1.966532e-09, -2.386044e-09, -2.988571e-09, -3.855255e-09,
  -4.22969e-09, -3.339729e-09, -2.868802e-09, -2.468017e-09, -2.11603e-09, 
    -1.797282e-09, -1.632524e-09, -1.606839e-09, -1.699576e-09, 
    -1.836428e-09, -2.027775e-09, -2.401303e-09, -2.87325e-09, -3.61875e-09, 
    -4.382427e-09,
  -5.698724e-09, -4.679124e-09, -3.999927e-09, -3.560823e-09, -3.236563e-09, 
    -2.942332e-09, -2.707608e-09, -2.395131e-09, -2.305626e-09, 
    -2.423224e-09, -2.66145e-09, -3.025131e-09, -3.517667e-09, -4.116315e-09, 
    -4.723647e-09,
  -6.99077e-09, -6.054269e-09, -5.169842e-09, -4.504325e-09, -4.085434e-09, 
    -3.762022e-09, -3.604173e-09, -3.57486e-09, -3.377588e-09, -3.241831e-09, 
    -3.313459e-09, -3.56606e-09, -3.966994e-09, -4.484367e-09, -5.135885e-09,
  -8.75924e-09, -7.421427e-09, -6.396078e-09, -5.494323e-09, -4.837025e-09, 
    -4.335497e-09, -4.111485e-09, -4.088045e-09, -4.143437e-09, 
    -4.180979e-09, -4.163526e-09, -4.286808e-09, -4.602211e-09, 
    -5.095942e-09, -5.711925e-09,
  -9.746416e-09, -9.526186e-09, -8.246148e-09, -7.017174e-09, -6.147491e-09, 
    -5.474061e-09, -5.00052e-09, -4.826641e-09, -4.90032e-09, -5.059833e-09, 
    -5.278758e-09, -5.426108e-09, -5.649989e-09, -5.96983e-09, -6.452899e-09,
  -1.09075e-08, -1.066852e-08, -1.010767e-08, -8.660781e-09, -7.35894e-09, 
    -6.609551e-09, -6.063976e-09, -5.798218e-09, -5.780652e-09, 
    -5.944542e-09, -6.221373e-09, -6.549607e-09, -6.828161e-09, 
    -7.130566e-09, -7.548989e-09,
  -3.42133e-10, -3.716333e-10, -4.102887e-10, -4.472418e-10, -4.881401e-10, 
    -5.230765e-10, -5.570051e-10, -6.126761e-10, -7.089024e-10, 
    -8.051803e-10, -8.584646e-10, -8.912976e-10, -9.414592e-10, -1.07894e-09, 
    -1.48326e-09,
  -3.575794e-10, -3.759837e-10, -4.15503e-10, -4.529008e-10, -5.011805e-10, 
    -5.490837e-10, -5.907422e-10, -6.539337e-10, -7.524829e-10, 
    -8.471313e-10, -8.943676e-10, -9.21748e-10, -9.55179e-10, -1.10542e-09, 
    -1.53457e-09,
  -4.177491e-10, -4.091614e-10, -4.432392e-10, -4.831183e-10, -5.362213e-10, 
    -5.848734e-10, -6.267211e-10, -6.807604e-10, -7.791441e-10, 
    -8.723888e-10, -9.249757e-10, -9.562056e-10, -9.905959e-10, 
    -1.147318e-09, -1.605335e-09,
  -4.910337e-10, -4.612461e-10, -4.831309e-10, -5.123288e-10, -5.632082e-10, 
    -6.116715e-10, -6.538002e-10, -7.075771e-10, -7.950687e-10, 
    -8.922661e-10, -9.450898e-10, -9.928502e-10, -1.033782e-09, 
    -1.207218e-09, -1.698051e-09,
  -5.908851e-10, -5.375554e-10, -5.494142e-10, -5.638598e-10, -6.118364e-10, 
    -6.543874e-10, -7.014862e-10, -7.518891e-10, -8.331625e-10, 
    -9.210539e-10, -9.75823e-10, -1.040338e-09, -1.10541e-09, -1.307468e-09, 
    -1.85168e-09,
  -7.276963e-10, -6.392601e-10, -6.399701e-10, -6.466892e-10, -6.802254e-10, 
    -7.090398e-10, -7.498181e-10, -7.996575e-10, -8.791595e-10, 
    -9.713362e-10, -1.034321e-09, -1.125334e-09, -1.213418e-09, 
    -1.453208e-09, -2.086155e-09,
  -9.145664e-10, -7.743088e-10, -7.557153e-10, -7.462296e-10, -7.641314e-10, 
    -7.788944e-10, -8.186887e-10, -8.68559e-10, -9.552042e-10, -1.040422e-09, 
    -1.123045e-09, -1.238659e-09, -1.36798e-09, -1.672688e-09, -2.403096e-09,
  -1.197479e-09, -9.828319e-10, -9.195587e-10, -8.801043e-10, -8.910053e-10, 
    -8.908714e-10, -9.307958e-10, -9.815669e-10, -1.076642e-09, 
    -1.157161e-09, -1.265339e-09, -1.41217e-09, -1.599552e-09, -1.982966e-09, 
    -2.807709e-09,
  -1.606758e-09, -1.330862e-09, -1.221597e-09, -1.116401e-09, -1.0845e-09, 
    -1.075817e-09, -1.110854e-09, -1.170589e-09, -1.257304e-09, 
    -1.342026e-09, -1.472685e-09, -1.658026e-09, -1.915368e-09, 
    -2.395289e-09, -3.355945e-09,
  -2.031475e-09, -1.750043e-09, -1.622261e-09, -1.472673e-09, -1.388328e-09, 
    -1.342069e-09, -1.346095e-09, -1.385752e-09, -1.477594e-09, 
    -1.580637e-09, -1.7377e-09, -1.95743e-09, -2.282124e-09, -2.866583e-09, 
    -3.953295e-09,
  -1.010846e-09, -9.15497e-10, -8.242364e-10, -7.962108e-10, -8.149792e-10, 
    -9.348031e-10, -1.145312e-09, -1.388054e-09, -1.701924e-09, 
    -2.271196e-09, -3.266762e-09, -4.860968e-09, -7.217172e-09, -1.015e-08, 
    -1.328226e-08,
  -9.89326e-10, -9.142992e-10, -8.401274e-10, -8.16272e-10, -8.466899e-10, 
    -9.75916e-10, -1.185771e-09, -1.441592e-09, -1.82107e-09, -2.524137e-09, 
    -3.708188e-09, -5.558351e-09, -8.159235e-09, -1.128866e-08, -1.445521e-08,
  -9.688977e-10, -9.131682e-10, -8.632104e-10, -8.413482e-10, -8.819725e-10, 
    -1.016669e-09, -1.229292e-09, -1.512005e-09, -1.982665e-09, 
    -2.832325e-09, -4.210517e-09, -6.275441e-09, -9.049856e-09, 
    -1.230928e-08, -1.572384e-08,
  -9.395688e-10, -9.059915e-10, -8.812022e-10, -8.633025e-10, -9.121302e-10, 
    -1.051081e-09, -1.271726e-09, -1.591203e-09, -2.1789e-09, -3.197343e-09, 
    -4.769474e-09, -7.028056e-09, -9.975149e-09, -1.335335e-08, -1.710594e-08,
  -9.211452e-10, -8.974024e-10, -8.914434e-10, -8.820945e-10, -9.397194e-10, 
    -1.085412e-09, -1.316741e-09, -1.694563e-09, -2.416581e-09, 
    -3.603029e-09, -5.360441e-09, -7.762084e-09, -1.084034e-08, 
    -1.452832e-08, -1.880322e-08,
  -9.19136e-10, -8.917098e-10, -9.072201e-10, -8.984856e-10, -9.657293e-10, 
    -1.117393e-09, -1.371362e-09, -1.817404e-09, -2.687474e-09, 
    -4.036607e-09, -5.947647e-09, -8.510725e-09, -1.181092e-08, -1.58872e-08, 
    -2.015748e-08,
  -9.256324e-10, -8.896623e-10, -9.21715e-10, -9.170654e-10, -9.902961e-10, 
    -1.149144e-09, -1.433179e-09, -1.964536e-09, -2.978669e-09, 
    -4.467056e-09, -6.511613e-09, -9.243387e-09, -1.28317e-08, -1.716341e-08, 
    -2.091654e-08,
  -9.300991e-10, -8.976453e-10, -9.384201e-10, -9.269979e-10, -1.012245e-09, 
    -1.181319e-09, -1.50736e-09, -2.130871e-09, -3.276215e-09, -4.885102e-09, 
    -7.06509e-09, -1.005712e-08, -1.391579e-08, -1.809981e-08, -2.052881e-08,
  -9.432731e-10, -9.213216e-10, -9.520538e-10, -9.397046e-10, -1.033598e-09, 
    -1.213881e-09, -1.586388e-09, -2.305308e-09, -3.567808e-09, 
    -5.269735e-09, -7.616825e-09, -1.083732e-08, -1.476627e-08, 
    -1.831656e-08, -1.9414e-08,
  -9.674276e-10, -9.508431e-10, -9.634256e-10, -9.531836e-10, -1.05287e-09, 
    -1.243453e-09, -1.664538e-09, -2.479908e-09, -3.836392e-09, 
    -5.621721e-09, -8.162536e-09, -1.15373e-08, -1.532602e-08, -1.795087e-08, 
    -1.826376e-08,
  -8.715486e-10, -9.713017e-10, -1.101328e-09, -1.269042e-09, -1.53471e-09, 
    -1.857503e-09, -2.295962e-09, -2.935981e-09, -3.974081e-09, 
    -5.459683e-09, -7.113753e-09, -8.733896e-09, -1.033559e-08, -1.19909e-08, 
    -1.36973e-08,
  -9.453999e-10, -1.036273e-09, -1.196695e-09, -1.40819e-09, -1.708225e-09, 
    -2.089685e-09, -2.644034e-09, -3.522518e-09, -4.864926e-09, -6.50005e-09, 
    -8.167634e-09, -9.889208e-09, -1.16126e-08, -1.337607e-08, -1.501987e-08,
  -9.919974e-10, -1.110684e-09, -1.316689e-09, -1.567354e-09, -1.91712e-09, 
    -2.391435e-09, -3.129206e-09, -4.279355e-09, -5.824609e-09, 
    -7.530307e-09, -9.296165e-09, -1.107717e-08, -1.291072e-08, 
    -1.472923e-08, -1.61819e-08,
  -1.031543e-09, -1.18799e-09, -1.437481e-09, -1.727922e-09, -2.156035e-09, 
    -2.780141e-09, -3.752666e-09, -5.143184e-09, -6.835939e-09, 
    -8.611702e-09, -1.044175e-08, -1.23743e-08, -1.435407e-08, -1.591364e-08, 
    -1.732704e-08,
  -1.08706e-09, -1.274558e-09, -1.563507e-09, -1.912783e-09, -2.462635e-09, 
    -3.28263e-09, -4.483394e-09, -6.060469e-09, -7.824312e-09, -9.694364e-09, 
    -1.169822e-08, -1.376007e-08, -1.553516e-08, -1.705729e-08, -1.843575e-08,
  -1.148625e-09, -1.364192e-09, -1.706137e-09, -2.140221e-09, -2.848655e-09, 
    -3.876296e-09, -5.277657e-09, -6.973015e-09, -8.842648e-09, 
    -1.085356e-08, -1.293857e-08, -1.496093e-08, -1.673901e-08, 
    -1.810328e-08, -1.938627e-08,
  -1.213317e-09, -1.461017e-09, -1.871203e-09, -2.411154e-09, -3.306807e-09, 
    -4.527034e-09, -6.07442e-09, -7.880149e-09, -9.865598e-09, -1.198104e-08, 
    -1.417406e-08, -1.625559e-08, -1.777501e-08, -1.902517e-08, -1.936949e-08,
  -1.280699e-09, -1.566493e-09, -2.06141e-09, -2.729244e-09, -3.822232e-09, 
    -5.202934e-09, -6.854147e-09, -8.793076e-09, -1.0911e-08, -1.317745e-08, 
    -1.54224e-08, -1.724241e-08, -1.853322e-08, -1.941959e-08, -1.85884e-08,
  -1.350355e-09, -1.684435e-09, -2.275568e-09, -3.092253e-09, -4.367054e-09, 
    -5.852343e-09, -7.627885e-09, -9.723875e-09, -1.195409e-08, 
    -1.429108e-08, -1.639835e-08, -1.810972e-08, -1.932986e-08, 
    -1.904783e-08, -1.781777e-08,
  -1.428201e-09, -1.812811e-09, -2.514827e-09, -3.487423e-09, -4.908924e-09, 
    -6.475794e-09, -8.418675e-09, -1.065739e-08, -1.300344e-08, 
    -1.532577e-08, -1.740803e-08, -1.896189e-08, -1.941359e-08, 
    -1.839101e-08, -1.742633e-08,
  -1.354949e-09, -1.499538e-09, -1.649032e-09, -1.97848e-09, -2.375087e-09, 
    -2.899448e-09, -3.478325e-09, -4.130323e-09, -4.834402e-09, 
    -5.588855e-09, -6.47889e-09, -7.556755e-09, -8.869653e-09, -1.04404e-08, 
    -1.218478e-08,
  -1.514236e-09, -1.665619e-09, -1.965851e-09, -2.419915e-09, -2.933431e-09, 
    -3.506554e-09, -4.087696e-09, -4.754913e-09, -5.470335e-09, 
    -6.286439e-09, -7.27177e-09, -8.476386e-09, -9.891713e-09, -1.149774e-08, 
    -1.322951e-08,
  -1.678958e-09, -1.934938e-09, -2.388717e-09, -2.910783e-09, -3.478094e-09, 
    -4.086266e-09, -4.728889e-09, -5.431351e-09, -6.169198e-09, 
    -7.042349e-09, -8.137604e-09, -9.434656e-09, -1.087373e-08, -1.24753e-08, 
    -1.44629e-08,
  -1.919384e-09, -2.276316e-09, -2.840381e-09, -3.388755e-09, -4.024129e-09, 
    -4.688447e-09, -5.367161e-09, -6.055228e-09, -6.856336e-09, 
    -7.888774e-09, -9.083398e-09, -1.036097e-08, -1.183577e-08, 
    -1.368433e-08, -1.596299e-08,
  -2.244051e-09, -2.692542e-09, -3.33216e-09, -3.929583e-09, -4.631525e-09, 
    -5.29487e-09, -5.980842e-09, -6.739252e-09, -7.704082e-09, -8.788123e-09, 
    -9.944642e-09, -1.129344e-08, -1.299133e-08, -1.507245e-08, -1.73859e-08,
  -2.617319e-09, -3.135271e-09, -3.847905e-09, -4.503522e-09, -5.238646e-09, 
    -5.917853e-09, -6.672529e-09, -7.545961e-09, -8.559417e-09, 
    -9.633918e-09, -1.088283e-08, -1.241728e-08, -1.427373e-08, 
    -1.654135e-08, -1.922229e-08,
  -3.010139e-09, -3.620591e-09, -4.409839e-09, -5.092352e-09, -5.86069e-09, 
    -6.571186e-09, -7.405748e-09, -8.359283e-09, -9.424238e-09, 
    -1.056712e-08, -1.194456e-08, -1.359922e-08, -1.575106e-08, 
    -1.852334e-08, -2.155065e-08,
  -3.452192e-09, -4.157645e-09, -4.977889e-09, -5.666743e-09, -6.484116e-09, 
    -7.234852e-09, -8.198398e-09, -9.234822e-09, -1.034055e-08, 
    -1.159938e-08, -1.311302e-08, -1.514458e-08, -1.780836e-08, 
    -2.094136e-08, -2.359103e-08,
  -3.91106e-09, -4.702236e-09, -5.509676e-09, -6.25282e-09, -7.115031e-09, 
    -7.981026e-09, -9.052936e-09, -1.013146e-08, -1.137438e-08, 
    -1.276946e-08, -1.471925e-08, -1.713553e-08, -2.024999e-08, 
    -2.324767e-08, -2.477896e-08,
  -4.39241e-09, -5.212833e-09, -6.020869e-09, -6.838934e-09, -7.780666e-09, 
    -8.769143e-09, -9.929391e-09, -1.114437e-08, -1.255991e-08, 
    -1.435393e-08, -1.66014e-08, -1.965686e-08, -2.28371e-08, -2.464622e-08, 
    -2.391648e-08,
  -1.128067e-09, -1.367369e-09, -1.630468e-09, -2.023095e-09, -2.478775e-09, 
    -3.34728e-09, -4.675347e-09, -6.575807e-09, -9.089346e-09, -1.162394e-08, 
    -1.405946e-08, -1.63522e-08, -1.826406e-08, -1.945663e-08, -2.066445e-08,
  -1.327006e-09, -1.592001e-09, -1.964282e-09, -2.364312e-09, -2.917974e-09, 
    -3.880622e-09, -5.385739e-09, -7.496512e-09, -9.993994e-09, 
    -1.245752e-08, -1.482761e-08, -1.698016e-08, -1.858042e-08, 
    -1.982769e-08, -2.130801e-08,
  -1.544171e-09, -1.820533e-09, -2.213284e-09, -2.639339e-09, -3.306336e-09, 
    -4.502979e-09, -6.193647e-09, -8.398746e-09, -1.087346e-08, 
    -1.326949e-08, -1.5502e-08, -1.743927e-08, -1.88503e-08, -2.026313e-08, 
    -2.117971e-08,
  -1.690349e-09, -1.985261e-09, -2.339418e-09, -2.860697e-09, -3.68942e-09, 
    -5.12355e-09, -6.953281e-09, -9.243228e-09, -1.17e-08, -1.397804e-08, 
    -1.62094e-08, -1.796742e-08, -1.928303e-08, -2.043693e-08, -2.078463e-08,
  -1.835381e-09, -2.189993e-09, -2.532891e-09, -3.144992e-09, -4.186032e-09, 
    -5.810004e-09, -7.738915e-09, -1.010809e-08, -1.252063e-08, 
    -1.472666e-08, -1.680425e-08, -1.834177e-08, -1.954336e-08, -2.04922e-08, 
    -2.054185e-08,
  -2.080407e-09, -2.378943e-09, -2.85017e-09, -3.544493e-09, -4.814651e-09, 
    -6.548638e-09, -8.589535e-09, -1.096144e-08, -1.330839e-08, -1.53768e-08, 
    -1.732124e-08, -1.874817e-08, -1.996649e-08, -2.064271e-08, -2.053404e-08,
  -2.342778e-09, -2.642466e-09, -3.195104e-09, -4.031608e-09, -5.494703e-09, 
    -7.338406e-09, -9.434537e-09, -1.178535e-08, -1.401619e-08, 
    -1.597309e-08, -1.781277e-08, -1.922112e-08, -2.039052e-08, 
    -2.084667e-08, -2.106326e-08,
  -2.55169e-09, -2.944739e-09, -3.601647e-09, -4.614336e-09, -6.222248e-09, 
    -8.142468e-09, -1.025765e-08, -1.257729e-08, -1.462992e-08, -1.65683e-08, 
    -1.836026e-08, -1.978731e-08, -2.082826e-08, -2.127825e-08, -2.176178e-08,
  -2.822117e-09, -3.291498e-09, -4.074103e-09, -5.260878e-09, -6.975205e-09, 
    -8.961491e-09, -1.107927e-08, -1.32822e-08, -1.523404e-08, -1.72046e-08, 
    -1.897274e-08, -2.038358e-08, -2.135319e-08, -2.183009e-08, -2.259267e-08,
  -3.1872e-09, -3.693041e-09, -4.617359e-09, -5.978264e-09, -7.789004e-09, 
    -9.777984e-09, -1.182091e-08, -1.392398e-08, -1.583328e-08, 
    -1.785213e-08, -1.960829e-08, -2.098935e-08, -2.195586e-08, 
    -2.250651e-08, -2.355134e-08,
  -1.957266e-09, -2.72471e-09, -3.575155e-09, -4.863765e-09, -6.456957e-09, 
    -8.686023e-09, -1.181991e-08, -1.620948e-08, -2.054404e-08, 
    -2.345177e-08, -2.460553e-08, -2.352708e-08, -2.20656e-08, -2.259993e-08, 
    -2.332787e-08,
  -2.091302e-09, -2.897896e-09, -3.778077e-09, -5.221555e-09, -6.947278e-09, 
    -9.403164e-09, -1.28531e-08, -1.766405e-08, -2.189027e-08, -2.43485e-08, 
    -2.451194e-08, -2.217189e-08, -2.200072e-08, -2.284651e-08, -2.287114e-08,
  -2.387417e-09, -3.197405e-09, -4.13245e-09, -5.730552e-09, -7.617056e-09, 
    -1.037387e-08, -1.431499e-08, -1.927078e-08, -2.302857e-08, 
    -2.479602e-08, -2.310281e-08, -2.18341e-08, -2.231664e-08, -2.242776e-08, 
    -2.310354e-08,
  -2.758244e-09, -3.551702e-09, -4.592292e-09, -6.384938e-09, -8.470207e-09, 
    -1.165195e-08, -1.616256e-08, -2.111629e-08, -2.407516e-08, 
    -2.414415e-08, -2.176668e-08, -2.214807e-08, -2.252201e-08, 
    -2.274608e-08, -2.433415e-08,
  -3.132158e-09, -3.9245e-09, -5.162376e-09, -7.170661e-09, -9.58748e-09, 
    -1.348163e-08, -1.853172e-08, -2.274362e-08, -2.437971e-08, 
    -2.249409e-08, -2.20728e-08, -2.282623e-08, -2.29036e-08, -2.409792e-08, 
    -2.504182e-08,
  -3.484648e-09, -4.376167e-09, -5.914347e-09, -8.205665e-09, -1.115801e-08, 
    -1.586211e-08, -2.072169e-08, -2.388673e-08, -2.316018e-08, 
    -2.212863e-08, -2.290135e-08, -2.339168e-08, -2.414641e-08, -2.53396e-08, 
    -2.559012e-08,
  -3.858579e-09, -4.976757e-09, -6.935444e-09, -9.49835e-09, -1.328436e-08, 
    -1.849829e-08, -2.247223e-08, -2.354625e-08, -2.245277e-08, 
    -2.320335e-08, -2.392012e-08, -2.452975e-08, -2.553504e-08, 
    -2.601601e-08, -2.517429e-08,
  -4.375242e-09, -5.814087e-09, -8.205222e-09, -1.133551e-08, -1.614116e-08, 
    -2.06161e-08, -2.331025e-08, -2.271693e-08, -2.321114e-08, -2.403396e-08, 
    -2.42353e-08, -2.5181e-08, -2.616286e-08, -2.583398e-08, -2.532381e-08,
  -5.150588e-09, -6.883919e-09, -9.853806e-09, -1.384359e-08, -1.8576e-08, 
    -2.214401e-08, -2.278153e-08, -2.299708e-08, -2.393729e-08, 
    -2.401322e-08, -2.527269e-08, -2.650798e-08, -2.659246e-08, 
    -2.594003e-08, -2.511064e-08,
  -6.112757e-09, -8.288903e-09, -1.214128e-08, -1.649597e-08, -2.054047e-08, 
    -2.230087e-08, -2.279862e-08, -2.387497e-08, -2.425137e-08, 
    -2.526021e-08, -2.66911e-08, -2.668467e-08, -2.608805e-08, -2.552894e-08, 
    -2.50606e-08,
  -8.446648e-09, -9.930397e-09, -1.125084e-08, -1.279481e-08, -1.398392e-08, 
    -1.548592e-08, -1.763565e-08, -1.971734e-08, -2.091901e-08, 
    -2.232905e-08, -2.286955e-08, -2.294812e-08, -2.468694e-08, 
    -2.447205e-08, -2.447826e-08,
  -8.53484e-09, -9.981895e-09, -1.134165e-08, -1.275563e-08, -1.395279e-08, 
    -1.578128e-08, -1.797669e-08, -1.982516e-08, -2.182312e-08, 
    -2.320072e-08, -2.318095e-08, -2.435054e-08, -2.552233e-08, 
    -2.566101e-08, -2.488936e-08,
  -8.982614e-09, -1.026957e-08, -1.142722e-08, -1.296364e-08, -1.420878e-08, 
    -1.613939e-08, -1.834492e-08, -2.066757e-08, -2.266885e-08, 
    -2.341277e-08, -2.372069e-08, -2.504794e-08, -2.628817e-08, 
    -2.656993e-08, -2.571634e-08,
  -9.546715e-09, -1.035991e-08, -1.161964e-08, -1.333955e-08, -1.473555e-08, 
    -1.685362e-08, -1.946324e-08, -2.148982e-08, -2.310233e-08, 
    -2.358526e-08, -2.385908e-08, -2.559484e-08, -2.709181e-08, 
    -2.578223e-08, -2.392613e-08,
  -9.661332e-09, -1.067488e-08, -1.204995e-08, -1.384325e-08, -1.540196e-08, 
    -1.762333e-08, -2.006492e-08, -2.218828e-08, -2.371478e-08, 
    -2.331344e-08, -2.434626e-08, -2.617547e-08, -2.483932e-08, 
    -2.345386e-08, -2.318376e-08,
  -9.989329e-09, -1.116985e-08, -1.260678e-08, -1.43555e-08, -1.598943e-08, 
    -1.863116e-08, -2.118411e-08, -2.315819e-08, -2.324004e-08, 
    -2.331243e-08, -2.458448e-08, -2.428031e-08, -2.247281e-08, 
    -2.286711e-08, -2.221776e-08,
  -1.070072e-08, -1.20139e-08, -1.346968e-08, -1.514394e-08, -1.719173e-08, 
    -2.017496e-08, -2.21336e-08, -2.291066e-08, -2.255504e-08, -2.322562e-08, 
    -2.359479e-08, -2.218058e-08, -2.212925e-08, -2.231894e-08, -2.169229e-08,
  -1.161753e-08, -1.295721e-08, -1.446997e-08, -1.635426e-08, -1.892981e-08, 
    -2.160033e-08, -2.278901e-08, -2.266833e-08, -2.191985e-08, -2.26678e-08, 
    -2.221492e-08, -2.183243e-08, -2.199172e-08, -2.193768e-08, -2.136117e-08,
  -1.268242e-08, -1.405333e-08, -1.573867e-08, -1.807072e-08, -2.090948e-08, 
    -2.281232e-08, -2.26351e-08, -2.103246e-08, -2.185114e-08, -2.253684e-08, 
    -2.28693e-08, -2.23434e-08, -2.183559e-08, -2.135081e-08, -2.089738e-08,
  -1.370224e-08, -1.52039e-08, -1.750867e-08, -2.031012e-08, -2.265685e-08, 
    -2.287003e-08, -2.069102e-08, -2.146188e-08, -2.303389e-08, 
    -2.388908e-08, -2.259643e-08, -2.180372e-08, -2.115098e-08, 
    -2.101264e-08, -2.102196e-08,
  -1.299832e-08, -1.41625e-08, -1.472153e-08, -1.581435e-08, -1.63737e-08, 
    -1.688919e-08, -1.726891e-08, -1.794648e-08, -1.849681e-08, 
    -1.895523e-08, -1.99636e-08, -2.099642e-08, -2.151276e-08, -2.204108e-08, 
    -2.152961e-08,
  -1.393814e-08, -1.481729e-08, -1.537918e-08, -1.637757e-08, -1.667417e-08, 
    -1.718331e-08, -1.780124e-08, -1.832789e-08, -1.864045e-08, 
    -1.897584e-08, -1.992432e-08, -2.095678e-08, -2.184498e-08, 
    -2.210748e-08, -2.200857e-08,
  -1.478069e-08, -1.547633e-08, -1.596251e-08, -1.686382e-08, -1.725792e-08, 
    -1.779421e-08, -1.822901e-08, -1.826699e-08, -1.848267e-08, 
    -1.874408e-08, -1.989893e-08, -2.126645e-08, -2.212712e-08, 
    -2.196607e-08, -2.212077e-08,
  -1.57723e-08, -1.589078e-08, -1.665846e-08, -1.752466e-08, -1.754226e-08, 
    -1.818252e-08, -1.844499e-08, -1.832221e-08, -1.847951e-08, 
    -1.887871e-08, -2.024968e-08, -2.170674e-08, -2.233245e-08, 
    -2.221606e-08, -2.215503e-08,
  -1.63985e-08, -1.634539e-08, -1.727955e-08, -1.812383e-08, -1.822639e-08, 
    -1.859047e-08, -1.866654e-08, -1.851003e-08, -1.864048e-08, 
    -1.918373e-08, -2.066616e-08, -2.225508e-08, -2.308935e-08, 
    -2.268444e-08, -2.196054e-08,
  -1.708769e-08, -1.69043e-08, -1.791904e-08, -1.84171e-08, -1.8797e-08, 
    -1.88724e-08, -1.876818e-08, -1.868139e-08, -1.908675e-08, -1.977417e-08, 
    -2.141542e-08, -2.299983e-08, -2.38403e-08, -2.258867e-08, -2.111983e-08,
  -1.713711e-08, -1.732608e-08, -1.796004e-08, -1.82204e-08, -1.886246e-08, 
    -1.878947e-08, -1.868139e-08, -1.912231e-08, -1.967111e-08, 
    -2.064581e-08, -2.215675e-08, -2.344483e-08, -2.344837e-08, 
    -2.191327e-08, -2.07611e-08,
  -1.709302e-08, -1.734943e-08, -1.762992e-08, -1.81422e-08, -1.856563e-08, 
    -1.858369e-08, -1.898692e-08, -1.939305e-08, -2.030038e-08, 
    -2.109257e-08, -2.25989e-08, -2.333207e-08, -2.277776e-08, -2.14822e-08, 
    -2.045379e-08,
  -1.647584e-08, -1.699495e-08, -1.738889e-08, -1.806602e-08, -1.840796e-08, 
    -1.859413e-08, -1.916014e-08, -1.96627e-08, -2.052974e-08, -2.165894e-08, 
    -2.267212e-08, -2.262155e-08, -2.190359e-08, -2.083995e-08, -1.984797e-08,
  -1.647813e-08, -1.684556e-08, -1.735795e-08, -1.789207e-08, -1.827767e-08, 
    -1.891011e-08, -1.952028e-08, -2.006931e-08, -2.100501e-08, -2.18214e-08, 
    -2.228637e-08, -2.205233e-08, -2.094518e-08, -2.01933e-08, -1.95093e-08,
  -8.726705e-09, -1.154359e-08, -1.350898e-08, -1.60064e-08, -1.851662e-08, 
    -2.018701e-08, -2.094229e-08, -2.11988e-08, -2.092725e-08, -1.989657e-08, 
    -1.857796e-08, -1.739273e-08, -1.632175e-08, -1.607813e-08, -1.663557e-08,
  -1.065328e-08, -1.290926e-08, -1.520832e-08, -1.77052e-08, -1.922075e-08, 
    -2.032252e-08, -2.082155e-08, -2.11113e-08, -2.04718e-08, -1.937031e-08, 
    -1.815967e-08, -1.714026e-08, -1.629137e-08, -1.673909e-08, -1.748769e-08,
  -1.21698e-08, -1.4285e-08, -1.66665e-08, -1.836194e-08, -1.938735e-08, 
    -2.017118e-08, -2.066307e-08, -2.091986e-08, -1.996132e-08, 
    -1.877364e-08, -1.787303e-08, -1.704906e-08, -1.705128e-08, 
    -1.769394e-08, -1.851325e-08,
  -1.35224e-08, -1.545892e-08, -1.765264e-08, -1.863897e-08, -1.946742e-08, 
    -2.000401e-08, -2.052501e-08, -2.047805e-08, -1.930352e-08, -1.84574e-08, 
    -1.78499e-08, -1.775224e-08, -1.809193e-08, -1.864796e-08, -1.919987e-08,
  -1.459685e-08, -1.648896e-08, -1.82621e-08, -1.87438e-08, -1.926645e-08, 
    -1.970113e-08, -2.009357e-08, -1.961735e-08, -1.86349e-08, -1.833708e-08, 
    -1.848504e-08, -1.892862e-08, -1.91121e-08, -1.933411e-08, -1.950622e-08,
  -1.550332e-08, -1.720651e-08, -1.856849e-08, -1.888774e-08, -1.904237e-08, 
    -1.935742e-08, -1.946666e-08, -1.872956e-08, -1.833546e-08, 
    -1.892507e-08, -1.96249e-08, -2.012646e-08, -1.967472e-08, -1.944162e-08, 
    -1.930854e-08,
  -1.62463e-08, -1.782725e-08, -1.870087e-08, -1.876608e-08, -1.887848e-08, 
    -1.903494e-08, -1.876958e-08, -1.82534e-08, -1.875793e-08, -1.976951e-08, 
    -2.053972e-08, -2.051178e-08, -1.957101e-08, -1.913326e-08, -1.893038e-08,
  -1.705939e-08, -1.803165e-08, -1.853708e-08, -1.865057e-08, -1.863128e-08, 
    -1.857397e-08, -1.843946e-08, -1.853644e-08, -1.943573e-08, 
    -2.047781e-08, -2.076795e-08, -2.032419e-08, -1.931209e-08, 
    -1.878162e-08, -1.834023e-08,
  -1.726986e-08, -1.804111e-08, -1.825391e-08, -1.852244e-08, -1.834367e-08, 
    -1.857613e-08, -1.876787e-08, -1.913708e-08, -2.005926e-08, 
    -2.067299e-08, -2.050041e-08, -1.999098e-08, -1.899117e-08, 
    -1.827303e-08, -1.787589e-08,
  -1.733182e-08, -1.777138e-08, -1.811442e-08, -1.840666e-08, -1.869476e-08, 
    -1.884777e-08, -1.898242e-08, -1.959671e-08, -2.023984e-08, 
    -2.063043e-08, -2.032023e-08, -1.96225e-08, -1.870636e-08, -1.791362e-08, 
    -1.760635e-08,
  -7.891961e-09, -1.000076e-08, -1.145553e-08, -1.271875e-08, -1.325159e-08, 
    -1.383087e-08, -1.392682e-08, -1.414568e-08, -1.522792e-08, 
    -1.704423e-08, -1.856408e-08, -1.934242e-08, -1.946337e-08, -1.91052e-08, 
    -1.843483e-08,
  -1.060168e-08, -1.195053e-08, -1.305451e-08, -1.372759e-08, -1.397566e-08, 
    -1.416848e-08, -1.425602e-08, -1.53532e-08, -1.712209e-08, -1.858351e-08, 
    -1.95377e-08, -1.992233e-08, -1.983794e-08, -1.905442e-08, -1.837304e-08,
  -1.276015e-08, -1.353696e-08, -1.411033e-08, -1.434635e-08, -1.438281e-08, 
    -1.458378e-08, -1.563368e-08, -1.734423e-08, -1.85274e-08, -1.952751e-08, 
    -2.017442e-08, -2.025778e-08, -1.947886e-08, -1.838812e-08, -1.698083e-08,
  -1.428388e-08, -1.475348e-08, -1.491647e-08, -1.48373e-08, -1.517782e-08, 
    -1.605992e-08, -1.729518e-08, -1.841926e-08, -1.939755e-08, 
    -2.044739e-08, -2.084709e-08, -2.014597e-08, -1.892351e-08, 
    -1.725366e-08, -1.624736e-08,
  -1.531488e-08, -1.572452e-08, -1.539284e-08, -1.57729e-08, -1.6413e-08, 
    -1.733931e-08, -1.839677e-08, -1.959754e-08, -2.082513e-08, 
    -2.138855e-08, -2.047067e-08, -1.897907e-08, -1.695549e-08, 
    -1.568771e-08, -1.570585e-08,
  -1.628375e-08, -1.639346e-08, -1.623086e-08, -1.679903e-08, -1.751092e-08, 
    -1.86447e-08, -1.992221e-08, -2.123496e-08, -2.143568e-08, -2.022922e-08, 
    -1.840279e-08, -1.653781e-08, -1.534389e-08, -1.53489e-08, -1.586596e-08,
  -1.690812e-08, -1.691781e-08, -1.710858e-08, -1.792869e-08, -1.901962e-08, 
    -2.035295e-08, -2.123818e-08, -2.102134e-08, -1.97422e-08, -1.788893e-08, 
    -1.623818e-08, -1.524685e-08, -1.533202e-08, -1.594887e-08, -1.672647e-08,
  -1.765982e-08, -1.783895e-08, -1.854224e-08, -1.954235e-08, -2.03874e-08, 
    -2.093193e-08, -2.046599e-08, -1.901002e-08, -1.741682e-08, 
    -1.610305e-08, -1.537548e-08, -1.569614e-08, -1.628653e-08, 
    -1.701084e-08, -1.780304e-08,
  -1.852197e-08, -1.879639e-08, -1.918814e-08, -1.98399e-08, -1.995324e-08, 
    -1.955427e-08, -1.842965e-08, -1.729661e-08, -1.629821e-08, -1.58061e-08, 
    -1.606977e-08, -1.655077e-08, -1.706724e-08, -1.76678e-08, -1.830139e-08,
  -1.854845e-08, -1.862708e-08, -1.870711e-08, -1.903573e-08, -1.867815e-08, 
    -1.807742e-08, -1.716745e-08, -1.633606e-08, -1.579214e-08, 
    -1.580169e-08, -1.604338e-08, -1.63339e-08, -1.671289e-08, -1.704457e-08, 
    -1.734682e-08,
  -7.429013e-09, -9.025185e-09, -1.063304e-08, -1.226621e-08, -1.400916e-08, 
    -1.50898e-08, -1.58834e-08, -1.598683e-08, -1.543374e-08, -1.465942e-08, 
    -1.438872e-08, -1.415385e-08, -1.431374e-08, -1.395233e-08, -1.314429e-08,
  -1.071273e-08, -1.155165e-08, -1.29802e-08, -1.400029e-08, -1.513814e-08, 
    -1.599703e-08, -1.62593e-08, -1.544225e-08, -1.486428e-08, -1.473435e-08, 
    -1.484874e-08, -1.499011e-08, -1.49948e-08, -1.435984e-08, -1.372094e-08,
  -1.277887e-08, -1.360633e-08, -1.467777e-08, -1.524984e-08, -1.615498e-08, 
    -1.600804e-08, -1.560606e-08, -1.50442e-08, -1.51755e-08, -1.530863e-08, 
    -1.549704e-08, -1.54932e-08, -1.545117e-08, -1.504894e-08, -1.460376e-08,
  -1.407691e-08, -1.503256e-08, -1.581826e-08, -1.604602e-08, -1.611916e-08, 
    -1.564492e-08, -1.553116e-08, -1.56878e-08, -1.586187e-08, -1.593523e-08, 
    -1.591002e-08, -1.608208e-08, -1.630076e-08, -1.608008e-08, -1.552428e-08,
  -1.513077e-08, -1.58643e-08, -1.611142e-08, -1.60448e-08, -1.595715e-08, 
    -1.600781e-08, -1.633408e-08, -1.646325e-08, -1.637357e-08, 
    -1.627281e-08, -1.665319e-08, -1.713669e-08, -1.749804e-08, 
    -1.720668e-08, -1.634538e-08,
  -1.594317e-08, -1.631967e-08, -1.639007e-08, -1.655058e-08, -1.677606e-08, 
    -1.711016e-08, -1.716956e-08, -1.684861e-08, -1.679175e-08, 
    -1.717998e-08, -1.790968e-08, -1.850581e-08, -1.873585e-08, 
    -1.810576e-08, -1.672742e-08,
  -1.700302e-08, -1.72241e-08, -1.750259e-08, -1.773395e-08, -1.781961e-08, 
    -1.759397e-08, -1.718479e-08, -1.718684e-08, -1.758155e-08, 
    -1.839927e-08, -1.908686e-08, -1.959444e-08, -1.947926e-08, 
    -1.848273e-08, -1.671636e-08,
  -1.830134e-08, -1.830379e-08, -1.808346e-08, -1.7966e-08, -1.764936e-08, 
    -1.75114e-08, -1.776132e-08, -1.82477e-08, -1.88406e-08, -1.931916e-08, 
    -1.992026e-08, -2.006701e-08, -1.9547e-08, -1.821236e-08, -1.683269e-08,
  -1.789835e-08, -1.782128e-08, -1.765857e-08, -1.79418e-08, -1.817244e-08, 
    -1.860185e-08, -1.905366e-08, -1.94579e-08, -1.997888e-08, -2.038437e-08, 
    -2.052619e-08, -2.030658e-08, -1.956794e-08, -1.833117e-08, -1.733397e-08,
  -1.831433e-08, -1.850348e-08, -1.896112e-08, -1.939025e-08, -1.988358e-08, 
    -2.025635e-08, -2.066237e-08, -2.099573e-08, -2.127173e-08, 
    -2.141673e-08, -2.133349e-08, -2.1043e-08, -2.005484e-08, -1.89077e-08, 
    -1.784145e-08,
  -4.805545e-09, -4.722585e-09, -4.837114e-09, -5.023673e-09, -5.153511e-09, 
    -5.432962e-09, -5.763483e-09, -5.420897e-09, -4.956922e-09, 
    -4.313739e-09, -4.05081e-09, -3.401456e-09, -3.634182e-09, -3.791647e-09, 
    -3.861794e-09,
  -6.895593e-09, -6.720999e-09, -6.949907e-09, -6.948036e-09, -7.059506e-09, 
    -6.999719e-09, -6.271103e-09, -5.680829e-09, -5.129071e-09, 
    -4.594795e-09, -4.357398e-09, -3.953425e-09, -3.859477e-09, 
    -3.789244e-09, -4.481848e-09,
  -7.388524e-09, -7.330151e-09, -7.946739e-09, -8.111314e-09, -8.302149e-09, 
    -7.356552e-09, -6.637999e-09, -5.899071e-09, -5.372096e-09, 
    -4.960867e-09, -4.692797e-09, -4.334151e-09, -4.16022e-09, -3.762579e-09, 
    -4.494257e-09,
  -1.063175e-08, -1.015209e-08, -1.031189e-08, -9.307192e-09, -8.482026e-09, 
    -7.43378e-09, -6.740455e-09, -6.113094e-09, -5.681003e-09, -5.468647e-09, 
    -5.03065e-09, -4.647489e-09, -4.357126e-09, -4.248833e-09, -4.710235e-09,
  -1.308499e-08, -1.157424e-08, -1.022663e-08, -8.912341e-09, -7.992334e-09, 
    -7.257761e-09, -6.767851e-09, -6.269245e-09, -6.014108e-09, 
    -5.800377e-09, -5.384682e-09, -5.037866e-09, -4.728789e-09, 
    -4.843566e-09, -4.990544e-09,
  -1.202829e-08, -1.095682e-08, -9.739506e-09, -8.905968e-09, -8.046158e-09, 
    -7.562083e-09, -7.049467e-09, -6.72846e-09, -6.468181e-09, -6.208648e-09, 
    -5.911883e-09, -5.690624e-09, -5.398454e-09, -5.468572e-09, -5.364392e-09,
  -1.285768e-08, -1.19709e-08, -1.094063e-08, -1.012483e-08, -9.130815e-09, 
    -8.447277e-09, -7.928015e-09, -7.572416e-09, -7.209416e-09, 
    -6.978279e-09, -6.878984e-09, -6.677224e-09, -6.149687e-09, 
    -5.838864e-09, -5.598959e-09,
  -1.384533e-08, -1.27444e-08, -1.169514e-08, -1.0933e-08, -1.004775e-08, 
    -9.374165e-09, -8.874316e-09, -8.432194e-09, -8.067704e-09, 
    -7.898935e-09, -7.693852e-09, -7.403703e-09, -6.493445e-09, 
    -6.025954e-09, -5.788765e-09,
  -1.488145e-08, -1.341629e-08, -1.219106e-08, -1.13701e-08, -1.067164e-08, 
    -1.009178e-08, -9.518563e-09, -9.058791e-09, -8.759287e-09, 
    -8.592021e-09, -8.350786e-09, -7.678356e-09, -6.693043e-09, 
    -6.185675e-09, -6.015108e-09,
  -1.543672e-08, -1.412873e-08, -1.286724e-08, -1.176336e-08, -1.099449e-08, 
    -1.040751e-08, -1.002326e-08, -9.606868e-09, -9.456635e-09, 
    -9.207996e-09, -8.675102e-09, -7.6557e-09, -6.833261e-09, -6.363972e-09, 
    -6.388014e-09,
  -3.506721e-09, -3.528217e-09, -3.359555e-09, -3.526146e-09, -3.586285e-09, 
    -3.176326e-09, -2.880709e-09, -2.855106e-09, -3.23111e-09, -4.015766e-09, 
    -5.2246e-09, -6.684722e-09, -8.576748e-09, -1.05287e-08, -1.251107e-08,
  -3.096994e-09, -3.671587e-09, -3.458234e-09, -3.256685e-09, -3.265029e-09, 
    -3.030068e-09, -2.78976e-09, -2.620437e-09, -3.034949e-09, -3.767822e-09, 
    -4.91694e-09, -6.385921e-09, -8.116603e-09, -1.004737e-08, -1.193147e-08,
  -2.677227e-09, -3.137917e-09, -3.750493e-09, -3.102656e-09, -3.016572e-09, 
    -2.910368e-09, -2.770727e-09, -2.527e-09, -2.775488e-09, -3.545023e-09, 
    -4.608392e-09, -5.773956e-09, -7.535981e-09, -9.497487e-09, -1.136239e-08,
  -2.530492e-09, -2.800913e-09, -3.680186e-09, -3.409842e-09, -3.021066e-09, 
    -2.856298e-09, -2.668602e-09, -2.405833e-09, -2.578451e-09, 
    -3.219614e-09, -4.245948e-09, -5.405878e-09, -6.97957e-09, -8.87606e-09, 
    -1.07432e-08,
  -2.305455e-09, -2.416717e-09, -3.243394e-09, -3.581223e-09, -3.147219e-09, 
    -2.893725e-09, -2.713483e-09, -2.398622e-09, -2.347215e-09, 
    -2.871646e-09, -3.898665e-09, -5.006763e-09, -6.352686e-09, 
    -8.284493e-09, -1.022168e-08,
  -2.049049e-09, -2.231889e-09, -2.763202e-09, -3.486984e-09, -3.313263e-09, 
    -2.911438e-09, -2.743136e-09, -2.381811e-09, -2.243744e-09, 
    -2.571146e-09, -3.598662e-09, -4.663149e-09, -5.702444e-09, 
    -7.618862e-09, -9.63857e-09,
  -1.891462e-09, -2.108427e-09, -2.432447e-09, -3.075168e-09, -3.277743e-09, 
    -2.986206e-09, -2.824822e-09, -2.46621e-09, -2.207614e-09, -2.445149e-09, 
    -3.380612e-09, -4.394749e-09, -5.216314e-09, -7.136285e-09, -9.009389e-09,
  -1.731567e-09, -2.02355e-09, -2.380713e-09, -2.678174e-09, -3.015577e-09, 
    -2.939931e-09, -2.897709e-09, -2.579628e-09, -2.241391e-09, 
    -2.423037e-09, -3.379738e-09, -4.35793e-09, -4.870628e-09, -6.660349e-09, 
    -8.410804e-09,
  -1.536058e-09, -1.7099e-09, -2.244866e-09, -2.512326e-09, -2.779028e-09, 
    -2.82102e-09, -2.909169e-09, -2.656051e-09, -2.260756e-09, -2.355238e-09, 
    -3.289614e-09, -4.203632e-09, -4.720061e-09, -6.143397e-09, -7.713991e-09,
  -1.307653e-09, -1.359892e-09, -1.885734e-09, -2.337407e-09, -2.744693e-09, 
    -2.775061e-09, -2.828949e-09, -2.715419e-09, -2.221279e-09, 
    -2.258659e-09, -3.153448e-09, -4.231469e-09, -4.754701e-09, 
    -5.761775e-09, -7.010796e-09,
  -2.242509e-09, -2.735056e-09, -3.315299e-09, -3.845387e-09, -4.883658e-09, 
    -6.307765e-09, -8.025572e-09, -1.005289e-08, -1.245923e-08, 
    -1.498594e-08, -1.709807e-08, -1.870459e-08, -1.986942e-08, 
    -2.079204e-08, -2.169567e-08,
  -2.208455e-09, -2.564466e-09, -3.150365e-09, -3.778674e-09, -4.782555e-09, 
    -6.179361e-09, -7.863512e-09, -9.889531e-09, -1.231919e-08, 
    -1.484877e-08, -1.69475e-08, -1.856626e-08, -1.969576e-08, -2.076533e-08, 
    -2.180001e-08,
  -2.163818e-09, -2.493919e-09, -2.977765e-09, -3.620792e-09, -4.648875e-09, 
    -6.03181e-09, -7.721306e-09, -9.733009e-09, -1.214589e-08, -1.469379e-08, 
    -1.677129e-08, -1.843966e-08, -1.968462e-08, -2.084748e-08, -2.188187e-08,
  -2.21079e-09, -2.431748e-09, -2.863984e-09, -3.461602e-09, -4.481209e-09, 
    -5.870799e-09, -7.547671e-09, -9.513219e-09, -1.190241e-08, 
    -1.442287e-08, -1.654796e-08, -1.8273e-08, -1.960158e-08, -2.08415e-08, 
    -2.196813e-08,
  -2.29703e-09, -2.413105e-09, -2.817627e-09, -3.325067e-09, -4.269648e-09, 
    -5.615978e-09, -7.306901e-09, -9.260816e-09, -1.162138e-08, 
    -1.414653e-08, -1.629811e-08, -1.807721e-08, -1.952379e-08, 
    -2.086132e-08, -2.203585e-08,
  -2.419388e-09, -2.493966e-09, -2.812406e-09, -3.266348e-09, -4.07309e-09, 
    -5.339247e-09, -7.006912e-09, -8.961184e-09, -1.130469e-08, -1.38355e-08, 
    -1.60429e-08, -1.788417e-08, -1.941177e-08, -2.081928e-08, -2.201353e-08,
  -2.538154e-09, -2.575186e-09, -2.81862e-09, -3.241686e-09, -3.958136e-09, 
    -5.065921e-09, -6.692197e-09, -8.634762e-09, -1.098011e-08, 
    -1.350835e-08, -1.57556e-08, -1.766917e-08, -1.931105e-08, -2.079868e-08, 
    -2.199761e-08,
  -2.781193e-09, -2.751438e-09, -2.825844e-09, -3.209404e-09, -3.885756e-09, 
    -4.85447e-09, -6.373966e-09, -8.294441e-09, -1.062536e-08, -1.316653e-08, 
    -1.545463e-08, -1.744883e-08, -1.91787e-08, -2.073723e-08, -2.193774e-08,
  -2.914695e-09, -2.999631e-09, -2.891832e-09, -3.184254e-09, -3.827205e-09, 
    -4.72262e-09, -6.105839e-09, -7.960212e-09, -1.028575e-08, -1.28182e-08, 
    -1.513591e-08, -1.722012e-08, -1.906327e-08, -2.06619e-08, -2.194346e-08,
  -3.054808e-09, -3.159634e-09, -3.17747e-09, -3.193464e-09, -3.763354e-09, 
    -4.60638e-09, -5.887921e-09, -7.633862e-09, -9.930011e-09, -1.248436e-08, 
    -1.482588e-08, -1.699487e-08, -1.889952e-08, -2.056902e-08, -2.197125e-08,
  -5.016546e-09, -6.979997e-09, -9.378773e-09, -1.174694e-08, -1.435463e-08, 
    -1.623244e-08, -1.816804e-08, -1.966211e-08, -2.074892e-08, 
    -2.149666e-08, -2.19068e-08, -2.209448e-08, -2.200683e-08, -2.144301e-08, 
    -2.079209e-08,
  -5.068405e-09, -7.248751e-09, -9.845864e-09, -1.23527e-08, -1.48995e-08, 
    -1.691915e-08, -1.901861e-08, -2.061534e-08, -2.172515e-08, 
    -2.231809e-08, -2.256127e-08, -2.263629e-08, -2.254962e-08, 
    -2.202172e-08, -2.113083e-08,
  -4.754549e-09, -7.168046e-09, -9.973652e-09, -1.261466e-08, -1.530605e-08, 
    -1.766688e-08, -1.990647e-08, -2.150765e-08, -2.25116e-08, -2.305448e-08, 
    -2.320497e-08, -2.306915e-08, -2.304376e-08, -2.239679e-08, -2.143363e-08,
  -4.76498e-09, -6.997043e-09, -9.909654e-09, -1.278933e-08, -1.572352e-08, 
    -1.82874e-08, -2.042313e-08, -2.208956e-08, -2.301964e-08, -2.339866e-08, 
    -2.335612e-08, -2.300955e-08, -2.294337e-08, -2.220249e-08, -2.120932e-08,
  -5.016553e-09, -6.96261e-09, -9.782959e-09, -1.285049e-08, -1.603072e-08, 
    -1.866972e-08, -2.077375e-08, -2.242644e-08, -2.330804e-08, -2.35234e-08, 
    -2.342804e-08, -2.300631e-08, -2.278058e-08, -2.206071e-08, -2.095841e-08,
  -5.245778e-09, -6.832821e-09, -9.640277e-09, -1.271563e-08, -1.621115e-08, 
    -1.886401e-08, -2.099747e-08, -2.260251e-08, -2.361385e-08, 
    -2.360262e-08, -2.324971e-08, -2.267739e-08, -2.260231e-08, 
    -2.172819e-08, -2.039318e-08,
  -5.522786e-09, -7.03863e-09, -9.46102e-09, -1.246099e-08, -1.624695e-08, 
    -1.889826e-08, -2.115097e-08, -2.271172e-08, -2.35535e-08, -2.338989e-08, 
    -2.28351e-08, -2.234072e-08, -2.204207e-08, -2.097983e-08, -1.971979e-08,
  -5.9539e-09, -7.203029e-09, -9.19804e-09, -1.219482e-08, -1.612301e-08, 
    -1.888072e-08, -2.120236e-08, -2.278668e-08, -2.341524e-08, 
    -2.321106e-08, -2.234712e-08, -2.183933e-08, -2.14756e-08, -2.044234e-08, 
    -1.910608e-08,
  -6.342168e-09, -7.404731e-09, -9.00527e-09, -1.201112e-08, -1.584592e-08, 
    -1.874655e-08, -2.121441e-08, -2.29452e-08, -2.324699e-08, -2.291102e-08, 
    -2.187862e-08, -2.140161e-08, -2.094934e-08, -1.9638e-08, -1.834145e-08,
  -6.69679e-09, -7.699224e-09, -9.011321e-09, -1.189141e-08, -1.540361e-08, 
    -1.851898e-08, -2.121332e-08, -2.305019e-08, -2.306517e-08, 
    -2.252859e-08, -2.149428e-08, -2.10343e-08, -2.040242e-08, -1.893032e-08, 
    -1.771032e-08,
  -1.572762e-08, -1.750434e-08, -1.785136e-08, -1.753965e-08, -1.679119e-08, 
    -1.667462e-08, -1.721132e-08, -1.799802e-08, -1.859294e-08, -1.85478e-08, 
    -1.840705e-08, -1.800099e-08, -1.754792e-08, -1.730844e-08, -1.685496e-08,
  -1.587376e-08, -1.771397e-08, -1.778722e-08, -1.710002e-08, -1.652388e-08, 
    -1.702784e-08, -1.777215e-08, -1.852073e-08, -1.902348e-08, 
    -1.882112e-08, -1.861277e-08, -1.814734e-08, -1.770577e-08, 
    -1.734065e-08, -1.694691e-08,
  -1.607589e-08, -1.78386e-08, -1.772157e-08, -1.673371e-08, -1.655437e-08, 
    -1.735434e-08, -1.810517e-08, -1.887681e-08, -1.916316e-08, 
    -1.895421e-08, -1.850714e-08, -1.800299e-08, -1.752e-08, -1.704616e-08, 
    -1.671837e-08,
  -1.616995e-08, -1.792584e-08, -1.762105e-08, -1.649293e-08, -1.678577e-08, 
    -1.795477e-08, -1.868919e-08, -1.906835e-08, -1.938971e-08, 
    -1.907903e-08, -1.852676e-08, -1.793648e-08, -1.749497e-08, 
    -1.704918e-08, -1.685779e-08,
  -1.633717e-08, -1.792714e-08, -1.756439e-08, -1.634011e-08, -1.714177e-08, 
    -1.848026e-08, -1.910458e-08, -1.916934e-08, -1.937074e-08, 
    -1.892354e-08, -1.845471e-08, -1.781632e-08, -1.741738e-08, 
    -1.705273e-08, -1.696926e-08,
  -1.645617e-08, -1.795205e-08, -1.744354e-08, -1.630301e-08, -1.761303e-08, 
    -1.887744e-08, -1.95513e-08, -1.944832e-08, -1.938646e-08, -1.886036e-08, 
    -1.846827e-08, -1.793173e-08, -1.749449e-08, -1.736281e-08, -1.712698e-08,
  -1.66621e-08, -1.789752e-08, -1.730121e-08, -1.637224e-08, -1.81077e-08, 
    -1.937911e-08, -1.994456e-08, -1.953178e-08, -1.906165e-08, 
    -1.880318e-08, -1.840903e-08, -1.819145e-08, -1.801143e-08, -1.79396e-08, 
    -1.762709e-08,
  -1.681985e-08, -1.784015e-08, -1.709522e-08, -1.651629e-08, -1.878014e-08, 
    -1.995785e-08, -1.996058e-08, -1.941347e-08, -1.8527e-08, -1.844599e-08, 
    -1.831502e-08, -1.826963e-08, -1.853757e-08, -1.861587e-08, -1.856647e-08,
  -1.701506e-08, -1.777013e-08, -1.693869e-08, -1.68715e-08, -1.934369e-08, 
    -2.03568e-08, -1.982111e-08, -1.893392e-08, -1.79333e-08, -1.81188e-08, 
    -1.820263e-08, -1.827716e-08, -1.86379e-08, -1.882331e-08, -1.869262e-08,
  -1.710196e-08, -1.768011e-08, -1.688109e-08, -1.740892e-08, -2.005617e-08, 
    -2.05851e-08, -1.955859e-08, -1.78781e-08, -1.764756e-08, -1.802997e-08, 
    -1.836889e-08, -1.865354e-08, -1.878694e-08, -1.88208e-08, -1.873478e-08,
  -1.80818e-08, -1.910914e-08, -1.94093e-08, -1.954898e-08, -1.944637e-08, 
    -1.92556e-08, -1.865099e-08, -1.799132e-08, -1.721349e-08, -1.668594e-08, 
    -1.645093e-08, -1.648124e-08, -1.669369e-08, -1.72025e-08, -1.790803e-08,
  -1.832663e-08, -1.886009e-08, -1.89878e-08, -1.958318e-08, -1.985303e-08, 
    -1.996292e-08, -1.97621e-08, -1.893009e-08, -1.815533e-08, -1.759952e-08, 
    -1.720048e-08, -1.707615e-08, -1.688997e-08, -1.715718e-08, -1.756926e-08,
  -1.84476e-08, -1.870808e-08, -1.888105e-08, -1.967324e-08, -2.004672e-08, 
    -2.038587e-08, -2.040946e-08, -1.96355e-08, -1.885891e-08, -1.843126e-08, 
    -1.806352e-08, -1.799647e-08, -1.767619e-08, -1.765973e-08, -1.77806e-08,
  -1.870336e-08, -1.872392e-08, -1.891066e-08, -1.970838e-08, -2.026484e-08, 
    -2.068458e-08, -2.085913e-08, -2.059842e-08, -1.942739e-08, 
    -1.919474e-08, -1.861285e-08, -1.870356e-08, -1.851588e-08, -1.85192e-08, 
    -1.847184e-08,
  -1.876298e-08, -1.88833e-08, -1.890035e-08, -1.970458e-08, -2.048633e-08, 
    -2.07514e-08, -2.103549e-08, -2.136844e-08, -2.047891e-08, -2.036397e-08, 
    -1.943075e-08, -1.912056e-08, -1.897245e-08, -1.901452e-08, -1.917765e-08,
  -1.871144e-08, -1.89934e-08, -1.880902e-08, -1.980176e-08, -2.062736e-08, 
    -2.097364e-08, -2.122814e-08, -2.16334e-08, -2.120765e-08, -2.135415e-08, 
    -2.088473e-08, -2.028932e-08, -1.949688e-08, -1.928581e-08, -1.943282e-08,
  -1.871652e-08, -1.905227e-08, -1.883808e-08, -1.972681e-08, -2.069117e-08, 
    -2.111978e-08, -2.180052e-08, -2.211681e-08, -2.163549e-08, 
    -2.153646e-08, -2.134057e-08, -2.15123e-08, -2.073745e-08, -2.010518e-08, 
    -1.965095e-08,
  -1.878279e-08, -1.909075e-08, -1.879198e-08, -1.966726e-08, -2.063631e-08, 
    -2.154486e-08, -2.274935e-08, -2.337652e-08, -2.297184e-08, 
    -2.223668e-08, -2.104084e-08, -2.13681e-08, -2.113356e-08, -2.104843e-08, 
    -2.047852e-08,
  -1.888831e-08, -1.913083e-08, -1.882366e-08, -1.953851e-08, -2.067125e-08, 
    -2.187532e-08, -2.334065e-08, -2.448067e-08, -2.435731e-08, 
    -2.409574e-08, -2.261825e-08, -2.134433e-08, -2.097781e-08, 
    -2.093559e-08, -2.08644e-08,
  -1.910607e-08, -1.920791e-08, -1.878329e-08, -1.943689e-08, -2.060447e-08, 
    -2.187561e-08, -2.374769e-08, -2.509368e-08, -2.528976e-08, 
    -2.562279e-08, -2.507462e-08, -2.371932e-08, -2.196393e-08, 
    -2.114581e-08, -2.102869e-08,
  -2.078293e-08, -2.174442e-08, -2.257618e-08, -2.269055e-08, -2.287622e-08, 
    -2.328546e-08, -2.438297e-08, -2.53458e-08, -2.583026e-08, -2.587808e-08, 
    -2.604477e-08, -2.542342e-08, -2.421541e-08, -2.256291e-08, -2.093483e-08,
  -2.063168e-08, -2.152566e-08, -2.212502e-08, -2.252481e-08, -2.262678e-08, 
    -2.250195e-08, -2.322832e-08, -2.377483e-08, -2.471417e-08, 
    -2.513748e-08, -2.541354e-08, -2.560848e-08, -2.532625e-08, -2.44071e-08, 
    -2.2726e-08,
  -2.032486e-08, -2.12814e-08, -2.199741e-08, -2.266123e-08, -2.335763e-08, 
    -2.285919e-08, -2.259804e-08, -2.327661e-08, -2.395577e-08, 
    -2.478226e-08, -2.510301e-08, -2.562828e-08, -2.603994e-08, 
    -2.595414e-08, -2.517685e-08,
  -1.995385e-08, -2.09234e-08, -2.155584e-08, -2.215248e-08, -2.314115e-08, 
    -2.406961e-08, -2.255973e-08, -2.249724e-08, -2.290478e-08, 
    -2.383576e-08, -2.432366e-08, -2.490549e-08, -2.536914e-08, 
    -2.590911e-08, -2.593509e-08,
  -1.947401e-08, -2.04376e-08, -2.131381e-08, -2.16697e-08, -2.266262e-08, 
    -2.467069e-08, -2.429915e-08, -2.241754e-08, -2.248905e-08, 
    -2.304589e-08, -2.350198e-08, -2.435426e-08, -2.481908e-08, -2.53396e-08, 
    -2.592679e-08,
  -1.913283e-08, -1.991621e-08, -2.081343e-08, -2.143792e-08, -2.198978e-08, 
    -2.449399e-08, -2.594071e-08, -2.363805e-08, -2.212794e-08, -2.2361e-08, 
    -2.277308e-08, -2.305438e-08, -2.394613e-08, -2.461316e-08, -2.532247e-08,
  -1.863944e-08, -1.934278e-08, -2.028538e-08, -2.109239e-08, -2.158996e-08, 
    -2.350377e-08, -2.638833e-08, -2.568376e-08, -2.281119e-08, 
    -2.179154e-08, -2.242001e-08, -2.256636e-08, -2.306221e-08, 
    -2.359017e-08, -2.423166e-08,
  -1.853146e-08, -1.895585e-08, -1.967428e-08, -2.055538e-08, -2.108688e-08, 
    -2.27482e-08, -2.575139e-08, -2.71315e-08, -2.472115e-08, -2.146858e-08, 
    -2.178352e-08, -2.186719e-08, -2.261368e-08, -2.277487e-08, -2.348658e-08,
  -1.837944e-08, -1.849338e-08, -1.909875e-08, -1.998946e-08, -2.064816e-08, 
    -2.207677e-08, -2.496445e-08, -2.738062e-08, -2.675254e-08, 
    -2.259199e-08, -2.141348e-08, -2.134261e-08, -2.190764e-08, 
    -2.246463e-08, -2.273852e-08,
  -1.851259e-08, -1.83181e-08, -1.855611e-08, -1.943177e-08, -2.037011e-08, 
    -2.151409e-08, -2.424893e-08, -2.717157e-08, -2.726041e-08, 
    -2.357229e-08, -2.180567e-08, -2.119832e-08, -2.143744e-08, 
    -2.216021e-08, -2.240417e-08,
  -2.431752e-08, -2.406747e-08, -2.44298e-08, -2.432775e-08, -2.460991e-08, 
    -2.462417e-08, -2.424443e-08, -2.266983e-08, -2.062153e-08, 
    -1.900209e-08, -1.784096e-08, -1.702944e-08, -1.693671e-08, 
    -1.711809e-08, -1.761482e-08,
  -2.354043e-08, -2.344273e-08, -2.343958e-08, -2.352485e-08, -2.375869e-08, 
    -2.386896e-08, -2.40483e-08, -2.34017e-08, -2.174364e-08, -1.973517e-08, 
    -1.849967e-08, -1.737815e-08, -1.682555e-08, -1.704723e-08, -1.767159e-08,
  -2.346492e-08, -2.353831e-08, -2.373541e-08, -2.378055e-08, -2.3884e-08, 
    -2.373802e-08, -2.384341e-08, -2.33281e-08, -2.239655e-08, -2.07359e-08, 
    -1.915569e-08, -1.83725e-08, -1.750443e-08, -1.728309e-08, -1.789232e-08,
  -2.320825e-08, -2.337118e-08, -2.356649e-08, -2.349295e-08, -2.376319e-08, 
    -2.3563e-08, -2.335164e-08, -2.330898e-08, -2.240331e-08, -2.139089e-08, 
    -1.984176e-08, -1.900516e-08, -1.849081e-08, -1.793765e-08, -1.804055e-08,
  -2.278678e-08, -2.313827e-08, -2.333874e-08, -2.365168e-08, -2.399434e-08, 
    -2.406631e-08, -2.344147e-08, -2.33666e-08, -2.269344e-08, -2.187927e-08, 
    -2.036331e-08, -1.959835e-08, -1.906383e-08, -1.869698e-08, -1.860026e-08,
  -2.247044e-08, -2.276396e-08, -2.293326e-08, -2.333392e-08, -2.354623e-08, 
    -2.395079e-08, -2.340698e-08, -2.29538e-08, -2.266219e-08, -2.204245e-08, 
    -2.084824e-08, -1.967724e-08, -1.934395e-08, -1.910054e-08, -1.941861e-08,
  -2.210222e-08, -2.251852e-08, -2.23807e-08, -2.295722e-08, -2.306144e-08, 
    -2.364475e-08, -2.358889e-08, -2.265161e-08, -2.233189e-08, 
    -2.184902e-08, -2.13457e-08, -1.998477e-08, -1.940114e-08, -1.939966e-08, 
    -1.986736e-08,
  -2.202182e-08, -2.230337e-08, -2.215901e-08, -2.25534e-08, -2.291297e-08, 
    -2.325883e-08, -2.368466e-08, -2.300992e-08, -2.197657e-08, 
    -2.171422e-08, -2.134432e-08, -2.039179e-08, -1.96406e-08, -1.938714e-08, 
    -2.003861e-08,
  -2.215563e-08, -2.223227e-08, -2.201273e-08, -2.219861e-08, -2.243973e-08, 
    -2.285775e-08, -2.351743e-08, -2.355264e-08, -2.191856e-08, 
    -2.153596e-08, -2.120576e-08, -2.079023e-08, -1.984501e-08, 
    -1.934041e-08, -2.005246e-08,
  -2.241092e-08, -2.212246e-08, -2.190705e-08, -2.193414e-08, -2.21433e-08, 
    -2.239423e-08, -2.294242e-08, -2.380274e-08, -2.229103e-08, 
    -2.142359e-08, -2.1219e-08, -2.103783e-08, -2.046359e-08, -1.968499e-08, 
    -2.00825e-08,
  -1.88532e-08, -1.827098e-08, -1.780569e-08, -1.746013e-08, -1.772138e-08, 
    -1.879719e-08, -2.006449e-08, -2.133204e-08, -2.179721e-08, 
    -2.236778e-08, -2.295623e-08, -2.395117e-08, -2.466515e-08, 
    -2.502681e-08, -2.511958e-08,
  -1.918268e-08, -1.850807e-08, -1.799385e-08, -1.745882e-08, -1.767603e-08, 
    -1.888744e-08, -2.035017e-08, -2.142645e-08, -2.174239e-08, 
    -2.239039e-08, -2.289605e-08, -2.372785e-08, -2.453511e-08, 
    -2.488284e-08, -2.497323e-08,
  -1.945254e-08, -1.865222e-08, -1.811067e-08, -1.743794e-08, -1.773511e-08, 
    -1.903881e-08, -2.051788e-08, -2.142526e-08, -2.173915e-08, 
    -2.242684e-08, -2.292813e-08, -2.401924e-08, -2.492028e-08, 
    -2.515381e-08, -2.520451e-08,
  -1.986478e-08, -1.881646e-08, -1.808878e-08, -1.743379e-08, -1.78653e-08, 
    -1.913693e-08, -2.048768e-08, -2.141696e-08, -2.183839e-08, -2.25743e-08, 
    -2.32232e-08, -2.43964e-08, -2.520285e-08, -2.538752e-08, -2.527311e-08,
  -2.045128e-08, -1.919439e-08, -1.809164e-08, -1.739806e-08, -1.788198e-08, 
    -1.916391e-08, -2.04767e-08, -2.143975e-08, -2.199176e-08, -2.283146e-08, 
    -2.359139e-08, -2.478279e-08, -2.561643e-08, -2.576199e-08, -2.56369e-08,
  -2.104389e-08, -1.968002e-08, -1.834398e-08, -1.748288e-08, -1.779462e-08, 
    -1.906211e-08, -2.046623e-08, -2.145005e-08, -2.213132e-08, -2.30313e-08, 
    -2.401351e-08, -2.525249e-08, -2.628132e-08, -2.662124e-08, -2.649626e-08,
  -2.162404e-08, -2.01874e-08, -1.867084e-08, -1.776482e-08, -1.779012e-08, 
    -1.899439e-08, -2.045596e-08, -2.148136e-08, -2.224719e-08, 
    -2.334855e-08, -2.452648e-08, -2.577286e-08, -2.703599e-08, 
    -2.748128e-08, -2.73723e-08,
  -2.216662e-08, -2.059945e-08, -1.896652e-08, -1.817152e-08, -1.796806e-08, 
    -1.889566e-08, -2.036926e-08, -2.153248e-08, -2.237607e-08, -2.355e-08, 
    -2.484833e-08, -2.61681e-08, -2.7511e-08, -2.811469e-08, -2.792893e-08,
  -2.269697e-08, -2.098542e-08, -1.919881e-08, -1.84334e-08, -1.830687e-08, 
    -1.886819e-08, -2.031527e-08, -2.154623e-08, -2.247906e-08, 
    -2.365744e-08, -2.503438e-08, -2.649407e-08, -2.803805e-08, 
    -2.880177e-08, -2.869051e-08,
  -2.327808e-08, -2.138879e-08, -1.945583e-08, -1.858864e-08, -1.854547e-08, 
    -1.91016e-08, -2.02487e-08, -2.155285e-08, -2.254189e-08, -2.368366e-08, 
    -2.517745e-08, -2.679546e-08, -2.83535e-08, -2.923562e-08, -2.932242e-08,
  -1.571384e-08, -1.820178e-08, -2.193822e-08, -2.474335e-08, -2.64381e-08, 
    -2.591943e-08, -2.340805e-08, -2.093311e-08, -1.943409e-08, 
    -1.824177e-08, -1.743182e-08, -1.7014e-08, -1.693997e-08, -1.697651e-08, 
    -1.710992e-08,
  -1.474064e-08, -1.724786e-08, -2.119056e-08, -2.452408e-08, -2.678763e-08, 
    -2.616793e-08, -2.32529e-08, -2.076331e-08, -1.903315e-08, -1.749983e-08, 
    -1.669042e-08, -1.627983e-08, -1.611537e-08, -1.612541e-08, -1.619672e-08,
  -1.388353e-08, -1.629967e-08, -2.042664e-08, -2.436337e-08, -2.689128e-08, 
    -2.608839e-08, -2.282038e-08, -1.997607e-08, -1.822204e-08, 
    -1.664616e-08, -1.609695e-08, -1.564356e-08, -1.529175e-08, -1.51963e-08, 
    -1.515204e-08,
  -1.318897e-08, -1.539514e-08, -1.970916e-08, -2.421862e-08, -2.712651e-08, 
    -2.624797e-08, -2.22844e-08, -1.955823e-08, -1.777108e-08, -1.629425e-08, 
    -1.594377e-08, -1.542789e-08, -1.504162e-08, -1.488947e-08, -1.47327e-08,
  -1.258873e-08, -1.460235e-08, -1.900678e-08, -2.414539e-08, -2.730163e-08, 
    -2.600532e-08, -2.17798e-08, -1.907462e-08, -1.731998e-08, -1.615745e-08, 
    -1.576725e-08, -1.537609e-08, -1.50472e-08, -1.488335e-08, -1.466013e-08,
  -1.209242e-08, -1.395514e-08, -1.840396e-08, -2.411003e-08, -2.749042e-08, 
    -2.570324e-08, -2.139681e-08, -1.883904e-08, -1.712441e-08, 
    -1.619797e-08, -1.581143e-08, -1.574233e-08, -1.524212e-08, 
    -1.508465e-08, -1.455149e-08,
  -1.161141e-08, -1.339089e-08, -1.794468e-08, -2.408682e-08, -2.756673e-08, 
    -2.527958e-08, -2.110171e-08, -1.873609e-08, -1.694041e-08, 
    -1.625323e-08, -1.611325e-08, -1.605782e-08, -1.548486e-08, 
    -1.519792e-08, -1.456989e-08,
  -1.122689e-08, -1.287997e-08, -1.757172e-08, -2.412463e-08, -2.760116e-08, 
    -2.488287e-08, -2.086925e-08, -1.864729e-08, -1.69084e-08, -1.675851e-08, 
    -1.682982e-08, -1.667022e-08, -1.622216e-08, -1.571359e-08, -1.50624e-08,
  -1.090338e-08, -1.244898e-08, -1.733789e-08, -2.412352e-08, -2.763199e-08, 
    -2.44596e-08, -2.074762e-08, -1.873033e-08, -1.732512e-08, -1.748155e-08, 
    -1.764198e-08, -1.735336e-08, -1.704835e-08, -1.637845e-08, -1.584782e-08,
  -1.070131e-08, -1.208374e-08, -1.714097e-08, -2.413786e-08, -2.758894e-08, 
    -2.408411e-08, -2.072007e-08, -1.889209e-08, -1.775858e-08, 
    -1.808901e-08, -1.818421e-08, -1.802493e-08, -1.782119e-08, -1.70958e-08, 
    -1.668544e-08,
  -2.581665e-08, -2.68559e-08, -2.591572e-08, -2.315337e-08, -1.887052e-08, 
    -1.624653e-08, -1.69499e-08, -1.851663e-08, -2.038255e-08, -2.183824e-08, 
    -2.317327e-08, -2.377373e-08, -2.4578e-08, -2.418233e-08, -2.27582e-08,
  -2.579111e-08, -2.6874e-08, -2.618133e-08, -2.353257e-08, -1.903851e-08, 
    -1.606176e-08, -1.633333e-08, -1.771641e-08, -1.944304e-08, 
    -2.094496e-08, -2.242747e-08, -2.326897e-08, -2.424335e-08, -2.45276e-08, 
    -2.339257e-08,
  -2.559833e-08, -2.658584e-08, -2.61565e-08, -2.374479e-08, -1.907465e-08, 
    -1.560619e-08, -1.601802e-08, -1.719691e-08, -1.913118e-08, 
    -2.059174e-08, -2.191194e-08, -2.26691e-08, -2.357062e-08, -2.425324e-08, 
    -2.366528e-08,
  -2.521184e-08, -2.622632e-08, -2.628643e-08, -2.410394e-08, -1.908012e-08, 
    -1.52713e-08, -1.562674e-08, -1.673181e-08, -1.860608e-08, -2.004363e-08, 
    -2.135819e-08, -2.211596e-08, -2.314133e-08, -2.397162e-08, -2.409572e-08,
  -2.488345e-08, -2.590044e-08, -2.635498e-08, -2.432581e-08, -1.884745e-08, 
    -1.482916e-08, -1.519961e-08, -1.634953e-08, -1.812328e-08, 
    -1.948303e-08, -2.062383e-08, -2.129127e-08, -2.226725e-08, -2.31997e-08, 
    -2.390538e-08,
  -2.455577e-08, -2.559917e-08, -2.636156e-08, -2.446797e-08, -1.836927e-08, 
    -1.461331e-08, -1.496656e-08, -1.62665e-08, -1.789208e-08, -1.905941e-08, 
    -2.009458e-08, -2.083397e-08, -2.178508e-08, -2.258513e-08, -2.339487e-08,
  -2.438774e-08, -2.539111e-08, -2.632303e-08, -2.443437e-08, -1.769635e-08, 
    -1.438995e-08, -1.466821e-08, -1.599825e-08, -1.731458e-08, 
    -1.832511e-08, -1.91476e-08, -1.998397e-08, -2.083422e-08, -2.164195e-08, 
    -2.247084e-08,
  -2.43533e-08, -2.526132e-08, -2.624914e-08, -2.424787e-08, -1.69159e-08, 
    -1.422912e-08, -1.457683e-08, -1.608093e-08, -1.724289e-08, 
    -1.813311e-08, -1.885839e-08, -1.989283e-08, -2.049967e-08, 
    -2.112304e-08, -2.180579e-08,
  -2.441727e-08, -2.523893e-08, -2.607604e-08, -2.35987e-08, -1.63074e-08, 
    -1.408544e-08, -1.458644e-08, -1.610582e-08, -1.696008e-08, 
    -1.784013e-08, -1.843216e-08, -1.961788e-08, -2.006336e-08, 
    -2.063043e-08, -2.096895e-08,
  -2.44662e-08, -2.52192e-08, -2.58843e-08, -2.277184e-08, -1.587976e-08, 
    -1.397603e-08, -1.477689e-08, -1.6301e-08, -1.704791e-08, -1.773812e-08, 
    -1.829948e-08, -1.939816e-08, -1.982753e-08, -2.034071e-08, -2.046372e-08,
  -1.746821e-08, -1.86062e-08, -1.923767e-08, -1.806631e-08, -1.786826e-08, 
    -2.402134e-08, -2.381923e-08, -2.209495e-08, -2.094771e-08, 
    -1.914919e-08, -1.839856e-08, -1.88187e-08, -1.955032e-08, -1.909798e-08, 
    -1.857894e-08,
  -1.750756e-08, -1.940257e-08, -1.948935e-08, -1.843524e-08, -2.003198e-08, 
    -2.264982e-08, -2.172055e-08, -2.067353e-08, -1.968441e-08, 
    -1.881859e-08, -1.834333e-08, -1.867457e-08, -1.93778e-08, -1.872552e-08, 
    -1.809323e-08,
  -1.843224e-08, -1.968336e-08, -1.940309e-08, -1.925184e-08, -2.086102e-08, 
    -2.145645e-08, -2.083504e-08, -1.948105e-08, -1.889986e-08, -1.87653e-08, 
    -1.855627e-08, -1.974719e-08, -2.000041e-08, -1.862707e-08, -1.802785e-08,
  -1.90778e-08, -2.012112e-08, -2.012188e-08, -1.971923e-08, -2.04179e-08, 
    -2.036074e-08, -1.976763e-08, -1.864202e-08, -1.829033e-08, 
    -1.876539e-08, -1.945734e-08, -2.056833e-08, -2.062702e-08, 
    -1.930029e-08, -1.827748e-08,
  -2.047762e-08, -2.105427e-08, -2.074685e-08, -1.936358e-08, -1.929183e-08, 
    -1.972894e-08, -1.900216e-08, -1.83828e-08, -1.841731e-08, -1.908681e-08, 
    -2.037027e-08, -2.093907e-08, -2.096349e-08, -1.97025e-08, -1.884765e-08,
  -2.211127e-08, -2.162526e-08, -2.011932e-08, -1.873134e-08, -1.902938e-08, 
    -1.876434e-08, -1.841875e-08, -1.816915e-08, -1.894884e-08, 
    -1.956094e-08, -2.071502e-08, -2.116183e-08, -2.105336e-08, -2.00768e-08, 
    -1.949867e-08,
  -2.280271e-08, -2.159166e-08, -1.92255e-08, -1.790022e-08, -1.856288e-08, 
    -1.766801e-08, -1.802642e-08, -1.783541e-08, -1.880939e-08, -1.93191e-08, 
    -2.012768e-08, -2.079156e-08, -2.104587e-08, -2.044429e-08, -1.984876e-08,
  -2.263897e-08, -2.056165e-08, -1.793597e-08, -1.727637e-08, -1.763498e-08, 
    -1.75518e-08, -1.777776e-08, -1.801045e-08, -1.858295e-08, -1.943815e-08, 
    -1.993256e-08, -2.027663e-08, -2.042652e-08, -2.053045e-08, -2.028309e-08,
  -2.211676e-08, -1.859575e-08, -1.679663e-08, -1.649396e-08, -1.689012e-08, 
    -1.718751e-08, -1.715696e-08, -1.734735e-08, -1.786787e-08, 
    -1.866307e-08, -1.930211e-08, -1.9817e-08, -1.999108e-08, -2.016789e-08, 
    -2.041755e-08,
  -1.965138e-08, -1.727717e-08, -1.619118e-08, -1.621554e-08, -1.699383e-08, 
    -1.723672e-08, -1.704261e-08, -1.73288e-08, -1.776811e-08, -1.837353e-08, 
    -1.873783e-08, -1.936798e-08, -1.97731e-08, -2.034249e-08, -2.078835e-08,
  -1.781869e-08, -1.923139e-08, -2.022997e-08, -2.079495e-08, -2.059594e-08, 
    -2.162568e-08, -2.020187e-08, -2.260054e-08, -2.540422e-08, 
    -2.101022e-08, -1.938708e-08, -1.561764e-08, -1.448127e-08, 
    -1.455612e-08, -1.41811e-08,
  -1.685751e-08, -1.88963e-08, -1.983024e-08, -2.015586e-08, -2.03015e-08, 
    -2.090523e-08, -2.079646e-08, -2.321809e-08, -2.257172e-08, 
    -1.891391e-08, -1.914747e-08, -1.536848e-08, -1.434308e-08, 
    -1.431987e-08, -1.442618e-08,
  -1.550023e-08, -1.837703e-08, -1.934386e-08, -1.931629e-08, -1.94092e-08, 
    -1.955237e-08, -2.18577e-08, -2.160358e-08, -2.094672e-08, -1.873268e-08, 
    -1.78515e-08, -1.486956e-08, -1.413778e-08, -1.399792e-08, -1.422683e-08,
  -1.71695e-08, -1.873444e-08, -1.834817e-08, -1.853332e-08, -1.963094e-08, 
    -1.819372e-08, -2.073637e-08, -2.089894e-08, -1.883087e-08, 
    -1.886804e-08, -1.664751e-08, -1.461985e-08, -1.361767e-08, 
    -1.343057e-08, -1.336838e-08,
  -1.711201e-08, -1.793122e-08, -1.787158e-08, -1.847986e-08, -1.888507e-08, 
    -1.834769e-08, -1.958155e-08, -2.002495e-08, -1.798881e-08, 
    -1.837224e-08, -1.581534e-08, -1.461286e-08, -1.359296e-08, 
    -1.342368e-08, -1.321937e-08,
  -1.72594e-08, -1.788166e-08, -1.82748e-08, -1.853819e-08, -1.85516e-08, 
    -1.853063e-08, -1.917583e-08, -1.877996e-08, -1.787831e-08, 
    -1.759863e-08, -1.570928e-08, -1.476684e-08, -1.42389e-08, -1.396552e-08, 
    -1.39885e-08,
  -1.843591e-08, -1.856181e-08, -1.85109e-08, -1.81832e-08, -1.763732e-08, 
    -1.836368e-08, -1.881793e-08, -1.8074e-08, -1.794125e-08, -1.696642e-08, 
    -1.59706e-08, -1.53015e-08, -1.474248e-08, -1.459454e-08, -1.47386e-08,
  -1.926757e-08, -1.83608e-08, -1.782615e-08, -1.695454e-08, -1.78034e-08, 
    -1.858684e-08, -1.80987e-08, -1.768389e-08, -1.760053e-08, -1.694273e-08, 
    -1.649979e-08, -1.564815e-08, -1.534558e-08, -1.514177e-08, -1.505969e-08,
  -1.864471e-08, -1.72577e-08, -1.669672e-08, -1.72241e-08, -1.85146e-08, 
    -1.794373e-08, -1.784185e-08, -1.809637e-08, -1.811205e-08, 
    -1.804495e-08, -1.747752e-08, -1.692331e-08, -1.66938e-08, -1.636042e-08, 
    -1.601629e-08,
  -1.669214e-08, -1.624058e-08, -1.705878e-08, -1.83462e-08, -1.835145e-08, 
    -1.822991e-08, -1.871534e-08, -1.859167e-08, -1.842629e-08, 
    -1.827977e-08, -1.790267e-08, -1.774617e-08, -1.738027e-08, 
    -1.674724e-08, -1.622909e-08,
  -2.20776e-08, -2.207565e-08, -2.253118e-08, -2.316947e-08, -2.294458e-08, 
    -2.274132e-08, -2.144704e-08, -1.893946e-08, -1.627928e-08, 
    -1.480677e-08, -1.330464e-08, -1.262928e-08, -1.283095e-08, 
    -1.260135e-08, -1.24495e-08,
  -2.180328e-08, -2.245253e-08, -2.237534e-08, -2.272464e-08, -2.282619e-08, 
    -2.322129e-08, -2.186856e-08, -1.950231e-08, -1.612781e-08, 
    -1.498583e-08, -1.331258e-08, -1.279726e-08, -1.301022e-08, 
    -1.285892e-08, -1.279817e-08,
  -2.065859e-08, -2.138481e-08, -2.2685e-08, -2.228332e-08, -2.2754e-08, 
    -2.339921e-08, -2.195644e-08, -1.996274e-08, -1.612191e-08, 
    -1.490293e-08, -1.262637e-08, -1.283744e-08, -1.324949e-08, 
    -1.322234e-08, -1.321345e-08,
  -1.949055e-08, -1.980665e-08, -2.180728e-08, -2.158959e-08, -2.215594e-08, 
    -2.282857e-08, -2.152504e-08, -1.999135e-08, -1.575646e-08, 
    -1.480463e-08, -1.249576e-08, -1.308196e-08, -1.355852e-08, 
    -1.374013e-08, -1.370534e-08,
  -2.004342e-08, -1.927515e-08, -2.037496e-08, -2.033293e-08, -2.134935e-08, 
    -2.167598e-08, -2.189295e-08, -2.01605e-08, -1.535919e-08, -1.382194e-08, 
    -1.288422e-08, -1.392857e-08, -1.401786e-08, -1.4376e-08, -1.420105e-08,
  -1.990542e-08, -1.924046e-08, -1.934508e-08, -1.958607e-08, -2.070598e-08, 
    -2.093014e-08, -2.147452e-08, -1.97446e-08, -1.5015e-08, -1.365934e-08, 
    -1.393747e-08, -1.418871e-08, -1.40814e-08, -1.449341e-08, -1.453677e-08,
  -1.889697e-08, -1.88017e-08, -1.898014e-08, -1.94516e-08, -2.045504e-08, 
    -2.100146e-08, -2.122128e-08, -1.848273e-08, -1.46312e-08, -1.380169e-08, 
    -1.420092e-08, -1.409792e-08, -1.420232e-08, -1.472542e-08, -1.51486e-08,
  -1.823463e-08, -1.904882e-08, -1.931059e-08, -1.934342e-08, -2.077395e-08, 
    -2.135325e-08, -2.013705e-08, -1.798316e-08, -1.467485e-08, 
    -1.411935e-08, -1.40765e-08, -1.381009e-08, -1.423557e-08, -1.470924e-08, 
    -1.532213e-08,
  -1.819559e-08, -1.89898e-08, -1.919646e-08, -2.02505e-08, -2.123971e-08, 
    -2.082518e-08, -1.964625e-08, -1.71116e-08, -1.467075e-08, -1.354729e-08, 
    -1.348929e-08, -1.391331e-08, -1.405365e-08, -1.464508e-08, -1.547122e-08,
  -1.812234e-08, -1.972652e-08, -2.056743e-08, -2.088476e-08, -2.078892e-08, 
    -1.994612e-08, -1.886784e-08, -1.626297e-08, -1.387878e-08, 
    -1.299558e-08, -1.372144e-08, -1.404374e-08, -1.389044e-08, 
    -1.479185e-08, -1.53656e-08,
  -1.436842e-08, -1.384247e-08, -1.327508e-08, -1.247353e-08, -1.180147e-08, 
    -1.173998e-08, -1.198264e-08, -1.225039e-08, -1.257377e-08, 
    -1.296226e-08, -1.346414e-08, -1.381352e-08, -1.414018e-08, -1.44747e-08, 
    -1.478426e-08,
  -1.485384e-08, -1.436538e-08, -1.379232e-08, -1.325394e-08, -1.262906e-08, 
    -1.2426e-08, -1.274912e-08, -1.304999e-08, -1.329128e-08, -1.371257e-08, 
    -1.42224e-08, -1.456296e-08, -1.496403e-08, -1.539867e-08, -1.575203e-08,
  -1.540662e-08, -1.479718e-08, -1.420259e-08, -1.403136e-08, -1.340167e-08, 
    -1.308434e-08, -1.325387e-08, -1.366285e-08, -1.397061e-08, 
    -1.447851e-08, -1.508077e-08, -1.559227e-08, -1.612893e-08, -1.67295e-08, 
    -1.723826e-08,
  -1.59509e-08, -1.5258e-08, -1.481177e-08, -1.475956e-08, -1.40141e-08, 
    -1.380735e-08, -1.367333e-08, -1.427207e-08, -1.473789e-08, 
    -1.543284e-08, -1.624609e-08, -1.704796e-08, -1.768326e-08, 
    -1.836086e-08, -1.897461e-08,
  -1.665267e-08, -1.588123e-08, -1.545032e-08, -1.547771e-08, -1.469269e-08, 
    -1.460732e-08, -1.417149e-08, -1.505328e-08, -1.580811e-08, 
    -1.674061e-08, -1.759601e-08, -1.836674e-08, -1.901155e-08, -1.95985e-08, 
    -2.01678e-08,
  -1.722314e-08, -1.631997e-08, -1.612239e-08, -1.612542e-08, -1.556138e-08, 
    -1.554334e-08, -1.510425e-08, -1.602931e-08, -1.699308e-08, 
    -1.796661e-08, -1.86037e-08, -1.935057e-08, -1.988337e-08, -2.046018e-08, 
    -2.092311e-08,
  -1.827202e-08, -1.701008e-08, -1.696457e-08, -1.673821e-08, -1.646317e-08, 
    -1.669268e-08, -1.623422e-08, -1.702625e-08, -1.798563e-08, 
    -1.873213e-08, -1.933685e-08, -2.007359e-08, -2.057674e-08, 
    -2.123603e-08, -2.163006e-08,
  -1.924438e-08, -1.774063e-08, -1.783422e-08, -1.760026e-08, -1.748461e-08, 
    -1.774419e-08, -1.731178e-08, -1.788517e-08, -1.861135e-08, -1.93364e-08, 
    -1.992116e-08, -2.064119e-08, -2.12404e-08, -2.197832e-08, -2.238177e-08,
  -1.983013e-08, -1.833984e-08, -1.836275e-08, -1.843712e-08, -1.837331e-08, 
    -1.873184e-08, -1.808842e-08, -1.846306e-08, -1.908631e-08, 
    -1.968916e-08, -2.033397e-08, -2.118297e-08, -2.212578e-08, -2.29717e-08, 
    -2.351599e-08,
  -1.966929e-08, -1.895795e-08, -1.908793e-08, -1.916583e-08, -1.924043e-08, 
    -1.949385e-08, -1.862658e-08, -1.884603e-08, -1.939745e-08, 
    -2.013418e-08, -2.097988e-08, -2.210894e-08, -2.330464e-08, 
    -2.407317e-08, -2.45011e-08,
  -1.269411e-08, -1.345779e-08, -1.33299e-08, -1.425924e-08, -1.490126e-08, 
    -1.562998e-08, -1.626369e-08, -1.689384e-08, -1.73476e-08, -1.765883e-08, 
    -1.794602e-08, -1.81846e-08, -1.840642e-08, -1.865682e-08, -1.891807e-08,
  -1.314864e-08, -1.348807e-08, -1.358034e-08, -1.452944e-08, -1.514642e-08, 
    -1.580961e-08, -1.65354e-08, -1.719292e-08, -1.767329e-08, -1.80916e-08, 
    -1.834403e-08, -1.862694e-08, -1.894032e-08, -1.929704e-08, -1.967141e-08,
  -1.362124e-08, -1.354559e-08, -1.389815e-08, -1.478068e-08, -1.535268e-08, 
    -1.613729e-08, -1.700138e-08, -1.7623e-08, -1.806846e-08, -1.839994e-08, 
    -1.881874e-08, -1.930699e-08, -1.979827e-08, -2.026435e-08, -2.076229e-08,
  -1.36591e-08, -1.361508e-08, -1.418594e-08, -1.50536e-08, -1.56751e-08, 
    -1.667073e-08, -1.741868e-08, -1.786099e-08, -1.847515e-08, 
    -1.915125e-08, -1.99073e-08, -2.048434e-08, -2.098616e-08, -2.150152e-08, 
    -2.206751e-08,
  -1.35799e-08, -1.379217e-08, -1.457629e-08, -1.541481e-08, -1.622956e-08, 
    -1.721236e-08, -1.780677e-08, -1.863411e-08, -1.964644e-08, 
    -2.059265e-08, -2.110351e-08, -2.152624e-08, -2.211605e-08, 
    -2.261799e-08, -2.313014e-08,
  -1.358397e-08, -1.41075e-08, -1.502839e-08, -1.585385e-08, -1.679671e-08, 
    -1.775441e-08, -1.855043e-08, -1.979546e-08, -2.080177e-08, 
    -2.142424e-08, -2.185728e-08, -2.253437e-08, -2.301351e-08, 
    -2.360255e-08, -2.397411e-08,
  -1.370619e-08, -1.452946e-08, -1.551154e-08, -1.642175e-08, -1.737936e-08, 
    -1.846449e-08, -1.958396e-08, -2.096567e-08, -2.169355e-08, -2.23472e-08, 
    -2.304765e-08, -2.366489e-08, -2.428979e-08, -2.471932e-08, -2.471775e-08,
  -1.393726e-08, -1.500411e-08, -1.597883e-08, -1.700288e-08, -1.802059e-08, 
    -1.934918e-08, -2.068754e-08, -2.185014e-08, -2.25249e-08, -2.327388e-08, 
    -2.403728e-08, -2.473447e-08, -2.525366e-08, -2.546043e-08, -2.534028e-08,
  -1.428611e-08, -1.547262e-08, -1.651116e-08, -1.760957e-08, -1.883607e-08, 
    -2.036517e-08, -2.165181e-08, -2.258872e-08, -2.326528e-08, 
    -2.428445e-08, -2.513805e-08, -2.585154e-08, -2.638061e-08, 
    -2.643187e-08, -2.649136e-08,
  -1.470386e-08, -1.595765e-08, -1.705226e-08, -1.834849e-08, -1.976869e-08, 
    -2.125258e-08, -2.227802e-08, -2.322698e-08, -2.419144e-08, 
    -2.523782e-08, -2.60823e-08, -2.674591e-08, -2.718007e-08, -2.72452e-08, 
    -2.738221e-08,
  -1.924198e-08, -1.982324e-08, -1.993289e-08, -2.044063e-08, -2.065844e-08, 
    -2.091832e-08, -2.113218e-08, -2.137197e-08, -2.156267e-08, -2.17234e-08, 
    -2.185132e-08, -2.195428e-08, -2.202655e-08, -2.209451e-08, -2.211832e-08,
  -1.975492e-08, -2.022783e-08, -2.041801e-08, -2.093411e-08, -2.108284e-08, 
    -2.137109e-08, -2.162768e-08, -2.185979e-08, -2.203452e-08, 
    -2.222621e-08, -2.239958e-08, -2.255358e-08, -2.267828e-08, 
    -2.278822e-08, -2.287686e-08,
  -2.052335e-08, -2.094257e-08, -2.112976e-08, -2.157214e-08, -2.167607e-08, 
    -2.199208e-08, -2.214761e-08, -2.233687e-08, -2.256457e-08, 
    -2.282805e-08, -2.308469e-08, -2.336469e-08, -2.362957e-08, 
    -2.388707e-08, -2.410318e-08,
  -2.095573e-08, -2.115994e-08, -2.138091e-08, -2.182656e-08, -2.194136e-08, 
    -2.230661e-08, -2.255231e-08, -2.286128e-08, -2.314317e-08, 
    -2.342303e-08, -2.370443e-08, -2.393667e-08, -2.416131e-08, 
    -2.433771e-08, -2.453654e-08,
  -2.115104e-08, -2.136233e-08, -2.171648e-08, -2.213887e-08, -2.228278e-08, 
    -2.279307e-08, -2.30182e-08, -2.330515e-08, -2.353983e-08, -2.375274e-08, 
    -2.390188e-08, -2.404731e-08, -2.412729e-08, -2.42327e-08, -2.439362e-08,
  -2.137573e-08, -2.162212e-08, -2.202265e-08, -2.234118e-08, -2.273714e-08, 
    -2.320689e-08, -2.345246e-08, -2.375404e-08, -2.391487e-08, 
    -2.411241e-08, -2.425277e-08, -2.441676e-08, -2.457131e-08, 
    -2.483142e-08, -2.504357e-08,
  -2.156558e-08, -2.178966e-08, -2.219721e-08, -2.262415e-08, -2.31411e-08, 
    -2.354806e-08, -2.385192e-08, -2.407667e-08, -2.42577e-08, -2.44806e-08, 
    -2.459085e-08, -2.483406e-08, -2.504094e-08, -2.526668e-08, -2.543024e-08,
  -2.160456e-08, -2.193475e-08, -2.239876e-08, -2.301652e-08, -2.359307e-08, 
    -2.397008e-08, -2.426044e-08, -2.435808e-08, -2.454503e-08, 
    -2.470611e-08, -2.496254e-08, -2.533351e-08, -2.555347e-08, 
    -2.570549e-08, -2.574701e-08,
  -2.167319e-08, -2.206323e-08, -2.265043e-08, -2.340959e-08, -2.393424e-08, 
    -2.425062e-08, -2.439647e-08, -2.461399e-08, -2.486888e-08, 
    -2.506472e-08, -2.542963e-08, -2.558163e-08, -2.558124e-08, 
    -2.561693e-08, -2.556735e-08,
  -2.164445e-08, -2.224361e-08, -2.303703e-08, -2.383086e-08, -2.433197e-08, 
    -2.454281e-08, -2.493279e-08, -2.524755e-08, -2.543163e-08, 
    -2.564886e-08, -2.587944e-08, -2.57771e-08, -2.563998e-08, -2.536775e-08, 
    -2.514615e-08,
  -1.658271e-08, -1.465193e-08, -1.396551e-08, -1.314239e-08, -1.243727e-08, 
    -1.17199e-08, -1.089577e-08, -9.953298e-09, -9.016279e-09, -8.270518e-09, 
    -7.662387e-09, -7.225936e-09, -6.818141e-09, -6.500378e-09, -6.218196e-09,
  -2.425644e-08, -2.193728e-08, -2.047202e-08, -1.892209e-08, -1.748145e-08, 
    -1.632633e-08, -1.528417e-08, -1.434402e-08, -1.345731e-08, 
    -1.264884e-08, -1.18107e-08, -1.107399e-08, -1.048156e-08, -1.007133e-08, 
    -9.703598e-09,
  -2.946952e-08, -2.814794e-08, -2.680074e-08, -2.588482e-08, -2.44915e-08, 
    -2.299807e-08, -2.116007e-08, -1.962537e-08, -1.837995e-08, 
    -1.742169e-08, -1.664656e-08, -1.593686e-08, -1.521735e-08, 
    -1.453071e-08, -1.384682e-08,
  -2.958422e-08, -3.0069e-08, -2.940792e-08, -2.832865e-08, -2.687011e-08, 
    -2.555551e-08, -2.447326e-08, -2.352684e-08, -2.268381e-08, 
    -2.194954e-08, -2.090606e-08, -1.993224e-08, -1.892901e-08, 
    -1.796682e-08, -1.713132e-08,
  -2.63788e-08, -2.666923e-08, -2.663266e-08, -2.687139e-08, -2.654936e-08, 
    -2.597194e-08, -2.513525e-08, -2.423093e-08, -2.320713e-08, 
    -2.221526e-08, -2.143929e-08, -2.092554e-08, -2.062038e-08, 
    -2.029034e-08, -1.987805e-08,
  -2.637e-08, -2.637669e-08, -2.61312e-08, -2.619682e-08, -2.614633e-08, 
    -2.629237e-08, -2.61815e-08, -2.574302e-08, -2.503048e-08, -2.423883e-08, 
    -2.323236e-08, -2.21469e-08, -2.113778e-08, -2.040826e-08, -1.996718e-08,
  -2.788068e-08, -2.735779e-08, -2.670477e-08, -2.633709e-08, -2.603963e-08, 
    -2.596236e-08, -2.602685e-08, -2.608841e-08, -2.604757e-08, 
    -2.574233e-08, -2.510559e-08, -2.422923e-08, -2.318796e-08, 
    -2.210887e-08, -2.106533e-08,
  -2.761504e-08, -2.770238e-08, -2.757118e-08, -2.724609e-08, -2.681787e-08, 
    -2.630338e-08, -2.581019e-08, -2.530547e-08, -2.497354e-08, 
    -2.487514e-08, -2.500288e-08, -2.490877e-08, -2.457464e-08, 
    -2.406097e-08, -2.320132e-08,
  -2.751744e-08, -2.748294e-08, -2.742819e-08, -2.73823e-08, -2.747956e-08, 
    -2.733666e-08, -2.6834e-08, -2.638376e-08, -2.568686e-08, -2.48764e-08, 
    -2.410638e-08, -2.384113e-08, -2.38119e-08, -2.387068e-08, -2.400926e-08,
  -2.747547e-08, -2.780127e-08, -2.782327e-08, -2.788463e-08, -2.78125e-08, 
    -2.797419e-08, -2.777586e-08, -2.730386e-08, -2.676473e-08, 
    -2.604122e-08, -2.510838e-08, -2.445499e-08, -2.398783e-08, 
    -2.372102e-08, -2.38916e-08,
  -2.763176e-09, -2.079386e-09, -2.154259e-09, -2.261673e-09, -2.427374e-09, 
    -2.54129e-09, -2.56744e-09, -2.394339e-09, -2.291235e-09, -2.297871e-09, 
    -2.35436e-09, -2.478854e-09, -2.755889e-09, -3.169331e-09, -3.658712e-09,
  -4.437662e-09, -3.02521e-09, -2.457003e-09, -2.038366e-09, -2.064259e-09, 
    -2.18003e-09, -2.222598e-09, -2.162784e-09, -1.94516e-09, -1.87703e-09, 
    -1.881596e-09, -2.044882e-09, -2.297147e-09, -2.868013e-09, -3.574575e-09,
  -7.533552e-09, -5.388306e-09, -4.048353e-09, -3.195976e-09, -2.303017e-09, 
    -1.846149e-09, -1.69554e-09, -1.78525e-09, -1.773753e-09, -1.730173e-09, 
    -1.788257e-09, -2.063287e-09, -2.461776e-09, -3.143181e-09, -3.882121e-09,
  -1.167211e-08, -8.9625e-09, -6.767521e-09, -5.33808e-09, -4.23539e-09, 
    -3.519886e-09, -2.781791e-09, -2.466977e-09, -2.284295e-09, 
    -2.348252e-09, -2.387408e-09, -2.533804e-09, -2.872671e-09, -3.51601e-09, 
    -4.203267e-09,
  -1.499061e-08, -1.303094e-08, -1.09217e-08, -8.830076e-09, -6.956261e-09, 
    -5.607331e-09, -4.667768e-09, -3.989064e-09, -3.429838e-09, 
    -3.393175e-09, -3.46804e-09, -3.683612e-09, -4.089928e-09, -4.511053e-09, 
    -4.709348e-09,
  -1.618414e-08, -1.509098e-08, -1.385559e-08, -1.264995e-08, -1.100284e-08, 
    -9.23785e-09, -7.628985e-09, -6.372755e-09, -5.582694e-09, -5.115833e-09, 
    -4.591739e-09, -4.420408e-09, -4.466221e-09, -4.593258e-09, -4.832708e-09,
  -1.674137e-08, -1.545802e-08, -1.440554e-08, -1.377484e-08, -1.293243e-08, 
    -1.188271e-08, -1.061086e-08, -9.211161e-09, -8.041182e-09, 
    -6.937669e-09, -6.222994e-09, -5.729846e-09, -5.613591e-09, 
    -5.723014e-09, -5.787742e-09,
  -1.917124e-08, -1.683639e-08, -1.504348e-08, -1.398666e-08, -1.336343e-08, 
    -1.279556e-08, -1.212089e-08, -1.136746e-08, -1.045584e-08, 
    -9.469967e-09, -8.500765e-09, -7.772348e-09, -7.282897e-09, 
    -7.050908e-09, -7.00406e-09,
  -2.186411e-08, -1.999282e-08, -1.785884e-08, -1.572337e-08, -1.406553e-08, 
    -1.318591e-08, -1.265145e-08, -1.218657e-08, -1.174455e-08, -1.13269e-08, 
    -1.072634e-08, -1.004835e-08, -9.382255e-09, -8.816655e-09, -8.447518e-09,
  -2.404178e-08, -2.265428e-08, -2.068717e-08, -1.926026e-08, -1.702626e-08, 
    -1.498099e-08, -1.346211e-08, -1.261451e-08, -1.200953e-08, 
    -1.150576e-08, -1.10219e-08, -1.060116e-08, -1.002565e-08, -9.574084e-09, 
    -9.050312e-09,
  -2.365796e-09, -2.430457e-09, -2.638189e-09, -2.954757e-09, -3.446594e-09, 
    -4.159624e-09, -5.03236e-09, -6.116013e-09, -7.373421e-09, -8.852112e-09, 
    -1.050488e-08, -1.219878e-08, -1.387944e-08, -1.529234e-08, -1.665616e-08,
  -3.073798e-09, -3.16479e-09, -3.396373e-09, -3.676119e-09, -4.180429e-09, 
    -4.946448e-09, -5.936066e-09, -7.182882e-09, -8.516769e-09, 
    -9.909915e-09, -1.127427e-08, -1.267936e-08, -1.416613e-08, 
    -1.563423e-08, -1.703643e-08,
  -4.011043e-09, -4.292604e-09, -4.665438e-09, -5.042224e-09, -5.587917e-09, 
    -6.266239e-09, -7.118492e-09, -8.115199e-09, -9.256348e-09, 
    -1.049866e-08, -1.175237e-08, -1.305689e-08, -1.444043e-08, 
    -1.571205e-08, -1.688193e-08,
  -5.296035e-09, -5.632483e-09, -6.221328e-09, -6.867419e-09, -7.554669e-09, 
    -8.232862e-09, -8.944603e-09, -9.773754e-09, -1.069561e-08, 
    -1.170789e-08, -1.276943e-08, -1.390887e-08, -1.498888e-08, -1.60879e-08, 
    -1.7197e-08,
  -6.966475e-09, -7.120221e-09, -7.618683e-09, -8.166338e-09, -8.864723e-09, 
    -9.62018e-09, -1.040518e-08, -1.119589e-08, -1.193995e-08, -1.275731e-08, 
    -1.365743e-08, -1.459088e-08, -1.547197e-08, -1.646138e-08, -1.750095e-08,
  -8.297212e-09, -8.554747e-09, -8.886998e-09, -9.270364e-09, -9.849327e-09, 
    -1.046719e-08, -1.12024e-08, -1.196203e-08, -1.278194e-08, -1.362569e-08, 
    -1.451782e-08, -1.541619e-08, -1.624722e-08, -1.704657e-08, -1.772358e-08,
  -9.321178e-09, -9.976409e-09, -1.04442e-08, -1.07911e-08, -1.119077e-08, 
    -1.155804e-08, -1.21029e-08, -1.27124e-08, -1.343559e-08, -1.412855e-08, 
    -1.482071e-08, -1.545241e-08, -1.607386e-08, -1.665398e-08, -1.725539e-08,
  -9.973012e-09, -1.050233e-08, -1.099072e-08, -1.154037e-08, -1.201944e-08, 
    -1.245958e-08, -1.293403e-08, -1.343607e-08, -1.404547e-08, 
    -1.465338e-08, -1.531946e-08, -1.595668e-08, -1.656633e-08, 
    -1.716577e-08, -1.772767e-08,
  -1.133878e-08, -1.121265e-08, -1.145613e-08, -1.173461e-08, -1.220006e-08, 
    -1.26973e-08, -1.326758e-08, -1.379159e-08, -1.427598e-08, -1.476969e-08, 
    -1.526181e-08, -1.576842e-08, -1.629695e-08, -1.683001e-08, -1.729389e-08,
  -1.331752e-08, -1.30862e-08, -1.31026e-08, -1.307957e-08, -1.330503e-08, 
    -1.35498e-08, -1.395363e-08, -1.438187e-08, -1.490024e-08, -1.538898e-08, 
    -1.589977e-08, -1.63675e-08, -1.683107e-08, -1.724267e-08, -1.76041e-08,
  -6.649632e-09, -7.831661e-09, -8.887141e-09, -1.035937e-08, -1.162773e-08, 
    -1.302609e-08, -1.445499e-08, -1.577568e-08, -1.674219e-08, 
    -1.745948e-08, -1.807711e-08, -1.853481e-08, -1.891636e-08, 
    -1.938553e-08, -1.97108e-08,
  -8.465686e-09, -9.696905e-09, -1.091913e-08, -1.227236e-08, -1.346343e-08, 
    -1.49462e-08, -1.620552e-08, -1.710021e-08, -1.778735e-08, -1.841185e-08, 
    -1.891882e-08, -1.932576e-08, -1.970731e-08, -1.998881e-08, -2.024979e-08,
  -1.030488e-08, -1.145814e-08, -1.263345e-08, -1.400981e-08, -1.529674e-08, 
    -1.658784e-08, -1.748269e-08, -1.820345e-08, -1.877525e-08, 
    -1.931601e-08, -1.975116e-08, -2.011448e-08, -2.036104e-08, 
    -2.066396e-08, -2.093437e-08,
  -1.190505e-08, -1.296736e-08, -1.422999e-08, -1.55598e-08, -1.663655e-08, 
    -1.762053e-08, -1.826794e-08, -1.886776e-08, -1.942669e-08, 
    -1.998104e-08, -2.036868e-08, -2.072093e-08, -2.10589e-08, -2.140835e-08, 
    -2.165085e-08,
  -1.374556e-08, -1.476502e-08, -1.608059e-08, -1.706423e-08, -1.780296e-08, 
    -1.859926e-08, -1.916726e-08, -1.979302e-08, -2.036127e-08, 
    -2.080209e-08, -2.11762e-08, -2.154328e-08, -2.184789e-08, -2.21212e-08, 
    -2.230018e-08,
  -1.553884e-08, -1.645501e-08, -1.75092e-08, -1.820891e-08, -1.893543e-08, 
    -1.949176e-08, -1.989728e-08, -2.042321e-08, -2.078395e-08, -2.11933e-08, 
    -2.15348e-08, -2.180728e-08, -2.210451e-08, -2.242122e-08, -2.261419e-08,
  -1.628649e-08, -1.717557e-08, -1.787151e-08, -1.845841e-08, -1.905431e-08, 
    -1.95116e-08, -1.999624e-08, -2.044677e-08, -2.079883e-08, -2.119897e-08, 
    -2.14844e-08, -2.182514e-08, -2.219502e-08, -2.243513e-08, -2.257002e-08,
  -1.67352e-08, -1.74108e-08, -1.79812e-08, -1.848049e-08, -1.907923e-08, 
    -1.956561e-08, -2.00943e-08, -2.054325e-08, -2.090846e-08, -2.126206e-08, 
    -2.150026e-08, -2.178575e-08, -2.194054e-08, -2.210961e-08, -2.223197e-08,
  -1.7057e-08, -1.7692e-08, -1.812038e-08, -1.872067e-08, -1.924428e-08, 
    -1.970279e-08, -2.020888e-08, -2.057849e-08, -2.084491e-08, 
    -2.109283e-08, -2.126452e-08, -2.144765e-08, -2.154515e-08, 
    -2.161591e-08, -2.160958e-08,
  -1.789795e-08, -1.845602e-08, -1.876632e-08, -1.93873e-08, -1.970873e-08, 
    -2.011037e-08, -2.046742e-08, -2.077584e-08, -2.089662e-08, 
    -2.106304e-08, -2.112144e-08, -2.116358e-08, -2.113409e-08, 
    -2.114519e-08, -2.116637e-08,
  -9.844918e-09, -1.167896e-08, -1.288655e-08, -1.448107e-08, -1.58102e-08, 
    -1.72024e-08, -1.822472e-08, -1.906939e-08, -1.971288e-08, -2.028557e-08, 
    -2.067623e-08, -2.108591e-08, -2.142127e-08, -2.183866e-08, -2.210371e-08,
  -1.039454e-08, -1.202123e-08, -1.33006e-08, -1.492952e-08, -1.622231e-08, 
    -1.75433e-08, -1.846687e-08, -1.92146e-08, -1.981543e-08, -2.035613e-08, 
    -2.069629e-08, -2.10569e-08, -2.131052e-08, -2.154361e-08, -2.163145e-08,
  -1.088104e-08, -1.240353e-08, -1.373921e-08, -1.533536e-08, -1.655341e-08, 
    -1.77886e-08, -1.850429e-08, -1.923092e-08, -1.982013e-08, -2.032416e-08, 
    -2.060103e-08, -2.092223e-08, -2.101647e-08, -2.109737e-08, -2.105689e-08,
  -1.140338e-08, -1.287246e-08, -1.42254e-08, -1.56932e-08, -1.686406e-08, 
    -1.793208e-08, -1.857182e-08, -1.92947e-08, -1.9856e-08, -2.029197e-08, 
    -2.048656e-08, -2.073744e-08, -2.079082e-08, -2.075038e-08, -2.065457e-08,
  -1.197064e-08, -1.336877e-08, -1.467149e-08, -1.605628e-08, -1.708192e-08, 
    -1.798461e-08, -1.855366e-08, -1.928232e-08, -1.972875e-08, 
    -2.007006e-08, -2.023731e-08, -2.049196e-08, -2.041314e-08, 
    -2.031064e-08, -2.019955e-08,
  -1.259315e-08, -1.394432e-08, -1.519253e-08, -1.637434e-08, -1.719361e-08, 
    -1.79479e-08, -1.845762e-08, -1.917829e-08, -1.956156e-08, -1.985057e-08, 
    -2.000972e-08, -2.018214e-08, -2.00469e-08, -1.994893e-08, -1.994199e-08,
  -1.330007e-08, -1.456047e-08, -1.564793e-08, -1.661164e-08, -1.730235e-08, 
    -1.796841e-08, -1.84968e-08, -1.916045e-08, -1.939776e-08, -1.955094e-08, 
    -1.964504e-08, -1.973652e-08, -1.947155e-08, -1.944478e-08, -1.957898e-08,
  -1.399206e-08, -1.506365e-08, -1.594484e-08, -1.678664e-08, -1.73693e-08, 
    -1.794926e-08, -1.83969e-08, -1.890286e-08, -1.905983e-08, -1.919576e-08, 
    -1.925388e-08, -1.926292e-08, -1.905075e-08, -1.914736e-08, -1.945289e-08,
  -1.444055e-08, -1.536986e-08, -1.617085e-08, -1.687958e-08, -1.734965e-08, 
    -1.787781e-08, -1.835161e-08, -1.882046e-08, -1.886392e-08, 
    -1.889568e-08, -1.887308e-08, -1.885929e-08, -1.875408e-08, 
    -1.893275e-08, -1.935018e-08,
  -1.489309e-08, -1.568978e-08, -1.638439e-08, -1.698293e-08, -1.745137e-08, 
    -1.79741e-08, -1.84055e-08, -1.87157e-08, -1.879873e-08, -1.895397e-08, 
    -1.903996e-08, -1.897611e-08, -1.894911e-08, -1.932568e-08, -1.986979e-08,
  -1.559251e-08, -1.711698e-08, -1.819081e-08, -1.944465e-08, -2.022427e-08, 
    -2.085112e-08, -2.108298e-08, -2.125293e-08, -2.127065e-08, 
    -2.153149e-08, -2.188125e-08, -2.230835e-08, -2.271904e-08, -2.33137e-08, 
    -2.385152e-08,
  -1.583871e-08, -1.738473e-08, -1.850977e-08, -1.975701e-08, -2.047653e-08, 
    -2.112731e-08, -2.131221e-08, -2.151386e-08, -2.168512e-08, 
    -2.208825e-08, -2.248624e-08, -2.291637e-08, -2.334656e-08, 
    -2.390343e-08, -2.442548e-08,
  -1.616523e-08, -1.76951e-08, -1.889721e-08, -2.009443e-08, -2.082391e-08, 
    -2.136735e-08, -2.145335e-08, -2.18307e-08, -2.215331e-08, -2.256338e-08, 
    -2.28375e-08, -2.317709e-08, -2.359724e-08, -2.40396e-08, -2.455954e-08,
  -1.644296e-08, -1.799467e-08, -1.924271e-08, -2.042668e-08, -2.10435e-08, 
    -2.143952e-08, -2.166078e-08, -2.233455e-08, -2.272592e-08, 
    -2.312121e-08, -2.326088e-08, -2.358948e-08, -2.386104e-08, 
    -2.410324e-08, -2.453095e-08,
  -1.672344e-08, -1.834393e-08, -1.967132e-08, -2.071537e-08, -2.117664e-08, 
    -2.151877e-08, -2.190899e-08, -2.275045e-08, -2.314132e-08, 
    -2.357697e-08, -2.364636e-08, -2.391645e-08, -2.401529e-08, 
    -2.418551e-08, -2.439761e-08,
  -1.701103e-08, -1.866127e-08, -1.993543e-08, -2.088905e-08, -2.118555e-08, 
    -2.151937e-08, -2.218376e-08, -2.300876e-08, -2.344686e-08, 
    -2.398209e-08, -2.403117e-08, -2.427204e-08, -2.429035e-08, 
    -2.437377e-08, -2.451857e-08,
  -1.728634e-08, -1.894191e-08, -2.019359e-08, -2.100455e-08, -2.124004e-08, 
    -2.1684e-08, -2.241841e-08, -2.312075e-08, -2.359402e-08, -2.411077e-08, 
    -2.420724e-08, -2.453763e-08, -2.454769e-08, -2.457409e-08, -2.463327e-08,
  -1.750871e-08, -1.914973e-08, -2.034955e-08, -2.106609e-08, -2.130785e-08, 
    -2.18578e-08, -2.268987e-08, -2.330696e-08, -2.378275e-08, -2.418466e-08, 
    -2.428689e-08, -2.45521e-08, -2.457293e-08, -2.469403e-08, -2.478793e-08,
  -1.767657e-08, -1.929288e-08, -2.046207e-08, -2.115388e-08, -2.146208e-08, 
    -2.214086e-08, -2.284257e-08, -2.340398e-08, -2.371151e-08, 
    -2.401106e-08, -2.403697e-08, -2.422478e-08, -2.413415e-08, 
    -2.422135e-08, -2.43702e-08,
  -1.782833e-08, -1.94014e-08, -2.052866e-08, -2.120013e-08, -2.156228e-08, 
    -2.228892e-08, -2.281947e-08, -2.331395e-08, -2.351709e-08, 
    -2.366199e-08, -2.354283e-08, -2.350435e-08, -2.321046e-08, 
    -2.317961e-08, -2.327089e-08,
  -1.729185e-08, -1.849151e-08, -1.895233e-08, -1.95671e-08, -1.965781e-08, 
    -1.98787e-08, -1.989662e-08, -2.005906e-08, -2.002804e-08, -2.031416e-08, 
    -2.09111e-08, -2.197303e-08, -2.306798e-08, -2.400478e-08, -2.487604e-08,
  -1.766326e-08, -1.86958e-08, -1.90812e-08, -1.964194e-08, -1.96814e-08, 
    -1.987253e-08, -1.984332e-08, -1.996425e-08, -2.001405e-08, 
    -2.030197e-08, -2.085005e-08, -2.1914e-08, -2.306358e-08, -2.415898e-08, 
    -2.517284e-08,
  -1.800232e-08, -1.887681e-08, -1.92734e-08, -1.975252e-08, -1.973916e-08, 
    -1.992053e-08, -1.985521e-08, -1.996535e-08, -2.000648e-08, 
    -2.027251e-08, -2.079805e-08, -2.18624e-08, -2.299047e-08, -2.420721e-08, 
    -2.524871e-08,
  -1.831202e-08, -1.908387e-08, -1.942415e-08, -1.98045e-08, -1.974841e-08, 
    -1.991521e-08, -1.987975e-08, -1.998488e-08, -2.001508e-08, 
    -2.026458e-08, -2.066993e-08, -2.160088e-08, -2.269206e-08, 
    -2.397536e-08, -2.520806e-08,
  -1.859587e-08, -1.922392e-08, -1.951429e-08, -1.982776e-08, -1.977425e-08, 
    -1.996165e-08, -1.988552e-08, -2.00296e-08, -2.007983e-08, -2.029616e-08, 
    -2.052778e-08, -2.132248e-08, -2.230748e-08, -2.357884e-08, -2.500964e-08,
  -1.881975e-08, -1.935476e-08, -1.961842e-08, -1.986709e-08, -1.977707e-08, 
    -1.994079e-08, -1.989661e-08, -2.009257e-08, -2.016404e-08, 
    -2.037418e-08, -2.059495e-08, -2.117674e-08, -2.196997e-08, -2.31466e-08, 
    -2.450425e-08,
  -1.90395e-08, -1.949964e-08, -1.970565e-08, -1.987973e-08, -1.974389e-08, 
    -1.987531e-08, -1.981526e-08, -2.003903e-08, -2.01286e-08, -2.036317e-08, 
    -2.054245e-08, -2.104325e-08, -2.174304e-08, -2.277415e-08, -2.405507e-08,
  -1.921537e-08, -1.961831e-08, -1.977058e-08, -1.989611e-08, -1.973585e-08, 
    -1.985296e-08, -1.982408e-08, -2.005064e-08, -2.015378e-08, 
    -2.044489e-08, -2.06661e-08, -2.111117e-08, -2.1654e-08, -2.251689e-08, 
    -2.358551e-08,
  -1.935737e-08, -1.974831e-08, -1.991238e-08, -1.994896e-08, -1.976018e-08, 
    -1.989092e-08, -1.992446e-08, -2.015795e-08, -2.0349e-08, -2.057584e-08, 
    -2.078094e-08, -2.118722e-08, -2.16462e-08, -2.235934e-08, -2.330662e-08,
  -1.948424e-08, -1.987974e-08, -2.003312e-08, -2.002071e-08, -1.987466e-08, 
    -2.023624e-08, -2.035073e-08, -2.06467e-08, -2.086253e-08, -2.109938e-08, 
    -2.131954e-08, -2.163259e-08, -2.193308e-08, -2.253614e-08, -2.327001e-08,
  -1.750226e-08, -1.951522e-08, -1.983392e-08, -2.063594e-08, -2.123542e-08, 
    -2.162113e-08, -2.236865e-08, -2.346372e-08, -2.326531e-08, 
    -2.306679e-08, -2.342293e-08, -2.482479e-08, -2.549711e-08, 
    -2.550368e-08, -2.554622e-08,
  -1.785708e-08, -1.969035e-08, -2.011715e-08, -2.091204e-08, -2.150895e-08, 
    -2.184877e-08, -2.263778e-08, -2.339883e-08, -2.299405e-08, 
    -2.342669e-08, -2.457442e-08, -2.567329e-08, -2.624097e-08, 
    -2.646912e-08, -2.661557e-08,
  -1.814606e-08, -1.975924e-08, -2.032995e-08, -2.106671e-08, -2.166277e-08, 
    -2.202439e-08, -2.267354e-08, -2.329746e-08, -2.299593e-08, 
    -2.376408e-08, -2.477315e-08, -2.563411e-08, -2.582475e-08, 
    -2.624805e-08, -2.628328e-08,
  -1.824501e-08, -1.974946e-08, -2.048412e-08, -2.116295e-08, -2.171778e-08, 
    -2.206895e-08, -2.277594e-08, -2.329686e-08, -2.296122e-08, 
    -2.388186e-08, -2.49127e-08, -2.546902e-08, -2.568558e-08, -2.595061e-08, 
    -2.601686e-08,
  -1.841793e-08, -1.975783e-08, -2.065187e-08, -2.123148e-08, -2.168127e-08, 
    -2.200972e-08, -2.259011e-08, -2.306149e-08, -2.291822e-08, 
    -2.398387e-08, -2.491779e-08, -2.536177e-08, -2.555934e-08, 
    -2.574795e-08, -2.591764e-08,
  -1.850957e-08, -1.984579e-08, -2.088709e-08, -2.129633e-08, -2.163694e-08, 
    -2.19513e-08, -2.23875e-08, -2.280796e-08, -2.279345e-08, -2.381516e-08, 
    -2.481857e-08, -2.528727e-08, -2.552694e-08, -2.604878e-08, -2.619537e-08,
  -1.85616e-08, -2.001753e-08, -2.122567e-08, -2.147212e-08, -2.163813e-08, 
    -2.190927e-08, -2.221467e-08, -2.265794e-08, -2.268073e-08, 
    -2.363895e-08, -2.472456e-08, -2.524052e-08, -2.549465e-08, 
    -2.604283e-08, -2.619776e-08,
  -1.857095e-08, -2.009159e-08, -2.160064e-08, -2.170971e-08, -2.170332e-08, 
    -2.190609e-08, -2.202061e-08, -2.236479e-08, -2.256723e-08, 
    -2.340829e-08, -2.44919e-08, -2.511607e-08, -2.53441e-08, -2.588305e-08, 
    -2.59736e-08,
  -1.844611e-08, -2.003388e-08, -2.189087e-08, -2.190529e-08, -2.174279e-08, 
    -2.190039e-08, -2.185589e-08, -2.218542e-08, -2.24117e-08, -2.30759e-08, 
    -2.420288e-08, -2.496222e-08, -2.510071e-08, -2.557201e-08, -2.581357e-08,
  -1.817565e-08, -1.984528e-08, -2.208657e-08, -2.197873e-08, -2.171927e-08, 
    -2.17966e-08, -2.175144e-08, -2.202119e-08, -2.221593e-08, -2.283621e-08, 
    -2.381913e-08, -2.467434e-08, -2.480544e-08, -2.516816e-08, -2.568303e-08,
  -1.255694e-08, -1.699512e-08, -2.028567e-08, -2.337722e-08, -2.332134e-08, 
    -2.218762e-08, -2.095953e-08, -2.057315e-08, -2.02155e-08, -1.987176e-08, 
    -1.959189e-08, -2.076541e-08, -2.166482e-08, -2.221488e-08, -2.24406e-08,
  -1.312977e-08, -1.805653e-08, -2.087727e-08, -2.413157e-08, -2.385021e-08, 
    -2.241619e-08, -2.133628e-08, -2.075778e-08, -1.998028e-08, 
    -1.973499e-08, -2.042988e-08, -2.172027e-08, -2.200065e-08, 
    -2.228985e-08, -2.264271e-08,
  -1.344279e-08, -1.858072e-08, -2.15845e-08, -2.500468e-08, -2.459159e-08, 
    -2.282316e-08, -2.157138e-08, -2.090981e-08, -1.992534e-08, 
    -2.054906e-08, -2.174714e-08, -2.249378e-08, -2.291612e-08, 
    -2.329758e-08, -2.348591e-08,
  -1.376459e-08, -1.884945e-08, -2.225718e-08, -2.593714e-08, -2.548639e-08, 
    -2.317336e-08, -2.184201e-08, -2.094121e-08, -2.034753e-08, 
    -2.174716e-08, -2.237762e-08, -2.292979e-08, -2.358414e-08, 
    -2.389414e-08, -2.415172e-08,
  -1.405343e-08, -1.915867e-08, -2.288396e-08, -2.685268e-08, -2.6144e-08, 
    -2.35063e-08, -2.207672e-08, -2.120771e-08, -2.119381e-08, -2.28169e-08, 
    -2.306208e-08, -2.376225e-08, -2.430516e-08, -2.470449e-08, -2.517805e-08,
  -1.440992e-08, -1.942707e-08, -2.317691e-08, -2.727531e-08, -2.676768e-08, 
    -2.356429e-08, -2.223802e-08, -2.145558e-08, -2.228618e-08, 
    -2.357291e-08, -2.375768e-08, -2.447343e-08, -2.479087e-08, 
    -2.508811e-08, -2.548114e-08,
  -1.470346e-08, -1.978981e-08, -2.310588e-08, -2.747112e-08, -2.709418e-08, 
    -2.355669e-08, -2.236012e-08, -2.183463e-08, -2.309947e-08, 
    -2.419435e-08, -2.445754e-08, -2.488409e-08, -2.502034e-08, 
    -2.532095e-08, -2.563844e-08,
  -1.511115e-08, -1.997411e-08, -2.288526e-08, -2.747873e-08, -2.733333e-08, 
    -2.338025e-08, -2.245004e-08, -2.217063e-08, -2.371509e-08, 
    -2.467993e-08, -2.489986e-08, -2.496062e-08, -2.499973e-08, 
    -2.531045e-08, -2.552268e-08,
  -1.554527e-08, -1.991627e-08, -2.262803e-08, -2.770315e-08, -2.747607e-08, 
    -2.319564e-08, -2.240437e-08, -2.24398e-08, -2.416351e-08, -2.497312e-08, 
    -2.49683e-08, -2.514396e-08, -2.500512e-08, -2.545042e-08, -2.538675e-08,
  -1.617131e-08, -1.973837e-08, -2.271371e-08, -2.804693e-08, -2.753171e-08, 
    -2.296266e-08, -2.23708e-08, -2.266098e-08, -2.427057e-08, -2.499637e-08, 
    -2.521155e-08, -2.542652e-08, -2.542483e-08, -2.553628e-08, -2.553082e-08,
  -9.281575e-09, -1.162519e-08, -1.403922e-08, -1.793353e-08, -2.172568e-08, 
    -2.438142e-08, -2.481181e-08, -2.356209e-08, -2.243538e-08, 
    -2.334625e-08, -2.35728e-08, -2.43226e-08, -2.477431e-08, -2.41267e-08, 
    -2.41985e-08,
  -9.091555e-09, -1.179376e-08, -1.367533e-08, -1.711707e-08, -2.109778e-08, 
    -2.44064e-08, -2.521358e-08, -2.361613e-08, -2.252657e-08, -2.345677e-08, 
    -2.324534e-08, -2.428433e-08, -2.500645e-08, -2.489276e-08, -2.499376e-08,
  -8.943059e-09, -1.198151e-08, -1.389698e-08, -1.690269e-08, -2.087536e-08, 
    -2.470249e-08, -2.552677e-08, -2.360564e-08, -2.263399e-08, -2.36274e-08, 
    -2.351368e-08, -2.521957e-08, -2.571583e-08, -2.582325e-08, -2.565457e-08,
  -9.074899e-09, -1.202475e-08, -1.436875e-08, -1.729977e-08, -2.109235e-08, 
    -2.527685e-08, -2.565768e-08, -2.353428e-08, -2.268104e-08, 
    -2.390999e-08, -2.39589e-08, -2.578551e-08, -2.575153e-08, -2.656736e-08, 
    -2.653439e-08,
  -9.362902e-09, -1.234897e-08, -1.50482e-08, -1.795546e-08, -2.148454e-08, 
    -2.577249e-08, -2.574949e-08, -2.347145e-08, -2.287242e-08, 
    -2.411326e-08, -2.416296e-08, -2.606489e-08, -2.600324e-08, 
    -2.686068e-08, -2.708565e-08,
  -9.564551e-09, -1.290781e-08, -1.590303e-08, -1.909831e-08, -2.246078e-08, 
    -2.616301e-08, -2.583273e-08, -2.338067e-08, -2.328467e-08, 
    -2.437879e-08, -2.469803e-08, -2.640984e-08, -2.644532e-08, 
    -2.723016e-08, -2.744993e-08,
  -1.001126e-08, -1.377578e-08, -1.678915e-08, -2.015469e-08, -2.407399e-08, 
    -2.644177e-08, -2.602123e-08, -2.348434e-08, -2.403836e-08, 
    -2.441345e-08, -2.568401e-08, -2.705729e-08, -2.675874e-08, 
    -2.747448e-08, -2.731809e-08,
  -1.077974e-08, -1.453889e-08, -1.745345e-08, -2.161364e-08, -2.519309e-08, 
    -2.720117e-08, -2.669615e-08, -2.353226e-08, -2.484806e-08, 
    -2.483906e-08, -2.714201e-08, -2.707431e-08, -2.729211e-08, 
    -2.758725e-08, -2.722373e-08,
  -1.162133e-08, -1.524628e-08, -1.880587e-08, -2.306639e-08, -2.652196e-08, 
    -2.895434e-08, -2.681296e-08, -2.383039e-08, -2.541844e-08, 
    -2.533747e-08, -2.753832e-08, -2.719823e-08, -2.777778e-08, 
    -2.757288e-08, -2.75904e-08,
  -1.254468e-08, -1.637919e-08, -2.039971e-08, -2.483434e-08, -2.866063e-08, 
    -3.052064e-08, -2.692346e-08, -2.425508e-08, -2.535048e-08, 
    -2.618564e-08, -2.756384e-08, -2.769024e-08, -2.801929e-08, 
    -2.785928e-08, -2.786989e-08,
  -1.63666e-08, -1.860944e-08, -2.080976e-08, -2.315575e-08, -2.336498e-08, 
    -2.317427e-08, -2.332953e-08, -2.345305e-08, -2.438472e-08, 
    -2.551835e-08, -2.500908e-08, -2.483232e-08, -2.393376e-08, -2.34142e-08, 
    -2.293985e-08,
  -1.459952e-08, -1.767738e-08, -2.007775e-08, -2.279077e-08, -2.357388e-08, 
    -2.3194e-08, -2.340201e-08, -2.395486e-08, -2.45435e-08, -2.582739e-08, 
    -2.575676e-08, -2.55423e-08, -2.506038e-08, -2.484893e-08, -2.472105e-08,
  -1.293607e-08, -1.649975e-08, -1.939772e-08, -2.245592e-08, -2.38308e-08, 
    -2.313538e-08, -2.343264e-08, -2.414545e-08, -2.445235e-08, 
    -2.624668e-08, -2.631787e-08, -2.601065e-08, -2.56066e-08, -2.556754e-08, 
    -2.573152e-08,
  -1.16353e-08, -1.537375e-08, -1.877254e-08, -2.21693e-08, -2.419056e-08, 
    -2.328208e-08, -2.320104e-08, -2.401171e-08, -2.446768e-08, 
    -2.625744e-08, -2.632661e-08, -2.598656e-08, -2.568809e-08, 
    -2.580938e-08, -2.604312e-08,
  -1.085295e-08, -1.427133e-08, -1.819444e-08, -2.200872e-08, -2.46141e-08, 
    -2.371314e-08, -2.32558e-08, -2.372428e-08, -2.420307e-08, -2.628899e-08, 
    -2.614081e-08, -2.651321e-08, -2.624681e-08, -2.663551e-08, -2.695303e-08,
  -1.043007e-08, -1.336814e-08, -1.75539e-08, -2.180845e-08, -2.509626e-08, 
    -2.428804e-08, -2.333362e-08, -2.354532e-08, -2.434884e-08, 
    -2.594618e-08, -2.643692e-08, -2.701139e-08, -2.6821e-08, -2.739802e-08, 
    -2.781172e-08,
  -1.012423e-08, -1.267649e-08, -1.703524e-08, -2.155597e-08, -2.559348e-08, 
    -2.484375e-08, -2.361337e-08, -2.345012e-08, -2.420929e-08, 
    -2.566349e-08, -2.662227e-08, -2.724299e-08, -2.727164e-08, 
    -2.772179e-08, -2.846208e-08,
  -9.980643e-09, -1.230369e-08, -1.66089e-08, -2.151312e-08, -2.62025e-08, 
    -2.538417e-08, -2.378098e-08, -2.352678e-08, -2.411778e-08, -2.53922e-08, 
    -2.679819e-08, -2.719216e-08, -2.74554e-08, -2.773103e-08, -2.849597e-08,
  -9.750885e-09, -1.21202e-08, -1.645604e-08, -2.17439e-08, -2.698974e-08, 
    -2.562848e-08, -2.397438e-08, -2.36721e-08, -2.418805e-08, -2.544377e-08, 
    -2.702317e-08, -2.709909e-08, -2.760228e-08, -2.774817e-08, -2.838344e-08,
  -9.689928e-09, -1.226752e-08, -1.654867e-08, -2.273105e-08, -2.794543e-08, 
    -2.586645e-08, -2.430999e-08, -2.378811e-08, -2.452502e-08, 
    -2.576537e-08, -2.698963e-08, -2.717918e-08, -2.757099e-08, 
    -2.765016e-08, -2.839214e-08,
  -1.827149e-08, -1.84027e-08, -1.834388e-08, -1.784087e-08, -1.69365e-08, 
    -1.591831e-08, -1.507377e-08, -1.439679e-08, -1.37445e-08, -1.275686e-08, 
    -1.191845e-08, -1.106394e-08, -1.016173e-08, -9.320034e-09, -8.654919e-09,
  -1.76811e-08, -1.797489e-08, -1.803514e-08, -1.797337e-08, -1.748692e-08, 
    -1.676193e-08, -1.610052e-08, -1.555959e-08, -1.488629e-08, 
    -1.397046e-08, -1.307553e-08, -1.233205e-08, -1.148601e-08, 
    -1.059678e-08, -9.809179e-09,
  -1.777896e-08, -1.7843e-08, -1.811781e-08, -1.817761e-08, -1.793572e-08, 
    -1.758768e-08, -1.717345e-08, -1.663849e-08, -1.596175e-08, 
    -1.517776e-08, -1.431227e-08, -1.355563e-08, -1.286822e-08, 
    -1.217177e-08, -1.13921e-08,
  -1.806657e-08, -1.786973e-08, -1.823649e-08, -1.863833e-08, -1.851499e-08, 
    -1.829875e-08, -1.793717e-08, -1.743112e-08, -1.684283e-08, 
    -1.606061e-08, -1.523316e-08, -1.435558e-08, -1.370978e-08, 
    -1.316567e-08, -1.262162e-08,
  -1.852821e-08, -1.809147e-08, -1.844331e-08, -1.911886e-08, -1.917433e-08, 
    -1.894556e-08, -1.870016e-08, -1.845859e-08, -1.797628e-08, 
    -1.745775e-08, -1.672348e-08, -1.586497e-08, -1.49997e-08, -1.429657e-08, 
    -1.376399e-08,
  -1.915696e-08, -1.869786e-08, -1.878672e-08, -1.963101e-08, -1.974805e-08, 
    -1.96893e-08, -1.952023e-08, -1.953735e-08, -1.928443e-08, -1.880955e-08, 
    -1.816105e-08, -1.729104e-08, -1.636947e-08, -1.550264e-08, -1.488834e-08,
  -1.980202e-08, -1.942137e-08, -1.921055e-08, -1.991577e-08, -2.016556e-08, 
    -2.036566e-08, -2.053976e-08, -2.088322e-08, -2.080456e-08, 
    -2.035255e-08, -1.977204e-08, -1.896719e-08, -1.795953e-08, 
    -1.699659e-08, -1.609019e-08,
  -2.021945e-08, -1.996167e-08, -1.968702e-08, -2.031044e-08, -2.076614e-08, 
    -2.102634e-08, -2.144313e-08, -2.174327e-08, -2.203205e-08, 
    -2.166459e-08, -2.096492e-08, -2.030643e-08, -1.944054e-08, 
    -1.856567e-08, -1.769271e-08,
  -2.032258e-08, -2.039047e-08, -2.021278e-08, -2.084158e-08, -2.141823e-08, 
    -2.161469e-08, -2.178795e-08, -2.212014e-08, -2.260973e-08, 
    -2.255434e-08, -2.18487e-08, -2.117653e-08, -2.03729e-08, -1.952863e-08, 
    -1.876131e-08,
  -2.044939e-08, -2.080152e-08, -2.079164e-08, -2.146235e-08, -2.209742e-08, 
    -2.21625e-08, -2.20281e-08, -2.2192e-08, -2.272394e-08, -2.298789e-08, 
    -2.252343e-08, -2.185348e-08, -2.105294e-08, -2.017615e-08, -1.943244e-08,
  -1.120998e-08, -9.947639e-09, -9.078742e-09, -8.249467e-09, -7.808837e-09, 
    -7.252304e-09, -6.815598e-09, -6.543671e-09, -6.396721e-09, 
    -6.269578e-09, -6.172899e-09, -6.230496e-09, -6.657596e-09, 
    -7.469525e-09, -8.484339e-09,
  -1.199475e-08, -1.08371e-08, -9.99324e-09, -8.979957e-09, -8.195353e-09, 
    -7.703985e-09, -7.100792e-09, -6.845474e-09, -6.694361e-09, 
    -6.721173e-09, -6.591468e-09, -6.494714e-09, -6.674065e-09, 
    -7.300877e-09, -8.326013e-09,
  -1.24521e-08, -1.141969e-08, -1.046376e-08, -9.625201e-09, -8.613549e-09, 
    -8.120397e-09, -7.392746e-09, -7.026617e-09, -6.823126e-09, 
    -6.743692e-09, -6.72967e-09, -6.792402e-09, -6.951355e-09, -7.510741e-09, 
    -8.259485e-09,
  -1.309408e-08, -1.220871e-08, -1.107614e-08, -1.011176e-08, -9.11165e-09, 
    -8.570893e-09, -7.993006e-09, -7.48068e-09, -7.266745e-09, -6.978483e-09, 
    -6.945054e-09, -7.137651e-09, -7.500686e-09, -8.007815e-09, -8.661071e-09,
  -1.338019e-08, -1.28307e-08, -1.164822e-08, -1.057029e-08, -9.437365e-09, 
    -8.540296e-09, -8.084608e-09, -7.728295e-09, -7.595201e-09, 
    -7.458572e-09, -7.430657e-09, -7.614448e-09, -8.00658e-09, -8.502301e-09, 
    -9.048794e-09,
  -1.385838e-08, -1.350891e-08, -1.248493e-08, -1.136072e-08, -1.025214e-08, 
    -9.147588e-09, -8.245605e-09, -7.779076e-09, -7.639312e-09, 
    -7.594698e-09, -7.698883e-09, -7.884402e-09, -8.373347e-09, 
    -8.852391e-09, -9.435e-09,
  -1.406436e-08, -1.380751e-08, -1.308348e-08, -1.200964e-08, -1.109181e-08, 
    -1.006721e-08, -9.025751e-09, -8.181325e-09, -7.740033e-09, 
    -7.628294e-09, -7.697961e-09, -7.92152e-09, -8.33004e-09, -8.935733e-09, 
    -9.681377e-09,
  -1.422117e-08, -1.38495e-08, -1.331971e-08, -1.248636e-08, -1.175244e-08, 
    -1.097454e-08, -9.939146e-09, -9.095559e-09, -8.39552e-09, -8.011583e-09, 
    -7.932091e-09, -8.062028e-09, -8.382827e-09, -8.893244e-09, -9.576307e-09,
  -1.44155e-08, -1.390587e-08, -1.342984e-08, -1.267028e-08, -1.216312e-08, 
    -1.165507e-08, -1.078858e-08, -9.927268e-09, -9.182773e-09, 
    -8.657828e-09, -8.435952e-09, -8.55104e-09, -8.877905e-09, -9.326661e-09, 
    -9.803462e-09,
  -1.430693e-08, -1.38783e-08, -1.334113e-08, -1.253523e-08, -1.225867e-08, 
    -1.207131e-08, -1.167708e-08, -1.094395e-08, -1.016166e-08, 
    -9.540646e-09, -9.21726e-09, -9.225251e-09, -9.501638e-09, -9.80449e-09, 
    -1.005884e-08,
  -5.739188e-09, -5.506595e-09, -5.275874e-09, -5.249856e-09, -5.33204e-09, 
    -5.50255e-09, -5.818935e-09, -6.287154e-09, -6.902624e-09, -7.621377e-09, 
    -8.480722e-09, -9.433937e-09, -1.072433e-08, -1.21959e-08, -1.386415e-08,
  -6.114133e-09, -5.828931e-09, -5.604499e-09, -5.463901e-09, -5.558062e-09, 
    -5.735882e-09, -6.057389e-09, -6.519718e-09, -7.168949e-09, 
    -7.877853e-09, -8.834014e-09, -9.838481e-09, -1.112452e-08, 
    -1.254681e-08, -1.421425e-08,
  -6.368976e-09, -6.12788e-09, -5.944861e-09, -5.701258e-09, -5.7788e-09, 
    -5.930484e-09, -6.249825e-09, -6.738987e-09, -7.366314e-09, 
    -8.103743e-09, -9.127928e-09, -1.017712e-08, -1.146413e-08, 
    -1.285865e-08, -1.444674e-08,
  -6.447451e-09, -6.360132e-09, -6.266315e-09, -6.022701e-09, -5.99396e-09, 
    -6.110213e-09, -6.430751e-09, -6.970032e-09, -7.611894e-09, 
    -8.329433e-09, -9.340737e-09, -1.046479e-08, -1.172166e-08, 
    -1.304204e-08, -1.46035e-08,
  -6.403057e-09, -6.506333e-09, -6.493357e-09, -6.371515e-09, -6.21628e-09, 
    -6.32387e-09, -6.672552e-09, -7.245418e-09, -7.92165e-09, -8.618643e-09, 
    -9.630594e-09, -1.077071e-08, -1.199827e-08, -1.324696e-08, -1.477902e-08,
  -6.40959e-09, -6.607798e-09, -6.667318e-09, -6.621759e-09, -6.460021e-09, 
    -6.602769e-09, -6.954497e-09, -7.545272e-09, -8.225137e-09, 
    -8.945301e-09, -9.988855e-09, -1.111968e-08, -1.227155e-08, 
    -1.346155e-08, -1.499853e-08,
  -6.312414e-09, -6.660084e-09, -6.839568e-09, -6.896973e-09, -6.756846e-09, 
    -6.861091e-09, -7.24319e-09, -7.829347e-09, -8.566651e-09, -9.350078e-09, 
    -1.044382e-08, -1.152273e-08, -1.259575e-08, -1.371068e-08, -1.524072e-08,
  -6.320615e-09, -6.688408e-09, -6.995796e-09, -7.019337e-09, -7.024429e-09, 
    -7.124004e-09, -7.525309e-09, -8.124013e-09, -8.928888e-09, 
    -9.805508e-09, -1.095702e-08, -1.192516e-08, -1.283935e-08, 
    -1.400474e-08, -1.554114e-08,
  -6.494452e-09, -6.756756e-09, -7.083387e-09, -7.208695e-09, -7.321719e-09, 
    -7.461732e-09, -7.848274e-09, -8.491656e-09, -9.348904e-09, 
    -1.036585e-08, -1.15118e-08, -1.235154e-08, -1.312634e-08, -1.437032e-08, 
    -1.575967e-08,
  -6.67104e-09, -6.903806e-09, -7.237152e-09, -7.46544e-09, -7.635879e-09, 
    -7.838814e-09, -8.186868e-09, -8.902042e-09, -9.826177e-09, 
    -1.096699e-08, -1.209308e-08, -1.280957e-08, -1.352477e-08, 
    -1.479406e-08, -1.599667e-08,
  -6.637292e-09, -7.155883e-09, -7.510709e-09, -7.948526e-09, -8.23422e-09, 
    -8.52109e-09, -8.650954e-09, -8.570446e-09, -8.655552e-09, -9.117636e-09, 
    -1.027804e-08, -1.334186e-08, -1.715233e-08, -2.025247e-08, -2.255834e-08,
  -6.793957e-09, -7.288659e-09, -7.70822e-09, -8.052484e-09, -8.294041e-09, 
    -8.476747e-09, -8.532522e-09, -8.531588e-09, -8.830306e-09, 
    -9.608973e-09, -1.156148e-08, -1.536393e-08, -1.885119e-08, 
    -2.145449e-08, -2.346099e-08,
  -6.813389e-09, -7.261388e-09, -7.601385e-09, -7.879338e-09, -8.083807e-09, 
    -8.260182e-09, -8.295916e-09, -8.459917e-09, -8.938994e-09, 
    -1.019894e-08, -1.295088e-08, -1.683805e-08, -1.978957e-08, 
    -2.223748e-08, -2.386321e-08,
  -6.736811e-09, -7.16912e-09, -7.433036e-09, -7.647265e-09, -7.837855e-09, 
    -8.017484e-09, -8.111928e-09, -8.411581e-09, -9.100853e-09, 
    -1.088678e-08, -1.409313e-08, -1.76381e-08, -2.034719e-08, -2.266168e-08, 
    -2.402832e-08,
  -6.678705e-09, -7.071522e-09, -7.324999e-09, -7.473084e-09, -7.655524e-09, 
    -7.822946e-09, -8.011279e-09, -8.409964e-09, -9.320416e-09, 
    -1.154267e-08, -1.492343e-08, -1.810574e-08, -2.066939e-08, 
    -2.283647e-08, -2.396035e-08,
  -6.630919e-09, -6.956019e-09, -7.232714e-09, -7.384391e-09, -7.57369e-09, 
    -7.716954e-09, -7.972337e-09, -8.449812e-09, -9.58414e-09, -1.208492e-08, 
    -1.544181e-08, -1.834521e-08, -2.07518e-08, -2.277884e-08, -2.373988e-08,
  -6.621701e-09, -6.898055e-09, -7.174736e-09, -7.330569e-09, -7.533088e-09, 
    -7.645428e-09, -7.956009e-09, -8.512597e-09, -9.835712e-09, 
    -1.252133e-08, -1.578064e-08, -1.847884e-08, -2.071696e-08, 
    -2.259332e-08, -2.35181e-08,
  -6.61254e-09, -6.870545e-09, -7.145986e-09, -7.301715e-09, -7.515525e-09, 
    -7.615435e-09, -7.974865e-09, -8.617309e-09, -1.007851e-08, 
    -1.284258e-08, -1.601263e-08, -1.853651e-08, -2.062723e-08, 
    -2.238487e-08, -2.331926e-08,
  -6.634372e-09, -6.891071e-09, -7.175102e-09, -7.319371e-09, -7.537372e-09, 
    -7.645756e-09, -8.040368e-09, -8.727318e-09, -1.028962e-08, -1.31045e-08, 
    -1.615106e-08, -1.852478e-08, -2.05269e-08, -2.22025e-08, -2.311946e-08,
  -6.6839e-09, -6.934005e-09, -7.217069e-09, -7.37356e-09, -7.583724e-09, 
    -7.711022e-09, -8.138532e-09, -8.847091e-09, -1.049046e-08, 
    -1.329858e-08, -1.621532e-08, -1.848874e-08, -2.043398e-08, 
    -2.207398e-08, -2.292143e-08,
  -1.282545e-08, -1.379658e-08, -1.408656e-08, -1.476762e-08, -1.529978e-08, 
    -1.580452e-08, -1.579154e-08, -1.533015e-08, -1.540944e-08, 
    -1.580369e-08, -1.642678e-08, -1.775824e-08, -1.953696e-08, 
    -2.115724e-08, -2.269434e-08,
  -1.341347e-08, -1.39727e-08, -1.441738e-08, -1.51861e-08, -1.56533e-08, 
    -1.593387e-08, -1.57438e-08, -1.563553e-08, -1.595745e-08, -1.668914e-08, 
    -1.852088e-08, -2.078625e-08, -2.252997e-08, -2.363603e-08, -2.458314e-08,
  -1.357932e-08, -1.410082e-08, -1.481811e-08, -1.555656e-08, -1.58062e-08, 
    -1.594404e-08, -1.564783e-08, -1.585374e-08, -1.659673e-08, -1.87874e-08, 
    -2.14385e-08, -2.335199e-08, -2.408432e-08, -2.458342e-08, -2.416854e-08,
  -1.35518e-08, -1.42681e-08, -1.509972e-08, -1.553774e-08, -1.567415e-08, 
    -1.569752e-08, -1.557387e-08, -1.631249e-08, -1.833273e-08, 
    -2.141361e-08, -2.361357e-08, -2.445395e-08, -2.455297e-08, 
    -2.416797e-08, -2.413321e-08,
  -1.36032e-08, -1.445179e-08, -1.518814e-08, -1.537897e-08, -1.554013e-08, 
    -1.55565e-08, -1.606386e-08, -1.782417e-08, -2.072754e-08, -2.35171e-08, 
    -2.46558e-08, -2.476045e-08, -2.438934e-08, -2.425906e-08, -2.437382e-08,
  -1.366771e-08, -1.453646e-08, -1.509484e-08, -1.521914e-08, -1.549423e-08, 
    -1.594935e-08, -1.723611e-08, -1.965092e-08, -2.252601e-08, 
    -2.449912e-08, -2.497366e-08, -2.484371e-08, -2.488921e-08, 
    -2.505404e-08, -2.510338e-08,
  -1.370884e-08, -1.451639e-08, -1.490337e-08, -1.517058e-08, -1.575321e-08, 
    -1.673311e-08, -1.856668e-08, -2.115403e-08, -2.374345e-08, 
    -2.498053e-08, -2.533342e-08, -2.554345e-08, -2.587336e-08, 
    -2.604153e-08, -2.611419e-08,
  -1.371575e-08, -1.432636e-08, -1.470494e-08, -1.528747e-08, -1.620549e-08, 
    -1.75645e-08, -1.970212e-08, -2.226037e-08, -2.423018e-08, -2.536428e-08, 
    -2.60728e-08, -2.638111e-08, -2.68018e-08, -2.703617e-08, -2.731987e-08,
  -1.360844e-08, -1.407121e-08, -1.45589e-08, -1.546592e-08, -1.665435e-08, 
    -1.827181e-08, -2.042354e-08, -2.260561e-08, -2.438616e-08, 
    -2.593182e-08, -2.67197e-08, -2.720342e-08, -2.768919e-08, -2.800042e-08, 
    -2.856927e-08,
  -1.343208e-08, -1.38038e-08, -1.444091e-08, -1.566764e-08, -1.706007e-08, 
    -1.882859e-08, -2.083427e-08, -2.282267e-08, -2.477286e-08, 
    -2.650612e-08, -2.730284e-08, -2.764539e-08, -2.77948e-08, -2.813115e-08, 
    -2.866513e-08,
  -2.055143e-08, -2.157909e-08, -2.15645e-08, -2.166089e-08, -2.174198e-08, 
    -2.199562e-08, -2.207808e-08, -2.210325e-08, -2.217233e-08, -2.22008e-08, 
    -2.226312e-08, -2.233603e-08, -2.244693e-08, -2.251602e-08, -2.259079e-08,
  -2.136247e-08, -2.136548e-08, -2.133777e-08, -2.192311e-08, -2.234409e-08, 
    -2.26323e-08, -2.291431e-08, -2.325985e-08, -2.342793e-08, -2.354645e-08, 
    -2.356949e-08, -2.353186e-08, -2.343264e-08, -2.329134e-08, -2.312758e-08,
  -2.09429e-08, -2.143224e-08, -2.230238e-08, -2.31693e-08, -2.38824e-08, 
    -2.430323e-08, -2.438686e-08, -2.402838e-08, -2.363669e-08, 
    -2.321856e-08, -2.294981e-08, -2.260118e-08, -2.232683e-08, 
    -2.203102e-08, -2.180539e-08,
  -2.136874e-08, -2.271239e-08, -2.400793e-08, -2.49626e-08, -2.496599e-08, 
    -2.442623e-08, -2.349238e-08, -2.277045e-08, -2.225173e-08, 
    -2.181235e-08, -2.143648e-08, -2.111082e-08, -2.086588e-08, 
    -2.069693e-08, -2.059368e-08,
  -2.26932e-08, -2.451212e-08, -2.55178e-08, -2.50512e-08, -2.411438e-08, 
    -2.294451e-08, -2.187035e-08, -2.126311e-08, -2.068276e-08, 
    -2.030188e-08, -1.990691e-08, -1.962998e-08, -1.943476e-08, 
    -1.937824e-08, -1.934995e-08,
  -2.418428e-08, -2.539952e-08, -2.48199e-08, -2.366557e-08, -2.215136e-08, 
    -2.04757e-08, -1.934045e-08, -1.865802e-08, -1.837339e-08, -1.81863e-08, 
    -1.808084e-08, -1.805275e-08, -1.81397e-08, -1.835071e-08, -1.849233e-08,
  -2.482327e-08, -2.488356e-08, -2.342414e-08, -2.14053e-08, -1.925313e-08, 
    -1.789199e-08, -1.75207e-08, -1.766271e-08, -1.800785e-08, -1.837346e-08, 
    -1.867122e-08, -1.902763e-08, -1.946813e-08, -1.990914e-08, -2.010651e-08,
  -2.450695e-08, -2.363933e-08, -2.102221e-08, -1.857108e-08, -1.74531e-08, 
    -1.755414e-08, -1.808334e-08, -1.883814e-08, -1.951303e-08, 
    -2.018618e-08, -2.082536e-08, -2.146826e-08, -2.202452e-08, 
    -2.245159e-08, -2.275581e-08,
  -2.342285e-08, -2.157686e-08, -1.875922e-08, -1.776326e-08, -1.816276e-08, 
    -1.908713e-08, -2.004669e-08, -2.120896e-08, -2.249253e-08, 
    -2.385589e-08, -2.489461e-08, -2.571261e-08, -2.621568e-08, 
    -2.657406e-08, -2.66603e-08,
  -2.17794e-08, -1.981517e-08, -1.806827e-08, -1.83826e-08, -1.930186e-08, 
    -2.061672e-08, -2.224964e-08, -2.420104e-08, -2.594029e-08, 
    -2.716006e-08, -2.789008e-08, -2.828337e-08, -2.855745e-08, 
    -2.889433e-08, -2.913272e-08,
  -2.44481e-08, -2.44383e-08, -2.429655e-08, -2.414868e-08, -2.382523e-08, 
    -2.365212e-08, -2.350569e-08, -2.329554e-08, -2.306293e-08, 
    -2.281616e-08, -2.247065e-08, -2.200735e-08, -2.139306e-08, 
    -2.059168e-08, -1.96416e-08,
  -2.445766e-08, -2.450261e-08, -2.415608e-08, -2.395318e-08, -2.376216e-08, 
    -2.38002e-08, -2.386131e-08, -2.402665e-08, -2.424638e-08, -2.434209e-08, 
    -2.433457e-08, -2.412988e-08, -2.375679e-08, -2.315596e-08, -2.228217e-08,
  -2.426784e-08, -2.418826e-08, -2.365813e-08, -2.349675e-08, -2.337866e-08, 
    -2.341605e-08, -2.363333e-08, -2.398871e-08, -2.441156e-08, 
    -2.487089e-08, -2.525963e-08, -2.549028e-08, -2.547482e-08, 
    -2.514453e-08, -2.456218e-08,
  -2.41525e-08, -2.39974e-08, -2.360028e-08, -2.351549e-08, -2.356527e-08, 
    -2.382211e-08, -2.423916e-08, -2.463261e-08, -2.488703e-08, 
    -2.508805e-08, -2.527511e-08, -2.549327e-08, -2.565666e-08, 
    -2.568927e-08, -2.547935e-08,
  -2.438792e-08, -2.414744e-08, -2.41042e-08, -2.436434e-08, -2.458349e-08, 
    -2.498207e-08, -2.539346e-08, -2.55164e-08, -2.562394e-08, -2.563577e-08, 
    -2.576391e-08, -2.58636e-08, -2.595086e-08, -2.59271e-08, -2.586951e-08,
  -2.526723e-08, -2.52153e-08, -2.552779e-08, -2.595082e-08, -2.645262e-08, 
    -2.696398e-08, -2.729691e-08, -2.734425e-08, -2.729129e-08, 
    -2.717882e-08, -2.689401e-08, -2.673823e-08, -2.638419e-08, 
    -2.600928e-08, -2.569731e-08,
  -2.552619e-08, -2.578093e-08, -2.624239e-08, -2.682967e-08, -2.7458e-08, 
    -2.784072e-08, -2.817519e-08, -2.832034e-08, -2.839405e-08, 
    -2.844497e-08, -2.830807e-08, -2.807394e-08, -2.747691e-08, 
    -2.672153e-08, -2.610905e-08,
  -2.615749e-08, -2.678534e-08, -2.736965e-08, -2.787683e-08, -2.824797e-08, 
    -2.847675e-08, -2.857246e-08, -2.862475e-08, -2.854068e-08, 
    -2.852344e-08, -2.825982e-08, -2.806717e-08, -2.778022e-08, 
    -2.726029e-08, -2.657853e-08,
  -2.644349e-08, -2.733519e-08, -2.814206e-08, -2.859842e-08, -2.867239e-08, 
    -2.879472e-08, -2.890414e-08, -2.898346e-08, -2.888808e-08, 
    -2.854229e-08, -2.821251e-08, -2.771973e-08, -2.740686e-08, 
    -2.714457e-08, -2.693627e-08,
  -2.646377e-08, -2.772946e-08, -2.873313e-08, -2.887533e-08, -2.869305e-08, 
    -2.858201e-08, -2.858306e-08, -2.863809e-08, -2.854395e-08, 
    -2.840003e-08, -2.828049e-08, -2.798453e-08, -2.749933e-08, 
    -2.697961e-08, -2.647202e-08,
  -2.308686e-08, -2.333118e-08, -2.340088e-08, -2.338072e-08, -2.33958e-08, 
    -2.343506e-08, -2.3464e-08, -2.350418e-08, -2.352271e-08, -2.345745e-08, 
    -2.307038e-08, -2.247737e-08, -2.16678e-08, -2.078188e-08, -1.997385e-08,
  -2.377021e-08, -2.415197e-08, -2.422952e-08, -2.423845e-08, -2.435014e-08, 
    -2.44515e-08, -2.459434e-08, -2.476187e-08, -2.499717e-08, -2.505865e-08, 
    -2.481093e-08, -2.431202e-08, -2.366533e-08, -2.275339e-08, -2.187507e-08,
  -2.421502e-08, -2.452793e-08, -2.45271e-08, -2.466464e-08, -2.484958e-08, 
    -2.500234e-08, -2.519965e-08, -2.546547e-08, -2.57662e-08, -2.585703e-08, 
    -2.568039e-08, -2.526978e-08, -2.485022e-08, -2.425887e-08, -2.351878e-08,
  -2.456433e-08, -2.471555e-08, -2.466351e-08, -2.498998e-08, -2.517516e-08, 
    -2.550321e-08, -2.575242e-08, -2.613481e-08, -2.651958e-08, 
    -2.672026e-08, -2.654691e-08, -2.608568e-08, -2.553145e-08, 
    -2.516795e-08, -2.47543e-08,
  -2.48121e-08, -2.473015e-08, -2.487887e-08, -2.512088e-08, -2.545489e-08, 
    -2.579265e-08, -2.602882e-08, -2.6379e-08, -2.682714e-08, -2.71157e-08, 
    -2.719252e-08, -2.699924e-08, -2.653121e-08, -2.607296e-08, -2.560634e-08,
  -2.490284e-08, -2.490106e-08, -2.523067e-08, -2.550502e-08, -2.602592e-08, 
    -2.635729e-08, -2.654836e-08, -2.67752e-08, -2.705699e-08, -2.734209e-08, 
    -2.75135e-08, -2.758458e-08, -2.751359e-08, -2.715807e-08, -2.679637e-08,
  -2.508368e-08, -2.532462e-08, -2.573207e-08, -2.611978e-08, -2.672643e-08, 
    -2.703367e-08, -2.710426e-08, -2.728348e-08, -2.75188e-08, -2.788519e-08, 
    -2.817019e-08, -2.824477e-08, -2.832398e-08, -2.826506e-08, -2.792155e-08,
  -2.556112e-08, -2.593343e-08, -2.644571e-08, -2.696611e-08, -2.753611e-08, 
    -2.781176e-08, -2.773087e-08, -2.774243e-08, -2.790226e-08, 
    -2.832324e-08, -2.885335e-08, -2.914006e-08, -2.929444e-08, 
    -2.922842e-08, -2.892839e-08,
  -2.657055e-08, -2.695972e-08, -2.743647e-08, -2.803211e-08, -2.84599e-08, 
    -2.871189e-08, -2.869411e-08, -2.864522e-08, -2.865369e-08, -2.8881e-08, 
    -2.93996e-08, -2.967827e-08, -2.992353e-08, -3.015186e-08, -3.006857e-08,
  -2.800759e-08, -2.852905e-08, -2.888809e-08, -2.926654e-08, -2.963272e-08, 
    -2.983709e-08, -3.006816e-08, -3.015683e-08, -3.017135e-08, 
    -3.010046e-08, -3.026594e-08, -3.046875e-08, -3.038906e-08, 
    -3.064608e-08, -3.082034e-08,
  -3.070679e-08, -3.013844e-08, -2.931571e-08, -2.859967e-08, -2.792967e-08, 
    -2.729394e-08, -2.694103e-08, -2.64378e-08, -2.592972e-08, -2.520841e-08, 
    -2.455606e-08, -2.391819e-08, -2.32842e-08, -2.272174e-08, -2.214288e-08,
  -3.138428e-08, -3.107753e-08, -3.028269e-08, -2.930316e-08, -2.862113e-08, 
    -2.788462e-08, -2.72592e-08, -2.661653e-08, -2.618227e-08, -2.560726e-08, 
    -2.522213e-08, -2.476162e-08, -2.422157e-08, -2.367756e-08, -2.314656e-08,
  -3.153622e-08, -3.183144e-08, -3.141412e-08, -3.008066e-08, -2.906642e-08, 
    -2.828379e-08, -2.756221e-08, -2.653693e-08, -2.563968e-08, 
    -2.498956e-08, -2.480654e-08, -2.473989e-08, -2.461026e-08, 
    -2.435459e-08, -2.391401e-08,
  -3.092105e-08, -3.166299e-08, -3.216362e-08, -3.126427e-08, -3.008038e-08, 
    -2.86844e-08, -2.789685e-08, -2.709302e-08, -2.618042e-08, -2.515618e-08, 
    -2.470068e-08, -2.457162e-08, -2.455906e-08, -2.459958e-08, -2.432644e-08,
  -3.010951e-08, -3.11045e-08, -3.204615e-08, -3.171369e-08, -3.097548e-08, 
    -2.989125e-08, -2.865936e-08, -2.754057e-08, -2.665842e-08, 
    -2.562687e-08, -2.492432e-08, -2.461999e-08, -2.443069e-08, 
    -2.436276e-08, -2.408991e-08,
  -2.933038e-08, -3.045472e-08, -3.144067e-08, -3.163854e-08, -3.104084e-08, 
    -3.04287e-08, -2.988395e-08, -2.863297e-08, -2.759012e-08, -2.635765e-08, 
    -2.534861e-08, -2.485495e-08, -2.457806e-08, -2.423898e-08, -2.386024e-08,
  -2.893441e-08, -2.989814e-08, -3.07569e-08, -3.123257e-08, -3.071209e-08, 
    -3.012633e-08, -3.001787e-08, -2.954792e-08, -2.857183e-08, 
    -2.751421e-08, -2.637439e-08, -2.549223e-08, -2.514615e-08, 
    -2.480467e-08, -2.422749e-08,
  -2.877191e-08, -2.964462e-08, -3.005802e-08, -3.050064e-08, -3.053061e-08, 
    -2.970951e-08, -2.944138e-08, -2.950467e-08, -2.92034e-08, -2.811277e-08, 
    -2.739977e-08, -2.671518e-08, -2.620482e-08, -2.563131e-08, -2.505267e-08,
  -2.888947e-08, -2.966251e-08, -2.980988e-08, -2.988623e-08, -3.00342e-08, 
    -2.976712e-08, -2.919572e-08, -2.881577e-08, -2.891413e-08, 
    -2.852846e-08, -2.77375e-08, -2.756857e-08, -2.746891e-08, -2.681002e-08, 
    -2.596547e-08,
  -2.925473e-08, -2.996664e-08, -2.9989e-08, -3.003948e-08, -2.993291e-08, 
    -2.970567e-08, -2.942107e-08, -2.872783e-08, -2.838734e-08, 
    -2.840779e-08, -2.81162e-08, -2.78628e-08, -2.80055e-08, -2.797395e-08, 
    -2.723152e-08,
  -2.901421e-08, -2.710518e-08, -2.576287e-08, -2.508039e-08, -2.488976e-08, 
    -2.488023e-08, -2.458778e-08, -2.385216e-08, -2.349239e-08, 
    -2.302146e-08, -2.233839e-08, -2.118702e-08, -2.01146e-08, -1.918018e-08, 
    -1.84677e-08,
  -2.776908e-08, -2.6009e-08, -2.525745e-08, -2.491754e-08, -2.482742e-08, 
    -2.478374e-08, -2.464089e-08, -2.400741e-08, -2.338611e-08, 
    -2.265627e-08, -2.189772e-08, -2.084921e-08, -1.986103e-08, 
    -1.895242e-08, -1.828099e-08,
  -2.688342e-08, -2.53162e-08, -2.470889e-08, -2.453424e-08, -2.432911e-08, 
    -2.425951e-08, -2.424769e-08, -2.346007e-08, -2.251066e-08, 
    -2.178106e-08, -2.111343e-08, -2.014606e-08, -1.912259e-08, 
    -1.828249e-08, -1.748896e-08,
  -2.605887e-08, -2.498437e-08, -2.44101e-08, -2.425911e-08, -2.429838e-08, 
    -2.410364e-08, -2.417883e-08, -2.330517e-08, -2.183473e-08, 
    -2.092072e-08, -2.018855e-08, -1.952659e-08, -1.875606e-08, 
    -1.772634e-08, -1.695508e-08,
  -2.505149e-08, -2.468196e-08, -2.427559e-08, -2.389974e-08, -2.397272e-08, 
    -2.400401e-08, -2.395419e-08, -2.295859e-08, -2.134818e-08, 
    -2.042446e-08, -1.970315e-08, -1.904156e-08, -1.827133e-08, 
    -1.751788e-08, -1.66697e-08,
  -2.452723e-08, -2.432692e-08, -2.416162e-08, -2.353051e-08, -2.344862e-08, 
    -2.375425e-08, -2.346999e-08, -2.258991e-08, -2.113693e-08, 
    -2.016317e-08, -1.940234e-08, -1.871623e-08, -1.794262e-08, 
    -1.727804e-08, -1.643971e-08,
  -2.445058e-08, -2.432858e-08, -2.401959e-08, -2.337383e-08, -2.313438e-08, 
    -2.345007e-08, -2.314201e-08, -2.252484e-08, -2.102225e-08, 
    -1.997449e-08, -1.925193e-08, -1.850916e-08, -1.758483e-08, 
    -1.677753e-08, -1.594321e-08,
  -2.460733e-08, -2.44972e-08, -2.410264e-08, -2.332901e-08, -2.299734e-08, 
    -2.323052e-08, -2.288016e-08, -2.227484e-08, -2.103617e-08, 
    -1.995839e-08, -1.913044e-08, -1.834617e-08, -1.73113e-08, -1.646416e-08, 
    -1.568157e-08,
  -2.484338e-08, -2.458745e-08, -2.433904e-08, -2.349999e-08, -2.294039e-08, 
    -2.309105e-08, -2.287789e-08, -2.236608e-08, -2.124368e-08, 
    -1.995935e-08, -1.910225e-08, -1.815267e-08, -1.715471e-08, 
    -1.627557e-08, -1.563348e-08,
  -2.51957e-08, -2.480214e-08, -2.471245e-08, -2.400031e-08, -2.321143e-08, 
    -2.292799e-08, -2.275777e-08, -2.245615e-08, -2.168136e-08, -2.03144e-08, 
    -1.906762e-08, -1.811381e-08, -1.708493e-08, -1.606482e-08, -1.546788e-08,
  -1.512072e-08, -1.470676e-08, -1.436655e-08, -1.383244e-08, -1.396655e-08, 
    -1.406241e-08, -1.478309e-08, -1.541665e-08, -1.55704e-08, -1.57831e-08, 
    -1.512995e-08, -1.444289e-08, -1.467623e-08, -1.498394e-08, -1.400962e-08,
  -1.45086e-08, -1.427652e-08, -1.373876e-08, -1.340249e-08, -1.394119e-08, 
    -1.429645e-08, -1.475472e-08, -1.493144e-08, -1.48488e-08, -1.490548e-08, 
    -1.426114e-08, -1.379623e-08, -1.388918e-08, -1.410614e-08, -1.330652e-08,
  -1.436475e-08, -1.379946e-08, -1.362151e-08, -1.384587e-08, -1.474162e-08, 
    -1.479737e-08, -1.492259e-08, -1.484076e-08, -1.470859e-08, 
    -1.429865e-08, -1.349792e-08, -1.309493e-08, -1.301994e-08, 
    -1.316585e-08, -1.253859e-08,
  -1.400599e-08, -1.384047e-08, -1.425915e-08, -1.460304e-08, -1.502353e-08, 
    -1.494772e-08, -1.487766e-08, -1.474907e-08, -1.472015e-08, -1.41461e-08, 
    -1.325641e-08, -1.279791e-08, -1.260468e-08, -1.252129e-08, -1.218607e-08,
  -1.447594e-08, -1.459965e-08, -1.486324e-08, -1.50212e-08, -1.521041e-08, 
    -1.476685e-08, -1.453571e-08, -1.449798e-08, -1.460532e-08, 
    -1.382783e-08, -1.306729e-08, -1.260366e-08, -1.242726e-08, 
    -1.226007e-08, -1.213509e-08,
  -1.469955e-08, -1.48501e-08, -1.52783e-08, -1.554173e-08, -1.541672e-08, 
    -1.441021e-08, -1.40084e-08, -1.413165e-08, -1.433509e-08, -1.360904e-08, 
    -1.287517e-08, -1.255359e-08, -1.232336e-08, -1.219797e-08, -1.236571e-08,
  -1.525355e-08, -1.527428e-08, -1.517329e-08, -1.528738e-08, -1.502372e-08, 
    -1.420623e-08, -1.375816e-08, -1.375891e-08, -1.368736e-08, 
    -1.313146e-08, -1.288237e-08, -1.254236e-08, -1.232946e-08, 
    -1.222431e-08, -1.237641e-08,
  -1.492588e-08, -1.461929e-08, -1.438387e-08, -1.452157e-08, -1.430781e-08, 
    -1.381941e-08, -1.342301e-08, -1.340274e-08, -1.308653e-08, 
    -1.263748e-08, -1.290123e-08, -1.254248e-08, -1.229769e-08, 
    -1.215562e-08, -1.226962e-08,
  -1.476158e-08, -1.448013e-08, -1.415623e-08, -1.416234e-08, -1.411172e-08, 
    -1.369298e-08, -1.306182e-08, -1.2733e-08, -1.274626e-08, -1.253442e-08, 
    -1.271433e-08, -1.218743e-08, -1.208381e-08, -1.196231e-08, -1.231369e-08,
  -1.468818e-08, -1.435438e-08, -1.412545e-08, -1.401443e-08, -1.376659e-08, 
    -1.332149e-08, -1.284397e-08, -1.261248e-08, -1.245303e-08, 
    -1.241347e-08, -1.239173e-08, -1.181386e-08, -1.185075e-08, 
    -1.189617e-08, -1.280265e-08,
  -2.147081e-08, -2.012757e-08, -1.91044e-08, -1.851124e-08, -1.702544e-08, 
    -1.543764e-08, -1.397001e-08, -1.43729e-08, -1.573472e-08, -1.630723e-08, 
    -1.510471e-08, -1.474643e-08, -1.534151e-08, -1.64231e-08, -1.788977e-08,
  -1.957759e-08, -1.878814e-08, -1.759618e-08, -1.648303e-08, -1.498745e-08, 
    -1.350892e-08, -1.331862e-08, -1.478437e-08, -1.577124e-08, -1.531e-08, 
    -1.443352e-08, -1.461412e-08, -1.548026e-08, -1.672333e-08, -1.825798e-08,
  -1.777448e-08, -1.661893e-08, -1.55327e-08, -1.453706e-08, -1.302442e-08, 
    -1.284208e-08, -1.398477e-08, -1.514939e-08, -1.519045e-08, 
    -1.434945e-08, -1.417172e-08, -1.489645e-08, -1.596892e-08, 
    -1.723219e-08, -1.891973e-08,
  -1.615643e-08, -1.499501e-08, -1.390015e-08, -1.285207e-08, -1.266632e-08, 
    -1.361757e-08, -1.468322e-08, -1.500892e-08, -1.436281e-08, 
    -1.405317e-08, -1.438043e-08, -1.546246e-08, -1.663056e-08, 
    -1.814149e-08, -1.977988e-08,
  -1.466783e-08, -1.344231e-08, -1.268147e-08, -1.276603e-08, -1.370496e-08, 
    -1.468689e-08, -1.486401e-08, -1.435172e-08, -1.397327e-08, 
    -1.415125e-08, -1.519572e-08, -1.630307e-08, -1.773843e-08, 
    -1.918251e-08, -2.057001e-08,
  -1.305524e-08, -1.274313e-08, -1.300938e-08, -1.390837e-08, -1.460103e-08, 
    -1.475218e-08, -1.427871e-08, -1.401349e-08, -1.430929e-08, 
    -1.510567e-08, -1.613576e-08, -1.749665e-08, -1.881801e-08, 
    -2.011768e-08, -2.119905e-08,
  -1.300827e-08, -1.336864e-08, -1.398572e-08, -1.451343e-08, -1.450106e-08, 
    -1.422058e-08, -1.405548e-08, -1.453329e-08, -1.515667e-08, 
    -1.595938e-08, -1.731172e-08, -1.850555e-08, -1.979024e-08, 
    -2.090729e-08, -2.1956e-08,
  -1.366713e-08, -1.407414e-08, -1.43254e-08, -1.434551e-08, -1.410564e-08, 
    -1.435002e-08, -1.470761e-08, -1.532554e-08, -1.60062e-08, -1.739315e-08, 
    -1.850087e-08, -1.971033e-08, -2.073805e-08, -2.1754e-08, -2.249762e-08,
  -1.414964e-08, -1.419621e-08, -1.413594e-08, -1.400081e-08, -1.435438e-08, 
    -1.484611e-08, -1.53419e-08, -1.605099e-08, -1.745573e-08, -1.866472e-08, 
    -1.97954e-08, -2.077721e-08, -2.163164e-08, -2.237005e-08, -2.270198e-08,
  -1.414508e-08, -1.383865e-08, -1.387742e-08, -1.439525e-08, -1.517159e-08, 
    -1.56809e-08, -1.641949e-08, -1.742529e-08, -1.88118e-08, -1.989258e-08, 
    -2.096686e-08, -2.156775e-08, -2.21958e-08, -2.263035e-08, -2.272155e-08,
  -1.555972e-08, -1.754251e-08, -1.936036e-08, -2.114692e-08, -2.184356e-08, 
    -2.280186e-08, -2.269867e-08, -2.131199e-08, -1.998879e-08, 
    -1.848059e-08, -1.762089e-08, -1.866783e-08, -1.989394e-08, 
    -1.919191e-08, -1.876093e-08,
  -1.623333e-08, -1.825518e-08, -2.011007e-08, -2.168752e-08, -2.235262e-08, 
    -2.249642e-08, -2.124631e-08, -2.060502e-08, -1.911848e-08, 
    -1.747997e-08, -1.723422e-08, -1.953611e-08, -2.032384e-08, 
    -1.935689e-08, -1.893432e-08,
  -1.716026e-08, -1.91809e-08, -2.093669e-08, -2.221869e-08, -2.208424e-08, 
    -2.094434e-08, -2.029727e-08, -1.992935e-08, -1.786718e-08, 
    -1.659452e-08, -1.793749e-08, -2.061815e-08, -2.044559e-08, 
    -1.960322e-08, -1.908747e-08,
  -1.833966e-08, -2.031891e-08, -2.164321e-08, -2.177426e-08, -2.033812e-08, 
    -2.013699e-08, -1.957862e-08, -1.818203e-08, -1.647832e-08, 
    -1.675934e-08, -2.00307e-08, -2.143879e-08, -2.074819e-08, -1.969619e-08, 
    -1.926299e-08,
  -1.965986e-08, -2.114724e-08, -2.109992e-08, -2.037141e-08, -1.972317e-08, 
    -1.911795e-08, -1.791534e-08, -1.668628e-08, -1.658002e-08, 
    -1.972632e-08, -2.186169e-08, -2.180006e-08, -2.043904e-08, -1.96777e-08, 
    -1.943843e-08,
  -2.032576e-08, -2.080341e-08, -2.002905e-08, -1.949158e-08, -1.851824e-08, 
    -1.775033e-08, -1.681338e-08, -1.737348e-08, -1.990836e-08, 
    -2.222528e-08, -2.241616e-08, -2.12077e-08, -2.02057e-08, -1.982023e-08, 
    -1.964725e-08,
  -2.010269e-08, -2.008603e-08, -1.896432e-08, -1.830566e-08, -1.741135e-08, 
    -1.74362e-08, -1.884322e-08, -2.1036e-08, -2.281621e-08, -2.285979e-08, 
    -2.200035e-08, -2.080762e-08, -2.032982e-08, -1.999505e-08, -1.993473e-08,
  -1.933984e-08, -1.884464e-08, -1.785189e-08, -1.783535e-08, -1.912751e-08, 
    -2.087157e-08, -2.254962e-08, -2.34498e-08, -2.324083e-08, -2.251071e-08, 
    -2.147765e-08, -2.086066e-08, -2.052739e-08, -2.025035e-08, -2.017438e-08,
  -1.845713e-08, -1.835262e-08, -1.95251e-08, -2.17401e-08, -2.308566e-08, 
    -2.388677e-08, -2.410166e-08, -2.371554e-08, -2.290618e-08, 
    -2.216588e-08, -2.144097e-08, -2.101511e-08, -2.066319e-08, 
    -2.046009e-08, -2.023223e-08,
  -1.970903e-08, -2.218263e-08, -2.412916e-08, -2.484722e-08, -2.496732e-08, 
    -2.464334e-08, -2.424285e-08, -2.339683e-08, -2.28127e-08, -2.207531e-08, 
    -2.161404e-08, -2.109085e-08, -2.082453e-08, -2.046391e-08, -2.030919e-08,
  -1.038291e-08, -1.13884e-08, -1.272126e-08, -1.356734e-08, -1.444527e-08, 
    -1.589472e-08, -1.717657e-08, -1.821145e-08, -1.793383e-08, 
    -1.781372e-08, -1.86246e-08, -1.969135e-08, -2.01683e-08, -2.00754e-08, 
    -1.988891e-08,
  -1.095519e-08, -1.210707e-08, -1.307111e-08, -1.363556e-08, -1.456767e-08, 
    -1.616842e-08, -1.727942e-08, -1.812685e-08, -1.79768e-08, -1.802731e-08, 
    -1.862084e-08, -1.932287e-08, -2.005874e-08, -1.9832e-08, -1.973038e-08,
  -1.163244e-08, -1.252673e-08, -1.339325e-08, -1.394039e-08, -1.480588e-08, 
    -1.631649e-08, -1.738489e-08, -1.807866e-08, -1.809953e-08, 
    -1.837335e-08, -1.873544e-08, -1.939979e-08, -1.989526e-08, 
    -1.961653e-08, -1.973349e-08,
  -1.205578e-08, -1.290262e-08, -1.385861e-08, -1.436229e-08, -1.518143e-08, 
    -1.648934e-08, -1.740586e-08, -1.80992e-08, -1.829877e-08, -1.870802e-08, 
    -1.897941e-08, -1.943533e-08, -1.958102e-08, -1.934828e-08, -1.975691e-08,
  -1.247164e-08, -1.338705e-08, -1.437544e-08, -1.481228e-08, -1.566371e-08, 
    -1.688871e-08, -1.784136e-08, -1.828683e-08, -1.858728e-08, 
    -1.897935e-08, -1.917738e-08, -1.944526e-08, -1.924695e-08, 
    -1.925584e-08, -2.002661e-08,
  -1.306613e-08, -1.412176e-08, -1.485799e-08, -1.541355e-08, -1.636467e-08, 
    -1.75772e-08, -1.816306e-08, -1.860796e-08, -1.87753e-08, -1.920986e-08, 
    -1.935641e-08, -1.933929e-08, -1.90246e-08, -1.927829e-08, -2.063845e-08,
  -1.384624e-08, -1.473073e-08, -1.54312e-08, -1.626374e-08, -1.734208e-08, 
    -1.823861e-08, -1.851578e-08, -1.877888e-08, -1.911312e-08, 
    -1.946261e-08, -1.948517e-08, -1.909151e-08, -1.906948e-08, 
    -1.971694e-08, -2.149381e-08,
  -1.436881e-08, -1.529972e-08, -1.637104e-08, -1.744569e-08, -1.824961e-08, 
    -1.860581e-08, -1.876963e-08, -1.917066e-08, -1.952161e-08, 
    -1.967506e-08, -1.926124e-08, -1.897458e-08, -1.933335e-08, 
    -2.058106e-08, -2.221875e-08,
  -1.530618e-08, -1.620047e-08, -1.759044e-08, -1.831292e-08, -1.866183e-08, 
    -1.89733e-08, -1.933778e-08, -1.96528e-08, -1.976216e-08, -1.942846e-08, 
    -1.907078e-08, -1.921497e-08, -2.00756e-08, -2.144118e-08, -2.276238e-08,
  -1.643584e-08, -1.725382e-08, -1.845721e-08, -1.895117e-08, -1.931147e-08, 
    -1.968281e-08, -1.985651e-08, -1.98891e-08, -1.950844e-08, -1.924542e-08, 
    -1.926996e-08, -1.981713e-08, -2.099695e-08, -2.198057e-08, -2.318004e-08,
  -1.109603e-08, -1.261941e-08, -1.447514e-08, -1.708823e-08, -1.542406e-08, 
    -1.227101e-08, -1.316805e-08, -1.533727e-08, -1.78841e-08, -1.996743e-08, 
    -2.038414e-08, -2.098095e-08, -2.064155e-08, -1.974897e-08, -1.976953e-08,
  -9.974468e-09, -1.091347e-08, -1.256785e-08, -1.400936e-08, -1.551291e-08, 
    -1.397673e-08, -1.275718e-08, -1.364959e-08, -1.571213e-08, 
    -1.828371e-08, -1.986889e-08, -2.068745e-08, -2.120333e-08, 
    -2.031486e-08, -1.992525e-08,
  -9.205265e-09, -9.732807e-09, -1.129974e-08, -1.212397e-08, -1.407298e-08, 
    -1.456653e-08, -1.325071e-08, -1.318958e-08, -1.44465e-08, -1.681182e-08, 
    -1.883005e-08, -2.033937e-08, -2.124113e-08, -2.084261e-08, -2.024766e-08,
  -9.520275e-09, -9.355753e-09, -1.067819e-08, -1.113903e-08, -1.190187e-08, 
    -1.406768e-08, -1.376938e-08, -1.295685e-08, -1.371049e-08, 
    -1.555728e-08, -1.771705e-08, -1.960182e-08, -2.108604e-08, 
    -2.130023e-08, -2.064941e-08,
  -9.645384e-09, -9.524145e-09, -1.037747e-08, -1.048029e-08, -1.053875e-08, 
    -1.247512e-08, -1.400242e-08, -1.294408e-08, -1.309671e-08, 
    -1.468872e-08, -1.672986e-08, -1.868321e-08, -2.040702e-08, 
    -2.151404e-08, -2.117201e-08,
  -9.231655e-09, -9.574658e-09, -1.014869e-08, -1.061023e-08, -1.007145e-08, 
    -1.11375e-08, -1.322291e-08, -1.287997e-08, -1.257506e-08, -1.401368e-08, 
    -1.585914e-08, -1.789736e-08, -1.959118e-08, -2.117863e-08, -2.146792e-08,
  -8.952033e-09, -9.585921e-09, -1.015015e-08, -1.05877e-08, -9.961454e-09, 
    -1.022119e-08, -1.246304e-08, -1.260714e-08, -1.225076e-08, 
    -1.351403e-08, -1.531753e-08, -1.730544e-08, -1.89053e-08, -2.053213e-08, 
    -2.144176e-08,
  -8.767874e-09, -9.447787e-09, -1.035104e-08, -1.079292e-08, -1.005813e-08, 
    -9.941198e-09, -1.168337e-08, -1.223963e-08, -1.186429e-08, 
    -1.311528e-08, -1.48496e-08, -1.683893e-08, -1.850763e-08, -1.989536e-08, 
    -2.108918e-08,
  -8.687117e-09, -9.451412e-09, -1.031784e-08, -1.080109e-08, -1.029912e-08, 
    -9.958568e-09, -1.121378e-08, -1.161496e-08, -1.16248e-08, -1.302115e-08, 
    -1.44992e-08, -1.66028e-08, -1.81884e-08, -1.94343e-08, -2.076579e-08,
  -8.58602e-09, -9.412088e-09, -1.031229e-08, -1.091033e-08, -1.025757e-08, 
    -9.923077e-09, -1.078467e-08, -1.116412e-08, -1.160775e-08, 
    -1.298713e-08, -1.43668e-08, -1.639712e-08, -1.808463e-08, -1.908539e-08, 
    -2.046488e-08,
  -1.851832e-08, -1.879505e-08, -1.882775e-08, -1.928398e-08, -1.948003e-08, 
    -2.008248e-08, -2.077783e-08, -2.110895e-08, -2.042505e-08, 
    -2.180713e-08, -2.294825e-08, -2.361613e-08, -2.412752e-08, 
    -2.391173e-08, -2.40686e-08,
  -1.834469e-08, -1.84788e-08, -1.847554e-08, -1.866908e-08, -1.861325e-08, 
    -1.917635e-08, -1.933248e-08, -2.064821e-08, -2.098032e-08, 
    -2.092457e-08, -2.205875e-08, -2.282032e-08, -2.35283e-08, -2.42222e-08, 
    -2.404134e-08,
  -1.810406e-08, -1.817159e-08, -1.799527e-08, -1.818011e-08, -1.805872e-08, 
    -1.824918e-08, -1.858166e-08, -1.915775e-08, -2.057713e-08, 
    -2.123033e-08, -2.118133e-08, -2.199621e-08, -2.287384e-08, 
    -2.331099e-08, -2.39187e-08,
  -1.787973e-08, -1.811937e-08, -1.817667e-08, -1.811584e-08, -1.78635e-08, 
    -1.768118e-08, -1.79479e-08, -1.84454e-08, -1.915693e-08, -2.035518e-08, 
    -2.111369e-08, -2.152352e-08, -2.203855e-08, -2.268131e-08, -2.31803e-08,
  -1.75193e-08, -1.773262e-08, -1.788546e-08, -1.783911e-08, -1.780781e-08, 
    -1.74272e-08, -1.739179e-08, -1.78915e-08, -1.803765e-08, -1.890016e-08, 
    -1.998173e-08, -2.04733e-08, -2.14336e-08, -2.189087e-08, -2.247779e-08,
  -1.702907e-08, -1.760448e-08, -1.784736e-08, -1.767008e-08, -1.758411e-08, 
    -1.719482e-08, -1.691619e-08, -1.749124e-08, -1.740324e-08, 
    -1.753413e-08, -1.869249e-08, -1.963215e-08, -2.015118e-08, 
    -2.104026e-08, -2.162382e-08,
  -1.625262e-08, -1.687954e-08, -1.77321e-08, -1.761898e-08, -1.742737e-08, 
    -1.678488e-08, -1.641529e-08, -1.690288e-08, -1.712176e-08, -1.6565e-08, 
    -1.736912e-08, -1.864477e-08, -1.94826e-08, -1.973511e-08, -2.074212e-08,
  -1.602608e-08, -1.65992e-08, -1.73652e-08, -1.763022e-08, -1.76543e-08, 
    -1.674428e-08, -1.577206e-08, -1.614703e-08, -1.677531e-08, 
    -1.615104e-08, -1.664285e-08, -1.75474e-08, -1.866828e-08, -1.89747e-08, 
    -1.954233e-08,
  -1.560249e-08, -1.634566e-08, -1.715948e-08, -1.757252e-08, -1.747769e-08, 
    -1.68663e-08, -1.560035e-08, -1.564926e-08, -1.606511e-08, -1.577593e-08, 
    -1.600399e-08, -1.704699e-08, -1.773533e-08, -1.828653e-08, -1.85611e-08,
  -1.546654e-08, -1.601459e-08, -1.697301e-08, -1.764942e-08, -1.735075e-08, 
    -1.675655e-08, -1.55827e-08, -1.557276e-08, -1.553186e-08, -1.542104e-08, 
    -1.558477e-08, -1.663468e-08, -1.717883e-08, -1.781031e-08, -1.79881e-08,
  -2.748552e-08, -2.73571e-08, -2.576628e-08, -2.517127e-08, -2.454391e-08, 
    -2.44094e-08, -2.426321e-08, -2.432317e-08, -2.431058e-08, -2.431054e-08, 
    -2.431141e-08, -2.425928e-08, -2.417755e-08, -2.400891e-08, -2.379908e-08,
  -2.6701e-08, -2.652972e-08, -2.564106e-08, -2.521329e-08, -2.471416e-08, 
    -2.467106e-08, -2.452432e-08, -2.455704e-08, -2.458475e-08, -2.46219e-08, 
    -2.44697e-08, -2.445482e-08, -2.435501e-08, -2.431474e-08, -2.425478e-08,
  -2.609152e-08, -2.61155e-08, -2.543124e-08, -2.482141e-08, -2.427375e-08, 
    -2.415733e-08, -2.396728e-08, -2.415612e-08, -2.411582e-08, 
    -2.408711e-08, -2.385105e-08, -2.376549e-08, -2.367298e-08, 
    -2.362624e-08, -2.357056e-08,
  -2.583372e-08, -2.575205e-08, -2.500101e-08, -2.418594e-08, -2.35921e-08, 
    -2.321826e-08, -2.315515e-08, -2.342168e-08, -2.366927e-08, 
    -2.375084e-08, -2.360098e-08, -2.343799e-08, -2.331974e-08, 
    -2.324244e-08, -2.317033e-08,
  -2.563217e-08, -2.537059e-08, -2.475782e-08, -2.393129e-08, -2.322442e-08, 
    -2.287551e-08, -2.286208e-08, -2.305876e-08, -2.334614e-08, 
    -2.341882e-08, -2.339678e-08, -2.335746e-08, -2.336827e-08, 
    -2.325289e-08, -2.318787e-08,
  -2.570995e-08, -2.540883e-08, -2.469629e-08, -2.401157e-08, -2.338514e-08, 
    -2.28763e-08, -2.280991e-08, -2.290654e-08, -2.31774e-08, -2.309653e-08, 
    -2.30397e-08, -2.299717e-08, -2.300465e-08, -2.290722e-08, -2.286043e-08,
  -2.579476e-08, -2.54588e-08, -2.480396e-08, -2.411349e-08, -2.352382e-08, 
    -2.312084e-08, -2.280894e-08, -2.282719e-08, -2.310159e-08, 
    -2.313534e-08, -2.318792e-08, -2.312442e-08, -2.289178e-08, 
    -2.287296e-08, -2.278161e-08,
  -2.589935e-08, -2.556474e-08, -2.504682e-08, -2.436464e-08, -2.373015e-08, 
    -2.325241e-08, -2.27989e-08, -2.28465e-08, -2.297679e-08, -2.296323e-08, 
    -2.288368e-08, -2.301763e-08, -2.298137e-08, -2.29883e-08, -2.28387e-08,
  -2.603806e-08, -2.562691e-08, -2.526551e-08, -2.461828e-08, -2.374833e-08, 
    -2.310927e-08, -2.271425e-08, -2.27936e-08, -2.286936e-08, -2.274306e-08, 
    -2.261962e-08, -2.277352e-08, -2.277507e-08, -2.28834e-08, -2.293299e-08,
  -2.605202e-08, -2.557669e-08, -2.547509e-08, -2.488792e-08, -2.391931e-08, 
    -2.310103e-08, -2.279892e-08, -2.266118e-08, -2.279267e-08, 
    -2.235832e-08, -2.242649e-08, -2.229013e-08, -2.256655e-08, 
    -2.267386e-08, -2.304759e-08,
  -1.966614e-08, -1.982747e-08, -2.013045e-08, -2.043602e-08, -2.058347e-08, 
    -2.061461e-08, -2.048833e-08, -2.036001e-08, -2.017323e-08, 
    -1.992876e-08, -1.966667e-08, -1.932748e-08, -1.901296e-08, 
    -1.871974e-08, -1.848369e-08,
  -2.070582e-08, -2.05109e-08, -2.066217e-08, -2.062898e-08, -2.070814e-08, 
    -2.073362e-08, -2.075871e-08, -2.076006e-08, -2.083109e-08, 
    -2.088642e-08, -2.092904e-08, -2.091041e-08, -2.086196e-08, 
    -2.078153e-08, -2.069995e-08,
  -2.161979e-08, -2.151774e-08, -2.153801e-08, -2.150843e-08, -2.152162e-08, 
    -2.144681e-08, -2.12941e-08, -2.115488e-08, -2.108283e-08, -2.110475e-08, 
    -2.121295e-08, -2.137928e-08, -2.154033e-08, -2.17035e-08, -2.181866e-08,
  -2.261678e-08, -2.246824e-08, -2.236656e-08, -2.228927e-08, -2.223099e-08, 
    -2.210423e-08, -2.18978e-08, -2.171494e-08, -2.147712e-08, -2.132554e-08, 
    -2.124846e-08, -2.120815e-08, -2.120967e-08, -2.120716e-08, -2.128022e-08,
  -2.2981e-08, -2.277647e-08, -2.259239e-08, -2.242706e-08, -2.229189e-08, 
    -2.205607e-08, -2.184018e-08, -2.158266e-08, -2.143785e-08, 
    -2.124556e-08, -2.112451e-08, -2.099868e-08, -2.09839e-08, -2.099279e-08, 
    -2.101357e-08,
  -2.271337e-08, -2.254465e-08, -2.232046e-08, -2.211637e-08, -2.192439e-08, 
    -2.170919e-08, -2.149098e-08, -2.125396e-08, -2.116735e-08, 
    -2.099153e-08, -2.093183e-08, -2.074148e-08, -2.064055e-08, 
    -2.054097e-08, -2.053164e-08,
  -2.253137e-08, -2.236491e-08, -2.226969e-08, -2.212442e-08, -2.200817e-08, 
    -2.180565e-08, -2.172068e-08, -2.156966e-08, -2.160349e-08, 
    -2.142085e-08, -2.136001e-08, -2.113139e-08, -2.097083e-08, 
    -2.078603e-08, -2.063347e-08,
  -2.235682e-08, -2.225886e-08, -2.224438e-08, -2.217801e-08, -2.216577e-08, 
    -2.215172e-08, -2.226797e-08, -2.233971e-08, -2.24554e-08, -2.244349e-08, 
    -2.236319e-08, -2.22515e-08, -2.208434e-08, -2.182328e-08, -2.159291e-08,
  -2.228536e-08, -2.232296e-08, -2.232702e-08, -2.231142e-08, -2.240197e-08, 
    -2.25395e-08, -2.283674e-08, -2.303071e-08, -2.319924e-08, -2.336702e-08, 
    -2.341935e-08, -2.340668e-08, -2.332399e-08, -2.317292e-08, -2.293732e-08,
  -2.229811e-08, -2.238877e-08, -2.237369e-08, -2.236817e-08, -2.248562e-08, 
    -2.275482e-08, -2.316865e-08, -2.345663e-08, -2.374823e-08, 
    -2.396754e-08, -2.419401e-08, -2.425388e-08, -2.436803e-08, 
    -2.430668e-08, -2.414645e-08,
  -2.139515e-08, -2.092572e-08, -2.057009e-08, -2.022146e-08, -1.991053e-08, 
    -1.961189e-08, -1.933746e-08, -1.904858e-08, -1.873753e-08, 
    -1.837802e-08, -1.798962e-08, -1.764562e-08, -1.737273e-08, 
    -1.720385e-08, -1.708187e-08,
  -2.244523e-08, -2.231122e-08, -2.216125e-08, -2.199351e-08, -2.182462e-08, 
    -2.166869e-08, -2.151911e-08, -2.133997e-08, -2.110035e-08, 
    -2.076966e-08, -2.043327e-08, -2.005603e-08, -1.974964e-08, 
    -1.944881e-08, -1.920235e-08,
  -2.284581e-08, -2.289007e-08, -2.293278e-08, -2.289978e-08, -2.286211e-08, 
    -2.278885e-08, -2.278449e-08, -2.278825e-08, -2.285112e-08, 
    -2.286344e-08, -2.278242e-08, -2.2535e-08, -2.219489e-08, -2.18055e-08, 
    -2.145961e-08,
  -2.183216e-08, -2.178781e-08, -2.190416e-08, -2.196876e-08, -2.210556e-08, 
    -2.217337e-08, -2.236924e-08, -2.248921e-08, -2.27029e-08, -2.285049e-08, 
    -2.299206e-08, -2.306e-08, -2.306685e-08, -2.29082e-08, -2.271545e-08,
  -2.11789e-08, -2.088241e-08, -2.090221e-08, -2.084918e-08, -2.095528e-08, 
    -2.101941e-08, -2.119081e-08, -2.134607e-08, -2.158308e-08, 
    -2.185005e-08, -2.2141e-08, -2.234977e-08, -2.25114e-08, -2.262374e-08, 
    -2.268811e-08,
  -2.110936e-08, -2.079339e-08, -2.063759e-08, -2.042996e-08, -2.036852e-08, 
    -2.024636e-08, -2.020126e-08, -2.014367e-08, -2.016493e-08, 
    -2.027775e-08, -2.052523e-08, -2.079786e-08, -2.102936e-08, 
    -2.120516e-08, -2.131005e-08,
  -2.162548e-08, -2.129393e-08, -2.116461e-08, -2.09747e-08, -2.097948e-08, 
    -2.0846e-08, -2.078745e-08, -2.059345e-08, -2.044461e-08, -2.030531e-08, 
    -2.025701e-08, -2.029401e-08, -2.041259e-08, -2.057361e-08, -2.071543e-08,
  -2.280331e-08, -2.252931e-08, -2.23973e-08, -2.22741e-08, -2.23114e-08, 
    -2.220606e-08, -2.208745e-08, -2.186891e-08, -2.172273e-08, 
    -2.155848e-08, -2.142169e-08, -2.130481e-08, -2.124439e-08, 
    -2.124806e-08, -2.127187e-08,
  -2.301055e-08, -2.28805e-08, -2.278503e-08, -2.2765e-08, -2.279696e-08, 
    -2.269392e-08, -2.257857e-08, -2.244069e-08, -2.229008e-08, 
    -2.209356e-08, -2.190627e-08, -2.175984e-08, -2.166984e-08, 
    -2.165186e-08, -2.164693e-08,
  -2.272467e-08, -2.270079e-08, -2.27214e-08, -2.269621e-08, -2.273924e-08, 
    -2.257186e-08, -2.241991e-08, -2.222478e-08, -2.204564e-08, 
    -2.183558e-08, -2.163778e-08, -2.148629e-08, -2.136917e-08, 
    -2.134506e-08, -2.142058e-08,
  -1.972104e-08, -1.90458e-08, -1.872784e-08, -1.823405e-08, -1.798914e-08, 
    -1.774129e-08, -1.757065e-08, -1.743777e-08, -1.742445e-08, 
    -1.750445e-08, -1.768957e-08, -1.801267e-08, -1.847354e-08, 
    -1.897374e-08, -1.952642e-08,
  -2.120748e-08, -2.050583e-08, -2.024268e-08, -1.975152e-08, -1.951588e-08, 
    -1.925383e-08, -1.923783e-08, -1.927045e-08, -1.946454e-08, 
    -1.957473e-08, -1.967913e-08, -1.97925e-08, -1.999582e-08, -2.020794e-08, 
    -2.046308e-08,
  -2.173278e-08, -2.110788e-08, -2.083284e-08, -2.045538e-08, -2.016461e-08, 
    -1.986618e-08, -1.952714e-08, -1.918278e-08, -1.886018e-08, 
    -1.873298e-08, -1.874412e-08, -1.891618e-08, -1.922706e-08, 
    -1.951196e-08, -1.972701e-08,
  -2.16623e-08, -2.160121e-08, -2.123844e-08, -2.100476e-08, -2.074292e-08, 
    -2.052638e-08, -2.030667e-08, -2.00645e-08, -1.978416e-08, -1.946725e-08, 
    -1.918876e-08, -1.902031e-08, -1.894594e-08, -1.897704e-08, -1.911459e-08,
  -2.130404e-08, -2.123863e-08, -2.114302e-08, -2.10093e-08, -2.090064e-08, 
    -2.073756e-08, -2.064847e-08, -2.055536e-08, -2.038989e-08, 
    -2.014166e-08, -1.985315e-08, -1.959008e-08, -1.941025e-08, 
    -1.930222e-08, -1.928206e-08,
  -2.09541e-08, -2.076724e-08, -2.063734e-08, -2.057442e-08, -2.060522e-08, 
    -2.052199e-08, -2.051777e-08, -2.048735e-08, -2.05338e-08, -2.049772e-08, 
    -2.028989e-08, -2.00143e-08, -1.974294e-08, -1.955158e-08, -1.946243e-08,
  -2.117392e-08, -2.094608e-08, -2.070581e-08, -2.047772e-08, -2.043742e-08, 
    -2.033902e-08, -2.027787e-08, -2.031769e-08, -2.035499e-08, 
    -2.043399e-08, -2.040468e-08, -2.025145e-08, -2.000347e-08, 
    -1.974471e-08, -1.951822e-08,
  -2.083593e-08, -2.087048e-08, -2.073352e-08, -2.053728e-08, -2.043143e-08, 
    -2.043356e-08, -2.043896e-08, -2.049519e-08, -2.05232e-08, -2.055574e-08, 
    -2.051924e-08, -2.04079e-08, -2.022722e-08, -1.997056e-08, -1.97394e-08,
  -2.076359e-08, -2.078328e-08, -2.084008e-08, -2.06444e-08, -2.041029e-08, 
    -2.02956e-08, -2.034858e-08, -2.045668e-08, -2.056326e-08, -2.064831e-08, 
    -2.063339e-08, -2.052133e-08, -2.034975e-08, -2.010411e-08, -1.988641e-08,
  -2.091228e-08, -2.105916e-08, -2.12016e-08, -2.113528e-08, -2.095087e-08, 
    -2.066345e-08, -2.052252e-08, -2.048476e-08, -2.052811e-08, 
    -2.054403e-08, -2.056068e-08, -2.048837e-08, -2.035721e-08, 
    -2.008365e-08, -1.976617e-08,
  -1.867052e-08, -1.951392e-08, -1.983235e-08, -2.048493e-08, -2.164935e-08, 
    -2.273213e-08, -2.346458e-08, -2.430741e-08, -2.492793e-08, -2.54171e-08, 
    -2.575741e-08, -2.597242e-08, -2.616525e-08, -2.619717e-08, -2.621194e-08,
  -2.003091e-08, -2.083723e-08, -2.132186e-08, -2.204663e-08, -2.293046e-08, 
    -2.349548e-08, -2.419742e-08, -2.473891e-08, -2.522248e-08, 
    -2.559788e-08, -2.588102e-08, -2.608414e-08, -2.626975e-08, 
    -2.617385e-08, -2.599462e-08,
  -2.098851e-08, -2.163128e-08, -2.214248e-08, -2.289383e-08, -2.370982e-08, 
    -2.414155e-08, -2.457261e-08, -2.495339e-08, -2.545578e-08, 
    -2.589177e-08, -2.61777e-08, -2.617774e-08, -2.608376e-08, -2.57312e-08, 
    -2.524356e-08,
  -2.134696e-08, -2.184607e-08, -2.224403e-08, -2.322773e-08, -2.406376e-08, 
    -2.435198e-08, -2.48091e-08, -2.517451e-08, -2.565135e-08, -2.608189e-08, 
    -2.61756e-08, -2.599882e-08, -2.567483e-08, -2.516396e-08, -2.48032e-08,
  -2.167601e-08, -2.1968e-08, -2.217627e-08, -2.305977e-08, -2.385572e-08, 
    -2.424453e-08, -2.480923e-08, -2.506486e-08, -2.56141e-08, -2.58962e-08, 
    -2.584268e-08, -2.558886e-08, -2.509808e-08, -2.467822e-08, -2.450264e-08,
  -2.128147e-08, -2.176085e-08, -2.220878e-08, -2.26997e-08, -2.330811e-08, 
    -2.410384e-08, -2.458602e-08, -2.495751e-08, -2.538788e-08, 
    -2.547853e-08, -2.539577e-08, -2.49551e-08, -2.452725e-08, -2.433814e-08, 
    -2.432517e-08,
  -2.098073e-08, -2.164363e-08, -2.215989e-08, -2.249258e-08, -2.315435e-08, 
    -2.384134e-08, -2.425005e-08, -2.462884e-08, -2.501056e-08, 
    -2.512224e-08, -2.498198e-08, -2.460941e-08, -2.424091e-08, 
    -2.407332e-08, -2.403018e-08,
  -2.075651e-08, -2.1345e-08, -2.181863e-08, -2.234237e-08, -2.311295e-08, 
    -2.374772e-08, -2.403815e-08, -2.435737e-08, -2.459522e-08, -2.46089e-08, 
    -2.447434e-08, -2.415305e-08, -2.386309e-08, -2.373623e-08, -2.391668e-08,
  -2.070182e-08, -2.121607e-08, -2.150049e-08, -2.200621e-08, -2.289862e-08, 
    -2.351211e-08, -2.386448e-08, -2.422356e-08, -2.439895e-08, 
    -2.435393e-08, -2.412941e-08, -2.3901e-08, -2.366586e-08, -2.358843e-08, 
    -2.380823e-08,
  -2.074955e-08, -2.108927e-08, -2.139596e-08, -2.17595e-08, -2.250629e-08, 
    -2.319713e-08, -2.375476e-08, -2.415215e-08, -2.431367e-08, 
    -2.426916e-08, -2.402196e-08, -2.378063e-08, -2.358694e-08, 
    -2.352375e-08, -2.364681e-08,
  -2.589313e-08, -2.616602e-08, -2.548349e-08, -2.63448e-08, -2.557942e-08, 
    -2.57041e-08, -2.514335e-08, -2.486918e-08, -2.435899e-08, -2.397304e-08, 
    -2.367644e-08, -2.335243e-08, -2.312198e-08, -2.27064e-08, -2.238279e-08,
  -2.725829e-08, -2.690136e-08, -2.657158e-08, -2.643658e-08, -2.611017e-08, 
    -2.604364e-08, -2.522379e-08, -2.496318e-08, -2.443114e-08, 
    -2.400303e-08, -2.374346e-08, -2.363113e-08, -2.342364e-08, 
    -2.314467e-08, -2.286761e-08,
  -2.749251e-08, -2.819803e-08, -2.726987e-08, -2.721471e-08, -2.665387e-08, 
    -2.644365e-08, -2.571519e-08, -2.512873e-08, -2.450666e-08, 
    -2.396668e-08, -2.376914e-08, -2.354536e-08, -2.344093e-08, -2.32163e-08, 
    -2.303225e-08,
  -2.747287e-08, -2.777714e-08, -2.796396e-08, -2.737731e-08, -2.725376e-08, 
    -2.685842e-08, -2.608133e-08, -2.524737e-08, -2.444452e-08, 
    -2.380947e-08, -2.350039e-08, -2.322186e-08, -2.331909e-08, 
    -2.313111e-08, -2.300565e-08,
  -2.788784e-08, -2.719649e-08, -2.711403e-08, -2.745798e-08, -2.776464e-08, 
    -2.725971e-08, -2.65266e-08, -2.567563e-08, -2.449711e-08, -2.361546e-08, 
    -2.332468e-08, -2.3208e-08, -2.337666e-08, -2.336624e-08, -2.315602e-08,
  -2.84728e-08, -2.771085e-08, -2.718086e-08, -2.802648e-08, -2.760771e-08, 
    -2.73151e-08, -2.701697e-08, -2.604239e-08, -2.476538e-08, -2.360489e-08, 
    -2.332602e-08, -2.320964e-08, -2.34873e-08, -2.372639e-08, -2.356536e-08,
  -2.856039e-08, -2.803346e-08, -2.737767e-08, -2.805099e-08, -2.731319e-08, 
    -2.721328e-08, -2.732969e-08, -2.644834e-08, -2.510513e-08, 
    -2.380372e-08, -2.325976e-08, -2.328465e-08, -2.373615e-08, 
    -2.408737e-08, -2.406886e-08,
  -2.930795e-08, -2.825137e-08, -2.743255e-08, -2.724014e-08, -2.654767e-08, 
    -2.733512e-08, -2.750718e-08, -2.676341e-08, -2.558658e-08, 
    -2.401555e-08, -2.335909e-08, -2.348533e-08, -2.392347e-08, 
    -2.431499e-08, -2.434097e-08,
  -3.005641e-08, -2.865598e-08, -2.682006e-08, -2.590655e-08, -2.628551e-08, 
    -2.728968e-08, -2.751102e-08, -2.696998e-08, -2.601525e-08, 
    -2.432486e-08, -2.364759e-08, -2.35787e-08, -2.399562e-08, -2.434568e-08, 
    -2.439522e-08,
  -3.047385e-08, -2.897889e-08, -2.666384e-08, -2.514314e-08, -2.559057e-08, 
    -2.720916e-08, -2.758969e-08, -2.720421e-08, -2.643211e-08, 
    -2.466549e-08, -2.394794e-08, -2.37301e-08, -2.403367e-08, -2.422181e-08, 
    -2.429491e-08,
  -2.169508e-08, -2.115349e-08, -2.064325e-08, -2.043132e-08, -2.014837e-08, 
    -1.999176e-08, -1.981339e-08, -1.971927e-08, -1.95366e-08, -1.937034e-08, 
    -1.91467e-08, -1.89998e-08, -1.887785e-08, -1.881082e-08, -1.877938e-08,
  -2.222204e-08, -2.190767e-08, -2.15422e-08, -2.106731e-08, -2.09711e-08, 
    -2.075824e-08, -2.073589e-08, -2.065374e-08, -2.060997e-08, 
    -2.051404e-08, -2.041482e-08, -2.028447e-08, -2.020181e-08, -2.01484e-08, 
    -2.009525e-08,
  -2.255224e-08, -2.247245e-08, -2.190056e-08, -2.142229e-08, -2.127809e-08, 
    -2.106534e-08, -2.102829e-08, -2.099892e-08, -2.09999e-08, -2.098322e-08, 
    -2.099231e-08, -2.097687e-08, -2.0931e-08, -2.090623e-08, -2.088525e-08,
  -2.361165e-08, -2.307846e-08, -2.240955e-08, -2.206977e-08, -2.162234e-08, 
    -2.154461e-08, -2.144409e-08, -2.144571e-08, -2.146748e-08, 
    -2.150878e-08, -2.15528e-08, -2.161189e-08, -2.153555e-08, -2.153563e-08, 
    -2.147581e-08,
  -2.483555e-08, -2.426226e-08, -2.355837e-08, -2.265951e-08, -2.244392e-08, 
    -2.217744e-08, -2.215108e-08, -2.224825e-08, -2.253307e-08, 
    -2.261113e-08, -2.292066e-08, -2.307452e-08, -2.313307e-08, 
    -2.314093e-08, -2.312187e-08,
  -2.557259e-08, -2.500418e-08, -2.412848e-08, -2.347599e-08, -2.302513e-08, 
    -2.277759e-08, -2.260095e-08, -2.272623e-08, -2.315011e-08, 
    -2.338717e-08, -2.386172e-08, -2.407258e-08, -2.434744e-08, 
    -2.439707e-08, -2.448101e-08,
  -2.544889e-08, -2.555916e-08, -2.47375e-08, -2.396541e-08, -2.378358e-08, 
    -2.350664e-08, -2.317715e-08, -2.320911e-08, -2.337521e-08, -2.36647e-08, 
    -2.388984e-08, -2.407351e-08, -2.399879e-08, -2.407784e-08, -2.395898e-08,
  -2.571417e-08, -2.599342e-08, -2.514431e-08, -2.4147e-08, -2.430873e-08, 
    -2.401242e-08, -2.355995e-08, -2.330522e-08, -2.316156e-08, -2.34175e-08, 
    -2.360129e-08, -2.356885e-08, -2.361119e-08, -2.34062e-08, -2.351346e-08,
  -2.580118e-08, -2.654877e-08, -2.591063e-08, -2.437181e-08, -2.462921e-08, 
    -2.427928e-08, -2.381262e-08, -2.361699e-08, -2.321577e-08, 
    -2.323708e-08, -2.341457e-08, -2.344282e-08, -2.336282e-08, 
    -2.323897e-08, -2.351318e-08,
  -2.666439e-08, -2.73224e-08, -2.713328e-08, -2.48419e-08, -2.435942e-08, 
    -2.480539e-08, -2.4524e-08, -2.393809e-08, -2.343688e-08, -2.317934e-08, 
    -2.326183e-08, -2.336119e-08, -2.318492e-08, -2.312753e-08, -2.356832e-08,
  -2.054163e-08, -2.029231e-08, -2.025059e-08, -2.017602e-08, -2.01571e-08, 
    -2.014522e-08, -2.017293e-08, -2.021047e-08, -2.028216e-08, 
    -2.036209e-08, -2.048679e-08, -2.067352e-08, -2.091762e-08, 
    -2.119592e-08, -2.151102e-08,
  -2.226973e-08, -2.217628e-08, -2.202809e-08, -2.205865e-08, -2.197992e-08, 
    -2.20832e-08, -2.207397e-08, -2.215469e-08, -2.221725e-08, -2.232395e-08, 
    -2.243874e-08, -2.259202e-08, -2.27467e-08, -2.292255e-08, -2.309896e-08,
  -2.336483e-08, -2.338021e-08, -2.348285e-08, -2.344226e-08, -2.34333e-08, 
    -2.348966e-08, -2.357421e-08, -2.361418e-08, -2.367361e-08, 
    -2.372905e-08, -2.380317e-08, -2.386108e-08, -2.393249e-08, -2.39986e-08, 
    -2.40809e-08,
  -2.399638e-08, -2.398018e-08, -2.425401e-08, -2.436242e-08, -2.453758e-08, 
    -2.462895e-08, -2.474855e-08, -2.486735e-08, -2.493608e-08, 
    -2.500157e-08, -2.504425e-08, -2.506366e-08, -2.506357e-08, 
    -2.507737e-08, -2.507986e-08,
  -2.449129e-08, -2.436742e-08, -2.468977e-08, -2.476174e-08, -2.507919e-08, 
    -2.529972e-08, -2.546088e-08, -2.566685e-08, -2.588241e-08, 
    -2.595718e-08, -2.599968e-08, -2.596641e-08, -2.592679e-08, 
    -2.589991e-08, -2.584031e-08,
  -2.478874e-08, -2.480613e-08, -2.507242e-08, -2.521084e-08, -2.545489e-08, 
    -2.566501e-08, -2.591923e-08, -2.617273e-08, -2.641556e-08, 
    -2.649884e-08, -2.646864e-08, -2.639543e-08, -2.642199e-08, 
    -2.632098e-08, -2.625601e-08,
  -2.47994e-08, -2.487207e-08, -2.516746e-08, -2.530315e-08, -2.558668e-08, 
    -2.577295e-08, -2.615782e-08, -2.643449e-08, -2.658854e-08, 
    -2.665704e-08, -2.651895e-08, -2.650114e-08, -2.644168e-08, 
    -2.655414e-08, -2.631309e-08,
  -2.45519e-08, -2.477486e-08, -2.494985e-08, -2.510677e-08, -2.544809e-08, 
    -2.562808e-08, -2.592184e-08, -2.633416e-08, -2.656587e-08, 
    -2.650234e-08, -2.649007e-08, -2.637487e-08, -2.641761e-08, 
    -2.658922e-08, -2.655596e-08,
  -2.437326e-08, -2.451779e-08, -2.489895e-08, -2.532594e-08, -2.538883e-08, 
    -2.557571e-08, -2.577615e-08, -2.623537e-08, -2.632994e-08, 
    -2.644667e-08, -2.635201e-08, -2.616615e-08, -2.638346e-08, 
    -2.661346e-08, -2.683249e-08,
  -2.434986e-08, -2.473157e-08, -2.526002e-08, -2.523871e-08, -2.540684e-08, 
    -2.535491e-08, -2.579662e-08, -2.604301e-08, -2.608713e-08, 
    -2.668589e-08, -2.619858e-08, -2.633835e-08, -2.623507e-08, 
    -2.657553e-08, -2.685492e-08,
  -2.515673e-08, -2.479596e-08, -2.472556e-08, -2.451918e-08, -2.445336e-08, 
    -2.420093e-08, -2.399216e-08, -2.373324e-08, -2.346367e-08, 
    -2.314007e-08, -2.28436e-08, -2.252929e-08, -2.222022e-08, -2.198517e-08, 
    -2.204358e-08,
  -2.531193e-08, -2.50124e-08, -2.493181e-08, -2.465135e-08, -2.452516e-08, 
    -2.429495e-08, -2.401399e-08, -2.371865e-08, -2.339292e-08, 
    -2.297636e-08, -2.262803e-08, -2.231321e-08, -2.202912e-08, 
    -2.177291e-08, -2.150346e-08,
  -2.544301e-08, -2.504091e-08, -2.488255e-08, -2.463275e-08, -2.452483e-08, 
    -2.431449e-08, -2.412759e-08, -2.388467e-08, -2.365317e-08, 
    -2.326384e-08, -2.282331e-08, -2.235089e-08, -2.199151e-08, 
    -2.173928e-08, -2.146781e-08,
  -2.643887e-08, -2.60095e-08, -2.566477e-08, -2.534429e-08, -2.509086e-08, 
    -2.489963e-08, -2.477064e-08, -2.466932e-08, -2.454969e-08, 
    -2.418783e-08, -2.376835e-08, -2.332858e-08, -2.294351e-08, 
    -2.267793e-08, -2.244216e-08,
  -2.748717e-08, -2.68844e-08, -2.639013e-08, -2.603066e-08, -2.571529e-08, 
    -2.542247e-08, -2.531963e-08, -2.52564e-08, -2.528046e-08, -2.503767e-08, 
    -2.462128e-08, -2.416964e-08, -2.360486e-08, -2.315387e-08, -2.299744e-08,
  -2.80501e-08, -2.770774e-08, -2.714746e-08, -2.673823e-08, -2.64481e-08, 
    -2.60864e-08, -2.59321e-08, -2.571774e-08, -2.573779e-08, -2.573387e-08, 
    -2.552495e-08, -2.525065e-08, -2.485756e-08, -2.423971e-08, -2.384805e-08,
  -2.807439e-08, -2.809187e-08, -2.752772e-08, -2.704159e-08, -2.682217e-08, 
    -2.658784e-08, -2.649914e-08, -2.629744e-08, -2.608381e-08, 
    -2.576883e-08, -2.559771e-08, -2.541847e-08, -2.520853e-08, -2.48324e-08, 
    -2.436873e-08,
  -2.741491e-08, -2.779679e-08, -2.794953e-08, -2.762785e-08, -2.700212e-08, 
    -2.665256e-08, -2.657808e-08, -2.670428e-08, -2.671362e-08, 
    -2.659855e-08, -2.624952e-08, -2.59841e-08, -2.56365e-08, -2.522065e-08, 
    -2.479791e-08,
  -2.659816e-08, -2.690266e-08, -2.743573e-08, -2.767119e-08, -2.747002e-08, 
    -2.688272e-08, -2.658812e-08, -2.660512e-08, -2.6859e-08, -2.703796e-08, 
    -2.695122e-08, -2.67693e-08, -2.650091e-08, -2.612099e-08, -2.561884e-08,
  -2.603071e-08, -2.647142e-08, -2.688176e-08, -2.715388e-08, -2.724591e-08, 
    -2.706875e-08, -2.671106e-08, -2.637352e-08, -2.66402e-08, -2.698409e-08, 
    -2.726861e-08, -2.722649e-08, -2.713782e-08, -2.692306e-08, -2.660765e-08,
  -2.087649e-08, -2.081257e-08, -2.082134e-08, -2.088435e-08, -2.089383e-08, 
    -2.085218e-08, -2.080461e-08, -2.07331e-08, -2.067822e-08, -2.054899e-08, 
    -2.036664e-08, -2.009598e-08, -1.98445e-08, -1.959389e-08, -1.931126e-08,
  -2.113528e-08, -2.086952e-08, -2.081615e-08, -2.075628e-08, -2.079904e-08, 
    -2.083035e-08, -2.087652e-08, -2.087616e-08, -2.095207e-08, 
    -2.097954e-08, -2.098606e-08, -2.09144e-08, -2.076706e-08, -2.061308e-08, 
    -2.042889e-08,
  -2.206696e-08, -2.157507e-08, -2.139694e-08, -2.111861e-08, -2.102201e-08, 
    -2.091698e-08, -2.078109e-08, -2.059057e-08, -2.043236e-08, 
    -2.046072e-08, -2.049675e-08, -2.061428e-08, -2.070365e-08, 
    -2.080032e-08, -2.087898e-08,
  -2.294696e-08, -2.27019e-08, -2.24569e-08, -2.225897e-08, -2.205417e-08, 
    -2.199305e-08, -2.190371e-08, -2.178151e-08, -2.160105e-08, 
    -2.152929e-08, -2.159605e-08, -2.174171e-08, -2.18988e-08, -2.208001e-08, 
    -2.220979e-08,
  -2.314763e-08, -2.325896e-08, -2.310305e-08, -2.306718e-08, -2.284851e-08, 
    -2.279699e-08, -2.278948e-08, -2.284156e-08, -2.279219e-08, 
    -2.270503e-08, -2.268565e-08, -2.274924e-08, -2.276258e-08, 
    -2.285784e-08, -2.297009e-08,
  -2.336895e-08, -2.329591e-08, -2.313955e-08, -2.296933e-08, -2.272546e-08, 
    -2.254197e-08, -2.245923e-08, -2.241974e-08, -2.242184e-08, 
    -2.239996e-08, -2.237064e-08, -2.24145e-08, -2.251664e-08, -2.262449e-08, 
    -2.274691e-08,
  -2.356979e-08, -2.343793e-08, -2.312687e-08, -2.300433e-08, -2.268191e-08, 
    -2.225762e-08, -2.2055e-08, -2.200299e-08, -2.203887e-08, -2.212936e-08, 
    -2.21993e-08, -2.224945e-08, -2.233151e-08, -2.249942e-08, -2.267689e-08,
  -2.357672e-08, -2.361677e-08, -2.319295e-08, -2.296094e-08, -2.279137e-08, 
    -2.252233e-08, -2.212491e-08, -2.185132e-08, -2.183218e-08, 
    -2.189783e-08, -2.196362e-08, -2.211351e-08, -2.219429e-08, 
    -2.230513e-08, -2.244727e-08,
  -2.391564e-08, -2.361403e-08, -2.329938e-08, -2.290242e-08, -2.265388e-08, 
    -2.251575e-08, -2.231066e-08, -2.210396e-08, -2.175709e-08, 
    -2.177257e-08, -2.187678e-08, -2.203257e-08, -2.219428e-08, 
    -2.231227e-08, -2.2423e-08,
  -2.415104e-08, -2.361131e-08, -2.331911e-08, -2.291157e-08, -2.269882e-08, 
    -2.250846e-08, -2.234425e-08, -2.219322e-08, -2.202361e-08, 
    -2.181227e-08, -2.187879e-08, -2.208833e-08, -2.234513e-08, 
    -2.260872e-08, -2.281258e-08,
  -2.344441e-08, -2.296623e-08, -2.247533e-08, -2.199967e-08, -2.165609e-08, 
    -2.146122e-08, -2.175673e-08, -2.209392e-08, -2.280448e-08, 
    -2.350124e-08, -2.38326e-08, -2.383597e-08, -2.351745e-08, -2.292484e-08, 
    -2.233132e-08,
  -2.551214e-08, -2.409393e-08, -2.374503e-08, -2.329394e-08, -2.33978e-08, 
    -2.361631e-08, -2.398342e-08, -2.425603e-08, -2.442761e-08, 
    -2.440459e-08, -2.413906e-08, -2.393533e-08, -2.354979e-08, 
    -2.335782e-08, -2.305468e-08,
  -2.339423e-08, -2.344552e-08, -2.380964e-08, -2.372512e-08, -2.415812e-08, 
    -2.418372e-08, -2.436609e-08, -2.435007e-08, -2.431007e-08, -2.42075e-08, 
    -2.406057e-08, -2.396245e-08, -2.390118e-08, -2.392167e-08, -2.394841e-08,
  -2.336925e-08, -2.39627e-08, -2.427011e-08, -2.429478e-08, -2.466451e-08, 
    -2.470018e-08, -2.472803e-08, -2.467327e-08, -2.464844e-08, 
    -2.469319e-08, -2.473573e-08, -2.484069e-08, -2.490885e-08, 
    -2.497426e-08, -2.506112e-08,
  -2.505879e-08, -2.563147e-08, -2.579928e-08, -2.588908e-08, -2.581235e-08, 
    -2.566814e-08, -2.554304e-08, -2.552442e-08, -2.548217e-08, 
    -2.553039e-08, -2.558513e-08, -2.570957e-08, -2.583998e-08, 
    -2.596522e-08, -2.610583e-08,
  -2.576324e-08, -2.600141e-08, -2.5616e-08, -2.561539e-08, -2.537977e-08, 
    -2.541972e-08, -2.542713e-08, -2.559531e-08, -2.572119e-08, 
    -2.583937e-08, -2.599614e-08, -2.607281e-08, -2.618285e-08, 
    -2.623427e-08, -2.621927e-08,
  -2.53876e-08, -2.559012e-08, -2.547522e-08, -2.561308e-08, -2.568131e-08, 
    -2.591901e-08, -2.634637e-08, -2.655764e-08, -2.673418e-08, -2.67861e-08, 
    -2.685423e-08, -2.694362e-08, -2.700357e-08, -2.685519e-08, -2.66591e-08,
  -2.527603e-08, -2.539154e-08, -2.557326e-08, -2.580498e-08, -2.611171e-08, 
    -2.648169e-08, -2.690203e-08, -2.704832e-08, -2.717361e-08, 
    -2.722233e-08, -2.727847e-08, -2.725359e-08, -2.722328e-08, 
    -2.698895e-08, -2.677348e-08,
  -2.508845e-08, -2.525911e-08, -2.563056e-08, -2.599338e-08, -2.643066e-08, 
    -2.683162e-08, -2.714449e-08, -2.722106e-08, -2.724491e-08, 
    -2.720045e-08, -2.717407e-08, -2.712267e-08, -2.69971e-08, -2.680216e-08, 
    -2.668966e-08,
  -2.475877e-08, -2.518104e-08, -2.573509e-08, -2.624301e-08, -2.676957e-08, 
    -2.703631e-08, -2.726118e-08, -2.727951e-08, -2.730171e-08, 
    -2.729078e-08, -2.723805e-08, -2.719143e-08, -2.712542e-08, 
    -2.706167e-08, -2.710037e-08,
  -2.242925e-08, -2.219793e-08, -2.200393e-08, -2.192262e-08, -2.220196e-08, 
    -2.287532e-08, -2.358058e-08, -2.423799e-08, -2.467132e-08, 
    -2.493235e-08, -2.505425e-08, -2.507435e-08, -2.500208e-08, 
    -2.485378e-08, -2.468605e-08,
  -2.260994e-08, -2.246071e-08, -2.293694e-08, -2.354689e-08, -2.433876e-08, 
    -2.501034e-08, -2.549321e-08, -2.564636e-08, -2.587088e-08, 
    -2.589627e-08, -2.606249e-08, -2.613793e-08, -2.613246e-08, -2.6009e-08, 
    -2.586334e-08,
  -2.354823e-08, -2.372035e-08, -2.449428e-08, -2.498088e-08, -2.556986e-08, 
    -2.573222e-08, -2.560027e-08, -2.538478e-08, -2.52077e-08, -2.515361e-08, 
    -2.510078e-08, -2.513596e-08, -2.523449e-08, -2.529863e-08, -2.530279e-08,
  -2.421495e-08, -2.463363e-08, -2.528092e-08, -2.5488e-08, -2.497937e-08, 
    -2.482628e-08, -2.4257e-08, -2.409279e-08, -2.377712e-08, -2.359061e-08, 
    -2.345206e-08, -2.341995e-08, -2.358195e-08, -2.379906e-08, -2.411023e-08,
  -2.470549e-08, -2.533917e-08, -2.564566e-08, -2.527002e-08, -2.500401e-08, 
    -2.457421e-08, -2.423307e-08, -2.369025e-08, -2.329237e-08, 
    -2.283408e-08, -2.261092e-08, -2.270935e-08, -2.302913e-08, 
    -2.346247e-08, -2.39048e-08,
  -2.560029e-08, -2.636314e-08, -2.605911e-08, -2.581805e-08, -2.550836e-08, 
    -2.509258e-08, -2.459205e-08, -2.423142e-08, -2.375512e-08, -2.34518e-08, 
    -2.370756e-08, -2.403575e-08, -2.449001e-08, -2.473156e-08, -2.484337e-08,
  -2.658239e-08, -2.661563e-08, -2.558324e-08, -2.559504e-08, -2.489874e-08, 
    -2.452524e-08, -2.402626e-08, -2.374676e-08, -2.386951e-08, 
    -2.435933e-08, -2.479399e-08, -2.516674e-08, -2.511645e-08, 
    -2.536046e-08, -2.519976e-08,
  -2.653407e-08, -2.578825e-08, -2.541287e-08, -2.50719e-08, -2.454444e-08, 
    -2.423881e-08, -2.403073e-08, -2.44601e-08, -2.490544e-08, -2.516557e-08, 
    -2.523015e-08, -2.504576e-08, -2.490487e-08, -2.496148e-08, -2.490287e-08,
  -2.628712e-08, -2.552331e-08, -2.553276e-08, -2.482417e-08, -2.485874e-08, 
    -2.452454e-08, -2.496791e-08, -2.522545e-08, -2.548879e-08, 
    -2.539972e-08, -2.525007e-08, -2.5144e-08, -2.512975e-08, -2.518333e-08, 
    -2.518866e-08,
  -2.609808e-08, -2.574068e-08, -2.546872e-08, -2.511127e-08, -2.517691e-08, 
    -2.518596e-08, -2.5615e-08, -2.57413e-08, -2.597725e-08, -2.589536e-08, 
    -2.583509e-08, -2.585985e-08, -2.589874e-08, -2.596094e-08, -2.598022e-08,
  -2.273945e-08, -2.279285e-08, -2.250094e-08, -2.237411e-08, -2.220334e-08, 
    -2.212038e-08, -2.208562e-08, -2.191016e-08, -2.172893e-08, 
    -2.156869e-08, -2.142316e-08, -2.134771e-08, -2.133293e-08, 
    -2.137404e-08, -2.144721e-08,
  -2.31851e-08, -2.310151e-08, -2.277089e-08, -2.279391e-08, -2.271693e-08, 
    -2.266569e-08, -2.253374e-08, -2.21891e-08, -2.183009e-08, -2.156004e-08, 
    -2.135418e-08, -2.119248e-08, -2.114566e-08, -2.115786e-08, -2.118907e-08,
  -2.354008e-08, -2.339784e-08, -2.316011e-08, -2.33732e-08, -2.351388e-08, 
    -2.35103e-08, -2.31476e-08, -2.283466e-08, -2.258829e-08, -2.241279e-08, 
    -2.225686e-08, -2.212144e-08, -2.2014e-08, -2.194665e-08, -2.192655e-08,
  -2.377484e-08, -2.37596e-08, -2.391145e-08, -2.418602e-08, -2.42414e-08, 
    -2.396408e-08, -2.350859e-08, -2.335272e-08, -2.309592e-08, 
    -2.299452e-08, -2.281863e-08, -2.264123e-08, -2.246566e-08, 
    -2.229278e-08, -2.217977e-08,
  -2.407498e-08, -2.399377e-08, -2.436508e-08, -2.441879e-08, -2.412136e-08, 
    -2.369545e-08, -2.364022e-08, -2.360039e-08, -2.341247e-08, 
    -2.333607e-08, -2.302741e-08, -2.286002e-08, -2.258893e-08, 
    -2.244533e-08, -2.217947e-08,
  -2.432499e-08, -2.434971e-08, -2.470143e-08, -2.451867e-08, -2.392057e-08, 
    -2.383089e-08, -2.377882e-08, -2.35891e-08, -2.33671e-08, -2.29249e-08, 
    -2.256128e-08, -2.226629e-08, -2.215096e-08, -2.200664e-08, -2.190791e-08,
  -2.465097e-08, -2.462528e-08, -2.485757e-08, -2.425235e-08, -2.359423e-08, 
    -2.366945e-08, -2.346994e-08, -2.332442e-08, -2.278573e-08, 
    -2.247216e-08, -2.237804e-08, -2.240881e-08, -2.249874e-08, -2.24976e-08, 
    -2.248252e-08,
  -2.497432e-08, -2.488984e-08, -2.473867e-08, -2.370325e-08, -2.331721e-08, 
    -2.340611e-08, -2.330978e-08, -2.275931e-08, -2.257197e-08, 
    -2.260385e-08, -2.286179e-08, -2.314817e-08, -2.335381e-08, -2.34536e-08, 
    -2.359319e-08,
  -2.511208e-08, -2.497273e-08, -2.437114e-08, -2.334261e-08, -2.314303e-08, 
    -2.307685e-08, -2.274922e-08, -2.260175e-08, -2.297179e-08, 
    -2.341617e-08, -2.383239e-08, -2.405308e-08, -2.414479e-08, 
    -2.421237e-08, -2.421641e-08,
  -2.505245e-08, -2.482311e-08, -2.393865e-08, -2.305731e-08, -2.284991e-08, 
    -2.270448e-08, -2.277658e-08, -2.322664e-08, -2.391134e-08, 
    -2.408387e-08, -2.411775e-08, -2.377076e-08, -2.349906e-08, 
    -2.311535e-08, -2.294046e-08,
  -2.260194e-08, -2.249369e-08, -2.255375e-08, -2.248941e-08, -2.237805e-08, 
    -2.23158e-08, -2.219567e-08, -2.210522e-08, -2.201651e-08, -2.197879e-08, 
    -2.193597e-08, -2.198548e-08, -2.199113e-08, -2.201911e-08, -2.203474e-08,
  -2.287728e-08, -2.263307e-08, -2.250973e-08, -2.228282e-08, -2.2208e-08, 
    -2.21018e-08, -2.201734e-08, -2.194101e-08, -2.183828e-08, -2.178593e-08, 
    -2.179842e-08, -2.184457e-08, -2.18938e-08, -2.193921e-08, -2.20509e-08,
  -2.298406e-08, -2.250757e-08, -2.21758e-08, -2.191359e-08, -2.180786e-08, 
    -2.173741e-08, -2.168356e-08, -2.163607e-08, -2.162828e-08, 
    -2.161917e-08, -2.175487e-08, -2.182671e-08, -2.196615e-08, 
    -2.194631e-08, -2.201125e-08,
  -2.280868e-08, -2.236183e-08, -2.185134e-08, -2.145019e-08, -2.155492e-08, 
    -2.154104e-08, -2.15859e-08, -2.151086e-08, -2.159811e-08, -2.182061e-08, 
    -2.207359e-08, -2.223693e-08, -2.224587e-08, -2.222358e-08, -2.21305e-08,
  -2.302299e-08, -2.221255e-08, -2.160369e-08, -2.132251e-08, -2.14742e-08, 
    -2.145551e-08, -2.147541e-08, -2.140052e-08, -2.164779e-08, 
    -2.190947e-08, -2.221383e-08, -2.228957e-08, -2.230369e-08, 
    -2.228572e-08, -2.222436e-08,
  -2.276232e-08, -2.221329e-08, -2.16494e-08, -2.14231e-08, -2.147701e-08, 
    -2.159412e-08, -2.149717e-08, -2.146361e-08, -2.172314e-08, -2.19146e-08, 
    -2.216466e-08, -2.232303e-08, -2.2327e-08, -2.236949e-08, -2.22205e-08,
  -2.285686e-08, -2.23134e-08, -2.164413e-08, -2.151293e-08, -2.175931e-08, 
    -2.170716e-08, -2.16163e-08, -2.150105e-08, -2.162796e-08, -2.187195e-08, 
    -2.219e-08, -2.236634e-08, -2.22812e-08, -2.223744e-08, -2.213766e-08,
  -2.299122e-08, -2.244243e-08, -2.177096e-08, -2.172128e-08, -2.200405e-08, 
    -2.190266e-08, -2.161656e-08, -2.144721e-08, -2.166565e-08, 
    -2.209255e-08, -2.243113e-08, -2.259698e-08, -2.240907e-08, 
    -2.234278e-08, -2.218425e-08,
  -2.33741e-08, -2.280968e-08, -2.195995e-08, -2.182556e-08, -2.224632e-08, 
    -2.20988e-08, -2.15783e-08, -2.148425e-08, -2.19081e-08, -2.238307e-08, 
    -2.267356e-08, -2.283647e-08, -2.253094e-08, -2.245909e-08, -2.2257e-08,
  -2.428969e-08, -2.320016e-08, -2.23217e-08, -2.190963e-08, -2.241327e-08, 
    -2.216722e-08, -2.166727e-08, -2.163975e-08, -2.218259e-08, 
    -2.263842e-08, -2.287281e-08, -2.303338e-08, -2.281224e-08, 
    -2.273417e-08, -2.257724e-08,
  -2.144198e-08, -2.151229e-08, -2.146608e-08, -2.150429e-08, -2.156908e-08, 
    -2.172103e-08, -2.182053e-08, -2.185155e-08, -2.180833e-08, 
    -2.176116e-08, -2.162725e-08, -2.151451e-08, -2.137353e-08, 
    -2.131151e-08, -2.125917e-08,
  -2.186628e-08, -2.171812e-08, -2.176776e-08, -2.177258e-08, -2.184514e-08, 
    -2.191817e-08, -2.197917e-08, -2.203227e-08, -2.206928e-08, 
    -2.210308e-08, -2.208355e-08, -2.202596e-08, -2.198207e-08, 
    -2.193168e-08, -2.183231e-08,
  -2.211991e-08, -2.185368e-08, -2.189723e-08, -2.180671e-08, -2.196214e-08, 
    -2.207993e-08, -2.223587e-08, -2.245663e-08, -2.257125e-08, 
    -2.269296e-08, -2.274454e-08, -2.267036e-08, -2.260507e-08, 
    -2.250153e-08, -2.240189e-08,
  -2.233396e-08, -2.226192e-08, -2.235773e-08, -2.230794e-08, -2.24404e-08, 
    -2.251772e-08, -2.270517e-08, -2.300117e-08, -2.312359e-08, 
    -2.314845e-08, -2.309134e-08, -2.299123e-08, -2.298356e-08, 
    -2.293101e-08, -2.283302e-08,
  -2.26865e-08, -2.268714e-08, -2.265901e-08, -2.261828e-08, -2.255158e-08, 
    -2.267022e-08, -2.290844e-08, -2.319948e-08, -2.332468e-08, -2.33265e-08, 
    -2.328818e-08, -2.324089e-08, -2.326474e-08, -2.313955e-08, -2.310766e-08,
  -2.295616e-08, -2.303449e-08, -2.295218e-08, -2.293634e-08, -2.292169e-08, 
    -2.292436e-08, -2.313574e-08, -2.345442e-08, -2.355677e-08, 
    -2.356845e-08, -2.344843e-08, -2.322575e-08, -2.321499e-08, 
    -2.309372e-08, -2.316994e-08,
  -2.297956e-08, -2.313163e-08, -2.307118e-08, -2.310501e-08, -2.306806e-08, 
    -2.299434e-08, -2.306817e-08, -2.338898e-08, -2.343377e-08, 
    -2.341917e-08, -2.318963e-08, -2.282892e-08, -2.286905e-08, 
    -2.284549e-08, -2.304334e-08,
  -2.290276e-08, -2.309569e-08, -2.316181e-08, -2.326387e-08, -2.311276e-08, 
    -2.296959e-08, -2.298652e-08, -2.332326e-08, -2.341644e-08, 
    -2.344663e-08, -2.309723e-08, -2.275062e-08, -2.278368e-08, 
    -2.288253e-08, -2.309064e-08,
  -2.274093e-08, -2.303024e-08, -2.312275e-08, -2.325642e-08, -2.289214e-08, 
    -2.285474e-08, -2.288841e-08, -2.335862e-08, -2.358544e-08, 
    -2.368061e-08, -2.344762e-08, -2.31957e-08, -2.338921e-08, -2.356285e-08, 
    -2.378466e-08,
  -2.266106e-08, -2.285927e-08, -2.308034e-08, -2.315512e-08, -2.294453e-08, 
    -2.284358e-08, -2.292845e-08, -2.354082e-08, -2.401455e-08, -2.42148e-08, 
    -2.415265e-08, -2.406374e-08, -2.436042e-08, -2.457585e-08, -2.477124e-08,
  -2.06621e-08, -2.052785e-08, -2.04996e-08, -2.053589e-08, -2.05639e-08, 
    -2.058901e-08, -2.065656e-08, -2.068776e-08, -2.071391e-08, 
    -2.068587e-08, -2.066361e-08, -2.060189e-08, -2.060554e-08, -2.05951e-08, 
    -2.063689e-08,
  -2.081297e-08, -2.080118e-08, -2.087504e-08, -2.094857e-08, -2.10273e-08, 
    -2.1102e-08, -2.113735e-08, -2.117759e-08, -2.118133e-08, -2.117297e-08, 
    -2.111639e-08, -2.101527e-08, -2.089083e-08, -2.073047e-08, -2.061125e-08,
  -2.11112e-08, -2.11957e-08, -2.148679e-08, -2.169286e-08, -2.192853e-08, 
    -2.20328e-08, -2.209415e-08, -2.204979e-08, -2.197546e-08, -2.18698e-08, 
    -2.173895e-08, -2.159211e-08, -2.144681e-08, -2.124768e-08, -2.104654e-08,
  -2.172174e-08, -2.205964e-08, -2.24885e-08, -2.276335e-08, -2.296028e-08, 
    -2.300646e-08, -2.299482e-08, -2.283779e-08, -2.2653e-08, -2.241058e-08, 
    -2.221901e-08, -2.202172e-08, -2.187446e-08, -2.172609e-08, -2.156452e-08,
  -2.249822e-08, -2.285613e-08, -2.316709e-08, -2.332606e-08, -2.340008e-08, 
    -2.336472e-08, -2.321458e-08, -2.304351e-08, -2.278958e-08, 
    -2.252833e-08, -2.231532e-08, -2.210412e-08, -2.203108e-08, 
    -2.198756e-08, -2.189105e-08,
  -2.31551e-08, -2.335238e-08, -2.350867e-08, -2.339249e-08, -2.318401e-08, 
    -2.29505e-08, -2.281868e-08, -2.270488e-08, -2.252035e-08, -2.22788e-08, 
    -2.205911e-08, -2.188446e-08, -2.185034e-08, -2.184406e-08, -2.183843e-08,
  -2.355431e-08, -2.346912e-08, -2.301591e-08, -2.270163e-08, -2.238188e-08, 
    -2.232777e-08, -2.229261e-08, -2.23579e-08, -2.218056e-08, -2.203317e-08, 
    -2.175696e-08, -2.166354e-08, -2.153122e-08, -2.161351e-08, -2.163806e-08,
  -2.336563e-08, -2.283096e-08, -2.240659e-08, -2.216331e-08, -2.207342e-08, 
    -2.21263e-08, -2.223298e-08, -2.228924e-08, -2.215342e-08, -2.191845e-08, 
    -2.165588e-08, -2.154853e-08, -2.1406e-08, -2.151538e-08, -2.156303e-08,
  -2.28582e-08, -2.246644e-08, -2.228087e-08, -2.212366e-08, -2.216987e-08, 
    -2.234225e-08, -2.248492e-08, -2.249212e-08, -2.230156e-08, 
    -2.190398e-08, -2.159819e-08, -2.140139e-08, -2.124573e-08, 
    -2.134642e-08, -2.135836e-08,
  -2.263014e-08, -2.248052e-08, -2.244208e-08, -2.236576e-08, -2.257406e-08, 
    -2.276453e-08, -2.287568e-08, -2.280097e-08, -2.251426e-08, 
    -2.199117e-08, -2.167907e-08, -2.134441e-08, -2.124587e-08, 
    -2.127228e-08, -2.120203e-08,
  -2.078586e-08, -2.078838e-08, -2.08457e-08, -2.08569e-08, -2.096334e-08, 
    -2.130209e-08, -2.143806e-08, -2.162359e-08, -2.181392e-08, 
    -2.205601e-08, -2.223122e-08, -2.237154e-08, -2.241057e-08, 
    -2.232358e-08, -2.226846e-08,
  -2.086356e-08, -2.121689e-08, -2.131419e-08, -2.158564e-08, -2.177781e-08, 
    -2.202427e-08, -2.217609e-08, -2.235572e-08, -2.24277e-08, -2.239362e-08, 
    -2.232467e-08, -2.219998e-08, -2.215838e-08, -2.212949e-08, -2.2182e-08,
  -2.139345e-08, -2.172256e-08, -2.173041e-08, -2.197725e-08, -2.200594e-08, 
    -2.21661e-08, -2.222077e-08, -2.225789e-08, -2.219617e-08, -2.211752e-08, 
    -2.196157e-08, -2.185147e-08, -2.180859e-08, -2.185712e-08, -2.198194e-08,
  -2.176957e-08, -2.164354e-08, -2.177883e-08, -2.18219e-08, -2.178608e-08, 
    -2.179753e-08, -2.172538e-08, -2.171731e-08, -2.163627e-08, -2.16334e-08, 
    -2.15987e-08, -2.163381e-08, -2.163831e-08, -2.168106e-08, -2.174941e-08,
  -2.18594e-08, -2.172471e-08, -2.179952e-08, -2.162843e-08, -2.15489e-08, 
    -2.143108e-08, -2.132266e-08, -2.125087e-08, -2.124102e-08, 
    -2.131776e-08, -2.137772e-08, -2.149326e-08, -2.150368e-08, 
    -2.152367e-08, -2.16516e-08,
  -2.194913e-08, -2.18037e-08, -2.173695e-08, -2.154442e-08, -2.143484e-08, 
    -2.128848e-08, -2.11361e-08, -2.10462e-08, -2.105881e-08, -2.116164e-08, 
    -2.129806e-08, -2.137995e-08, -2.147156e-08, -2.160387e-08, -2.174499e-08,
  -2.209092e-08, -2.180791e-08, -2.167055e-08, -2.149025e-08, -2.136077e-08, 
    -2.118431e-08, -2.101833e-08, -2.090624e-08, -2.09247e-08, -2.100979e-08, 
    -2.115472e-08, -2.128196e-08, -2.154925e-08, -2.171421e-08, -2.192228e-08,
  -2.199387e-08, -2.17286e-08, -2.160219e-08, -2.141342e-08, -2.127053e-08, 
    -2.108237e-08, -2.091796e-08, -2.079543e-08, -2.078747e-08, 
    -2.093434e-08, -2.1066e-08, -2.130018e-08, -2.162045e-08, -2.190262e-08, 
    -2.216873e-08,
  -2.189009e-08, -2.166108e-08, -2.149848e-08, -2.12827e-08, -2.110981e-08, 
    -2.092049e-08, -2.077985e-08, -2.065363e-08, -2.069486e-08, 
    -2.089086e-08, -2.117364e-08, -2.155862e-08, -2.192708e-08, 
    -2.225431e-08, -2.249563e-08,
  -2.172659e-08, -2.151699e-08, -2.132915e-08, -2.109977e-08, -2.094001e-08, 
    -2.076245e-08, -2.067253e-08, -2.057768e-08, -2.0721e-08, -2.104604e-08, 
    -2.141947e-08, -2.182616e-08, -2.218543e-08, -2.246486e-08, -2.277532e-08,
  -2.168895e-08, -2.240803e-08, -2.241899e-08, -2.305448e-08, -2.319148e-08, 
    -2.361831e-08, -2.295458e-08, -2.250488e-08, -2.168798e-08, 
    -2.161749e-08, -2.163026e-08, -2.209173e-08, -2.239849e-08, 
    -2.268548e-08, -2.298098e-08,
  -2.199131e-08, -2.227737e-08, -2.248782e-08, -2.299866e-08, -2.320755e-08, 
    -2.280223e-08, -2.153704e-08, -2.156103e-08, -2.148838e-08, 
    -2.181825e-08, -2.206997e-08, -2.242264e-08, -2.242698e-08, 
    -2.255735e-08, -2.261276e-08,
  -2.241074e-08, -2.240131e-08, -2.257922e-08, -2.274937e-08, -2.279141e-08, 
    -2.185695e-08, -2.187276e-08, -2.22113e-08, -2.215423e-08, -2.235483e-08, 
    -2.226717e-08, -2.229823e-08, -2.22377e-08, -2.240916e-08, -2.258614e-08,
  -2.295169e-08, -2.293928e-08, -2.340021e-08, -2.337909e-08, -2.295931e-08, 
    -2.222865e-08, -2.290271e-08, -2.301103e-08, -2.304659e-08, 
    -2.312359e-08, -2.3012e-08, -2.309315e-08, -2.313234e-08, -2.308113e-08, 
    -2.307652e-08,
  -2.357798e-08, -2.380392e-08, -2.417841e-08, -2.359511e-08, -2.290122e-08, 
    -2.324574e-08, -2.412405e-08, -2.388291e-08, -2.388144e-08, 
    -2.346036e-08, -2.327634e-08, -2.322875e-08, -2.312434e-08, -2.30619e-08, 
    -2.289325e-08,
  -2.387248e-08, -2.40803e-08, -2.405258e-08, -2.339433e-08, -2.340858e-08, 
    -2.43299e-08, -2.42441e-08, -2.385156e-08, -2.352731e-08, -2.325866e-08, 
    -2.322447e-08, -2.310961e-08, -2.29705e-08, -2.29111e-08, -2.287003e-08,
  -2.390907e-08, -2.394343e-08, -2.387462e-08, -2.352411e-08, -2.401486e-08, 
    -2.414602e-08, -2.371131e-08, -2.359561e-08, -2.342623e-08, 
    -2.326803e-08, -2.314779e-08, -2.302467e-08, -2.302282e-08, 
    -2.303047e-08, -2.303791e-08,
  -2.401017e-08, -2.376057e-08, -2.391335e-08, -2.373465e-08, -2.393654e-08, 
    -2.362921e-08, -2.354205e-08, -2.355912e-08, -2.331386e-08, 
    -2.309953e-08, -2.314627e-08, -2.322422e-08, -2.32939e-08, -2.332505e-08, 
    -2.339144e-08,
  -2.391586e-08, -2.37071e-08, -2.386156e-08, -2.360447e-08, -2.361251e-08, 
    -2.344006e-08, -2.352929e-08, -2.329701e-08, -2.313448e-08, 
    -2.326382e-08, -2.3413e-08, -2.355221e-08, -2.371231e-08, -2.384644e-08, 
    -2.382184e-08,
  -2.375709e-08, -2.350903e-08, -2.35788e-08, -2.33816e-08, -2.343947e-08, 
    -2.334616e-08, -2.331336e-08, -2.318195e-08, -2.339839e-08, 
    -2.358734e-08, -2.377678e-08, -2.399935e-08, -2.415298e-08, 
    -2.407005e-08, -2.396924e-08,
  -2.168534e-08, -2.097635e-08, -2.040306e-08, -1.961551e-08, -2.021837e-08, 
    -2.020283e-08, -2.010017e-08, -2.036996e-08, -2.016282e-08, 
    -2.014468e-08, -2.023002e-08, -2.035428e-08, -2.074116e-08, 
    -2.103534e-08, -2.127353e-08,
  -2.164927e-08, -2.098986e-08, -2.050111e-08, -1.954321e-08, -2.004412e-08, 
    -2.087435e-08, -2.077077e-08, -2.071126e-08, -2.039643e-08, 
    -2.063685e-08, -2.048525e-08, -2.060245e-08, -2.074682e-08, -2.09005e-08, 
    -2.117348e-08,
  -2.118167e-08, -2.123656e-08, -2.084829e-08, -2.007212e-08, -1.99627e-08, 
    -2.098277e-08, -2.118796e-08, -2.095281e-08, -2.079719e-08, 
    -2.080898e-08, -2.049907e-08, -2.061319e-08, -2.067632e-08, 
    -2.081427e-08, -2.084271e-08,
  -2.073159e-08, -2.127926e-08, -2.133267e-08, -2.040664e-08, -2.009793e-08, 
    -2.140109e-08, -2.175172e-08, -2.110839e-08, -2.084787e-08, 
    -2.082186e-08, -2.048873e-08, -2.080513e-08, -2.078494e-08, 
    -2.097067e-08, -2.08871e-08,
  -2.075588e-08, -2.143104e-08, -2.200791e-08, -2.098359e-08, -2.059838e-08, 
    -2.20088e-08, -2.192658e-08, -2.111808e-08, -2.101014e-08, -2.083e-08, 
    -2.082845e-08, -2.112252e-08, -2.119752e-08, -2.151557e-08, -2.118237e-08,
  -2.093848e-08, -2.200549e-08, -2.245299e-08, -2.125018e-08, -2.091022e-08, 
    -2.241172e-08, -2.223959e-08, -2.121179e-08, -2.122891e-08, 
    -2.117161e-08, -2.169738e-08, -2.202637e-08, -2.219215e-08, -2.22118e-08, 
    -2.172192e-08,
  -2.186892e-08, -2.224828e-08, -2.243685e-08, -2.148617e-08, -2.15652e-08, 
    -2.303755e-08, -2.232854e-08, -2.134829e-08, -2.173281e-08, 
    -2.177894e-08, -2.230412e-08, -2.217473e-08, -2.221594e-08, 
    -2.207901e-08, -2.155055e-08,
  -2.260256e-08, -2.235152e-08, -2.201873e-08, -2.177563e-08, -2.183965e-08, 
    -2.295916e-08, -2.222388e-08, -2.185825e-08, -2.212656e-08, 
    -2.197434e-08, -2.221444e-08, -2.189936e-08, -2.209227e-08, 
    -2.183511e-08, -2.148307e-08,
  -2.260069e-08, -2.231491e-08, -2.176698e-08, -2.188356e-08, -2.21137e-08, 
    -2.29067e-08, -2.250607e-08, -2.235406e-08, -2.226045e-08, -2.183803e-08, 
    -2.192876e-08, -2.175896e-08, -2.200711e-08, -2.174675e-08, -2.148886e-08,
  -2.259188e-08, -2.225254e-08, -2.161061e-08, -2.200886e-08, -2.226629e-08, 
    -2.299593e-08, -2.279714e-08, -2.262881e-08, -2.222976e-08, 
    -2.180396e-08, -2.176027e-08, -2.175884e-08, -2.198247e-08, 
    -2.172354e-08, -2.145563e-08,
  -2.22475e-08, -2.101856e-08, -2.046981e-08, -1.992552e-08, -1.983965e-08, 
    -1.953909e-08, -1.940037e-08, -1.906514e-08, -1.857035e-08, 
    -1.813978e-08, -1.770683e-08, -1.743584e-08, -1.705257e-08, 
    -1.669795e-08, -1.636607e-08,
  -2.225565e-08, -2.189919e-08, -2.126316e-08, -2.105429e-08, -2.079104e-08, 
    -2.056572e-08, -2.053723e-08, -2.028183e-08, -1.991767e-08, 
    -1.966542e-08, -1.926491e-08, -1.90622e-08, -1.891004e-08, -1.872677e-08, 
    -1.854112e-08,
  -2.341626e-08, -2.294078e-08, -2.231828e-08, -2.19098e-08, -2.195407e-08, 
    -2.196772e-08, -2.176431e-08, -2.180251e-08, -2.132191e-08, -2.09982e-08, 
    -2.06917e-08, -2.040019e-08, -2.036909e-08, -2.034478e-08, -2.034133e-08,
  -2.432633e-08, -2.362899e-08, -2.31548e-08, -2.233898e-08, -2.218359e-08, 
    -2.23694e-08, -2.242269e-08, -2.230561e-08, -2.225944e-08, -2.211322e-08, 
    -2.207474e-08, -2.198505e-08, -2.200768e-08, -2.222465e-08, -2.237572e-08,
  -2.56161e-08, -2.380616e-08, -2.378214e-08, -2.320567e-08, -2.234239e-08, 
    -2.266714e-08, -2.312158e-08, -2.31167e-08, -2.2926e-08, -2.290677e-08, 
    -2.279277e-08, -2.293665e-08, -2.313451e-08, -2.346967e-08, -2.384134e-08,
  -2.641371e-08, -2.469458e-08, -2.410722e-08, -2.408923e-08, -2.274887e-08, 
    -2.238866e-08, -2.312513e-08, -2.355964e-08, -2.354689e-08, 
    -2.361367e-08, -2.354341e-08, -2.377887e-08, -2.401918e-08, 
    -2.439257e-08, -2.474558e-08,
  -2.530859e-08, -2.512357e-08, -2.478499e-08, -2.414669e-08, -2.329242e-08, 
    -2.242251e-08, -2.286931e-08, -2.337459e-08, -2.345215e-08, 
    -2.373319e-08, -2.372752e-08, -2.39851e-08, -2.428816e-08, -2.446414e-08, 
    -2.473757e-08,
  -2.540139e-08, -2.504319e-08, -2.535841e-08, -2.44028e-08, -2.346559e-08, 
    -2.265333e-08, -2.282848e-08, -2.307435e-08, -2.3258e-08, -2.365427e-08, 
    -2.366716e-08, -2.407351e-08, -2.411294e-08, -2.423359e-08, -2.436055e-08,
  -2.488081e-08, -2.486376e-08, -2.55332e-08, -2.456622e-08, -2.356241e-08, 
    -2.264991e-08, -2.296446e-08, -2.30074e-08, -2.307392e-08, -2.332143e-08, 
    -2.350434e-08, -2.387453e-08, -2.380036e-08, -2.386679e-08, -2.379385e-08,
  -2.395543e-08, -2.425109e-08, -2.539672e-08, -2.440876e-08, -2.335398e-08, 
    -2.274279e-08, -2.317724e-08, -2.302614e-08, -2.292159e-08, 
    -2.301312e-08, -2.331729e-08, -2.35977e-08, -2.346243e-08, -2.35014e-08, 
    -2.338907e-08,
  -6.166879e-09, -4.905987e-09, -4.199285e-09, -3.530302e-09, -3.006124e-09, 
    -2.563273e-09, -2.427906e-09, -2.363268e-09, -2.288415e-09, -2.39702e-09, 
    -2.896216e-09, -3.703554e-09, -4.439633e-09, -5.209385e-09, -6.22053e-09,
  -7.373889e-09, -6.312534e-09, -5.460159e-09, -4.715541e-09, -4.115026e-09, 
    -3.547474e-09, -3.191139e-09, -2.966064e-09, -2.840752e-09, 
    -2.955821e-09, -3.460254e-09, -4.349336e-09, -5.14293e-09, -5.941252e-09, 
    -6.977015e-09,
  -8.733365e-09, -7.715133e-09, -6.882011e-09, -5.973512e-09, -5.245315e-09, 
    -4.869356e-09, -4.459435e-09, -4.185359e-09, -3.980614e-09, 
    -4.048979e-09, -4.432003e-09, -5.317777e-09, -5.995341e-09, -6.73305e-09, 
    -7.733313e-09,
  -9.916119e-09, -9.064101e-09, -8.363411e-09, -7.541201e-09, -6.750623e-09, 
    -6.068904e-09, -5.778097e-09, -5.551171e-09, -5.467248e-09, 
    -5.470691e-09, -5.768766e-09, -6.471888e-09, -7.032977e-09, 
    -7.718139e-09, -8.679685e-09,
  -1.158718e-08, -1.069506e-08, -1.006339e-08, -9.444431e-09, -8.853939e-09, 
    -8.20084e-09, -7.588588e-09, -7.251193e-09, -7.169149e-09, -7.123705e-09, 
    -7.247554e-09, -7.707009e-09, -8.124306e-09, -8.781504e-09, -9.660527e-09,
  -1.328685e-08, -1.22962e-08, -1.158851e-08, -1.09186e-08, -1.042741e-08, 
    -1.002399e-08, -9.510013e-09, -9.051887e-09, -8.835185e-09, -8.64886e-09, 
    -8.582012e-09, -8.960335e-09, -9.417429e-09, -1.00516e-08, -1.076164e-08,
  -1.473707e-08, -1.385986e-08, -1.328188e-08, -1.252221e-08, -1.18958e-08, 
    -1.146488e-08, -1.106621e-08, -1.062881e-08, -1.038037e-08, 
    -1.018719e-08, -1.007146e-08, -1.037983e-08, -1.081375e-08, 
    -1.147517e-08, -1.209713e-08,
  -1.641162e-08, -1.554583e-08, -1.485535e-08, -1.41592e-08, -1.354324e-08, 
    -1.311861e-08, -1.280584e-08, -1.244456e-08, -1.217199e-08, 
    -1.190084e-08, -1.171588e-08, -1.186388e-08, -1.229496e-08, 
    -1.290841e-08, -1.345575e-08,
  -1.783401e-08, -1.685917e-08, -1.654843e-08, -1.573519e-08, -1.525608e-08, 
    -1.464215e-08, -1.428362e-08, -1.408044e-08, -1.395199e-08, 
    -1.361245e-08, -1.333151e-08, -1.335592e-08, -1.380567e-08, 
    -1.432823e-08, -1.481702e-08,
  -2.03657e-08, -1.856883e-08, -1.797201e-08, -1.756023e-08, -1.673948e-08, 
    -1.634991e-08, -1.587623e-08, -1.553057e-08, -1.539039e-08, 
    -1.504107e-08, -1.47268e-08, -1.473383e-08, -1.520981e-08, -1.560921e-08, 
    -1.61092e-08,
  -1.692056e-09, -1.783279e-09, -1.712288e-09, -1.575836e-09, -1.646916e-09, 
    -2.074115e-09, -2.727401e-09, -3.4755e-09, -4.366946e-09, -5.593288e-09, 
    -7.199228e-09, -9.175976e-09, -1.1213e-08, -1.354824e-08, -1.635295e-08,
  -1.824737e-09, -1.884608e-09, -1.942376e-09, -1.82266e-09, -1.835097e-09, 
    -2.275005e-09, -3.011027e-09, -3.783405e-09, -4.667661e-09, 
    -5.875894e-09, -7.435354e-09, -9.355295e-09, -1.141929e-08, 
    -1.385453e-08, -1.673987e-08,
  -2.088911e-09, -2.126236e-09, -2.21282e-09, -2.032114e-09, -2.121799e-09, 
    -2.608176e-09, -3.317423e-09, -4.048231e-09, -4.957482e-09, 
    -6.146768e-09, -7.655598e-09, -9.511257e-09, -1.15478e-08, -1.408661e-08, 
    -1.700832e-08,
  -2.157491e-09, -2.283235e-09, -2.30672e-09, -2.068495e-09, -2.191761e-09, 
    -2.758412e-09, -3.502608e-09, -4.253435e-09, -5.202537e-09, 
    -6.420911e-09, -7.941479e-09, -9.760071e-09, -1.180113e-08, 
    -1.440585e-08, -1.731163e-08,
  -2.254499e-09, -2.362363e-09, -2.25957e-09, -1.9699e-09, -2.128122e-09, 
    -2.842858e-09, -3.572822e-09, -4.412759e-09, -5.432055e-09, 
    -6.707642e-09, -8.246977e-09, -1.005847e-08, -1.209575e-08, 
    -1.475935e-08, -1.757313e-08,
  -2.334057e-09, -2.382601e-09, -2.159884e-09, -1.851026e-09, -2.120452e-09, 
    -2.969142e-09, -3.70439e-09, -4.627359e-09, -5.680497e-09, -7.000303e-09, 
    -8.55774e-09, -1.036428e-08, -1.24235e-08, -1.512016e-08, -1.783774e-08,
  -2.228354e-09, -2.399405e-09, -2.125522e-09, -1.858147e-09, -2.348431e-09, 
    -3.250479e-09, -3.955392e-09, -4.949973e-09, -5.990296e-09, 
    -7.311069e-09, -8.880524e-09, -1.069983e-08, -1.279451e-08, 
    -1.549372e-08, -1.807804e-08,
  -2.272232e-09, -2.561587e-09, -2.162819e-09, -2.052167e-09, -2.750995e-09, 
    -3.618698e-09, -4.313971e-09, -5.313762e-09, -6.341834e-09, 
    -7.675468e-09, -9.222403e-09, -1.106755e-08, -1.321081e-08, 
    -1.586802e-08, -1.833473e-08,
  -2.459918e-09, -2.66381e-09, -2.292855e-09, -2.452888e-09, -3.204259e-09, 
    -3.985605e-09, -4.729497e-09, -5.715772e-09, -6.722684e-09, 
    -8.065438e-09, -9.623349e-09, -1.148475e-08, -1.367349e-08, 
    -1.624285e-08, -1.858564e-08,
  -2.795646e-09, -2.823905e-09, -2.648408e-09, -2.962544e-09, -3.603491e-09, 
    -4.353296e-09, -5.176346e-09, -6.109324e-09, -7.123559e-09, 
    -8.469713e-09, -1.001604e-08, -1.190897e-08, -1.413966e-08, 
    -1.657527e-08, -1.885424e-08,
  -3.36065e-09, -4.270468e-09, -5.136724e-09, -6.136457e-09, -7.220853e-09, 
    -8.19371e-09, -9.341621e-09, -1.077633e-08, -1.239372e-08, -1.500803e-08, 
    -1.880802e-08, -2.254818e-08, -2.496761e-08, -2.581046e-08, -2.580703e-08,
  -3.36985e-09, -4.26286e-09, -5.087253e-09, -6.011618e-09, -6.984478e-09, 
    -8.001118e-09, -9.244848e-09, -1.077056e-08, -1.245449e-08, 
    -1.521627e-08, -1.918338e-08, -2.294935e-08, -2.519833e-08, 
    -2.601733e-08, -2.553721e-08,
  -3.374489e-09, -4.25376e-09, -5.079578e-09, -5.879417e-09, -6.783197e-09, 
    -7.808984e-09, -9.118683e-09, -1.073845e-08, -1.249188e-08, 
    -1.540741e-08, -1.952966e-08, -2.333428e-08, -2.546744e-08, 
    -2.597094e-08, -2.514818e-08,
  -3.307227e-09, -4.155837e-09, -5.029619e-09, -5.841682e-09, -6.633952e-09, 
    -7.67896e-09, -9.059057e-09, -1.070176e-08, -1.24821e-08, -1.55657e-08, 
    -1.983414e-08, -2.364389e-08, -2.561043e-08, -2.583071e-08, -2.455676e-08,
  -3.219426e-09, -4.073009e-09, -5.005076e-09, -5.850592e-09, -6.623079e-09, 
    -7.619429e-09, -8.988443e-09, -1.06745e-08, -1.25283e-08, -1.578401e-08, 
    -2.014028e-08, -2.393277e-08, -2.560988e-08, -2.530798e-08, -2.395681e-08,
  -3.176045e-09, -4.052657e-09, -5.022241e-09, -5.843653e-09, -6.652106e-09, 
    -7.629339e-09, -8.957583e-09, -1.063735e-08, -1.256744e-08, 
    -1.602566e-08, -2.047024e-08, -2.415136e-08, -2.537528e-08, 
    -2.469361e-08, -2.358141e-08,
  -3.167605e-09, -4.054035e-09, -5.041732e-09, -5.803477e-09, -6.675617e-09, 
    -7.684719e-09, -8.96382e-09, -1.059716e-08, -1.263988e-08, -1.630537e-08, 
    -2.078625e-08, -2.429732e-08, -2.493975e-08, -2.401372e-08, -2.338449e-08,
  -3.171232e-09, -4.073931e-09, -5.057701e-09, -5.757135e-09, -6.678055e-09, 
    -7.742996e-09, -9.007236e-09, -1.060524e-08, -1.277405e-08, -1.66292e-08, 
    -2.112394e-08, -2.426923e-08, -2.437358e-08, -2.350646e-08, -2.351929e-08,
  -3.167321e-09, -4.122084e-09, -5.069551e-09, -5.686386e-09, -6.665865e-09, 
    -7.798101e-09, -9.063513e-09, -1.066149e-08, -1.299005e-08, 
    -1.699758e-08, -2.145875e-08, -2.40238e-08, -2.367211e-08, -2.325339e-08, 
    -2.37538e-08,
  -3.150716e-09, -4.173991e-09, -5.072195e-09, -5.624202e-09, -6.639822e-09, 
    -7.844874e-09, -9.137499e-09, -1.07883e-08, -1.328257e-08, -1.738626e-08, 
    -2.163642e-08, -2.357296e-08, -2.312605e-08, -2.320642e-08, -2.411751e-08,
  -1.057436e-08, -1.213625e-08, -1.361176e-08, -1.516334e-08, -1.635405e-08, 
    -1.726733e-08, -1.79441e-08, -1.841011e-08, -1.858822e-08, -1.875128e-08, 
    -1.889535e-08, -1.901476e-08, -1.927046e-08, -1.979484e-08, -2.041795e-08,
  -1.057192e-08, -1.208215e-08, -1.352309e-08, -1.505784e-08, -1.624484e-08, 
    -1.712766e-08, -1.778578e-08, -1.821102e-08, -1.837115e-08, 
    -1.848906e-08, -1.86275e-08, -1.870918e-08, -1.902594e-08, -1.953501e-08, 
    -2.009e-08,
  -1.043677e-08, -1.197756e-08, -1.342267e-08, -1.498964e-08, -1.621474e-08, 
    -1.709898e-08, -1.776374e-08, -1.807993e-08, -1.822043e-08, 
    -1.838545e-08, -1.849709e-08, -1.849797e-08, -1.881828e-08, 
    -1.936224e-08, -1.988668e-08,
  -1.032375e-08, -1.189879e-08, -1.334528e-08, -1.49495e-08, -1.616374e-08, 
    -1.704405e-08, -1.770464e-08, -1.802752e-08, -1.814335e-08, 
    -1.831413e-08, -1.842308e-08, -1.837658e-08, -1.866195e-08, 
    -1.925052e-08, -1.986552e-08,
  -1.021295e-08, -1.178725e-08, -1.322685e-08, -1.486767e-08, -1.614606e-08, 
    -1.705051e-08, -1.76771e-08, -1.794116e-08, -1.812949e-08, -1.837626e-08, 
    -1.844022e-08, -1.837962e-08, -1.86154e-08, -1.91987e-08, -1.986179e-08,
  -1.00745e-08, -1.163065e-08, -1.306303e-08, -1.475393e-08, -1.608287e-08, 
    -1.700585e-08, -1.763377e-08, -1.791149e-08, -1.81106e-08, -1.849896e-08, 
    -1.858102e-08, -1.846217e-08, -1.865766e-08, -1.913125e-08, -1.978919e-08,
  -9.930664e-09, -1.146673e-08, -1.290808e-08, -1.463344e-08, -1.599402e-08, 
    -1.690818e-08, -1.750695e-08, -1.787402e-08, -1.818785e-08, -1.86815e-08, 
    -1.877606e-08, -1.864537e-08, -1.871691e-08, -1.910172e-08, -1.970574e-08,
  -9.779996e-09, -1.131782e-08, -1.276961e-08, -1.45148e-08, -1.586111e-08, 
    -1.678234e-08, -1.736771e-08, -1.779105e-08, -1.824457e-08, 
    -1.893287e-08, -1.903465e-08, -1.882434e-08, -1.884276e-08, 
    -1.907869e-08, -1.962109e-08,
  -9.653786e-09, -1.118909e-08, -1.266903e-08, -1.443472e-08, -1.570663e-08, 
    -1.661543e-08, -1.721569e-08, -1.773165e-08, -1.831267e-08, 
    -1.917647e-08, -1.929066e-08, -1.907947e-08, -1.90532e-08, -1.908962e-08, 
    -1.957136e-08,
  -9.555818e-09, -1.109067e-08, -1.262585e-08, -1.437651e-08, -1.556582e-08, 
    -1.647156e-08, -1.706969e-08, -1.768543e-08, -1.843266e-08, 
    -1.941224e-08, -1.950546e-08, -1.924878e-08, -1.927829e-08, 
    -1.919902e-08, -1.952547e-08,
  -1.427132e-08, -1.679635e-08, -1.846119e-08, -1.99591e-08, -2.117042e-08, 
    -2.229194e-08, -2.308522e-08, -2.382986e-08, -2.44553e-08, -2.495837e-08, 
    -2.530689e-08, -2.548716e-08, -2.569125e-08, -2.565186e-08, -2.565617e-08,
  -1.422983e-08, -1.67399e-08, -1.836819e-08, -1.983702e-08, -2.101225e-08, 
    -2.219809e-08, -2.308392e-08, -2.381042e-08, -2.440063e-08, 
    -2.486513e-08, -2.522151e-08, -2.554256e-08, -2.575587e-08, 
    -2.580824e-08, -2.594328e-08,
  -1.422364e-08, -1.670427e-08, -1.830951e-08, -1.983944e-08, -2.100507e-08, 
    -2.219237e-08, -2.311453e-08, -2.386028e-08, -2.429761e-08, 
    -2.476466e-08, -2.521272e-08, -2.569218e-08, -2.604648e-08, 
    -2.612655e-08, -2.625202e-08,
  -1.425398e-08, -1.675008e-08, -1.843753e-08, -2.005574e-08, -2.117927e-08, 
    -2.229541e-08, -2.324292e-08, -2.388377e-08, -2.426794e-08, -2.47966e-08, 
    -2.537248e-08, -2.596485e-08, -2.628611e-08, -2.633275e-08, -2.628068e-08,
  -1.426938e-08, -1.675494e-08, -1.848619e-08, -2.019011e-08, -2.134861e-08, 
    -2.242864e-08, -2.33272e-08, -2.389202e-08, -2.423578e-08, -2.482732e-08, 
    -2.546538e-08, -2.60586e-08, -2.638028e-08, -2.641595e-08, -2.635895e-08,
  -1.429672e-08, -1.677886e-08, -1.850819e-08, -2.027807e-08, -2.143093e-08, 
    -2.250397e-08, -2.335354e-08, -2.387755e-08, -2.429994e-08, 
    -2.494367e-08, -2.563231e-08, -2.627265e-08, -2.652053e-08, 
    -2.652147e-08, -2.649129e-08,
  -1.43155e-08, -1.682205e-08, -1.85616e-08, -2.031728e-08, -2.148144e-08, 
    -2.25727e-08, -2.343557e-08, -2.387982e-08, -2.437321e-08, -2.511594e-08, 
    -2.581428e-08, -2.638703e-08, -2.664943e-08, -2.664403e-08, -2.666504e-08,
  -1.434709e-08, -1.686127e-08, -1.862669e-08, -2.037367e-08, -2.150006e-08, 
    -2.263349e-08, -2.34291e-08, -2.397413e-08, -2.450616e-08, -2.527324e-08, 
    -2.595369e-08, -2.652883e-08, -2.674312e-08, -2.687045e-08, -2.686625e-08,
  -1.437446e-08, -1.685847e-08, -1.866433e-08, -2.03982e-08, -2.15406e-08, 
    -2.263526e-08, -2.341381e-08, -2.394196e-08, -2.454596e-08, 
    -2.538528e-08, -2.602178e-08, -2.661021e-08, -2.683121e-08, 
    -2.700875e-08, -2.706282e-08,
  -1.440728e-08, -1.681806e-08, -1.864485e-08, -2.040577e-08, -2.154463e-08, 
    -2.259772e-08, -2.332327e-08, -2.387265e-08, -2.455202e-08, 
    -2.532704e-08, -2.607444e-08, -2.666111e-08, -2.682133e-08, 
    -2.710115e-08, -2.729007e-08,
  -2.385426e-08, -2.42691e-08, -2.411288e-08, -2.386173e-08, -2.358714e-08, 
    -2.356226e-08, -2.363906e-08, -2.368967e-08, -2.374644e-08, 
    -2.377754e-08, -2.388054e-08, -2.389526e-08, -2.392365e-08, -2.38715e-08, 
    -2.382862e-08,
  -2.37564e-08, -2.424858e-08, -2.395989e-08, -2.369348e-08, -2.355695e-08, 
    -2.364228e-08, -2.379616e-08, -2.40498e-08, -2.438051e-08, -2.457953e-08, 
    -2.4723e-08, -2.482762e-08, -2.481831e-08, -2.473687e-08, -2.46205e-08,
  -2.379175e-08, -2.431232e-08, -2.403187e-08, -2.398104e-08, -2.390611e-08, 
    -2.413845e-08, -2.434569e-08, -2.461674e-08, -2.492913e-08, 
    -2.501237e-08, -2.527947e-08, -2.543734e-08, -2.543874e-08, 
    -2.539505e-08, -2.526182e-08,
  -2.376579e-08, -2.437127e-08, -2.421249e-08, -2.420378e-08, -2.414114e-08, 
    -2.416908e-08, -2.402977e-08, -2.411279e-08, -2.415788e-08, 
    -2.417663e-08, -2.441053e-08, -2.45368e-08, -2.468702e-08, -2.481904e-08, 
    -2.49561e-08,
  -2.370344e-08, -2.446678e-08, -2.447355e-08, -2.447523e-08, -2.414183e-08, 
    -2.37958e-08, -2.363835e-08, -2.361099e-08, -2.358628e-08, -2.367268e-08, 
    -2.374784e-08, -2.386514e-08, -2.401969e-08, -2.409253e-08, -2.422757e-08,
  -2.360562e-08, -2.454557e-08, -2.464369e-08, -2.446716e-08, -2.390068e-08, 
    -2.353271e-08, -2.339462e-08, -2.342053e-08, -2.350292e-08, 
    -2.351152e-08, -2.365983e-08, -2.382773e-08, -2.391418e-08, 
    -2.393151e-08, -2.397035e-08,
  -2.350153e-08, -2.458014e-08, -2.478122e-08, -2.44741e-08, -2.381455e-08, 
    -2.339616e-08, -2.337616e-08, -2.347204e-08, -2.361523e-08, 
    -2.369532e-08, -2.399062e-08, -2.413851e-08, -2.417947e-08, 
    -2.425157e-08, -2.42208e-08,
  -2.337915e-08, -2.452957e-08, -2.478662e-08, -2.441775e-08, -2.38239e-08, 
    -2.342973e-08, -2.351167e-08, -2.362794e-08, -2.389161e-08, 
    -2.407866e-08, -2.434314e-08, -2.449222e-08, -2.454095e-08, -2.45382e-08, 
    -2.452304e-08,
  -2.326641e-08, -2.446118e-08, -2.480449e-08, -2.451811e-08, -2.390763e-08, 
    -2.358678e-08, -2.361221e-08, -2.381549e-08, -2.409818e-08, 
    -2.429465e-08, -2.458134e-08, -2.471895e-08, -2.476345e-08, 
    -2.484028e-08, -2.488601e-08,
  -2.312957e-08, -2.435668e-08, -2.47734e-08, -2.456648e-08, -2.40388e-08, 
    -2.375349e-08, -2.369901e-08, -2.389559e-08, -2.417138e-08, 
    -2.444106e-08, -2.475026e-08, -2.490566e-08, -2.503643e-08, 
    -2.499234e-08, -2.51022e-08,
  -2.277492e-08, -2.324458e-08, -2.34799e-08, -2.347891e-08, -2.356997e-08, 
    -2.317573e-08, -2.304685e-08, -2.257675e-08, -2.228664e-08, 
    -2.194945e-08, -2.175365e-08, -2.158346e-08, -2.138355e-08, 
    -2.112244e-08, -2.082075e-08,
  -2.268339e-08, -2.303599e-08, -2.342805e-08, -2.344314e-08, -2.365422e-08, 
    -2.34287e-08, -2.331763e-08, -2.288198e-08, -2.256496e-08, -2.222781e-08, 
    -2.19927e-08, -2.17282e-08, -2.16046e-08, -2.143934e-08, -2.123754e-08,
  -2.293116e-08, -2.35494e-08, -2.403133e-08, -2.408617e-08, -2.424703e-08, 
    -2.408133e-08, -2.388659e-08, -2.345863e-08, -2.292054e-08, 
    -2.244663e-08, -2.204715e-08, -2.173077e-08, -2.139434e-08, 
    -2.126614e-08, -2.122048e-08,
  -2.324532e-08, -2.41185e-08, -2.484421e-08, -2.49508e-08, -2.488056e-08, 
    -2.467696e-08, -2.443498e-08, -2.416313e-08, -2.373655e-08, 
    -2.319529e-08, -2.268862e-08, -2.232855e-08, -2.194782e-08, 
    -2.157934e-08, -2.140571e-08,
  -2.344412e-08, -2.418024e-08, -2.47245e-08, -2.46515e-08, -2.445916e-08, 
    -2.437594e-08, -2.423952e-08, -2.403545e-08, -2.383377e-08, 
    -2.346327e-08, -2.301792e-08, -2.263651e-08, -2.238513e-08, -2.20738e-08, 
    -2.181736e-08,
  -2.341081e-08, -2.389537e-08, -2.401761e-08, -2.38476e-08, -2.382589e-08, 
    -2.398188e-08, -2.41105e-08, -2.415995e-08, -2.394251e-08, -2.368253e-08, 
    -2.329534e-08, -2.284466e-08, -2.259806e-08, -2.236597e-08, -2.216733e-08,
  -2.341115e-08, -2.364881e-08, -2.349745e-08, -2.330348e-08, -2.343415e-08, 
    -2.372019e-08, -2.394173e-08, -2.419694e-08, -2.417792e-08, 
    -2.395585e-08, -2.372808e-08, -2.327213e-08, -2.285543e-08, 
    -2.264214e-08, -2.246387e-08,
  -2.339106e-08, -2.340162e-08, -2.305524e-08, -2.292907e-08, -2.314497e-08, 
    -2.351392e-08, -2.374733e-08, -2.400063e-08, -2.421939e-08, -2.40108e-08, 
    -2.382583e-08, -2.355664e-08, -2.311223e-08, -2.277035e-08, -2.258952e-08,
  -2.326999e-08, -2.314083e-08, -2.282412e-08, -2.28015e-08, -2.324321e-08, 
    -2.371857e-08, -2.40325e-08, -2.412803e-08, -2.421147e-08, -2.428897e-08, 
    -2.398803e-08, -2.370956e-08, -2.332506e-08, -2.289232e-08, -2.258429e-08,
  -2.31365e-08, -2.29695e-08, -2.279782e-08, -2.299999e-08, -2.357694e-08, 
    -2.407353e-08, -2.444133e-08, -2.446676e-08, -2.45351e-08, -2.458045e-08, 
    -2.453235e-08, -2.40929e-08, -2.374982e-08, -2.328462e-08, -2.288017e-08,
  -1.790244e-08, -1.789387e-08, -1.765121e-08, -1.76497e-08, -1.759458e-08, 
    -1.763636e-08, -1.765304e-08, -1.775962e-08, -1.789675e-08, 
    -1.799486e-08, -1.808915e-08, -1.823908e-08, -1.852803e-08, 
    -1.880698e-08, -1.903786e-08,
  -1.845645e-08, -1.842752e-08, -1.816177e-08, -1.813026e-08, -1.803386e-08, 
    -1.795188e-08, -1.787419e-08, -1.797295e-08, -1.810239e-08, 
    -1.819831e-08, -1.825532e-08, -1.84532e-08, -1.859808e-08, -1.890498e-08, 
    -1.916286e-08,
  -1.903819e-08, -1.901901e-08, -1.885127e-08, -1.88103e-08, -1.852556e-08, 
    -1.837409e-08, -1.827966e-08, -1.831473e-08, -1.840104e-08, -1.84733e-08, 
    -1.855833e-08, -1.858041e-08, -1.877694e-08, -1.906525e-08, -1.92667e-08,
  -1.98176e-08, -1.991106e-08, -1.954868e-08, -1.949946e-08, -1.920653e-08, 
    -1.905883e-08, -1.884468e-08, -1.876932e-08, -1.871671e-08, -1.87474e-08, 
    -1.870124e-08, -1.863516e-08, -1.871058e-08, -1.900636e-08, -1.939578e-08,
  -2.067543e-08, -2.066044e-08, -2.03396e-08, -2.01547e-08, -1.984789e-08, 
    -1.967121e-08, -1.940598e-08, -1.923882e-08, -1.900035e-08, 
    -1.886155e-08, -1.879627e-08, -1.87379e-08, -1.87157e-08, -1.89953e-08, 
    -1.941682e-08,
  -2.138063e-08, -2.122375e-08, -2.110373e-08, -2.069226e-08, -2.037435e-08, 
    -2.009858e-08, -1.974672e-08, -1.948315e-08, -1.928502e-08, 
    -1.904422e-08, -1.89228e-08, -1.891638e-08, -1.896442e-08, -1.915877e-08, 
    -1.960853e-08,
  -2.179687e-08, -2.172402e-08, -2.16276e-08, -2.115121e-08, -2.077217e-08, 
    -2.043642e-08, -2.015171e-08, -1.972637e-08, -1.944704e-08, 
    -1.933308e-08, -1.917863e-08, -1.923836e-08, -1.93221e-08, -1.951198e-08, 
    -1.98738e-08,
  -2.237712e-08, -2.219929e-08, -2.215957e-08, -2.171336e-08, -2.130467e-08, 
    -2.090608e-08, -2.05062e-08, -2.010809e-08, -1.960635e-08, -1.946399e-08, 
    -1.941397e-08, -1.95038e-08, -1.974393e-08, -2.011414e-08, -2.040513e-08,
  -2.302371e-08, -2.258126e-08, -2.261069e-08, -2.217099e-08, -2.178077e-08, 
    -2.142465e-08, -2.097182e-08, -2.055854e-08, -2.00141e-08, -1.962868e-08, 
    -1.969349e-08, -1.987029e-08, -2.001817e-08, -2.043839e-08, -2.071898e-08,
  -2.337909e-08, -2.285879e-08, -2.283538e-08, -2.250867e-08, -2.217693e-08, 
    -2.188276e-08, -2.150142e-08, -2.116501e-08, -2.075415e-08, 
    -2.027385e-08, -2.002652e-08, -2.016318e-08, -2.036841e-08, 
    -2.072994e-08, -2.102482e-08,
  -2.122117e-08, -2.218508e-08, -2.26934e-08, -2.294434e-08, -2.295136e-08, 
    -2.287279e-08, -2.276585e-08, -2.258612e-08, -2.234224e-08, -2.21275e-08, 
    -2.195409e-08, -2.187041e-08, -2.184981e-08, -2.207644e-08, -2.237386e-08,
  -2.054586e-08, -2.159499e-08, -2.262365e-08, -2.312811e-08, -2.340526e-08, 
    -2.359916e-08, -2.374596e-08, -2.379851e-08, -2.372467e-08, 
    -2.376546e-08, -2.389032e-08, -2.409354e-08, -2.443101e-08, -2.50111e-08, 
    -2.577941e-08,
  -1.966671e-08, -2.058561e-08, -2.176814e-08, -2.265464e-08, -2.32298e-08, 
    -2.352771e-08, -2.396757e-08, -2.439936e-08, -2.480281e-08, 
    -2.527793e-08, -2.603918e-08, -2.688225e-08, -2.779075e-08, 
    -2.852821e-08, -2.918965e-08,
  -1.942146e-08, -1.989265e-08, -2.084447e-08, -2.211377e-08, -2.302479e-08, 
    -2.386117e-08, -2.4561e-08, -2.523074e-08, -2.606096e-08, -2.712078e-08, 
    -2.81272e-08, -2.885154e-08, -2.888513e-08, -2.860381e-08, -2.844848e-08,
  -1.939276e-08, -1.950056e-08, -1.975166e-08, -2.044231e-08, -2.16196e-08, 
    -2.278964e-08, -2.368616e-08, -2.452005e-08, -2.519059e-08, 
    -2.568611e-08, -2.605723e-08, -2.638567e-08, -2.691207e-08, 
    -2.742506e-08, -2.795569e-08,
  -1.92841e-08, -1.941683e-08, -1.946756e-08, -1.965941e-08, -2.024916e-08, 
    -2.093827e-08, -2.150936e-08, -2.189046e-08, -2.239193e-08, 
    -2.304867e-08, -2.375571e-08, -2.43256e-08, -2.488583e-08, -2.536468e-08, 
    -2.590591e-08,
  -1.917904e-08, -1.935155e-08, -1.943625e-08, -1.963561e-08, -2.01057e-08, 
    -2.061805e-08, -2.11191e-08, -2.155859e-08, -2.219301e-08, -2.2804e-08, 
    -2.345343e-08, -2.402781e-08, -2.45809e-08, -2.505764e-08, -2.551294e-08,
  -1.906799e-08, -1.926759e-08, -1.95197e-08, -1.979529e-08, -2.012734e-08, 
    -2.054352e-08, -2.099514e-08, -2.150216e-08, -2.216168e-08, 
    -2.282267e-08, -2.339183e-08, -2.386463e-08, -2.44132e-08, -2.494578e-08, 
    -2.538988e-08,
  -1.890492e-08, -1.921231e-08, -1.960454e-08, -1.986494e-08, -2.013699e-08, 
    -2.044233e-08, -2.093426e-08, -2.147863e-08, -2.216965e-08, 
    -2.282965e-08, -2.340102e-08, -2.391151e-08, -2.451267e-08, 
    -2.506559e-08, -2.547255e-08,
  -1.88255e-08, -1.916995e-08, -1.962328e-08, -1.9892e-08, -2.022283e-08, 
    -2.048134e-08, -2.084773e-08, -2.139867e-08, -2.207303e-08, 
    -2.269937e-08, -2.336559e-08, -2.404701e-08, -2.46334e-08, -2.505574e-08, 
    -2.528456e-08,
  -2.253514e-08, -2.125396e-08, -2.028204e-08, -1.930652e-08, -1.872559e-08, 
    -1.826112e-08, -1.776646e-08, -1.729973e-08, -1.709839e-08, 
    -1.685858e-08, -1.65738e-08, -1.588232e-08, -1.497903e-08, -1.407471e-08, 
    -1.331007e-08,
  -2.469499e-08, -2.373963e-08, -2.274373e-08, -2.174112e-08, -2.101262e-08, 
    -2.05972e-08, -2.005815e-08, -1.931695e-08, -1.87977e-08, -1.860464e-08, 
    -1.85695e-08, -1.829408e-08, -1.766693e-08, -1.65763e-08, -1.532263e-08,
  -2.658471e-08, -2.582015e-08, -2.483747e-08, -2.420267e-08, -2.394475e-08, 
    -2.367806e-08, -2.286425e-08, -2.176382e-08, -2.087632e-08, 
    -2.027895e-08, -2.000603e-08, -1.977384e-08, -1.970834e-08, -1.91114e-08, 
    -1.796528e-08,
  -2.863998e-08, -2.900518e-08, -2.853852e-08, -2.720741e-08, -2.631369e-08, 
    -2.568133e-08, -2.528173e-08, -2.475079e-08, -2.39569e-08, -2.297477e-08, 
    -2.201044e-08, -2.122399e-08, -2.07841e-08, -2.066606e-08, -2.029791e-08,
  -2.972937e-08, -3.10725e-08, -3.161276e-08, -3.173054e-08, -3.104043e-08, 
    -2.947286e-08, -2.822641e-08, -2.745507e-08, -2.702747e-08, 
    -2.644349e-08, -2.585575e-08, -2.491645e-08, -2.372083e-08, 
    -2.275072e-08, -2.209983e-08,
  -2.897244e-08, -3.064118e-08, -3.122152e-08, -3.130365e-08, -3.132221e-08, 
    -3.091931e-08, -3.030012e-08, -2.978026e-08, -2.903253e-08, 
    -2.833319e-08, -2.75405e-08, -2.701474e-08, -2.644787e-08, -2.552321e-08, 
    -2.443104e-08,
  -2.768509e-08, -2.901831e-08, -2.989371e-08, -3.030619e-08, -3.039581e-08, 
    -3.014975e-08, -3.010259e-08, -2.993205e-08, -2.956159e-08, 
    -2.876613e-08, -2.802206e-08, -2.75493e-08, -2.71494e-08, -2.667077e-08, 
    -2.558637e-08,
  -2.661692e-08, -2.805838e-08, -2.93129e-08, -2.996151e-08, -3.040291e-08, 
    -3.041156e-08, -3.013829e-08, -2.980728e-08, -2.937224e-08, 
    -2.878003e-08, -2.802248e-08, -2.726151e-08, -2.665517e-08, -2.63232e-08, 
    -2.594238e-08,
  -2.584753e-08, -2.674622e-08, -2.786875e-08, -2.897438e-08, -2.985946e-08, 
    -3.029934e-08, -3.031811e-08, -2.996339e-08, -2.97123e-08, -2.927672e-08, 
    -2.892378e-08, -2.843887e-08, -2.764703e-08, -2.67464e-08, -2.602936e-08,
  -2.534797e-08, -2.584422e-08, -2.660096e-08, -2.737592e-08, -2.865893e-08, 
    -2.948894e-08, -3.023556e-08, -3.053486e-08, -3.022741e-08, 
    -2.982696e-08, -2.955728e-08, -2.894399e-08, -2.836236e-08, 
    -2.784977e-08, -2.714803e-08,
  -7.147642e-09, -6.995977e-09, -6.586874e-09, -6.191249e-09, -6.093882e-09, 
    -6.163083e-09, -6.200481e-09, -5.970055e-09, -5.583859e-09, 
    -5.211545e-09, -5.026106e-09, -4.926138e-09, -4.885574e-09, 
    -4.838822e-09, -4.799847e-09,
  -7.782659e-09, -7.690248e-09, -7.174417e-09, -6.434567e-09, -6.016486e-09, 
    -5.830799e-09, -5.892254e-09, -5.93262e-09, -5.800332e-09, -5.573356e-09, 
    -5.472678e-09, -5.46806e-09, -5.37955e-09, -5.290913e-09, -5.177516e-09,
  -8.616944e-09, -8.405992e-09, -8.104861e-09, -7.416009e-09, -6.810631e-09, 
    -6.304202e-09, -6.098122e-09, -6.081221e-09, -6.070848e-09, 
    -5.804317e-09, -5.419828e-09, -5.092127e-09, -4.839286e-09, 
    -4.594383e-09, -4.400747e-09,
  -9.586218e-09, -8.987167e-09, -8.503765e-09, -7.962143e-09, -7.587039e-09, 
    -7.063191e-09, -6.588308e-09, -6.363346e-09, -6.265159e-09, 
    -6.121748e-09, -5.646665e-09, -5.121195e-09, -4.695914e-09, 
    -4.284821e-09, -4.117918e-09,
  -1.149675e-08, -1.04972e-08, -9.765474e-09, -8.879572e-09, -8.290201e-09, 
    -7.624424e-09, -7.023357e-09, -6.592679e-09, -6.361596e-09, 
    -6.267613e-09, -5.941925e-09, -5.397493e-09, -4.930432e-09, 
    -4.743403e-09, -4.769127e-09,
  -1.349521e-08, -1.238133e-08, -1.141618e-08, -1.060983e-08, -9.79204e-09, 
    -9.046536e-09, -8.174885e-09, -7.330893e-09, -6.718019e-09, 
    -6.368104e-09, -6.18895e-09, -5.930033e-09, -5.53419e-09, -5.438801e-09, 
    -5.768271e-09,
  -1.554228e-08, -1.471545e-08, -1.33063e-08, -1.212692e-08, -1.139002e-08, 
    -1.063309e-08, -9.878818e-09, -9.045319e-09, -8.129165e-09, 
    -7.340097e-09, -6.880395e-09, -6.635934e-09, -6.423815e-09, 
    -6.437487e-09, -6.845882e-09,
  -1.718593e-08, -1.666083e-08, -1.544534e-08, -1.410724e-08, -1.308182e-08, 
    -1.226069e-08, -1.165403e-08, -1.103213e-08, -1.032038e-08, 
    -9.433467e-09, -8.553844e-09, -7.97109e-09, -7.653733e-09, -7.522432e-09, 
    -7.516359e-09,
  -1.87603e-08, -1.822862e-08, -1.712704e-08, -1.583291e-08, -1.485347e-08, 
    -1.380001e-08, -1.28741e-08, -1.233928e-08, -1.194023e-08, -1.145802e-08, 
    -1.082665e-08, -1.008323e-08, -9.577268e-09, -9.222432e-09, -8.856375e-09,
  -2.038223e-08, -1.987414e-08, -1.895985e-08, -1.779158e-08, -1.652172e-08, 
    -1.556274e-08, -1.449065e-08, -1.353758e-08, -1.297339e-08, 
    -1.267542e-08, -1.244168e-08, -1.214904e-08, -1.172457e-08, 
    -1.126418e-08, -1.07331e-08,
  -3.622805e-09, -3.654681e-09, -3.719376e-09, -3.906911e-09, -4.015661e-09, 
    -4.13816e-09, -4.371298e-09, -4.726124e-09, -5.267482e-09, -5.959329e-09, 
    -6.721501e-09, -7.59742e-09, -8.53481e-09, -9.602768e-09, -1.072128e-08,
  -4.175188e-09, -4.204913e-09, -4.284179e-09, -4.394173e-09, -4.511567e-09, 
    -4.711829e-09, -4.966965e-09, -5.371354e-09, -5.950983e-09, 
    -6.633254e-09, -7.389618e-09, -8.243465e-09, -9.221052e-09, 
    -1.027064e-08, -1.136542e-08,
  -4.517311e-09, -4.577092e-09, -4.678619e-09, -4.775631e-09, -4.920115e-09, 
    -5.131388e-09, -5.43805e-09, -5.909178e-09, -6.55268e-09, -7.257468e-09, 
    -8.042231e-09, -8.960601e-09, -9.95905e-09, -1.098182e-08, -1.202531e-08,
  -4.71703e-09, -4.843498e-09, -4.905718e-09, -5.022005e-09, -5.214483e-09, 
    -5.479646e-09, -5.875044e-09, -6.418762e-09, -7.109434e-09, 
    -7.849559e-09, -8.713719e-09, -9.684928e-09, -1.068711e-08, 
    -1.165198e-08, -1.267075e-08,
  -4.943119e-09, -5.131901e-09, -5.169573e-09, -5.301152e-09, -5.527345e-09, 
    -5.894706e-09, -6.36086e-09, -6.949209e-09, -7.635417e-09, -8.430446e-09, 
    -9.348661e-09, -1.03868e-08, -1.1389e-08, -1.235443e-08, -1.341953e-08,
  -5.400052e-09, -5.553859e-09, -5.592018e-09, -5.788759e-09, -6.062693e-09, 
    -6.425454e-09, -6.868467e-09, -7.485164e-09, -8.246861e-09, 
    -9.121158e-09, -1.007583e-08, -1.109065e-08, -1.209371e-08, 
    -1.308709e-08, -1.418065e-08,
  -6.017784e-09, -6.042377e-09, -6.158371e-09, -6.432779e-09, -6.698558e-09, 
    -7.00238e-09, -7.467245e-09, -8.205829e-09, -9.024259e-09, -9.925186e-09, 
    -1.084433e-08, -1.186251e-08, -1.285819e-08, -1.390776e-08, -1.511576e-08,
  -6.80461e-09, -6.769687e-09, -6.852237e-09, -7.04716e-09, -7.258812e-09, 
    -7.630319e-09, -8.239887e-09, -9.030759e-09, -9.848912e-09, 
    -1.074362e-08, -1.164279e-08, -1.265868e-08, -1.367804e-08, 
    -1.482923e-08, -1.609635e-08,
  -7.571452e-09, -7.60823e-09, -7.685197e-09, -7.739287e-09, -8.000586e-09, 
    -8.439978e-09, -9.091513e-09, -9.874904e-09, -1.070456e-08, 
    -1.158725e-08, -1.248117e-08, -1.34938e-08, -1.455021e-08, -1.57079e-08, 
    -1.691984e-08,
  -8.262996e-09, -8.311198e-09, -8.469415e-09, -8.662647e-09, -8.976808e-09, 
    -9.416406e-09, -9.982822e-09, -1.066826e-08, -1.14628e-08, -1.232278e-08, 
    -1.327322e-08, -1.430693e-08, -1.533825e-08, -1.642602e-08, -1.753195e-08,
  -5.883045e-09, -6.554195e-09, -7.181643e-09, -7.883264e-09, -8.653881e-09, 
    -9.661032e-09, -1.072372e-08, -1.181981e-08, -1.312632e-08, 
    -1.459621e-08, -1.602731e-08, -1.740377e-08, -1.860801e-08, 
    -1.933548e-08, -1.972843e-08,
  -6.575545e-09, -7.079838e-09, -7.695477e-09, -8.433457e-09, -9.357537e-09, 
    -1.041978e-08, -1.145472e-08, -1.271571e-08, -1.413689e-08, 
    -1.553083e-08, -1.683998e-08, -1.80947e-08, -1.890877e-08, -1.934899e-08, 
    -2.008615e-08,
  -6.973337e-09, -7.485726e-09, -8.293769e-09, -9.187239e-09, -1.015543e-08, 
    -1.1141e-08, -1.229596e-08, -1.369351e-08, -1.508242e-08, -1.640161e-08, 
    -1.764029e-08, -1.851127e-08, -1.891967e-08, -1.960992e-08, -2.071284e-08,
  -7.281354e-09, -8.082184e-09, -8.998817e-09, -9.759942e-09, -1.07208e-08, 
    -1.187702e-08, -1.317605e-08, -1.456576e-08, -1.585133e-08, 
    -1.707988e-08, -1.797312e-08, -1.853581e-08, -1.919913e-08, 
    -2.032779e-08, -2.128296e-08,
  -7.866017e-09, -8.709103e-09, -9.547228e-09, -1.041927e-08, -1.159779e-08, 
    -1.278558e-08, -1.410769e-08, -1.544947e-08, -1.66543e-08, -1.762213e-08, 
    -1.82336e-08, -1.887469e-08, -1.98052e-08, -2.079294e-08, -2.1562e-08,
  -8.534024e-09, -9.399513e-09, -1.043355e-08, -1.137727e-08, -1.254691e-08, 
    -1.380025e-08, -1.522022e-08, -1.639639e-08, -1.733093e-08, 
    -1.790649e-08, -1.849358e-08, -1.932394e-08, -2.044605e-08, 
    -2.148142e-08, -2.251902e-08,
  -9.427838e-09, -1.028281e-08, -1.134082e-08, -1.233813e-08, -1.37663e-08, 
    -1.511048e-08, -1.62808e-08, -1.701794e-08, -1.759824e-08, -1.819277e-08, 
    -1.901419e-08, -2.029188e-08, -2.138226e-08, -2.222179e-08, -2.305591e-08,
  -1.026925e-08, -1.11661e-08, -1.253018e-08, -1.379751e-08, -1.515098e-08, 
    -1.604059e-08, -1.670235e-08, -1.722502e-08, -1.794102e-08, 
    -1.876455e-08, -2.005518e-08, -2.107573e-08, -2.185704e-08, 
    -2.278739e-08, -2.400638e-08,
  -1.133774e-08, -1.257951e-08, -1.409107e-08, -1.496345e-08, -1.58211e-08, 
    -1.638821e-08, -1.705557e-08, -1.772984e-08, -1.865305e-08, -1.9856e-08, 
    -2.095235e-08, -2.181834e-08, -2.291062e-08, -2.416646e-08, -2.551779e-08,
  -1.299532e-08, -1.403961e-08, -1.508708e-08, -1.565708e-08, -1.638684e-08, 
    -1.694741e-08, -1.771377e-08, -1.86147e-08, -1.983796e-08, -2.081627e-08, 
    -2.181818e-08, -2.295552e-08, -2.42013e-08, -2.533007e-08, -2.52515e-08,
  -1.298636e-08, -1.367544e-08, -1.441115e-08, -1.543876e-08, -1.63307e-08, 
    -1.740346e-08, -1.839926e-08, -1.932732e-08, -2.009128e-08, 
    -2.057509e-08, -2.09423e-08, -2.119539e-08, -2.143309e-08, -2.154443e-08, 
    -2.166873e-08,
  -1.426231e-08, -1.492901e-08, -1.57941e-08, -1.664883e-08, -1.753757e-08, 
    -1.855608e-08, -1.935505e-08, -2.007652e-08, -2.049128e-08, 
    -2.090016e-08, -2.123597e-08, -2.154156e-08, -2.17843e-08, -2.19297e-08, 
    -2.212271e-08,
  -1.487244e-08, -1.566625e-08, -1.665558e-08, -1.76511e-08, -1.866435e-08, 
    -1.954679e-08, -2.024897e-08, -2.079957e-08, -2.115777e-08, 
    -2.144133e-08, -2.161954e-08, -2.173411e-08, -2.181265e-08, 
    -2.200694e-08, -2.235475e-08,
  -1.553065e-08, -1.659235e-08, -1.782e-08, -1.873257e-08, -1.95972e-08, 
    -2.028431e-08, -2.084984e-08, -2.12346e-08, -2.151916e-08, -2.168888e-08, 
    -2.180481e-08, -2.195774e-08, -2.218198e-08, -2.260463e-08, -2.296265e-08,
  -1.662987e-08, -1.777649e-08, -1.893623e-08, -1.965459e-08, -2.039981e-08, 
    -2.093871e-08, -2.136668e-08, -2.163275e-08, -2.180418e-08, 
    -2.197884e-08, -2.226543e-08, -2.261931e-08, -2.301722e-08, 
    -2.345072e-08, -2.40772e-08,
  -1.799e-08, -1.890312e-08, -1.994766e-08, -2.049085e-08, -2.109001e-08, 
    -2.144776e-08, -2.180174e-08, -2.204714e-08, -2.235245e-08, 
    -2.275883e-08, -2.315374e-08, -2.360133e-08, -2.399196e-08, 
    -2.466163e-08, -2.523031e-08,
  -1.891107e-08, -1.968351e-08, -2.070117e-08, -2.097224e-08, -2.151099e-08, 
    -2.184652e-08, -2.234548e-08, -2.27651e-08, -2.322725e-08, -2.364094e-08, 
    -2.406794e-08, -2.45314e-08, -2.514249e-08, -2.566186e-08, -2.573015e-08,
  -1.963993e-08, -2.037461e-08, -2.130224e-08, -2.155706e-08, -2.225589e-08, 
    -2.269174e-08, -2.321527e-08, -2.365926e-08, -2.406468e-08, 
    -2.455216e-08, -2.499828e-08, -2.549081e-08, -2.576438e-08, 
    -2.565939e-08, -2.534387e-08,
  -2.014569e-08, -2.092083e-08, -2.1829e-08, -2.216914e-08, -2.282605e-08, 
    -2.31176e-08, -2.359379e-08, -2.396053e-08, -2.458092e-08, -2.513447e-08, 
    -2.551228e-08, -2.561449e-08, -2.557424e-08, -2.538787e-08, -2.514283e-08,
  -2.097824e-08, -2.174265e-08, -2.258327e-08, -2.281046e-08, -2.325574e-08, 
    -2.359475e-08, -2.407642e-08, -2.463091e-08, -2.507633e-08, 
    -2.517021e-08, -2.51956e-08, -2.529298e-08, -2.537062e-08, -2.518259e-08, 
    -2.481104e-08,
  -1.831286e-08, -1.861384e-08, -1.813957e-08, -1.739917e-08, -1.659535e-08, 
    -1.625587e-08, -1.594632e-08, -1.568901e-08, -1.545409e-08, 
    -1.525269e-08, -1.496789e-08, -1.46881e-08, -1.459507e-08, -1.462927e-08, 
    -1.475196e-08,
  -1.875125e-08, -1.856694e-08, -1.835752e-08, -1.827481e-08, -1.800422e-08, 
    -1.791328e-08, -1.767833e-08, -1.753165e-08, -1.754696e-08, 
    -1.764862e-08, -1.773219e-08, -1.779772e-08, -1.770144e-08, 
    -1.751354e-08, -1.737574e-08,
  -1.922126e-08, -1.899367e-08, -1.898552e-08, -1.884533e-08, -1.873407e-08, 
    -1.863944e-08, -1.849305e-08, -1.825019e-08, -1.79918e-08, -1.794311e-08, 
    -1.803078e-08, -1.810986e-08, -1.829312e-08, -1.834539e-08, -1.828588e-08,
  -1.999896e-08, -1.9816e-08, -1.987117e-08, -1.968059e-08, -1.951514e-08, 
    -1.946745e-08, -1.943416e-08, -1.935127e-08, -1.90727e-08, -1.889416e-08, 
    -1.894844e-08, -1.922891e-08, -1.94738e-08, -1.978559e-08, -2.013034e-08,
  -2.081589e-08, -2.077744e-08, -2.098802e-08, -2.075829e-08, -2.056348e-08, 
    -2.0393e-08, -2.057017e-08, -2.083194e-08, -2.10439e-08, -2.107043e-08, 
    -2.112202e-08, -2.126276e-08, -2.152555e-08, -2.177353e-08, -2.193778e-08,
  -2.143953e-08, -2.143017e-08, -2.194203e-08, -2.182677e-08, -2.186401e-08, 
    -2.164947e-08, -2.169863e-08, -2.195246e-08, -2.232503e-08, 
    -2.243815e-08, -2.24456e-08, -2.2383e-08, -2.242808e-08, -2.250402e-08, 
    -2.263755e-08,
  -2.206577e-08, -2.239115e-08, -2.269745e-08, -2.257877e-08, -2.265529e-08, 
    -2.255527e-08, -2.258331e-08, -2.269162e-08, -2.289486e-08, 
    -2.309859e-08, -2.313951e-08, -2.314101e-08, -2.323521e-08, 
    -2.349489e-08, -2.414588e-08,
  -2.364022e-08, -2.378888e-08, -2.451278e-08, -2.42812e-08, -2.433128e-08, 
    -2.419374e-08, -2.42055e-08, -2.415925e-08, -2.435384e-08, -2.46492e-08, 
    -2.50127e-08, -2.538716e-08, -2.573611e-08, -2.610797e-08, -2.645049e-08,
  -2.477572e-08, -2.538261e-08, -2.607551e-08, -2.638892e-08, -2.660495e-08, 
    -2.642022e-08, -2.626823e-08, -2.611764e-08, -2.606497e-08, 
    -2.619352e-08, -2.647409e-08, -2.669237e-08, -2.675514e-08, 
    -2.659398e-08, -2.625886e-08,
  -2.456871e-08, -2.498383e-08, -2.528576e-08, -2.531445e-08, -2.567719e-08, 
    -2.580254e-08, -2.594366e-08, -2.587917e-08, -2.588242e-08, 
    -2.581207e-08, -2.577229e-08, -2.550334e-08, -2.516033e-08, 
    -2.475111e-08, -2.44403e-08,
  -1.006792e-08, -1.005117e-08, -9.580691e-09, -8.767195e-09, -8.11636e-09, 
    -7.499954e-09, -7.106306e-09, -6.823931e-09, -6.643919e-09, 
    -6.454606e-09, -6.013363e-09, -5.620551e-09, -5.359283e-09, 
    -5.792859e-09, -7.022313e-09,
  -1.053043e-08, -1.093056e-08, -1.093101e-08, -1.038038e-08, -9.998835e-09, 
    -9.711881e-09, -9.360556e-09, -9.023779e-09, -8.542766e-09, 
    -7.966104e-09, -7.270365e-09, -6.819081e-09, -6.841301e-09, 
    -7.569652e-09, -8.868246e-09,
  -1.232015e-08, -1.310967e-08, -1.266771e-08, -1.218748e-08, -1.179621e-08, 
    -1.151446e-08, -1.102125e-08, -1.05421e-08, -9.886191e-09, -9.213453e-09, 
    -8.575976e-09, -8.253269e-09, -8.575839e-09, -9.61716e-09, -1.117036e-08,
  -1.35591e-08, -1.621358e-08, -1.567145e-08, -1.534065e-08, -1.48273e-08, 
    -1.426688e-08, -1.34958e-08, -1.250471e-08, -1.160074e-08, -1.081115e-08, 
    -1.023502e-08, -1.022458e-08, -1.079564e-08, -1.194974e-08, -1.327584e-08,
  -1.550716e-08, -1.818214e-08, -1.755679e-08, -1.718089e-08, -1.652259e-08, 
    -1.58715e-08, -1.495751e-08, -1.406875e-08, -1.320793e-08, -1.245244e-08, 
    -1.214617e-08, -1.236318e-08, -1.292758e-08, -1.375435e-08, -1.457817e-08,
  -1.808534e-08, -1.83895e-08, -1.807589e-08, -1.863322e-08, -1.852663e-08, 
    -1.814703e-08, -1.716683e-08, -1.624347e-08, -1.526633e-08, 
    -1.479599e-08, -1.467293e-08, -1.468054e-08, -1.502372e-08, 
    -1.536624e-08, -1.573947e-08,
  -1.971953e-08, -1.886706e-08, -1.845888e-08, -1.847356e-08, -1.871575e-08, 
    -1.875373e-08, -1.847428e-08, -1.823341e-08, -1.768351e-08, 
    -1.729515e-08, -1.683071e-08, -1.664542e-08, -1.659301e-08, -1.65281e-08, 
    -1.650071e-08,
  -2.106464e-08, -2.017032e-08, -1.966509e-08, -1.921306e-08, -1.906688e-08, 
    -1.87527e-08, -1.869502e-08, -1.860802e-08, -1.846768e-08, -1.832635e-08, 
    -1.808017e-08, -1.775289e-08, -1.742719e-08, -1.715717e-08, -1.703395e-08,
  -2.267846e-08, -2.170086e-08, -2.124045e-08, -2.075108e-08, -2.046523e-08, 
    -2.000249e-08, -1.961098e-08, -1.918467e-08, -1.887935e-08, 
    -1.849591e-08, -1.810528e-08, -1.775234e-08, -1.746895e-08, 
    -1.732539e-08, -1.723807e-08,
  -2.491244e-08, -2.424415e-08, -2.369696e-08, -2.31298e-08, -2.269172e-08, 
    -2.228358e-08, -2.18728e-08, -2.137285e-08, -2.071619e-08, -1.998765e-08, 
    -1.926785e-08, -1.866215e-08, -1.837311e-08, -1.815103e-08, -1.816769e-08,
  -5.350913e-09, -4.461898e-09, -3.981165e-09, -4.139495e-09, -4.868193e-09, 
    -6.073644e-09, -7.266558e-09, -8.321753e-09, -9.411852e-09, 
    -1.079297e-08, -1.239517e-08, -1.39656e-08, -1.56901e-08, -1.754875e-08, 
    -1.904204e-08,
  -5.312017e-09, -4.693663e-09, -4.467612e-09, -4.717797e-09, -5.281297e-09, 
    -5.884575e-09, -6.568637e-09, -7.058794e-09, -8.120971e-09, 
    -9.884098e-09, -1.171756e-08, -1.318877e-08, -1.45474e-08, -1.619429e-08, 
    -1.796179e-08,
  -5.003078e-09, -5.105797e-09, -5.377224e-09, -5.636696e-09, -6.192788e-09, 
    -6.421019e-09, -6.649227e-09, -6.910504e-09, -7.995228e-09, 
    -9.559458e-09, -1.092035e-08, -1.231556e-08, -1.365077e-08, 
    -1.514802e-08, -1.702953e-08,
  -4.231662e-09, -5.038375e-09, -5.393774e-09, -5.907546e-09, -6.649002e-09, 
    -7.127691e-09, -7.414313e-09, -7.780106e-09, -8.716063e-09, 
    -9.725432e-09, -1.080314e-08, -1.182946e-08, -1.291166e-08, 
    -1.456183e-08, -1.663173e-08,
  -4.421476e-09, -5.516943e-09, -5.355371e-09, -5.655386e-09, -6.313248e-09, 
    -6.764627e-09, -7.262159e-09, -7.93632e-09, -8.987077e-09, -1.019842e-08, 
    -1.155949e-08, -1.245692e-08, -1.307073e-08, -1.432421e-08, -1.632281e-08,
  -6.46695e-09, -7.412792e-09, -6.623841e-09, -6.21068e-09, -6.369314e-09, 
    -6.581033e-09, -6.754707e-09, -7.172833e-09, -8.211589e-09, 
    -9.679558e-09, -1.144558e-08, -1.28426e-08, -1.342425e-08, -1.435752e-08, 
    -1.590705e-08,
  -7.371397e-09, -8.864732e-09, -7.949044e-09, -6.976719e-09, -6.574174e-09, 
    -6.370994e-09, -6.317653e-09, -6.453287e-09, -7.336105e-09, 
    -9.157918e-09, -1.095747e-08, -1.208096e-08, -1.273804e-08, 
    -1.367752e-08, -1.492359e-08,
  -7.342926e-09, -9.53075e-09, -8.756196e-09, -8.341517e-09, -7.804963e-09, 
    -7.337741e-09, -7.079454e-09, -6.95906e-09, -7.295128e-09, -8.490991e-09, 
    -1.003053e-08, -1.120932e-08, -1.196197e-08, -1.309061e-08, -1.42561e-08,
  -8.099376e-09, -9.728663e-09, -9.127874e-09, -8.955247e-09, -8.832505e-09, 
    -8.245197e-09, -7.844285e-09, -7.626123e-09, -7.778995e-09, 
    -8.383363e-09, -9.193581e-09, -1.024861e-08, -1.094882e-08, 
    -1.198644e-08, -1.321855e-08,
  -1.046679e-08, -1.028234e-08, -9.580595e-09, -9.676159e-09, -1.012024e-08, 
    -9.162904e-09, -8.29238e-09, -7.620002e-09, -7.334198e-09, -7.709084e-09, 
    -8.337643e-09, -9.042485e-09, -9.80201e-09, -1.096406e-08, -1.280211e-08,
  -1.538743e-08, -1.709515e-08, -1.889705e-08, -2.173129e-08, -2.475068e-08, 
    -2.773365e-08, -2.955666e-08, -2.967762e-08, -2.84249e-08, -2.667157e-08, 
    -2.601914e-08, -2.589778e-08, -2.600149e-08, -2.590505e-08, -2.583846e-08,
  -1.575964e-08, -1.774595e-08, -1.9921e-08, -2.305688e-08, -2.62158e-08, 
    -2.891589e-08, -3.015749e-08, -2.959317e-08, -2.80853e-08, -2.674583e-08, 
    -2.639835e-08, -2.630061e-08, -2.640008e-08, -2.635955e-08, -2.641976e-08,
  -1.589828e-08, -1.794652e-08, -2.058838e-08, -2.38745e-08, -2.686988e-08, 
    -2.907929e-08, -2.971506e-08, -2.841008e-08, -2.71732e-08, -2.627073e-08, 
    -2.617975e-08, -2.632179e-08, -2.655758e-08, -2.672664e-08, -2.691773e-08,
  -1.584766e-08, -1.784015e-08, -2.069903e-08, -2.4173e-08, -2.665068e-08, 
    -2.836761e-08, -2.854613e-08, -2.726633e-08, -2.622748e-08, 
    -2.574127e-08, -2.582368e-08, -2.592957e-08, -2.617464e-08, 
    -2.630928e-08, -2.642136e-08,
  -1.580128e-08, -1.788329e-08, -2.060387e-08, -2.393767e-08, -2.614883e-08, 
    -2.736372e-08, -2.733167e-08, -2.637372e-08, -2.581168e-08, 
    -2.562896e-08, -2.566305e-08, -2.570092e-08, -2.578564e-08, 
    -2.587902e-08, -2.596155e-08,
  -1.584518e-08, -1.780172e-08, -2.049267e-08, -2.360649e-08, -2.547945e-08, 
    -2.640765e-08, -2.636441e-08, -2.579429e-08, -2.565116e-08, 
    -2.571926e-08, -2.609221e-08, -2.616615e-08, -2.610482e-08, 
    -2.617918e-08, -2.602675e-08,
  -1.565907e-08, -1.767761e-08, -2.026871e-08, -2.305216e-08, -2.461923e-08, 
    -2.566822e-08, -2.574363e-08, -2.539184e-08, -2.553862e-08, 
    -2.594845e-08, -2.660571e-08, -2.693351e-08, -2.671737e-08, -2.64398e-08, 
    -2.638243e-08,
  -1.549957e-08, -1.753502e-08, -1.991596e-08, -2.241692e-08, -2.389151e-08, 
    -2.507391e-08, -2.523838e-08, -2.499106e-08, -2.52457e-08, -2.585661e-08, 
    -2.657995e-08, -2.718982e-08, -2.727854e-08, -2.693475e-08, -2.67174e-08,
  -1.531059e-08, -1.737325e-08, -1.96293e-08, -2.191985e-08, -2.341083e-08, 
    -2.477071e-08, -2.49693e-08, -2.477061e-08, -2.50247e-08, -2.551367e-08, 
    -2.63945e-08, -2.674315e-08, -2.69098e-08, -2.693754e-08, -2.691426e-08,
  -1.520615e-08, -1.72072e-08, -1.929833e-08, -2.143679e-08, -2.300706e-08, 
    -2.44346e-08, -2.490468e-08, -2.491929e-08, -2.517442e-08, -2.550304e-08, 
    -2.604831e-08, -2.633047e-08, -2.634177e-08, -2.659435e-08, -2.692272e-08,
  -1.730827e-08, -1.736552e-08, -1.693338e-08, -1.675327e-08, -1.653738e-08, 
    -1.668123e-08, -1.692404e-08, -1.714919e-08, -1.722436e-08, 
    -1.723037e-08, -1.731561e-08, -1.742448e-08, -1.74456e-08, -1.752963e-08, 
    -1.759984e-08,
  -1.738563e-08, -1.72472e-08, -1.676977e-08, -1.66383e-08, -1.669027e-08, 
    -1.708954e-08, -1.732876e-08, -1.726555e-08, -1.713852e-08, 
    -1.721517e-08, -1.73411e-08, -1.74335e-08, -1.753036e-08, -1.761001e-08, 
    -1.770007e-08,
  -1.736188e-08, -1.709244e-08, -1.665247e-08, -1.68088e-08, -1.733205e-08, 
    -1.778674e-08, -1.771506e-08, -1.770454e-08, -1.782858e-08, 
    -1.805034e-08, -1.811008e-08, -1.816905e-08, -1.822662e-08, -1.82662e-08, 
    -1.843179e-08,
  -1.733176e-08, -1.697176e-08, -1.688956e-08, -1.771378e-08, -1.824825e-08, 
    -1.855235e-08, -1.866884e-08, -1.900364e-08, -1.934088e-08, 
    -1.959234e-08, -1.979994e-08, -1.997428e-08, -2.007193e-08, 
    -2.004586e-08, -2.00176e-08,
  -1.733958e-08, -1.71043e-08, -1.756825e-08, -1.833576e-08, -1.878918e-08, 
    -1.906156e-08, -1.94277e-08, -1.982266e-08, -2.019187e-08, -2.062324e-08, 
    -2.092685e-08, -2.121419e-08, -2.131631e-08, -2.139527e-08, -2.137626e-08,
  -1.733643e-08, -1.744099e-08, -1.813915e-08, -1.892647e-08, -1.94192e-08, 
    -1.984646e-08, -2.035611e-08, -2.078358e-08, -2.119901e-08, 
    -2.148843e-08, -2.175153e-08, -2.199033e-08, -2.218294e-08, 
    -2.227836e-08, -2.237948e-08,
  -1.754119e-08, -1.787028e-08, -1.875857e-08, -1.967998e-08, -2.019835e-08, 
    -2.065503e-08, -2.109723e-08, -2.154993e-08, -2.192649e-08, 
    -2.232721e-08, -2.25424e-08, -2.275249e-08, -2.27667e-08, -2.28492e-08, 
    -2.30312e-08,
  -1.76627e-08, -1.824012e-08, -1.938197e-08, -2.04947e-08, -2.100469e-08, 
    -2.159291e-08, -2.213603e-08, -2.26118e-08, -2.307402e-08, -2.316802e-08, 
    -2.320346e-08, -2.32378e-08, -2.342559e-08, -2.362808e-08, -2.379763e-08,
  -1.78578e-08, -1.873126e-08, -2.018871e-08, -2.141681e-08, -2.188502e-08, 
    -2.271214e-08, -2.32605e-08, -2.371709e-08, -2.3842e-08, -2.404069e-08, 
    -2.420099e-08, -2.450305e-08, -2.467421e-08, -2.485533e-08, -2.508393e-08,
  -1.810221e-08, -1.934049e-08, -2.104271e-08, -2.23996e-08, -2.304605e-08, 
    -2.367665e-08, -2.396379e-08, -2.403645e-08, -2.44813e-08, -2.483331e-08, 
    -2.511293e-08, -2.54545e-08, -2.552128e-08, -2.593703e-08, -2.599216e-08,
  -2.089344e-08, -2.078322e-08, -2.064305e-08, -2.063775e-08, -2.061032e-08, 
    -2.073774e-08, -2.120165e-08, -2.193153e-08, -2.219428e-08, -2.27265e-08, 
    -2.223457e-08, -2.194178e-08, -2.1713e-08, -2.160979e-08, -2.163664e-08,
  -2.104958e-08, -2.096326e-08, -2.072339e-08, -2.059561e-08, -2.049072e-08, 
    -2.062075e-08, -2.106655e-08, -2.15815e-08, -2.221426e-08, -2.229179e-08, 
    -2.171154e-08, -2.151818e-08, -2.132698e-08, -2.117739e-08, -2.163539e-08,
  -2.144148e-08, -2.113283e-08, -2.066113e-08, -2.033632e-08, -2.027956e-08, 
    -2.057328e-08, -2.097796e-08, -2.156873e-08, -2.195475e-08, 
    -2.175435e-08, -2.152563e-08, -2.138303e-08, -2.108713e-08, -2.12236e-08, 
    -2.197153e-08,
  -2.160066e-08, -2.081111e-08, -2.028724e-08, -1.999588e-08, -2.006488e-08, 
    -2.038331e-08, -2.075419e-08, -2.122572e-08, -2.139284e-08, 
    -2.116635e-08, -2.120271e-08, -2.106022e-08, -2.105946e-08, 
    -2.141249e-08, -2.215752e-08,
  -2.151551e-08, -2.066365e-08, -2.032333e-08, -2.001392e-08, -2.002955e-08, 
    -2.035493e-08, -2.060565e-08, -2.086987e-08, -2.085705e-08, 
    -2.091602e-08, -2.119453e-08, -2.09229e-08, -2.100511e-08, -2.146124e-08, 
    -2.203459e-08,
  -2.143126e-08, -2.069984e-08, -2.039863e-08, -2.003897e-08, -2.012697e-08, 
    -2.01278e-08, -2.044922e-08, -2.055164e-08, -2.064466e-08, -2.094356e-08, 
    -2.112789e-08, -2.077563e-08, -2.101078e-08, -2.149065e-08, -2.19458e-08,
  -2.111569e-08, -2.072386e-08, -2.047272e-08, -2.019115e-08, -2.022728e-08, 
    -2.020423e-08, -2.049603e-08, -2.057357e-08, -2.073638e-08, -2.09386e-08, 
    -2.089664e-08, -2.081851e-08, -2.112538e-08, -2.165597e-08, -2.210335e-08,
  -2.08262e-08, -2.077718e-08, -2.056281e-08, -2.032086e-08, -2.032342e-08, 
    -2.022262e-08, -2.038474e-08, -2.041782e-08, -2.064474e-08, 
    -2.072531e-08, -2.061235e-08, -2.080825e-08, -2.117431e-08, 
    -2.171526e-08, -2.201781e-08,
  -2.082321e-08, -2.083418e-08, -2.06889e-08, -2.044148e-08, -2.022829e-08, 
    -2.004963e-08, -2.013516e-08, -2.03249e-08, -2.067893e-08, -2.074124e-08, 
    -2.080362e-08, -2.10597e-08, -2.140907e-08, -2.175637e-08, -2.188031e-08,
  -2.055361e-08, -2.070933e-08, -2.084262e-08, -2.038327e-08, -2.014943e-08, 
    -1.999808e-08, -2.006351e-08, -2.057314e-08, -2.106289e-08, 
    -2.130861e-08, -2.140044e-08, -2.148991e-08, -2.167687e-08, 
    -2.188741e-08, -2.178024e-08,
  -2.241732e-08, -2.298637e-08, -2.345379e-08, -2.383804e-08, -2.413319e-08, 
    -2.415528e-08, -2.410648e-08, -2.434245e-08, -2.412208e-08, 
    -2.395262e-08, -2.39585e-08, -2.398332e-08, -2.409146e-08, -2.431103e-08, 
    -2.4529e-08,
  -2.272732e-08, -2.32228e-08, -2.369783e-08, -2.401822e-08, -2.408134e-08, 
    -2.40309e-08, -2.401361e-08, -2.413337e-08, -2.4117e-08, -2.40764e-08, 
    -2.403204e-08, -2.417126e-08, -2.439124e-08, -2.453072e-08, -2.469288e-08,
  -2.291435e-08, -2.337049e-08, -2.390126e-08, -2.420493e-08, -2.412834e-08, 
    -2.41101e-08, -2.413679e-08, -2.440328e-08, -2.426617e-08, -2.430765e-08, 
    -2.415586e-08, -2.431984e-08, -2.451707e-08, -2.46685e-08, -2.479791e-08,
  -2.30326e-08, -2.34847e-08, -2.404304e-08, -2.426995e-08, -2.409871e-08, 
    -2.419858e-08, -2.413206e-08, -2.448589e-08, -2.434765e-08, 
    -2.430163e-08, -2.406251e-08, -2.432178e-08, -2.453873e-08, 
    -2.462701e-08, -2.469195e-08,
  -2.306362e-08, -2.354043e-08, -2.40876e-08, -2.42113e-08, -2.4096e-08, 
    -2.408834e-08, -2.410314e-08, -2.4436e-08, -2.434208e-08, -2.422233e-08, 
    -2.39537e-08, -2.424047e-08, -2.441611e-08, -2.44345e-08, -2.447589e-08,
  -2.307594e-08, -2.355929e-08, -2.398328e-08, -2.39899e-08, -2.386809e-08, 
    -2.403428e-08, -2.402751e-08, -2.425729e-08, -2.426256e-08, 
    -2.414563e-08, -2.384377e-08, -2.409936e-08, -2.427576e-08, 
    -2.431605e-08, -2.425969e-08,
  -2.304501e-08, -2.343349e-08, -2.379849e-08, -2.371957e-08, -2.366162e-08, 
    -2.378386e-08, -2.389122e-08, -2.412019e-08, -2.405615e-08, 
    -2.395004e-08, -2.377917e-08, -2.40361e-08, -2.426824e-08, -2.430811e-08, 
    -2.415882e-08,
  -2.307063e-08, -2.332203e-08, -2.347911e-08, -2.338162e-08, -2.353163e-08, 
    -2.355232e-08, -2.365055e-08, -2.375788e-08, -2.387163e-08, 
    -2.388191e-08, -2.375386e-08, -2.406881e-08, -2.438074e-08, 
    -2.433275e-08, -2.423214e-08,
  -2.301495e-08, -2.31211e-08, -2.324941e-08, -2.325386e-08, -2.333769e-08, 
    -2.345027e-08, -2.351282e-08, -2.367721e-08, -2.370946e-08, 
    -2.366469e-08, -2.37751e-08, -2.41611e-08, -2.442179e-08, -2.433288e-08, 
    -2.42043e-08,
  -2.318107e-08, -2.308713e-08, -2.304461e-08, -2.299161e-08, -2.321238e-08, 
    -2.312949e-08, -2.333605e-08, -2.345439e-08, -2.380125e-08, 
    -2.383504e-08, -2.389689e-08, -2.427571e-08, -2.435254e-08, -2.41817e-08, 
    -2.420876e-08,
  -2.295304e-08, -2.294734e-08, -2.285281e-08, -2.26034e-08, -2.245867e-08, 
    -2.233532e-08, -2.23197e-08, -2.226347e-08, -2.222483e-08, -2.218708e-08, 
    -2.212097e-08, -2.203024e-08, -2.199737e-08, -2.203059e-08, -2.216175e-08,
  -2.262918e-08, -2.233459e-08, -2.222131e-08, -2.216653e-08, -2.223202e-08, 
    -2.229225e-08, -2.234987e-08, -2.236381e-08, -2.23905e-08, -2.246819e-08, 
    -2.256902e-08, -2.272542e-08, -2.293114e-08, -2.318765e-08, -2.339189e-08,
  -2.245209e-08, -2.221567e-08, -2.223612e-08, -2.229494e-08, -2.233367e-08, 
    -2.235503e-08, -2.245552e-08, -2.264752e-08, -2.292184e-08, 
    -2.319003e-08, -2.346157e-08, -2.372373e-08, -2.400926e-08, 
    -2.427129e-08, -2.441796e-08,
  -2.250153e-08, -2.231671e-08, -2.24493e-08, -2.25557e-08, -2.276788e-08, 
    -2.300615e-08, -2.333556e-08, -2.364153e-08, -2.401909e-08, 
    -2.434087e-08, -2.466338e-08, -2.490668e-08, -2.510293e-08, 
    -2.521603e-08, -2.527385e-08,
  -2.286873e-08, -2.294355e-08, -2.321284e-08, -2.326671e-08, -2.363479e-08, 
    -2.392596e-08, -2.434881e-08, -2.464625e-08, -2.497704e-08, 
    -2.523543e-08, -2.543276e-08, -2.552486e-08, -2.559424e-08, 
    -2.560559e-08, -2.560568e-08,
  -2.331965e-08, -2.346503e-08, -2.37084e-08, -2.399195e-08, -2.440193e-08, 
    -2.477102e-08, -2.515258e-08, -2.546827e-08, -2.579491e-08, 
    -2.599973e-08, -2.60757e-08, -2.607664e-08, -2.600773e-08, -2.588841e-08, 
    -2.581264e-08,
  -2.36521e-08, -2.403955e-08, -2.46648e-08, -2.49102e-08, -2.520179e-08, 
    -2.554683e-08, -2.592403e-08, -2.617943e-08, -2.634216e-08, -2.63054e-08, 
    -2.623747e-08, -2.607888e-08, -2.592716e-08, -2.576903e-08, -2.562661e-08,
  -2.410089e-08, -2.455556e-08, -2.523896e-08, -2.550018e-08, -2.582569e-08, 
    -2.604514e-08, -2.627033e-08, -2.644188e-08, -2.649179e-08, 
    -2.646358e-08, -2.639847e-08, -2.620072e-08, -2.600978e-08, -2.56991e-08, 
    -2.53856e-08,
  -2.436578e-08, -2.50154e-08, -2.578828e-08, -2.615076e-08, -2.629357e-08, 
    -2.637372e-08, -2.651643e-08, -2.661058e-08, -2.649075e-08, 
    -2.648401e-08, -2.632097e-08, -2.613387e-08, -2.583457e-08, 
    -2.555252e-08, -2.518579e-08,
  -2.450975e-08, -2.523742e-08, -2.605578e-08, -2.62445e-08, -2.631414e-08, 
    -2.65183e-08, -2.662736e-08, -2.669403e-08, -2.650878e-08, -2.623486e-08, 
    -2.599898e-08, -2.572954e-08, -2.542065e-08, -2.51414e-08, -2.486229e-08,
  -2.209734e-08, -2.188663e-08, -2.17265e-08, -2.153701e-08, -2.134567e-08, 
    -2.113609e-08, -2.094074e-08, -2.070286e-08, -2.049276e-08, -2.0302e-08, 
    -2.015632e-08, -2.003584e-08, -1.996492e-08, -1.991032e-08, -1.991313e-08,
  -2.216497e-08, -2.207074e-08, -2.193688e-08, -2.176213e-08, -2.150456e-08, 
    -2.129307e-08, -2.112483e-08, -2.098044e-08, -2.087334e-08, 
    -2.075899e-08, -2.064029e-08, -2.055816e-08, -2.051029e-08, 
    -2.052824e-08, -2.060271e-08,
  -2.163186e-08, -2.172102e-08, -2.162932e-08, -2.162895e-08, -2.150903e-08, 
    -2.146525e-08, -2.1367e-08, -2.133556e-08, -2.128198e-08, -2.126246e-08, 
    -2.123409e-08, -2.120929e-08, -2.120668e-08, -2.120191e-08, -2.124701e-08,
  -2.149151e-08, -2.158972e-08, -2.158641e-08, -2.167212e-08, -2.168475e-08, 
    -2.175117e-08, -2.172337e-08, -2.171759e-08, -2.165631e-08, -2.16464e-08, 
    -2.164002e-08, -2.167217e-08, -2.172284e-08, -2.1803e-08, -2.196791e-08,
  -2.192625e-08, -2.198726e-08, -2.20291e-08, -2.21151e-08, -2.21773e-08, 
    -2.225088e-08, -2.224204e-08, -2.222601e-08, -2.217815e-08, 
    -2.217064e-08, -2.217736e-08, -2.223345e-08, -2.229845e-08, 
    -2.246673e-08, -2.264281e-08,
  -2.214264e-08, -2.235047e-08, -2.245691e-08, -2.258765e-08, -2.264356e-08, 
    -2.272708e-08, -2.27604e-08, -2.278326e-08, -2.274731e-08, -2.275e-08, 
    -2.278479e-08, -2.281797e-08, -2.291653e-08, -2.303792e-08, -2.318946e-08,
  -2.215924e-08, -2.23968e-08, -2.257432e-08, -2.279744e-08, -2.297346e-08, 
    -2.310308e-08, -2.321964e-08, -2.327558e-08, -2.32775e-08, -2.322309e-08, 
    -2.319817e-08, -2.319177e-08, -2.32319e-08, -2.321562e-08, -2.320927e-08,
  -2.234578e-08, -2.249461e-08, -2.28477e-08, -2.30063e-08, -2.323913e-08, 
    -2.344663e-08, -2.359281e-08, -2.369924e-08, -2.368418e-08, 
    -2.359778e-08, -2.345279e-08, -2.342889e-08, -2.330566e-08, 
    -2.331599e-08, -2.333925e-08,
  -2.258105e-08, -2.281859e-08, -2.303145e-08, -2.325925e-08, -2.366216e-08, 
    -2.36972e-08, -2.389313e-08, -2.403167e-08, -2.419302e-08, -2.420435e-08, 
    -2.402324e-08, -2.387728e-08, -2.373375e-08, -2.358333e-08, -2.349075e-08,
  -2.30087e-08, -2.309745e-08, -2.319287e-08, -2.36402e-08, -2.371499e-08, 
    -2.392787e-08, -2.397684e-08, -2.409214e-08, -2.407108e-08, 
    -2.417679e-08, -2.412408e-08, -2.413e-08, -2.402246e-08, -2.38266e-08, 
    -2.363178e-08,
  -1.469143e-08, -1.41244e-08, -1.378521e-08, -1.351482e-08, -1.333088e-08, 
    -1.315009e-08, -1.305332e-08, -1.304866e-08, -1.314056e-08, 
    -1.335878e-08, -1.371117e-08, -1.418213e-08, -1.465396e-08, 
    -1.506429e-08, -1.546961e-08,
  -1.594204e-08, -1.52873e-08, -1.490747e-08, -1.457406e-08, -1.434571e-08, 
    -1.411891e-08, -1.400188e-08, -1.395956e-08, -1.401791e-08, 
    -1.419308e-08, -1.451367e-08, -1.488836e-08, -1.527231e-08, 
    -1.566077e-08, -1.610761e-08,
  -1.707644e-08, -1.644221e-08, -1.598368e-08, -1.563759e-08, -1.535964e-08, 
    -1.509556e-08, -1.491857e-08, -1.480978e-08, -1.480197e-08, 
    -1.491477e-08, -1.51631e-08, -1.547803e-08, -1.5785e-08, -1.623698e-08, 
    -1.679456e-08,
  -1.819008e-08, -1.749932e-08, -1.700243e-08, -1.659308e-08, -1.629421e-08, 
    -1.601048e-08, -1.579687e-08, -1.565978e-08, -1.562119e-08, -1.56731e-08, 
    -1.583548e-08, -1.607475e-08, -1.637724e-08, -1.680779e-08, -1.74172e-08,
  -1.928978e-08, -1.852295e-08, -1.804744e-08, -1.755948e-08, -1.728897e-08, 
    -1.696377e-08, -1.674733e-08, -1.657903e-08, -1.652154e-08, 
    -1.654788e-08, -1.668385e-08, -1.690796e-08, -1.717101e-08, -1.75391e-08, 
    -1.807544e-08,
  -2.057422e-08, -1.971049e-08, -1.926437e-08, -1.871348e-08, -1.833645e-08, 
    -1.796843e-08, -1.774401e-08, -1.757735e-08, -1.74979e-08, -1.746493e-08, 
    -1.755221e-08, -1.772515e-08, -1.797014e-08, -1.830122e-08, -1.883605e-08,
  -2.16657e-08, -2.100227e-08, -2.052984e-08, -2.000589e-08, -1.950938e-08, 
    -1.911652e-08, -1.879705e-08, -1.858552e-08, -1.8472e-08, -1.8446e-08, 
    -1.847268e-08, -1.856232e-08, -1.869776e-08, -1.899973e-08, -1.952779e-08,
  -2.233393e-08, -2.198917e-08, -2.164732e-08, -2.115595e-08, -2.075323e-08, 
    -2.028121e-08, -2.004305e-08, -1.972643e-08, -1.95627e-08, -1.94645e-08, 
    -1.944882e-08, -1.948678e-08, -1.958637e-08, -1.982399e-08, -2.011435e-08,
  -2.289013e-08, -2.281676e-08, -2.258014e-08, -2.227546e-08, -2.190963e-08, 
    -2.154042e-08, -2.116274e-08, -2.087638e-08, -2.061257e-08, 
    -2.040095e-08, -2.024315e-08, -2.023226e-08, -2.030626e-08, 
    -2.046918e-08, -2.065214e-08,
  -2.330533e-08, -2.331202e-08, -2.322231e-08, -2.305342e-08, -2.28697e-08, 
    -2.264916e-08, -2.237519e-08, -2.201638e-08, -2.167027e-08, 
    -2.143939e-08, -2.123228e-08, -2.105881e-08, -2.100146e-08, 
    -2.101006e-08, -2.118037e-08 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
