netcdf atmos_daily.00010101-00010701.pr.tile2 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float pr(time, grid_yt, grid_xt) ;
		pr:_FillValue = 1.e+20f ;
		pr:missing_value = 1.e+20f ;
		pr:units = "kg m-2 s-1" ;
		pr:long_name = "Precipitation" ;
		pr:cell_methods = "time: mean" ;
		pr:cell_measures = "area: area" ;
		pr:time_avg_info = "average_T1,average_T2,average_DT" ;
		pr:standard_name = "precipitation_flux" ;
		pr:interp_method = "conserve_order1" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:53:56 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile2.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile2.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 pr =
  1.161729e-05, 1.691405e-05, 1.638349e-05, 1.908949e-05, 2.157779e-05, 
    2.62694e-05, 2.886319e-05, 3.286671e-05, 3.166102e-05, 3.123579e-05, 
    5.729376e-05, 7.38681e-05, 5.774912e-05, 4.89551e-05, 5.128553e-05,
  1.25271e-05, 1.325042e-05, 1.642345e-05, 1.832482e-05, 1.983746e-05, 
    2.074077e-05, 2.384928e-05, 2.674543e-05, 2.576235e-05, 3.212753e-05, 
    3.604858e-05, 3.744663e-05, 4.725956e-05, 4.675364e-05, 3.297852e-05,
  8.096754e-06, 1.100705e-05, 1.702678e-05, 1.494308e-05, 1.735297e-05, 
    1.95243e-05, 2.20908e-05, 2.221207e-05, 2.531315e-05, 2.533537e-05, 
    2.68388e-05, 2.95811e-05, 3.252202e-05, 3.361184e-05, 2.419308e-05,
  5.124451e-06, 5.991461e-06, 1.243942e-05, 1.59606e-05, 1.669228e-05, 
    1.866712e-05, 1.901583e-05, 2.079517e-05, 2.026773e-05, 2.275752e-05, 
    2.341321e-05, 2.058888e-05, 1.77624e-05, 1.514094e-05, 1.195226e-05,
  2.73727e-05, 6.932391e-06, 7.833943e-06, 7.460317e-06, 1.262667e-05, 
    1.684751e-05, 1.616481e-05, 1.394697e-05, 1.520678e-05, 1.415674e-05, 
    1.360939e-05, 1.113266e-05, 1.083183e-05, 9.524561e-06, 9.838932e-06,
  9.419558e-05, 6.635887e-05, 2.026926e-05, 7.443448e-06, 7.670113e-06, 
    1.088731e-05, 8.680609e-06, 9.464618e-06, 9.851902e-06, 7.267643e-06, 
    7.461239e-06, 5.438018e-06, 6.557515e-06, 5.459541e-06, 5.319988e-06,
  0.0001101841, 0.0001169144, 9.56929e-05, 2.533108e-05, 3.243794e-06, 
    4.233695e-06, 5.491492e-06, 5.892324e-06, 5.115023e-06, 3.527996e-06, 
    3.232419e-06, 1.735499e-06, 2.121616e-06, 3.225198e-06, 4.002029e-06,
  0.0001608843, 0.0001230568, 0.0001256996, 7.375111e-05, 8.613373e-06, 
    6.602568e-07, 1.882308e-06, 3.386407e-06, 4.918399e-06, 2.694105e-06, 
    2.603405e-06, 1.032967e-06, 2.363221e-06, 3.010267e-06, 4.379255e-06,
  0.0002236797, 0.0001567304, 7.000624e-05, 4.795725e-05, 1.582928e-05, 
    2.166598e-06, 3.368054e-06, 4.026913e-06, 3.008117e-06, 2.137669e-06, 
    1.639845e-06, 2.18388e-06, 2.998048e-06, 5.334242e-06, 1.038257e-05,
  8.43892e-05, 7.462402e-05, 4.140318e-05, 2.627085e-05, 2.237191e-05, 
    1.300372e-05, 3.515723e-06, 2.505172e-06, 2.019738e-06, 1.633171e-06, 
    4.039902e-06, 2.075866e-06, 5.677262e-06, 1.404849e-05, 3.011666e-05,
  1.762383e-06, 2.36441e-06, 3.308956e-06, 5.368666e-06, 5.589327e-06, 
    7.921484e-06, 8.895505e-06, 1.197609e-05, 1.336903e-05, 1.513996e-05, 
    1.741214e-05, 1.909757e-05, 1.660041e-05, 1.500468e-05, 1.631331e-05,
  1.575226e-06, 1.177028e-06, 1.927537e-06, 2.328655e-06, 2.479722e-06, 
    4.320089e-06, 5.116291e-06, 6.542308e-06, 7.293909e-06, 7.903625e-06, 
    7.926939e-06, 7.627533e-06, 8.897496e-06, 1.031578e-05, 2.857368e-05,
  8.698723e-07, 1.145568e-06, 1.324162e-06, 1.455282e-06, 1.966147e-06, 
    2.990517e-06, 4.451485e-06, 3.641481e-06, 3.354548e-06, 5.206269e-06, 
    5.794736e-06, 8.435684e-06, 8.145939e-06, 1.130537e-05, 1.925593e-05,
  1.974582e-06, 1.435795e-06, 2.408525e-06, 1.604121e-06, 9.814516e-07, 
    1.461023e-06, 2.327216e-06, 2.806721e-06, 2.870065e-06, 2.636827e-06, 
    3.574821e-06, 8.751943e-06, 1.187878e-05, 1.81033e-05, 2.329342e-05,
  4.066411e-06, 2.999151e-06, 3.909696e-06, 4.796967e-06, 4.293325e-06, 
    3.69763e-06, 3.213311e-06, 4.536147e-06, 3.874054e-06, 5.667584e-06, 
    7.848234e-06, 9.237056e-06, 1.133333e-05, 1.363421e-05, 1.412673e-05,
  3.909884e-06, 2.583783e-06, 3.159113e-06, 3.87686e-06, 4.763878e-06, 
    5.050102e-06, 5.733659e-06, 6.780832e-06, 6.753802e-06, 6.818446e-06, 
    7.956594e-06, 1.017428e-05, 1.135897e-05, 1.077168e-05, 9.796132e-06,
  2.603891e-06, 1.926644e-06, 1.451241e-06, 2.098363e-06, 3.046049e-06, 
    4.657358e-06, 6.663771e-06, 8.998886e-06, 1.002371e-05, 1.054478e-05, 
    8.460161e-06, 1.069278e-05, 8.771702e-06, 7.272037e-06, 4.031264e-06,
  1.491636e-06, 1.273118e-05, 7.75864e-06, 3.948282e-06, 4.005991e-06, 
    4.046918e-06, 5.869841e-06, 7.163429e-06, 1.010696e-05, 8.768746e-06, 
    9.915009e-06, 7.913999e-06, 5.347454e-06, 4.591527e-06, 2.469481e-06,
  1.066892e-05, 2.243374e-05, 4.328568e-05, 3.493839e-05, 1.698216e-05, 
    4.080326e-06, 5.032727e-06, 7.828149e-06, 7.284579e-06, 8.013233e-06, 
    9.732737e-06, 5.975433e-06, 3.690671e-06, 2.606685e-06, 2.550634e-06,
  1.813638e-05, 5.725259e-05, 0.0001131333, 6.662159e-05, 3.125816e-05, 
    1.10207e-05, 4.584308e-06, 5.06709e-06, 5.535086e-06, 4.212909e-06, 
    3.659449e-06, 3.180579e-06, 2.243436e-06, 2.155381e-06, 2.472514e-06,
  5.333446e-06, 9.545482e-06, 9.527655e-06, 1.18347e-05, 1.346291e-05, 
    1.210652e-05, 1.38228e-05, 1.801451e-05, 1.651634e-05, 1.946675e-05, 
    1.454241e-05, 9.383085e-06, 7.569353e-06, 8.723363e-06, 1.300281e-05,
  4.775596e-06, 5.650654e-06, 7.180218e-06, 9.960591e-06, 1.313199e-05, 
    1.054423e-05, 1.30682e-05, 1.19334e-05, 1.565062e-05, 1.539624e-05, 
    2.030749e-05, 1.804458e-05, 1.574238e-05, 1.651573e-05, 1.465147e-05,
  3.258471e-06, 2.97571e-06, 5.751221e-06, 7.42369e-06, 1.030489e-05, 
    8.249031e-06, 1.430043e-05, 1.256109e-05, 1.089605e-05, 1.407541e-05, 
    1.617889e-05, 1.803271e-05, 2.33032e-05, 2.123457e-05, 2.113821e-05,
  2.221935e-06, 3.240792e-06, 3.013796e-06, 4.425149e-06, 5.109761e-06, 
    7.599896e-06, 9.584363e-06, 1.148191e-05, 1.353002e-05, 1.054295e-05, 
    1.081748e-05, 1.475674e-05, 1.597393e-05, 1.83217e-05, 1.902551e-05,
  1.719231e-06, 2.415078e-06, 2.417012e-06, 1.727454e-06, 3.444857e-06, 
    5.59015e-06, 6.880432e-06, 8.11486e-06, 1.117236e-05, 1.109941e-05, 
    1.084242e-05, 9.76675e-06, 1.081475e-05, 1.067768e-05, 1.288274e-05,
  4.342964e-06, 2.682163e-06, 1.756717e-06, 3.265477e-06, 2.093108e-06, 
    3.044194e-06, 3.903638e-06, 3.911591e-06, 4.979398e-06, 4.404352e-06, 
    7.573501e-06, 7.195499e-06, 7.585663e-06, 5.949825e-06, 6.50982e-06,
  2.402371e-06, 4.868076e-06, 4.74062e-06, 4.891233e-06, 3.806239e-06, 
    3.888773e-06, 4.072929e-06, 3.513869e-06, 3.738864e-06, 5.379482e-06, 
    4.619132e-06, 3.85677e-06, 4.638858e-06, 2.811288e-06, 2.169594e-06,
  5.483751e-06, 4.219946e-06, 5.610208e-06, 3.305419e-06, 6.484638e-06, 
    5.076728e-06, 5.109236e-06, 4.435145e-06, 3.422964e-06, 3.845312e-06, 
    3.849208e-06, 3.376936e-06, 2.70139e-06, 3.020176e-06, 3.643966e-06,
  9.018742e-06, 7.806046e-06, 4.049586e-06, 5.124555e-06, 5.339355e-06, 
    8.23859e-06, 7.191591e-06, 7.484635e-06, 5.303164e-06, 3.131624e-06, 
    3.90733e-06, 3.458953e-06, 5.199756e-06, 4.529644e-06, 4.132579e-06,
  4.852282e-06, 8.447524e-06, 5.207195e-06, 5.926567e-06, 7.821715e-06, 
    6.871259e-06, 9.841346e-06, 8.663387e-06, 5.250335e-06, 5.173093e-06, 
    6.626219e-06, 6.648645e-06, 6.250187e-06, 4.310292e-06, 5.162629e-06,
  4.113192e-06, 5.122034e-06, 7.787023e-06, 8.406569e-06, 9.485972e-06, 
    5.498837e-06, 4.041851e-06, 3.194109e-06, 7.958876e-07, 5.194572e-07, 
    7.787187e-07, 1.717527e-06, 2.174162e-06, 2.927592e-06, 5.17507e-06,
  7.011364e-06, 4.416693e-06, 4.217417e-06, 5.335227e-06, 7.718942e-06, 
    1.042801e-05, 6.756301e-06, 4.452386e-06, 2.116621e-06, 4.896918e-08, 
    9.901947e-08, 6.594531e-08, 1.960993e-07, 1.791115e-06, 3.318553e-06,
  5.711537e-06, 4.926861e-06, 3.294143e-06, 3.383363e-06, 4.945586e-06, 
    7.900102e-06, 6.660354e-06, 5.148081e-06, 2.614468e-06, 2.394247e-07, 
    5.668431e-07, 8.864809e-08, 9.130057e-08, 2.378534e-07, 6.061284e-07,
  6.68131e-06, 4.982141e-06, 2.291666e-06, 2.142856e-06, 3.054678e-06, 
    4.523653e-06, 7.516993e-06, 6.451444e-06, 2.794925e-06, 8.268484e-07, 
    2.363611e-07, 1.560586e-07, 9.680618e-08, 7.545106e-08, 1.364658e-07,
  5.217485e-06, 5.254973e-06, 2.466124e-06, 2.33748e-06, 1.584508e-06, 
    3.320929e-06, 4.707857e-06, 7.074599e-06, 5.180226e-06, 3.502855e-06, 
    1.756911e-06, 5.880646e-07, 1.205496e-07, 4.2075e-07, 4.741851e-08,
  4.835652e-06, 5.560567e-06, 4.443205e-06, 2.054647e-06, 3.373759e-06, 
    2.788015e-06, 4.373658e-06, 4.766961e-06, 6.196147e-06, 6.205556e-06, 
    5.834204e-06, 3.162541e-06, 1.726227e-06, 3.712625e-07, 9.703388e-08,
  5.924977e-06, 5.001574e-06, 5.091302e-06, 2.96902e-06, 3.519411e-06, 
    2.665059e-06, 3.838902e-06, 5.134516e-06, 6.284945e-06, 6.720647e-06, 
    5.882934e-06, 6.840804e-06, 4.229988e-06, 3.512616e-06, 2.393808e-06,
  6.164057e-06, 5.725035e-06, 7.156517e-06, 3.512005e-06, 3.374666e-06, 
    3.989916e-06, 3.244555e-06, 4.257578e-06, 5.721292e-06, 6.753886e-06, 
    7.086722e-06, 4.934699e-06, 4.795424e-06, 5.999069e-06, 7.257336e-06,
  6.732395e-06, 5.4554e-06, 4.0881e-06, 6.435231e-06, 4.799153e-06, 
    3.725788e-06, 3.932257e-06, 5.992259e-06, 4.583966e-06, 6.694808e-06, 
    6.782401e-06, 7.73894e-06, 5.008565e-06, 5.465544e-06, 4.726729e-06,
  5.848838e-06, 4.607046e-06, 3.982923e-06, 4.893005e-06, 2.262674e-06, 
    3.041054e-06, 3.869164e-06, 4.898465e-06, 5.283214e-06, 5.398772e-06, 
    4.636017e-06, 4.296802e-06, 4.746151e-06, 4.305907e-06, 3.555525e-06,
  1.342609e-06, 2.891465e-06, 4.227094e-06, 3.994607e-06, 4.49023e-06, 
    3.090478e-06, 5.445569e-06, 5.819451e-06, 2.317007e-06, 5.652239e-06, 
    3.342366e-06, 2.476726e-06, 2.459408e-06, 6.371035e-07, 1.397292e-06,
  1.221278e-05, 7.042825e-06, 3.704447e-06, 5.771453e-06, 3.626923e-06, 
    5.190987e-06, 4.019309e-06, 5.699018e-06, 3.924801e-06, 1.361644e-06, 
    2.848241e-06, 2.066287e-06, 1.241418e-06, 2.350323e-06, 1.477471e-06,
  1.278811e-05, 8.043646e-06, 8.824355e-06, 6.486276e-06, 6.464908e-06, 
    8.448308e-06, 4.782712e-06, 3.00939e-06, 3.099962e-06, 2.917675e-06, 
    1.693696e-06, 3.304785e-06, 2.862976e-06, 3.296479e-06, 2.590326e-06,
  1.429115e-05, 7.373927e-06, 1.053621e-05, 6.894718e-06, 9.916724e-06, 
    9.793825e-06, 4.476181e-06, 5.183161e-06, 4.353082e-06, 1.194439e-06, 
    1.065951e-06, 1.457524e-06, 2.74649e-06, 4.477355e-06, 2.592402e-06,
  1.405856e-05, 1.186093e-05, 6.33993e-06, 7.519558e-06, 1.068512e-05, 
    1.273772e-05, 1.266447e-05, 1.110316e-05, 8.654293e-06, 5.752043e-06, 
    2.049998e-06, 3.07973e-06, 1.858006e-06, 2.026664e-06, 3.54193e-06,
  1.347033e-05, 2.0151e-05, 8.539193e-06, 8.355951e-06, 1.432469e-05, 
    1.384067e-05, 1.11481e-05, 1.299705e-05, 1.2823e-05, 8.702502e-06, 
    9.542977e-06, 2.648022e-06, 1.726682e-06, 1.209705e-06, 1.611863e-06,
  1.532346e-05, 1.138435e-05, 1.232356e-05, 7.355154e-06, 9.438128e-06, 
    1.040981e-05, 1.426339e-05, 1.280474e-05, 2.361302e-05, 2.869684e-05, 
    4.698555e-06, 6.800948e-06, 4.209091e-06, 2.207501e-06, 2.229921e-06,
  2.099372e-05, 1.417081e-05, 7.04341e-06, 8.422967e-06, 7.760439e-06, 
    7.748574e-06, 1.168717e-05, 1.578807e-05, 1.420368e-05, 2.114527e-05, 
    1.160593e-05, 1.136796e-05, 3.931579e-06, 3.385106e-06, 4.196645e-06,
  3.958919e-05, 2.755242e-05, 1.328989e-05, 7.147687e-06, 8.498236e-06, 
    6.481941e-06, 9.701476e-06, 1.428146e-05, 1.755035e-05, 2.092305e-05, 
    2.651669e-05, 1.244422e-05, 1.023066e-05, 5.454449e-06, 2.893167e-06,
  5.251264e-05, 4.393631e-05, 3.358985e-05, 1.426403e-05, 8.241571e-06, 
    7.649867e-06, 6.749403e-06, 9.250525e-06, 1.690771e-05, 1.847042e-05, 
    2.495507e-05, 3.555007e-05, 2.612147e-05, 3.019079e-05, 1.521466e-05,
  0.0001243473, 9.543275e-05, 6.40217e-05, 6.216601e-05, 3.558188e-05, 
    4.967156e-05, 6.183756e-05, 7.514517e-05, 9.379534e-05, 0.0001005586, 
    9.720169e-05, 0.0001103927, 0.0001114969, 0.00010846, 0.0001188194,
  0.000209258, 0.0001978646, 0.0001664, 0.0001386634, 0.0001263745, 
    0.000118421, 0.0001166595, 0.0001299955, 0.0001195555, 0.0001052309, 
    7.663662e-05, 5.802595e-05, 5.044041e-05, 6.496925e-05, 8.331338e-05,
  0.0003165553, 0.0003273086, 0.0003350158, 0.0003317555, 0.0002823462, 
    0.0002129017, 0.000162058, 0.0001162707, 8.583158e-05, 6.221914e-05, 
    3.02599e-05, 1.537493e-05, 2.267845e-05, 3.924002e-05, 6.967713e-05,
  0.0003877175, 0.0003995951, 0.0004693849, 0.0004416555, 0.0003175515, 
    0.0002217881, 0.0001526948, 7.827505e-05, 5.655954e-05, 3.772476e-05, 
    1.884842e-05, 1.429557e-05, 1.833531e-05, 5.074536e-05, 7.236251e-05,
  0.0003401712, 0.0004057798, 0.00042815, 0.0004027254, 0.0003074079, 
    0.0001927435, 0.000101177, 6.101246e-05, 4.212643e-05, 3.051147e-05, 
    1.776625e-05, 2.215896e-05, 3.758251e-05, 5.791733e-05, 4.335747e-05,
  0.0002453577, 0.0002839639, 0.0003174684, 0.0002746508, 0.0002219532, 
    0.0001487982, 8.349738e-05, 5.557051e-05, 4.690511e-05, 4.131695e-05, 
    2.979793e-05, 2.546176e-05, 2.447138e-05, 1.971597e-05, 4.608674e-06,
  0.0001436311, 0.0001558331, 0.0001677762, 0.0001672022, 0.0001451684, 
    0.000148005, 9.378131e-05, 4.597781e-05, 4.469301e-05, 3.148423e-05, 
    1.578046e-05, 3.942178e-06, 3.826235e-06, 1.429987e-06, 1.183247e-07,
  9.927939e-05, 8.520929e-05, 6.046115e-05, 9.34547e-05, 0.0001480222, 
    9.903718e-05, 8.487461e-05, 9.88587e-05, 1.418264e-05, 8.097127e-06, 
    1.938887e-06, 9.593576e-08, 6.569388e-08, 1.923846e-08, 5.400506e-08,
  8.931409e-05, 9.545085e-05, 6.814074e-05, 7.218985e-05, 8.126489e-05, 
    5.82279e-05, 4.6747e-05, 8.174587e-05, 7.417222e-06, 2.032902e-07, 
    7.093328e-06, 7.802393e-06, 1.133844e-05, 8.236238e-06, 8.85457e-08,
  9.57747e-05, 7.881346e-05, 7.126619e-05, 7.307583e-05, 6.609364e-05, 
    4.18893e-05, 4.320336e-05, 2.256345e-05, 1.394597e-05, 1.721938e-06, 
    6.479645e-06, 3.905932e-06, 2.826451e-08, 1.309423e-08, 3.816852e-06,
  2.853481e-06, 1.928149e-06, 1.151994e-06, 1.06741e-06, 9.565198e-07, 
    7.783239e-07, 1.838488e-06, 7.440287e-06, 2.515335e-05, 2.252503e-05, 
    5.271224e-06, 5.130114e-06, 4.771409e-06, 7.399789e-06, 2.602419e-06,
  5.823397e-06, 6.000228e-06, 2.7075e-06, 2.849842e-06, 3.547123e-06, 
    3.983089e-06, 7.588409e-06, 1.907581e-05, 5.603591e-05, 6.436338e-05, 
    1.977947e-05, 1.600275e-05, 6.760681e-06, 4.585822e-07, 3.550058e-07,
  1.190607e-05, 1.250139e-05, 1.480493e-05, 1.711966e-05, 2.62701e-05, 
    3.186138e-05, 6.976614e-05, 0.0001183667, 0.0002038343, 0.0002917146, 
    0.0001983197, 5.999255e-05, 4.437658e-06, 3.525047e-07, 7.479306e-07,
  1.297433e-05, 1.727906e-05, 2.669919e-05, 4.947614e-05, 8.290088e-05, 
    0.0001298297, 0.000213896, 0.000317176, 0.0005225295, 0.0008220266, 
    0.0009363128, 0.0007480115, 0.0003763893, 5.918662e-05, 2.189799e-05,
  1.567121e-05, 1.761192e-05, 2.676783e-05, 5.251317e-05, 7.341146e-05, 
    0.0001068966, 0.0001386162, 0.0001723202, 0.0003436873, 0.000620447, 
    0.0006254644, 0.0003525675, 0.0002051692, 9.561483e-05, 0.000113829,
  1.493075e-05, 1.860123e-05, 1.989399e-05, 1.702061e-05, 2.296731e-05, 
    3.183845e-05, 1.454163e-05, 2.161636e-05, 5.966633e-05, 7.0749e-05, 
    4.282353e-05, 2.880343e-05, 2.610613e-05, 5.243632e-05, 0.0001046152,
  1.818571e-05, 1.420779e-05, 1.461073e-05, 5.030655e-05, 5.113631e-05, 
    4.697115e-05, 6.545788e-05, 2.423566e-05, 2.214724e-05, 9.446989e-06, 
    2.375014e-05, 1.689565e-05, 2.325325e-05, 2.007562e-05, 2.491213e-05,
  2.46082e-05, 1.480511e-05, 1.579784e-05, 1.30172e-05, 5.322135e-05, 
    4.279557e-05, 6.986412e-05, 5.327563e-05, 2.136746e-05, 2.762528e-05, 
    3.086066e-05, 2.875124e-05, 1.270809e-05, 1.279653e-05, 1.527833e-05,
  2.004876e-05, 1.731834e-05, 9.20797e-06, 4.235366e-06, 2.493497e-05, 
    2.365251e-05, 5.82104e-05, 4.303588e-05, 4.67631e-05, 9.469187e-05, 
    6.404895e-05, 5.392346e-05, 1.884397e-05, 5.638914e-06, 3.942806e-05,
  1.579172e-05, 2.021222e-05, 5.663755e-06, 7.656411e-07, 2.910962e-05, 
    4.445883e-05, 2.333939e-05, 5.044859e-05, 0.0001237152, 0.0001237563, 
    0.0001286606, 7.050238e-05, 5.527287e-05, 1.862681e-05, 1.533812e-05,
  1.575171e-05, 1.667818e-05, 1.282156e-05, 1.135109e-05, 7.518226e-06, 
    4.399122e-06, 7.20085e-06, 2.69767e-05, 0.0001114763, 0.0001858298, 
    0.0001077895, 3.08137e-05, 3.272049e-05, 4.788338e-05, 5.585541e-05,
  9.521708e-06, 1.553387e-05, 1.4252e-05, 1.255896e-05, 1.12928e-05, 
    7.353899e-06, 7.306594e-06, 1.892386e-05, 9.26689e-05, 0.0001179978, 
    3.392306e-05, 2.579477e-05, 3.313426e-05, 4.749003e-05, 3.898676e-05,
  8.638573e-06, 7.017216e-06, 6.470422e-06, 8.713733e-06, 9.360716e-06, 
    7.543759e-06, 6.796386e-06, 1.824424e-05, 5.602374e-05, 4.924712e-05, 
    2.041112e-05, 2.663081e-05, 2.824781e-05, 2.824128e-05, 1.571069e-05,
  5.867203e-06, 5.088057e-06, 9.159259e-06, 1.052789e-05, 9.859918e-06, 
    6.768584e-06, 9.282897e-06, 1.305159e-05, 1.486803e-05, 1.031734e-05, 
    1.542805e-05, 2.522077e-05, 1.627909e-05, 9.293565e-06, 7.103191e-06,
  2.813749e-06, 5.606627e-06, 8.923863e-06, 7.492527e-06, 7.39906e-06, 
    9.943924e-06, 9.928731e-06, 9.077628e-06, 6.072236e-06, 7.655862e-06, 
    1.178479e-05, 1.937442e-05, 2.143431e-05, 1.114195e-05, 5.967924e-06,
  2.842532e-06, 5.890319e-06, 5.847802e-06, 9.020008e-06, 1.177742e-05, 
    1.663221e-05, 6.080606e-06, 1.879864e-05, 9.447266e-06, 8.962784e-06, 
    5.422207e-06, 1.047879e-05, 1.891387e-05, 1.363489e-05, 7.631094e-06,
  3.688052e-06, 8.264418e-06, 8.946832e-06, 9.475092e-06, 1.45068e-05, 
    2.248526e-05, 3.818972e-05, 3.172688e-05, 2.308774e-05, 2.79208e-05, 
    1.43118e-05, 1.237187e-05, 1.388165e-05, 1.201344e-05, 2.202809e-05,
  3.584424e-06, 5.456965e-06, 7.013729e-06, 8.255803e-06, 1.977183e-05, 
    1.667972e-05, 2.680368e-05, 3.58975e-05, 2.551693e-05, 3.52765e-05, 
    2.747312e-05, 6.283725e-06, 7.087475e-06, 8.905024e-06, 8.516351e-06,
  4.234576e-06, 4.968654e-06, 6.476573e-06, 7.807413e-06, 2.031038e-05, 
    2.361641e-06, 9.619345e-06, 2.669788e-05, 3.427296e-05, 3.773398e-05, 
    2.544171e-05, 1.967156e-05, 1.498303e-05, 6.988245e-06, 5.90055e-06,
  4.116394e-06, 2.871177e-06, 3.184105e-06, 3.004116e-05, 3.673511e-05, 
    1.468655e-05, 2.181909e-05, 2.896032e-05, 4.136302e-05, 2.977741e-05, 
    3.78035e-05, 1.011506e-05, 3.372736e-06, 2.63649e-06, 1.950256e-06,
  2.059377e-06, 1.864687e-06, 2.430435e-06, 2.716812e-06, 3.19327e-06, 
    3.487023e-06, 3.58824e-06, 3.499961e-06, 2.624733e-06, 1.566925e-06, 
    1.200381e-06, 5.319451e-07, 7.318752e-07, 6.867966e-07, 2.191711e-06,
  1.53304e-06, 3.625658e-07, 3.180661e-07, 4.002251e-07, 7.680908e-07, 
    1.42082e-06, 1.469916e-06, 8.848545e-07, 1.257526e-06, 3.497998e-07, 
    7.60534e-07, 1.172583e-06, 7.027148e-07, 2.247984e-06, 7.360146e-06,
  2.151571e-07, 7.610628e-08, 7.048715e-08, 1.322841e-07, 1.822774e-07, 
    2.24504e-08, 5.419026e-07, 9.783881e-07, 4.549343e-07, 1.396362e-06, 
    1.096539e-06, 2.173114e-06, 7.323729e-06, 9.260558e-06, 8.036314e-06,
  1.404735e-07, 2.657536e-07, 3.56812e-07, 7.296757e-07, 1.749205e-06, 
    1.993872e-06, 2.009179e-06, 9.975089e-07, 2.121211e-06, 9.209859e-07, 
    1.158203e-06, 8.536121e-06, 1.213709e-05, 1.374055e-05, 1.004251e-05,
  1.354902e-06, 9.852268e-07, 9.514719e-07, 2.595902e-06, 2.313305e-06, 
    4.474817e-06, 4.360994e-06, 2.755071e-06, 2.504102e-06, 4.028409e-06, 
    6.990042e-06, 5.639361e-06, 9.331457e-06, 1.183858e-05, 7.400222e-06,
  2.324522e-06, 2.944793e-06, 2.465399e-06, 2.742529e-06, 2.827109e-06, 
    3.490822e-06, 4.335067e-06, 3.74661e-06, 3.36518e-06, 2.232996e-06, 
    5.555013e-06, 1.211192e-05, 1.472586e-05, 1.318173e-05, 1.490038e-05,
  3.720145e-06, 3.593598e-06, 2.320261e-06, 3.86034e-06, 3.970821e-06, 
    3.309995e-06, 5.600072e-06, 6.501549e-06, 4.749385e-06, 1.082537e-05, 
    8.914546e-06, 2.027807e-05, 1.691951e-05, 1.789133e-05, 1.728268e-05,
  2.518628e-06, 2.726591e-06, 5.429191e-06, 3.979879e-06, 5.069288e-06, 
    6.63965e-06, 5.614749e-06, 6.734433e-06, 9.912868e-06, 1.906404e-05, 
    2.302296e-05, 1.704699e-05, 1.524425e-05, 1.172724e-05, 2.034181e-05,
  2.108422e-06, 2.462014e-06, 5.70758e-06, 6.844914e-06, 7.700363e-06, 
    8.637399e-06, 1.12643e-05, 1.070667e-05, 1.489433e-05, 2.990774e-05, 
    2.787693e-05, 1.725671e-05, 1.32519e-05, 1.426418e-05, 1.400309e-05,
  2.965139e-06, 4.285485e-06, 7.199109e-06, 1.317068e-05, 1.423831e-05, 
    7.878512e-06, 1.372689e-05, 1.84984e-05, 2.742029e-05, 1.971007e-05, 
    2.061307e-05, 2.266992e-05, 1.433733e-05, 1.29473e-05, 1.68438e-05,
  1.134641e-06, 1.102003e-06, 2.190507e-06, 2.478974e-06, 2.703674e-06, 
    5.678582e-06, 9.830968e-06, 1.345213e-05, 1.30196e-05, 8.137374e-06, 
    3.809344e-06, 3.531291e-06, 2.837915e-06, 4.217831e-07, 1.92367e-06,
  2.447286e-07, 7.584308e-07, 5.546547e-07, 7.633671e-07, 1.601261e-06, 
    2.299848e-06, 3.536491e-06, 4.448776e-06, 2.836273e-06, 1.256639e-06, 
    1.571784e-08, 4.096256e-07, 3.467484e-07, 3.818695e-07, 8.407925e-07,
  1.326358e-06, 4.14604e-07, 7.272756e-07, 1.730695e-07, 7.855978e-08, 
    6.114193e-07, 1.168965e-06, 1.147927e-06, 1.067856e-08, 1.249837e-07, 
    4.54114e-07, 3.041932e-08, 1.5437e-07, 2.759574e-06, 1.129326e-05,
  8.954345e-07, 8.619389e-07, 2.834244e-08, 4.275523e-08, 1.322463e-07, 
    1.76007e-08, 4.105464e-07, 4.341309e-08, 1.533135e-07, 3.708172e-07, 
    9.412683e-07, 4.271175e-06, 1.556448e-05, 1.900855e-05, 3.076283e-05,
  2.200603e-06, 4.996159e-07, 4.055119e-07, 6.434138e-07, 3.654309e-08, 
    8.578668e-08, 1.17947e-07, 1.740419e-07, 7.74257e-07, 2.522188e-06, 
    6.769842e-06, 1.73103e-05, 2.357789e-05, 2.211185e-05, 3.089256e-05,
  1.082835e-06, 1.438345e-06, 5.898322e-07, 6.327045e-07, 8.475435e-07, 
    6.354939e-07, 2.861476e-07, 1.502467e-06, 6.063848e-07, 3.26672e-06, 
    1.258464e-05, 2.455636e-05, 3.019372e-05, 2.333936e-05, 2.201066e-05,
  2.880915e-06, 9.951927e-07, 1.318654e-06, 9.001952e-07, 6.370901e-07, 
    1.928512e-07, 7.21593e-07, 1.377148e-06, 2.211023e-06, 3.264413e-06, 
    1.484139e-05, 3.01085e-05, 2.589162e-05, 2.670029e-05, 2.850818e-05,
  4.142839e-06, 3.090016e-06, 3.081464e-06, 2.704594e-06, 8.394774e-07, 
    8.178144e-07, 2.119761e-06, 2.099017e-06, 3.899429e-06, 3.815077e-06, 
    1.041117e-05, 1.832975e-05, 2.15065e-05, 4.023321e-05, 3.068606e-05,
  5.817046e-06, 5.469352e-06, 3.868143e-06, 4.235509e-06, 4.458721e-06, 
    3.835744e-06, 4.910743e-06, 5.961148e-06, 6.368439e-06, 1.032474e-05, 
    1.014292e-05, 1.27983e-05, 2.004541e-05, 2.978049e-05, 3.655215e-05,
  7.298193e-06, 8.118331e-06, 6.374895e-06, 5.811081e-06, 6.162535e-06, 
    6.073885e-06, 8.440844e-06, 9.853052e-06, 1.080679e-05, 1.054006e-05, 
    9.51474e-06, 1.32173e-05, 2.957587e-05, 1.885415e-05, 2.500447e-05,
  5.548873e-06, 5.73845e-06, 6.458576e-06, 6.149727e-06, 4.93673e-06, 
    5.150008e-06, 3.793205e-06, 6.325801e-06, 7.928155e-06, 1.180318e-05, 
    1.080581e-05, 1.152677e-05, 8.139848e-06, 8.52471e-06, 9.315871e-06,
  1.598699e-06, 4.885116e-06, 5.419593e-06, 4.588045e-06, 5.667439e-06, 
    4.347645e-06, 4.025426e-06, 3.844052e-06, 6.01694e-06, 5.788327e-06, 
    7.641753e-06, 6.984309e-06, 4.714158e-06, 4.323709e-06, 3.932093e-06,
  1.719108e-06, 1.783021e-06, 1.288541e-06, 3.409178e-06, 4.905648e-06, 
    4.821921e-06, 4.476277e-06, 3.766361e-06, 4.246802e-06, 4.463446e-06, 
    2.83999e-06, 3.513664e-06, 2.64889e-06, 5.660121e-06, 2.724302e-05,
  6.012424e-07, 2.789372e-06, 5.191004e-07, 2.076007e-06, 1.906311e-06, 
    1.328462e-06, 2.843897e-06, 2.968893e-06, 2.3278e-06, 2.146834e-06, 
    2.20693e-06, 3.583024e-06, 4.545494e-06, 1.236284e-05, 4.742062e-05,
  2.721364e-07, 5.493436e-07, 3.380001e-07, 7.495498e-07, 6.156725e-07, 
    7.292093e-07, 4.553475e-07, 2.084647e-06, 2.454647e-06, 3.1542e-06, 
    3.773635e-06, 5.460362e-06, 6.932178e-06, 9.113135e-06, 1.913086e-05,
  5.943105e-07, 3.429612e-07, 1.183281e-06, 6.886815e-08, 1.676995e-07, 
    3.666188e-07, 2.86893e-07, 1.864814e-06, 1.687119e-06, 3.728839e-06, 
    9.557062e-06, 1.111357e-05, 7.135328e-06, 4.440573e-06, 4.934116e-06,
  5.443302e-07, 1.110275e-07, 6.459719e-07, 1.175998e-06, 2.12749e-06, 
    1.565184e-06, 9.840543e-07, 8.526459e-07, 3.132233e-06, 8.497383e-06, 
    1.034076e-05, 1.192034e-05, 5.737467e-06, 7.784466e-06, 8.755361e-06,
  4.236774e-07, 6.214903e-08, 5.088938e-07, 1.339753e-06, 1.169089e-06, 
    9.859486e-07, 1.023414e-06, 2.293809e-06, 4.057544e-06, 5.809469e-06, 
    1.158728e-05, 1.327588e-05, 1.72424e-05, 2.526666e-05, 2.714122e-05,
  6.068556e-07, 2.950007e-07, 1.758088e-07, 1.437202e-07, 1.780239e-07, 
    5.504624e-07, 1.150467e-06, 2.320285e-06, 4.537138e-06, 7.344612e-06, 
    9.216816e-06, 1.016633e-05, 2.05234e-05, 4.513134e-05, 9.824186e-05,
  6.265918e-07, 1.222493e-06, 1.037553e-06, 3.962722e-07, 1.070747e-06, 
    1.515785e-06, 2.82013e-06, 5.012278e-06, 8.036743e-06, 7.62794e-06, 
    9.710438e-06, 2.211605e-05, 6.96569e-05, 0.0001406407, 9.69686e-05,
  8.292755e-05, 0.0002480442, 0.0003997856, 0.0003923131, 0.0003686263, 
    0.000300457, 0.0002362459, 0.0002282047, 0.000186916, 0.0001275684, 
    6.004698e-05, 2.783627e-05, 1.892912e-05, 1.734424e-05, 2.080958e-05,
  8.978693e-06, 5.243507e-05, 0.0001454762, 0.000213785, 0.0001980761, 
    0.0001600237, 0.0001452349, 0.0001522417, 0.0001625882, 0.0001318402, 
    7.931185e-05, 4.102477e-05, 2.140541e-05, 1.635969e-05, 1.595604e-05,
  4.146613e-06, 6.915279e-06, 7.060267e-06, 5.494332e-05, 0.0001158182, 
    0.0001345474, 0.0001200304, 0.0001119875, 0.0001099561, 8.471129e-05, 
    4.865783e-05, 2.425405e-05, 1.531031e-05, 1.114145e-05, 1.161927e-05,
  1.34605e-06, 2.770367e-06, 5.430068e-06, 5.838558e-06, 6.466063e-06, 
    3.111042e-05, 7.169792e-05, 9.077469e-05, 7.977364e-05, 5.779621e-05, 
    2.449611e-05, 1.139694e-05, 9.203944e-06, 8.240385e-06, 6.994958e-06,
  3.989608e-07, 1.326739e-06, 2.990918e-06, 4.416105e-06, 4.903626e-06, 
    4.770935e-06, 7.688051e-06, 1.149619e-05, 1.844363e-05, 2.330383e-05, 
    1.969917e-05, 1.855398e-05, 1.54093e-05, 1.224407e-05, 9.185994e-06,
  4.008294e-07, 4.894505e-07, 1.617834e-06, 1.666752e-06, 2.711548e-06, 
    3.847086e-06, 4.100283e-06, 6.353073e-06, 1.148527e-05, 1.444794e-05, 
    1.665349e-05, 2.455736e-05, 2.448117e-05, 2.281924e-05, 1.813589e-05,
  3.081569e-07, 1.754567e-07, 1.071752e-06, 3.395007e-06, 4.325887e-06, 
    6.046502e-06, 5.228355e-06, 5.673246e-06, 8.777984e-06, 9.659057e-06, 
    2.968819e-05, 3.427818e-05, 5.725801e-05, 5.137728e-05, 4.648926e-05,
  4.188746e-07, 3.612561e-07, 2.371609e-07, 1.665389e-06, 2.885721e-06, 
    2.686232e-06, 4.205129e-06, 3.88734e-06, 5.621529e-06, 1.645396e-05, 
    1.936525e-05, 4.759856e-06, 1.475623e-05, 2.573952e-05, 4.236163e-05,
  1.174266e-08, 4.498022e-08, 5.281891e-07, 1.757738e-06, 2.288956e-06, 
    1.588883e-06, 2.821852e-06, 3.273403e-06, 6.523544e-06, 1.86576e-05, 
    2.963231e-05, 1.634967e-05, 4.763571e-05, 8.155569e-05, 0.0001167018,
  3.92408e-07, 4.275228e-07, 7.326188e-07, 1.059156e-06, 1.169073e-06, 
    1.544496e-06, 2.154518e-06, 2.197023e-06, 4.002498e-06, 1.481251e-05, 
    2.227843e-05, 5.065705e-05, 0.0001015469, 0.0001151921, 0.0001529434,
  4.468975e-06, 6.465677e-06, 1.392336e-05, 3.058264e-05, 3.225932e-05, 
    1.754558e-05, 9.771762e-06, 7.630045e-06, 1.16212e-05, 1.433729e-05, 
    2.809553e-05, 4.064842e-05, 4.309114e-05, 3.184687e-05, 1.822605e-05,
  6.34914e-06, 8.178185e-06, 2.109245e-05, 4.471541e-05, 7.879052e-05, 
    8.152066e-05, 5.545357e-05, 4.405997e-05, 2.791331e-05, 2.255628e-05, 
    3.27806e-05, 3.723763e-05, 3.55641e-05, 3.788603e-05, 4.733571e-05,
  6.425951e-06, 3.183438e-05, 2.170082e-05, 2.811523e-05, 5.617531e-05, 
    0.0001046326, 0.0001114938, 9.872381e-05, 9.489145e-05, 9.728815e-05, 
    0.0001023005, 9.146191e-05, 8.714781e-05, 7.587152e-05, 0.0001138978,
  2.675884e-05, 5.512992e-05, 2.699177e-05, 9.56646e-07, 2.313848e-06, 
    3.303818e-05, 0.0001237943, 0.0001564453, 0.0001417038, 0.0001619143, 
    0.0002112603, 0.0002542092, 0.0002468997, 0.0002383143, 0.0002225871,
  2.918503e-05, 2.670196e-05, 1.887531e-05, 1.050458e-05, 1.098726e-06, 
    1.275873e-05, 8.996734e-05, 5.332572e-05, 7.828686e-05, 8.816799e-05, 
    0.0001129799, 0.0001386812, 0.00017088, 0.0001922768, 0.0002047164,
  3.343145e-06, 7.379817e-06, 5.950013e-06, 4.295041e-06, 2.85119e-06, 
    6.935329e-06, 1.219562e-05, 2.668908e-05, 1.977398e-05, 4.906468e-05, 
    6.067578e-05, 4.356011e-05, 6.530798e-05, 3.338558e-05, 6.940692e-05,
  2.481987e-05, 1.298243e-06, 5.721055e-07, 6.718247e-07, 3.017584e-06, 
    2.281967e-06, 4.917308e-06, 4.933317e-06, 5.678045e-06, 5.17836e-05, 
    5.583745e-05, 2.380629e-05, 1.602729e-05, 2.753041e-05, 2.124812e-06,
  2.769198e-05, 1.642964e-05, 7.969246e-06, 3.276171e-06, 5.331301e-06, 
    4.516283e-06, 1.050439e-05, 1.185497e-05, 2.564125e-05, 4.664112e-05, 
    4.88912e-05, 3.580083e-05, 6.462596e-06, 7.191225e-06, 9.830113e-06,
  4.411665e-06, 3.44425e-06, 3.672639e-06, 4.384918e-06, 2.606571e-06, 
    5.700153e-06, 6.481481e-06, 8.552217e-06, 1.893526e-05, 6.263327e-05, 
    6.814823e-05, 4.222144e-05, 7.5603e-05, 6.640705e-05, 6.877381e-05,
  5.33234e-06, 2.077181e-06, 2.223981e-06, 2.148682e-06, 2.016049e-06, 
    2.200293e-06, 2.367762e-06, 3.194444e-05, 3.060342e-05, 4.976626e-05, 
    4.577396e-05, 5.483953e-05, 6.45841e-05, 4.726817e-05, 3.426545e-05,
  2.882877e-06, 2.963998e-06, 2.998888e-06, 2.995326e-06, 3.868511e-06, 
    2.790518e-06, 2.357749e-06, 2.822501e-06, 2.189325e-06, 1.861477e-06, 
    1.031706e-06, 1.433852e-06, 4.59041e-07, 8.32286e-07, 2.855562e-06,
  7.224959e-06, 7.212272e-06, 6.396511e-06, 5.946554e-06, 4.781508e-06, 
    3.516432e-06, 3.350404e-06, 3.173015e-06, 2.901245e-06, 1.590753e-06, 
    7.802569e-07, 3.721408e-07, 8.696479e-07, 8.929619e-07, 3.252056e-06,
  7.044076e-06, 7.742013e-06, 9.579248e-06, 6.063794e-06, 5.846262e-06, 
    3.876342e-06, 2.559828e-06, 3.213439e-06, 3.682346e-06, 2.620167e-06, 
    1.164643e-06, 8.153451e-07, 7.965886e-07, 3.436324e-07, 2.85752e-06,
  2.634235e-06, 3.741603e-06, 2.095589e-06, 1.445672e-06, 1.12094e-06, 
    1.681193e-06, 1.911375e-06, 2.394883e-06, 2.729414e-06, 1.770216e-06, 
    7.930698e-07, 8.165637e-08, 7.570815e-07, 6.264015e-07, 1.707788e-06,
  3.246767e-06, 2.219601e-06, 9.106076e-07, 5.701102e-07, 5.78534e-07, 
    4.153279e-07, 4.696306e-07, 4.559404e-07, 2.003632e-07, 3.301596e-07, 
    2.956444e-07, 3.418082e-07, 8.706549e-07, 8.989222e-07, 1.982451e-06,
  2.833011e-06, 1.147652e-06, 4.319246e-07, 6.318944e-07, 7.389417e-07, 
    1.09191e-06, 9.766933e-07, 6.72953e-07, 1.236022e-07, 8.288844e-08, 
    7.309974e-08, 9.123254e-07, 1.521814e-06, 7.362985e-06, 2.820922e-06,
  4.270323e-07, 2.836049e-07, 1.157449e-08, 4.449375e-08, 3.17766e-07, 
    4.370793e-07, 6.268895e-07, 5.39733e-07, 3.742398e-07, 2.349003e-07, 
    9.502768e-07, 8.795048e-06, 1.321781e-05, 1.412279e-05, 2.135214e-05,
  6.147832e-07, 4.518589e-07, 2.705229e-06, 1.597155e-06, 1.053778e-06, 
    2.608838e-06, 1.026317e-06, 8.565081e-07, 1.073494e-06, 1.415023e-06, 
    9.64138e-06, 1.700703e-05, 1.844856e-05, 4.777277e-05, 1.733403e-05,
  1.933123e-06, 1.17207e-06, 8.88438e-07, 1.462072e-06, 1.064039e-06, 
    1.690994e-06, 3.800185e-06, 6.428505e-06, 1.723434e-05, 2.112752e-05, 
    1.88752e-05, 4.16045e-05, 5.700414e-05, 7.280372e-05, 0.0001014504,
  6.272766e-06, 4.433399e-06, 3.465731e-06, 1.656668e-06, 2.49152e-06, 
    2.428782e-06, 3.257735e-06, 3.292603e-06, 6.425704e-06, 2.199844e-05, 
    3.772305e-05, 6.30113e-05, 7.749636e-05, 6.808185e-05, 7.467295e-05,
  5.535883e-06, 4.009628e-06, 4.756906e-06, 4.921129e-06, 5.800899e-06, 
    5.304969e-06, 3.336326e-06, 4.18498e-06, 4.6884e-06, 5.228599e-06, 
    3.460887e-06, 1.468429e-06, 1.754553e-06, 9.56677e-07, 5.859427e-07,
  2.325369e-06, 3.484522e-06, 3.585194e-06, 4.285925e-06, 3.584574e-06, 
    2.797007e-06, 3.14144e-06, 2.811053e-06, 1.927358e-06, 1.734377e-06, 
    1.753403e-06, 4.749298e-07, 2.0793e-08, 1.063851e-08, 9.659837e-09,
  1.560406e-06, 7.179221e-07, 8.660124e-07, 1.391941e-06, 2.056511e-06, 
    1.836795e-06, 1.686133e-06, 2.185898e-06, 1.909354e-06, 1.261875e-06, 
    1.174352e-06, 1.358103e-06, 8.581756e-07, 8.615019e-07, 3.919166e-07,
  3.436987e-08, 2.125246e-08, 5.97417e-08, 1.948088e-07, 4.782344e-07, 
    2.473898e-06, 1.913033e-06, 1.630907e-06, 2.683e-06, 2.305098e-06, 
    3.079474e-06, 5.907882e-06, 8.005821e-06, 5.199807e-06, 3.713079e-06,
  1.631933e-09, 1.211569e-08, 3.946316e-08, 1.360491e-07, 6.274175e-07, 
    2.686013e-06, 1.755455e-06, 3.268717e-06, 4.536585e-06, 4.652048e-06, 
    4.616758e-06, 3.96578e-06, 8.415983e-06, 1.144649e-05, 9.708483e-06,
  1.603626e-08, 1.034622e-07, 1.085601e-07, 2.794944e-07, 1.043172e-06, 
    1.32569e-06, 3.366731e-06, 4.500581e-06, 5.027939e-06, 6.187502e-06, 
    6.487639e-06, 4.325889e-06, 5.638191e-06, 3.194198e-06, 4.405743e-06,
  2.295978e-07, 5.328851e-07, 3.097322e-07, 4.456502e-07, 1.308946e-06, 
    2.531322e-06, 3.89778e-06, 5.5354e-06, 5.970294e-06, 5.195628e-06, 
    5.20356e-06, 4.586323e-06, 2.257737e-06, 1.261456e-05, 8.728332e-06,
  6.29894e-08, 3.803701e-07, 4.365407e-07, 1.02417e-06, 5.962531e-07, 
    3.483229e-06, 4.151695e-06, 5.586975e-06, 7.024096e-06, 5.635668e-06, 
    7.827614e-06, 8.02069e-06, 1.389367e-05, 2.746919e-05, 3.130723e-05,
  9.893564e-08, 2.67492e-07, 9.844008e-07, 7.57872e-07, 1.476874e-06, 
    1.459969e-06, 2.047364e-06, 4.208492e-06, 7.461896e-06, 8.272321e-06, 
    2.727841e-05, 1.896286e-05, 3.444121e-05, 2.460873e-05, 3.228849e-05,
  2.737815e-07, 1.130623e-06, 7.865927e-07, 9.144023e-07, 1.525449e-06, 
    2.460052e-06, 3.110166e-06, 5.009921e-06, 9.256081e-06, 2.711839e-05, 
    3.273205e-05, 4.198033e-05, 3.315497e-05, 3.503516e-05, 4.047089e-05,
  2.299595e-05, 2.490396e-05, 1.515205e-05, 8.33e-06, 5.751887e-06, 
    2.12334e-06, 1.279295e-06, 2.784102e-06, 6.63463e-06, 1.699497e-05, 
    2.163862e-05, 2.790818e-05, 1.927255e-05, 8.100252e-06, 2.913613e-06,
  6.92368e-06, 1.61005e-05, 2.674412e-05, 1.31382e-05, 6.315114e-06, 
    6.021811e-07, 1.202466e-06, 4.577956e-06, 7.102666e-06, 8.463828e-06, 
    1.048451e-05, 6.985538e-06, 5.227941e-06, 3.190994e-06, 2.607245e-06,
  3.175846e-05, 2.226381e-05, 9.189303e-06, 4.095715e-06, 2.351903e-06, 
    1.902252e-06, 4.424275e-06, 7.255655e-06, 8.388224e-06, 7.560142e-06, 
    6.147531e-06, 6.664955e-06, 4.788927e-06, 6.04419e-06, 5.776236e-06,
  1.889449e-05, 1.987169e-06, 1.405896e-07, 5.094611e-07, 3.282846e-06, 
    2.220826e-06, 7.13218e-06, 6.163159e-06, 6.133323e-06, 4.923005e-06, 
    3.590592e-06, 5.570172e-06, 4.670717e-06, 5.292497e-06, 6.159364e-06,
  7.961054e-06, 4.252169e-07, 1.908425e-07, 1.270586e-06, 3.139818e-06, 
    2.200952e-06, 5.45081e-06, 5.132283e-06, 1.192481e-05, 4.635747e-06, 
    2.823315e-07, 1.791198e-06, 2.360325e-06, 2.22028e-06, 3.72194e-06,
  5.912147e-07, 3.529578e-07, 1.324043e-07, 2.103171e-06, 2.392917e-06, 
    2.52962e-06, 2.163935e-06, 9.509816e-06, 7.565409e-06, 7.732776e-06, 
    1.989415e-07, 1.367795e-07, 1.344481e-07, 2.127436e-07, 4.076395e-06,
  5.726343e-07, 4.722635e-07, 1.013137e-06, 1.531131e-06, 2.051012e-06, 
    2.513866e-06, 5.020913e-06, 1.153374e-05, 1.56475e-05, 1.20195e-05, 
    1.259323e-05, 1.705601e-05, 1.917405e-05, 1.318833e-05, 3.608835e-06,
  2.288258e-07, 3.759685e-07, 2.296864e-06, 3.55397e-06, 5.522535e-06, 
    4.402995e-06, 6.190707e-06, 1.263313e-05, 2.076683e-05, 3.04444e-05, 
    1.963981e-05, 2.365511e-05, 1.882535e-05, 6.088339e-06, 2.599934e-05,
  1.83853e-07, 4.341763e-07, 1.909088e-06, 3.352722e-06, 3.769914e-06, 
    4.698425e-06, 6.270265e-06, 1.938871e-05, 2.485262e-05, 2.239204e-05, 
    2.910804e-05, 1.710214e-05, 1.562939e-05, 2.110134e-05, 1.679231e-05,
  3.023977e-07, 1.715443e-06, 3.488163e-06, 3.453257e-06, 4.540534e-06, 
    5.026059e-06, 9.623012e-06, 2.106385e-05, 3.561874e-05, 2.484923e-05, 
    3.535375e-05, 2.772282e-05, 2.369097e-05, 2.393033e-05, 2.015836e-05,
  3.649561e-09, 1.195311e-07, 5.309734e-06, 2.68839e-05, 5.22933e-05, 
    6.757941e-05, 3.879375e-05, 1.552877e-05, 1.65159e-05, 1.091892e-05, 
    1.59253e-05, 2.252423e-05, 3.336406e-05, 3.624056e-05, 1.794218e-05,
  4.331067e-07, 4.034403e-06, 2.19398e-05, 2.852726e-05, 3.216053e-05, 
    2.003216e-05, 1.247408e-05, 1.660518e-05, 3.203053e-05, 1.166184e-05, 
    1.491171e-05, 1.249804e-05, 1.313088e-05, 6.679953e-06, 5.976231e-06,
  2.361828e-06, 1.969098e-05, 4.07111e-05, 3.214662e-05, 1.98143e-05, 
    9.854172e-06, 1.003848e-05, 1.987852e-05, 2.869791e-05, 1.989725e-05, 
    4.885799e-06, 2.527366e-06, 2.693434e-06, 3.128366e-06, 4.087806e-06,
  1.175617e-05, 3.475002e-05, 2.010349e-05, 1.538917e-05, 1.21595e-05, 
    6.912942e-06, 1.082167e-05, 1.863339e-05, 2.644379e-05, 1.865407e-05, 
    4.595814e-06, 2.11287e-07, 1.292997e-07, 2.532492e-06, 2.217023e-06,
  9.01196e-06, 9.465636e-06, 9.276339e-06, 8.909484e-06, 7.785566e-06, 
    1.298834e-05, 1.222088e-05, 2.559549e-05, 3.062791e-05, 3.522778e-05, 
    8.897352e-06, 5.505804e-06, 4.272012e-06, 3.632457e-06, 2.096783e-06,
  6.572435e-06, 6.271458e-06, 3.897045e-06, 5.461639e-06, 6.590623e-06, 
    8.196364e-06, 1.221944e-05, 1.675116e-05, 1.820276e-05, 1.255224e-05, 
    6.014189e-06, 1.049662e-05, 4.024445e-06, 5.483918e-06, 4.346966e-06,
  2.007927e-06, 8.792056e-07, 1.595211e-06, 1.687532e-06, 5.26815e-06, 
    1.211175e-05, 9.617902e-06, 9.606059e-06, 6.449252e-06, 4.729873e-06, 
    5.540548e-06, 2.455737e-06, 8.60711e-06, 6.710756e-06, 8.04907e-06,
  9.396946e-07, 1.759763e-06, 1.498373e-06, 3.205069e-06, 5.399659e-06, 
    6.205869e-06, 6.240526e-06, 3.665137e-06, 5.748736e-06, 5.861737e-06, 
    9.961709e-06, 4.235302e-06, 1.993853e-06, 4.45818e-06, 5.563557e-06,
  6.91257e-07, 1.683072e-06, 3.755954e-06, 5.325667e-06, 7.208233e-06, 
    3.751996e-06, 2.860893e-06, 2.812702e-06, 3.684403e-06, 1.955404e-06, 
    2.446267e-06, 3.783657e-06, 3.778134e-06, 4.381636e-06, 4.472784e-06,
  2.13282e-06, 4.05416e-06, 6.390685e-06, 4.443931e-06, 3.585675e-06, 
    2.592797e-06, 2.260665e-06, 2.363817e-06, 4.816657e-06, 3.360781e-06, 
    3.015181e-06, 4.931433e-06, 3.116119e-06, 3.191313e-06, 4.323259e-06,
  1.229173e-06, 1.087035e-06, 1.851681e-06, 8.545762e-07, 3.810089e-07, 
    1.193323e-06, 1.33689e-06, 2.102801e-06, 3.9185e-06, 1.676428e-05, 
    1.143762e-05, 1.65669e-05, 2.388591e-05, 2.87277e-05, 2.855371e-05,
  1.460697e-07, 9.135201e-07, 5.822027e-07, 1.706139e-06, 2.448823e-06, 
    1.963111e-06, 3.017336e-06, 5.959067e-06, 1.724467e-05, 1.847981e-05, 
    1.501489e-05, 1.338788e-05, 2.058526e-05, 1.860515e-05, 2.07639e-05,
  1.396208e-09, 6.836519e-09, 3.953209e-08, 6.410052e-08, 1.240616e-06, 
    3.112155e-06, 2.123112e-06, 3.126546e-06, 2.267297e-05, 4.286432e-05, 
    1.162507e-05, 1.603129e-05, 3.764281e-05, 1.141984e-05, 1.736676e-05,
  1.068421e-07, 6.99202e-08, 1.087216e-06, 1.710256e-06, 8.215232e-07, 
    2.427406e-06, 3.229491e-06, 1.145354e-05, 2.956329e-05, 1.958626e-05, 
    2.215301e-05, 4.056681e-05, 3.639096e-05, 3.252332e-05, 1.662229e-05,
  1.365146e-06, 1.139275e-06, 1.998086e-06, 2.000271e-06, 1.41948e-06, 
    2.387126e-06, 4.478393e-06, 2.216576e-05, 3.455409e-05, 2.644593e-05, 
    3.670042e-05, 5.475003e-05, 4.447668e-05, 2.850314e-05, 1.92967e-05,
  1.056119e-06, 1.556942e-06, 1.632031e-06, 1.877741e-06, 2.8278e-06, 
    4.914047e-06, 1.673722e-05, 2.595785e-05, 2.835061e-05, 5.915193e-05, 
    7.60016e-05, 6.346328e-05, 5.654318e-05, 3.119067e-05, 1.614628e-05,
  2.977079e-06, 3.761638e-06, 2.251794e-06, 2.274855e-06, 3.345151e-06, 
    1.298488e-05, 1.483961e-05, 2.587051e-05, 5.163705e-05, 5.649734e-05, 
    4.783608e-05, 1.493822e-05, 1.05803e-05, 6.486892e-06, 3.929264e-06,
  3.408555e-06, 3.589092e-06, 4.05533e-06, 3.155599e-06, 3.812921e-06, 
    3.762109e-06, 2.619626e-05, 2.735872e-05, 2.878136e-05, 1.69792e-05, 
    5.649772e-06, 1.688993e-06, 1.740322e-06, 1.334493e-06, 1.571479e-06,
  2.943867e-06, 3.573212e-06, 4.093861e-06, 3.287374e-06, 4.711233e-06, 
    7.883154e-06, 1.18571e-05, 2.015115e-05, 4.523507e-06, 1.981289e-06, 
    1.026197e-06, 1.775359e-06, 1.41909e-06, 1.463114e-06, 1.285604e-06,
  2.393767e-06, 2.52029e-06, 3.206794e-06, 3.176096e-06, 4.340334e-06, 
    4.798947e-06, 4.418874e-06, 2.932518e-06, 7.065099e-07, 7.0941e-07, 
    1.00539e-06, 1.061109e-06, 1.917142e-06, 1.688081e-06, 3.111704e-06,
  3.955189e-06, 4.571747e-06, 5.584393e-06, 1.144494e-05, 5.133496e-06, 
    3.570633e-06, 5.235511e-06, 9.768319e-06, 1.434157e-05, 1.060637e-05, 
    1.424263e-05, 3.379158e-06, 2.860621e-06, 8.53673e-07, 2.64726e-07,
  4.537842e-06, 6.7329e-06, 8.564536e-06, 8.014612e-06, 1.162215e-05, 
    1.494511e-05, 1.382782e-05, 1.368436e-05, 1.273961e-05, 1.288306e-05, 
    6.386158e-06, 4.23684e-07, 1.152729e-07, 6.886646e-08, 1.378028e-06,
  9.897423e-06, 8.798874e-06, 1.347169e-05, 1.701508e-05, 1.87668e-05, 
    2.317488e-05, 1.336746e-05, 1.415098e-05, 7.512501e-06, 4.484492e-06, 
    1.293528e-06, 3.721513e-09, 9.013274e-08, 1.589663e-06, 3.855907e-06,
  1.817143e-05, 1.761399e-05, 1.549181e-05, 2.068511e-05, 1.645383e-05, 
    1.283508e-05, 7.656809e-06, 2.628609e-06, 1.859719e-06, 7.136694e-07, 
    2.601555e-07, 8.560739e-08, 9.005607e-07, 1.042845e-05, 9.973519e-06,
  1.350047e-05, 1.950221e-05, 1.790816e-05, 1.483539e-05, 7.82187e-06, 
    1.568507e-06, 4.027873e-07, 5.036859e-07, 1.513192e-07, 8.219836e-09, 
    2.405787e-08, 3.709547e-06, 6.676393e-06, 8.065872e-06, 5.028963e-06,
  7.040039e-06, 4.703757e-06, 7.92232e-06, 7.16352e-06, 2.039956e-06, 
    1.19559e-06, 1.764651e-07, 5.774132e-09, 1.620101e-08, 3.140139e-07, 
    4.093901e-06, 8.067978e-06, 4.288473e-06, 2.451608e-06, 7.531554e-07,
  2.13213e-05, 4.003359e-06, 5.204413e-06, 4.949994e-06, 3.530463e-06, 
    1.198596e-06, 4.309058e-07, 6.922967e-07, 2.029559e-06, 4.553091e-06, 
    3.442969e-06, 2.598102e-06, 7.588719e-07, 1.732807e-07, 6.069258e-07,
  4.29846e-06, 3.204052e-06, 3.819385e-06, 4.267884e-06, 3.245801e-06, 
    2.084288e-06, 2.815925e-06, 1.36961e-06, 2.287909e-06, 2.381263e-06, 
    1.621486e-06, 4.331044e-07, 3.459994e-07, 3.555971e-08, 8.667263e-07,
  1.550333e-06, 2.674569e-06, 3.127658e-06, 3.504411e-06, 3.167453e-06, 
    2.19679e-06, 2.97597e-06, 1.938755e-06, 2.431073e-06, 4.786575e-06, 
    1.256404e-07, 1.572189e-07, 3.135223e-08, 4.593183e-07, 2.813766e-06,
  2.383188e-06, 3.165072e-06, 2.575609e-06, 2.927999e-06, 2.421782e-06, 
    2.408006e-06, 1.540004e-06, 1.819279e-06, 4.034986e-06, 1.964932e-06, 
    6.532231e-07, 3.33529e-07, 1.280371e-06, 2.65079e-06, 1.343212e-05,
  1.868257e-07, 1.100655e-07, 2.093117e-07, 1.458007e-07, 6.657758e-08, 
    3.452757e-08, 1.535136e-09, 3.250273e-09, 1.555395e-08, 2.574112e-07, 
    1.00226e-06, 1.379996e-06, 3.079294e-06, 7.786806e-06, 1.194441e-05,
  3.9158e-07, 8.984306e-08, 9.863546e-09, 5.668961e-10, 1.415552e-08, 
    4.422608e-08, 4.531742e-08, 3.370375e-08, 4.147765e-07, 5.310309e-07, 
    1.964104e-06, 6.650874e-06, 7.421542e-06, 1.100041e-05, 1.162942e-05,
  6.213175e-07, 7.466523e-07, 1.409289e-07, 4.651722e-08, 1.452744e-07, 
    1.048933e-07, 1.736801e-06, 1.318862e-06, 3.268251e-06, 3.916758e-06, 
    5.666668e-06, 5.803888e-06, 9.309045e-06, 5.653243e-06, 5.252022e-06,
  2.538419e-06, 1.475673e-06, 2.236524e-06, 3.015712e-06, 4.426422e-06, 
    4.881429e-06, 6.356851e-06, 8.763735e-06, 7.840872e-06, 6.684516e-06, 
    6.506593e-06, 8.357295e-06, 7.571427e-06, 7.855439e-06, 9.19784e-06,
  1.385788e-05, 1.712649e-05, 1.236993e-05, 1.089907e-05, 1.381834e-05, 
    8.67686e-06, 9.473603e-06, 1.463477e-05, 1.299161e-05, 1.173269e-05, 
    1.123042e-05, 1.191517e-05, 9.906133e-06, 6.547658e-06, 7.595914e-06,
  2.684216e-05, 2.953598e-05, 2.487376e-05, 2.327192e-05, 2.003638e-05, 
    1.630215e-05, 1.458562e-05, 1.639279e-05, 1.516889e-05, 1.101492e-05, 
    8.611553e-06, 7.475963e-06, 5.489615e-06, 6.513371e-06, 4.525377e-06,
  1.592986e-05, 1.952861e-05, 2.147795e-05, 2.123814e-05, 1.49777e-05, 
    1.329275e-05, 1.018842e-05, 1.10313e-05, 1.051565e-05, 8.933108e-06, 
    8.024654e-06, 4.611467e-06, 3.474775e-06, 5.441003e-06, 9.415123e-06,
  1.128988e-05, 1.3674e-05, 1.934181e-05, 1.435651e-05, 1.155608e-05, 
    8.515038e-06, 1.007487e-05, 8.005012e-06, 8.009972e-06, 6.138852e-06, 
    4.488817e-06, 4.013349e-06, 4.885596e-06, 1.042061e-05, 1.777557e-05,
  7.173921e-06, 1.057275e-05, 1.717097e-05, 1.228458e-05, 8.916423e-06, 
    6.676957e-06, 7.855927e-06, 7.579326e-06, 6.129296e-06, 5.048561e-06, 
    3.803569e-06, 4.302071e-06, 8.838745e-06, 1.484675e-05, 2.449442e-05,
  5.883079e-06, 9.695459e-06, 9.615403e-06, 1.073088e-05, 8.796038e-06, 
    6.582891e-06, 6.063046e-06, 5.43552e-06, 4.653222e-06, 3.730862e-06, 
    3.469682e-06, 8.217959e-06, 1.206301e-05, 1.828665e-05, 3.946284e-05,
  1.052885e-06, 5.958576e-07, 1.84098e-06, 2.475667e-06, 3.107519e-06, 
    3.681113e-06, 4.467698e-06, 7.360792e-06, 1.01059e-05, 1.157386e-05, 
    1.223443e-05, 1.29248e-05, 1.018847e-05, 1.003447e-05, 1.223278e-05,
  2.27617e-06, 3.608401e-07, 1.337549e-06, 4.248695e-06, 6.833502e-06, 
    7.311179e-06, 8.84811e-06, 1.3888e-05, 1.469423e-05, 1.384261e-05, 
    1.274481e-05, 1.292073e-05, 1.051479e-05, 1.317062e-05, 2.105953e-05,
  3.510017e-06, 7.278752e-06, 6.968728e-06, 7.332967e-06, 1.005171e-05, 
    9.65153e-06, 1.040884e-05, 1.137693e-05, 1.148951e-05, 1.048954e-05, 
    1.123185e-05, 2.148914e-05, 3.697873e-05, 5.711581e-05, 7.610422e-05,
  5.514042e-07, 1.485709e-06, 3.091306e-06, 7.430022e-06, 1.001447e-05, 
    1.674925e-05, 1.481381e-05, 1.578334e-05, 1.677408e-05, 1.436108e-05, 
    2.593557e-05, 4.128112e-05, 5.449302e-05, 6.739141e-05, 7.453281e-05,
  1.924924e-07, 3.581092e-06, 5.008021e-06, 4.140003e-06, 9.838048e-06, 
    1.191618e-05, 1.309891e-05, 1.011421e-05, 1.232368e-05, 1.895021e-05, 
    3.05367e-05, 4.187157e-05, 5.031534e-05, 6.137552e-05, 7.059343e-05,
  4.782208e-07, 2.036069e-06, 3.360479e-06, 5.779774e-06, 1.060923e-05, 
    1.251943e-05, 9.825866e-06, 8.539135e-06, 1.186822e-05, 1.658585e-05, 
    1.887258e-05, 2.609615e-05, 4.154194e-05, 5.954782e-05, 7.168557e-05,
  1.756991e-06, 2.237771e-06, 3.990026e-06, 6.170165e-06, 1.219482e-05, 
    1.354589e-05, 8.611399e-06, 1.068879e-05, 1.524162e-05, 1.505678e-05, 
    1.637578e-05, 2.492256e-05, 3.704002e-05, 4.410058e-05, 4.196279e-05,
  5.313067e-06, 2.220997e-06, 2.922568e-06, 6.735232e-06, 9.50271e-06, 
    1.317717e-05, 1.084456e-05, 1.466552e-05, 2.469263e-05, 2.493274e-05, 
    2.734976e-05, 3.090904e-05, 2.546967e-05, 2.43485e-05, 1.264525e-05,
  8.792748e-06, 4.11829e-06, 3.720917e-06, 5.285092e-06, 7.448163e-06, 
    1.521207e-05, 1.485564e-05, 1.900178e-05, 2.460823e-05, 3.93646e-05, 
    6.351872e-05, 6.906112e-05, 3.950515e-05, 1.251713e-05, 5.388149e-06,
  8.704028e-06, 1.097278e-05, 3.586783e-06, 3.829573e-06, 7.236929e-06, 
    1.04936e-05, 1.641898e-05, 1.583087e-05, 2.26478e-05, 3.875937e-05, 
    7.863879e-05, 0.0001257261, 0.0001531898, 9.509363e-05, 6.857664e-06,
  8.944747e-06, 4.757368e-06, 4.057656e-06, 5.018642e-06, 9.038888e-06, 
    1.259636e-05, 1.950011e-05, 1.815183e-05, 1.031096e-05, 1.471167e-05, 
    3.61635e-05, 7.866146e-05, 0.0001773236, 0.0003190755, 0.0004390563,
  7.524529e-06, 4.16339e-06, 5.581562e-06, 6.477594e-06, 9.418603e-06, 
    1.031156e-05, 8.597463e-06, 7.328023e-06, 1.094447e-05, 4.710147e-05, 
    0.000159068, 0.0002680773, 0.0004313058, 0.0005960062, 0.0007295539,
  4.044843e-06, 4.083378e-06, 6.043758e-06, 1.054611e-05, 9.987853e-06, 
    6.882306e-06, 7.250452e-06, 8.709107e-06, 3.826959e-05, 0.000254595, 
    0.0004267179, 0.0004450613, 0.0004949161, 0.0006186816, 0.000681219,
  3.28106e-06, 6.236698e-06, 8.047488e-06, 1.289002e-05, 1.067234e-05, 
    8.151046e-06, 9.817874e-06, 2.073369e-05, 0.0002128555, 0.0005094401, 
    0.0004538209, 0.0003203193, 0.0003588672, 0.0004323248, 0.0004206507,
  4.041962e-06, 6.238824e-06, 1.073528e-05, 2.246556e-05, 1.605589e-05, 
    8.995184e-06, 8.647719e-06, 3.732651e-05, 0.000295572, 0.000373459, 
    0.0002776204, 0.000260889, 0.0001934781, 0.0001893462, 0.0001814498,
  5.184795e-06, 7.458047e-06, 2.152719e-05, 3.11993e-05, 1.861216e-05, 
    1.112424e-05, 1.13954e-05, 4.089795e-05, 0.0001238906, 0.0001667244, 
    0.000237915, 0.0001923103, 7.436997e-05, 9.482834e-05, 0.0001307422,
  1.06555e-05, 1.503823e-05, 2.50718e-05, 3.053771e-05, 2.357036e-05, 
    1.629583e-05, 1.813447e-05, 3.114398e-05, 3.272217e-05, 8.190193e-05, 
    0.0001602662, 0.0001442793, 2.920688e-05, 6.481271e-05, 8.841007e-05,
  1.141713e-05, 1.713619e-05, 2.644527e-05, 2.958135e-05, 2.198511e-05, 
    1.834851e-05, 2.353363e-05, 3.133152e-05, 1.599879e-05, 3.288694e-05, 
    8.107639e-05, 0.000121973, 7.427747e-05, 3.275153e-05, 7.327135e-05,
  1.233377e-05, 1.937521e-05, 2.739453e-05, 2.372875e-05, 1.967605e-05, 
    1.950171e-05, 2.839841e-05, 2.91319e-05, 2.560389e-05, 2.536285e-05, 
    5.542659e-05, 0.0001049986, 0.0001207097, 2.44656e-05, 4.553868e-05,
  1.427444e-05, 1.736524e-05, 2.408254e-05, 2.213438e-05, 1.890529e-05, 
    2.318415e-05, 3.82478e-05, 4.017452e-05, 2.92757e-05, 4.120759e-05, 
    3.256326e-05, 0.0001129501, 0.0001522576, 7.314964e-06, 2.371138e-05,
  1.600752e-06, 1.626167e-06, 5.299262e-07, 2.225331e-07, 1.890064e-07, 
    7.128224e-08, 6.301777e-08, 6.834261e-08, 6.952268e-08, 1.377595e-07, 
    1.232725e-07, 8.748401e-08, 7.401673e-08, 2.053163e-08, 1.047433e-07,
  1.882656e-06, 6.553083e-07, 3.661278e-07, 1.650622e-07, 8.237019e-08, 
    3.475878e-08, 7.394888e-08, 5.77013e-07, 1.766199e-07, 1.230392e-08, 
    8.503358e-08, 6.43923e-07, 8.469036e-07, 4.43321e-07, 3.181509e-06,
  5.830884e-07, 5.468211e-07, 1.841982e-07, 8.243367e-08, 2.638979e-07, 
    6.104349e-07, 4.690411e-07, 4.368625e-07, 2.886818e-08, 8.564935e-07, 
    1.775913e-06, 4.197227e-06, 1.035599e-05, 2.037417e-05, 7.991629e-05,
  2.005167e-06, 1.279595e-06, 3.932058e-07, 2.980671e-07, 3.140755e-07, 
    8.348993e-07, 4.38974e-07, 4.177523e-07, 6.283387e-07, 1.479001e-06, 
    5.004273e-06, 3.942714e-05, 0.0002271645, 0.0005220466, 0.0006443706,
  3.131936e-06, 2.094628e-06, 5.5676e-07, 1.431309e-06, 1.875879e-06, 
    2.19407e-06, 1.311109e-06, 7.216083e-07, 1.599422e-06, 2.245653e-06, 
    9.252628e-05, 0.0004826667, 0.000885198, 0.001186546, 0.001150001,
  5.724816e-06, 5.652763e-06, 2.873411e-06, 1.976612e-06, 2.459948e-06, 
    4.418567e-06, 5.029022e-06, 5.850908e-06, 9.575758e-06, 4.871347e-05, 
    0.0003399267, 0.0005940303, 0.0008754538, 0.001063882, 0.0008321953,
  8.820265e-06, 8.503404e-06, 5.269665e-06, 4.301955e-06, 6.668005e-06, 
    7.844974e-06, 1.32999e-05, 1.982175e-05, 3.173688e-05, 0.0001181794, 
    0.0002594609, 0.0004161614, 0.0004764894, 0.0003014023, 3.764651e-05,
  8.598667e-06, 8.084166e-06, 9.441429e-06, 1.070107e-05, 1.385487e-05, 
    2.289802e-05, 3.51221e-05, 4.459812e-05, 5.764273e-05, 8.80147e-05, 
    0.0001129594, 0.0001343266, 5.566004e-05, 8.51341e-07, 3.634286e-08,
  1.253182e-05, 1.01845e-05, 1.22454e-05, 1.56323e-05, 1.732751e-05, 
    3.186127e-05, 4.911521e-05, 6.240468e-05, 7.489515e-05, 5.345793e-05, 
    2.893546e-05, 2.124172e-05, 1.588772e-06, 5.437783e-08, 2.823014e-07,
  1.995273e-05, 1.681396e-05, 1.32785e-05, 1.554925e-05, 2.68835e-05, 
    3.743673e-05, 4.798737e-05, 5.526502e-05, 5.391224e-05, 2.96205e-05, 
    9.200923e-05, 1.025982e-05, 5.252686e-06, 1.221854e-07, 5.086499e-08,
  9.35868e-06, 4.152331e-06, 1.478146e-06, 8.79767e-07, 4.569739e-07, 
    1.60146e-07, 2.189176e-07, 1.581777e-07, 5.765008e-08, 5.170428e-08, 
    6.010929e-08, 6.207182e-08, 2.602691e-06, 1.913751e-05, 5.351647e-05,
  1.140335e-05, 1.215153e-05, 5.286172e-06, 1.640008e-06, 2.86311e-06, 
    7.37935e-06, 7.016725e-06, 2.996994e-06, 3.90335e-07, 6.894577e-09, 
    9.967814e-08, 5.364414e-07, 4.348188e-06, 4.442546e-05, 0.000134851,
  1.362799e-05, 1.408848e-05, 1.057684e-05, 8.087185e-06, 2.276606e-05, 
    4.111189e-05, 5.697056e-05, 4.385348e-05, 1.576297e-05, 3.584726e-06, 
    9.214018e-08, 1.113794e-06, 5.186339e-06, 6.340371e-05, 0.0002515524,
  1.840772e-05, 1.739453e-05, 1.013341e-05, 1.452069e-05, 2.868934e-05, 
    5.651022e-05, 7.431744e-05, 5.12419e-05, 2.305969e-05, 1.401016e-05, 
    6.745762e-06, 4.869702e-06, 1.60505e-05, 0.0001654355, 0.0005444211,
  1.503564e-05, 9.940578e-06, 1.138774e-05, 1.025187e-05, 2.135534e-05, 
    4.035312e-05, 4.745522e-05, 3.56782e-05, 2.585243e-05, 1.745322e-05, 
    1.755423e-05, 1.627317e-05, 6.109008e-05, 0.0003279042, 0.0007059841,
  1.050874e-05, 1.073471e-05, 1.249026e-05, 1.279641e-05, 1.526845e-05, 
    2.639741e-05, 3.711884e-05, 3.599996e-05, 3.228211e-05, 3.441433e-05, 
    3.924762e-05, 4.49154e-05, 0.0001065805, 0.0002754229, 0.0003824615,
  1.17633e-05, 1.142364e-05, 1.135874e-05, 1.512626e-05, 1.856308e-05, 
    2.650865e-05, 2.710393e-05, 2.689497e-05, 2.66264e-05, 3.279084e-05, 
    4.476466e-05, 4.996457e-05, 3.213162e-05, 2.867657e-06, 5.952456e-07,
  7.473647e-06, 1.13265e-05, 1.05275e-05, 2.058357e-05, 2.153012e-05, 
    1.992076e-05, 1.747258e-05, 1.637948e-05, 1.961467e-05, 1.934731e-05, 
    2.186124e-05, 9.769575e-06, 1.814852e-06, 1.914491e-06, 1.076886e-06,
  6.076608e-06, 5.105847e-06, 1.183839e-05, 1.945559e-05, 1.970523e-05, 
    1.428035e-05, 1.434688e-05, 1.70977e-05, 2.06714e-05, 2.49671e-05, 
    1.606107e-05, 2.050259e-06, 5.440631e-07, 5.679443e-07, 1.490269e-06,
  4.227851e-06, 3.203502e-06, 7.977102e-06, 1.99296e-05, 1.711554e-05, 
    1.399911e-05, 1.890443e-05, 2.209416e-05, 7.474539e-05, 7.184791e-05, 
    1.943856e-05, 1.348089e-06, 2.163655e-06, 2.840995e-07, 7.860821e-07,
  1.189232e-06, 2.612066e-06, 2.198577e-06, 3.23684e-06, 3.573757e-06, 
    8.93325e-06, 0.0001136342, 0.00026577, 0.0004060779, 0.0005296196, 
    0.0006139955, 0.0006464259, 0.0006326772, 0.0005774418, 0.0004720916,
  1.865357e-06, 5.316339e-06, 5.460674e-06, 7.971245e-06, 2.015137e-05, 
    7.424656e-05, 0.0001558144, 0.0002175234, 0.0002588119, 0.0002913626, 
    0.0003542537, 0.0004140016, 0.0004651595, 0.0004699754, 0.000379428,
  3.213731e-06, 5.131905e-06, 4.861567e-06, 5.516025e-06, 2.550527e-05, 
    7.209725e-05, 9.984914e-05, 8.127152e-05, 6.804709e-05, 6.67089e-05, 
    5.749236e-05, 4.659953e-05, 3.049347e-05, 2.107714e-05, 1.425208e-05,
  3.348984e-06, 4.633822e-06, 8.755739e-06, 8.120694e-06, 2.344668e-05, 
    4.095314e-05, 4.204174e-05, 4.488907e-05, 4.522732e-05, 3.684679e-05, 
    2.459572e-05, 1.317357e-05, 6.488783e-06, 4.264577e-06, 4.271674e-06,
  8.002097e-07, 3.478767e-06, 7.829711e-06, 9.179632e-06, 1.559819e-05, 
    1.990833e-05, 2.862325e-05, 3.262067e-05, 1.359928e-05, 3.274354e-06, 
    1.778474e-06, 2.124753e-06, 2.182848e-06, 7.469231e-07, 3.519695e-07,
  2.257406e-07, 2.416946e-06, 4.848427e-06, 8.014808e-06, 9.019996e-06, 
    1.308215e-05, 1.899352e-05, 1.637836e-05, 9.6314e-07, 7.487126e-08, 
    3.285229e-07, 3.276705e-07, 5.800277e-08, 4.42708e-08, 1.187608e-07,
  1.780651e-06, 1.121283e-06, 5.90331e-06, 8.438773e-06, 1.67214e-05, 
    9.742564e-06, 1.592523e-05, 9.195724e-06, 2.082727e-07, 9.838816e-08, 
    9.503749e-08, 3.243774e-06, 1.117754e-06, 1.797215e-06, 8.944806e-07,
  1.307494e-06, 1.874785e-06, 5.498936e-06, 1.051347e-05, 1.983874e-05, 
    1.395539e-05, 3.8354e-05, 8.300806e-07, 1.149613e-07, 2.430609e-06, 
    9.70473e-06, 6.053882e-06, 2.442627e-06, 9.481313e-07, 7.058169e-07,
  2.851576e-06, 2.044622e-06, 4.702973e-06, 1.420926e-05, 1.570431e-05, 
    1.982899e-05, 1.872183e-05, 5.622487e-06, 1.768646e-06, 8.088507e-06, 
    5.247422e-06, 3.199114e-06, 1.745708e-06, 9.825804e-07, 1.141953e-06,
  1.464069e-06, 4.040852e-06, 3.712399e-06, 1.526313e-05, 2.087773e-05, 
    1.762042e-05, 2.844754e-05, 7.14445e-06, 1.037957e-05, 8.269089e-06, 
    3.356768e-06, 1.474258e-06, 8.921615e-07, 1.053344e-06, 8.217729e-07,
  4.907976e-07, 9.006725e-07, 7.202053e-07, 2.746036e-06, 1.657321e-06, 
    2.932991e-06, 3.089454e-06, 5.367854e-06, 2.311221e-06, 2.984471e-06, 
    1.926585e-06, 3.047202e-06, 3.30142e-06, 8.261973e-06, 5.292086e-05,
  1.630765e-06, 1.257294e-06, 2.105977e-06, 1.77166e-06, 4.229558e-06, 
    3.821471e-06, 5.694244e-06, 4.556894e-06, 1.461505e-06, 2.381121e-06, 
    1.756642e-06, 3.415739e-06, 7.471499e-06, 4.1546e-05, 0.0001439053,
  5.435514e-06, 5.664266e-06, 4.522802e-06, 2.995124e-06, 3.602926e-06, 
    6.274473e-06, 6.020155e-06, 3.808948e-06, 3.929933e-06, 5.811599e-06, 
    1.447187e-05, 2.75035e-05, 4.888272e-05, 9.475881e-05, 0.0001488892,
  3.940129e-06, 4.717457e-06, 3.653803e-06, 6.680594e-06, 4.898087e-06, 
    6.843954e-06, 6.180931e-06, 8.641982e-06, 6.894451e-06, 1.703998e-05, 
    3.074109e-05, 5.221812e-05, 6.914286e-05, 8.635064e-05, 0.0001018338,
  3.166791e-06, 3.376633e-06, 3.489216e-06, 4.711544e-06, 3.128959e-06, 
    7.113179e-06, 6.888397e-06, 8.199419e-06, 1.684036e-05, 3.118192e-05, 
    5.169928e-05, 6.210709e-05, 6.790303e-05, 7.471184e-05, 7.651086e-05,
  3.271925e-06, 1.916392e-06, 2.572949e-06, 3.002802e-06, 5.46578e-06, 
    8.232472e-06, 8.022163e-06, 2.156965e-05, 3.554186e-05, 5.424365e-05, 
    7.439453e-05, 7.508864e-05, 7.357579e-05, 6.234609e-05, 6.07404e-05,
  5.437634e-06, 4.957346e-07, 2.097981e-06, 3.024111e-06, 4.856908e-06, 
    1.10888e-05, 1.435934e-05, 3.588111e-05, 3.967573e-05, 2.605751e-05, 
    8.679056e-06, 3.233195e-05, 2.022636e-05, 9.430521e-06, 3.641302e-06,
  2.69498e-06, 2.841944e-06, 1.755235e-06, 2.720752e-06, 9.015345e-06, 
    1.734304e-05, 6.183996e-05, 7.554893e-05, 3.229762e-05, 2.810762e-05, 
    3.713221e-06, 3.063941e-06, 1.211246e-06, 1.061835e-06, 1.133445e-06,
  3.028887e-06, 1.762278e-06, 1.672488e-06, 6.099523e-06, 1.671869e-05, 
    3.799639e-05, 0.0001663399, 8.357505e-05, 1.010247e-05, 2.568695e-06, 
    1.575399e-06, 7.864218e-07, 6.600793e-07, 3.995162e-07, 1.965929e-07,
  2.112602e-06, 2.502831e-06, 2.673227e-06, 9.237763e-06, 1.942739e-05, 
    0.0001132539, 9.245561e-05, 1.081717e-05, 1.481703e-06, 8.816287e-07, 
    3.721947e-07, 1.823682e-08, 4.48519e-08, 2.088628e-07, 6.321648e-08,
  5.570319e-06, 5.84566e-06, 4.595167e-06, 3.62596e-06, 1.298013e-05, 
    2.933531e-05, 3.460305e-05, 3.037422e-05, 1.813177e-05, 1.015122e-05, 
    8.574978e-06, 9.641481e-06, 7.44047e-06, 5.967574e-06, 8.927331e-06,
  6.15751e-06, 5.605926e-06, 4.948874e-06, 8.093451e-06, 1.454925e-05, 
    2.797556e-05, 2.231278e-05, 1.397242e-05, 6.842752e-06, 6.57977e-06, 
    4.566387e-06, 4.180758e-06, 2.759496e-06, 2.724679e-06, 4.298405e-06,
  6.217304e-06, 6.71405e-06, 7.551466e-06, 1.205312e-05, 1.304457e-05, 
    1.733827e-05, 1.032797e-05, 7.250406e-06, 5.342596e-06, 4.353438e-06, 
    4.314282e-06, 2.697257e-06, 1.885312e-06, 1.220639e-06, 1.983984e-06,
  5.731536e-06, 8.223621e-06, 9.767986e-06, 1.190441e-05, 7.562066e-06, 
    9.673253e-06, 8.780111e-06, 9.707257e-06, 8.833103e-06, 4.097006e-06, 
    2.569284e-06, 2.370124e-06, 1.448313e-06, 9.069673e-07, 1.416359e-07,
  2.239327e-06, 8.36236e-06, 8.049999e-06, 1.337685e-05, 1.442837e-05, 
    9.648836e-06, 8.862909e-06, 9.395234e-06, 8.653251e-06, 6.749605e-06, 
    6.951997e-06, 9.528206e-06, 1.422814e-05, 1.691678e-05, 1.81082e-05,
  5.685126e-06, 9.693394e-06, 9.818612e-06, 3.21278e-05, 1.99259e-05, 
    1.551819e-05, 8.161759e-06, 4.984509e-06, 3.421569e-06, 1.671585e-06, 
    6.117008e-07, 3.187346e-06, 7.985816e-06, 2.579224e-05, 2.558848e-05,
  5.753852e-06, 5.995885e-06, 1.254112e-05, 3.924784e-05, 2.574824e-05, 
    1.886504e-05, 1.392452e-05, 4.269065e-06, 1.0067e-05, 1.849473e-05, 
    1.853603e-05, 1.113088e-05, 5.452796e-06, 5.827834e-06, 4.203617e-06,
  4.616437e-06, 1.20147e-05, 1.656141e-05, 7.751182e-05, 6.101387e-05, 
    5.577457e-05, 3.650597e-05, 2.282967e-05, 4.44865e-05, 3.318436e-05, 
    7.652267e-06, 2.547919e-06, 1.792925e-06, 2.379786e-06, 2.204285e-06,
  2.430806e-06, 7.987283e-06, 2.695153e-05, 6.217559e-05, 6.639441e-05, 
    3.432071e-05, 1.80637e-06, 3.990362e-06, 6.908539e-06, 6.503045e-06, 
    7.486713e-06, 2.788687e-06, 1.607464e-06, 2.017714e-06, 2.575623e-06,
  1.282656e-06, 1.003128e-05, 2.151799e-05, 4.317189e-05, 2.786288e-05, 
    4.433098e-06, 4.627545e-07, 1.562249e-06, 3.332654e-06, 7.74872e-06, 
    7.632133e-06, 4.472005e-06, 2.096083e-06, 2.235125e-06, 3.359662e-06,
  5.396131e-05, 3.881418e-05, 0.0001351227, 0.0001161812, 0.0001284415, 
    0.0001340612, 0.0001292992, 0.0001001318, 0.0001081991, 0.000127515, 
    0.0001658184, 0.0002003809, 0.0001962945, 0.0001597942, 0.0001235048,
  2.818466e-05, 8.770279e-05, 7.476473e-05, 0.0001699043, 0.0001425014, 
    0.0001160847, 0.0001102093, 0.0001016408, 7.995968e-05, 0.0001025317, 
    0.0001363813, 0.0001415497, 0.0001488124, 0.0001369856, 0.0001177177,
  3.431803e-05, 4.24846e-05, 0.0001399725, 9.689628e-05, 0.0001105714, 
    8.65515e-05, 8.521532e-05, 7.777357e-05, 6.678605e-05, 7.564443e-05, 
    0.0001097679, 0.00012566, 0.0001318085, 0.0001184364, 0.0001131913,
  3.386289e-05, 4.409329e-05, 4.293221e-05, 5.179796e-05, 4.516757e-05, 
    5.237813e-05, 4.624695e-05, 3.947699e-05, 5.355348e-05, 6.712322e-05, 
    7.827977e-05, 9.681815e-05, 9.75114e-05, 8.969256e-05, 8.236521e-05,
  1.529615e-05, 3.562275e-05, 2.503226e-05, 2.834096e-05, 3.746073e-05, 
    2.548232e-05, 2.793004e-05, 3.053503e-05, 4.466608e-05, 5.87725e-05, 
    6.133803e-05, 6.435056e-05, 6.697796e-05, 6.335065e-05, 5.908165e-05,
  2.130576e-05, 1.7959e-05, 1.74089e-05, 2.696191e-05, 3.228518e-05, 
    4.672615e-05, 5.507566e-05, 2.902479e-05, 3.660101e-05, 3.597143e-05, 
    4.930985e-05, 4.937394e-05, 5.862182e-05, 5.074419e-05, 7.58992e-05,
  1.549809e-05, 1.849512e-05, 2.203686e-05, 4.692556e-05, 6.157572e-05, 
    3.42989e-05, 2.315296e-05, 2.863924e-05, 2.099654e-05, 2.908953e-05, 
    5.040293e-05, 0.0001302754, 0.0001064102, 6.236933e-05, 7.883547e-05,
  2.352174e-05, 1.654285e-05, 4.12385e-05, 6.944522e-05, 6.547159e-05, 
    4.831762e-05, 3.643869e-05, 3.048659e-05, 4.46134e-05, 7.332356e-05, 
    0.000103865, 5.853601e-05, 3.846671e-05, 4.362961e-05, 5.090614e-05,
  4.292303e-05, 2.069267e-05, 4.069244e-05, 6.922825e-05, 4.796192e-05, 
    4.589213e-05, 4.265751e-05, 3.502318e-05, 4.9086e-05, 5.361174e-05, 
    5.906068e-05, 2.987335e-05, 2.029506e-05, 4.422575e-05, 3.858405e-05,
  3.418271e-05, 3.057437e-05, 3.953677e-05, 6.346941e-05, 5.274118e-05, 
    4.792151e-05, 5.173595e-05, 3.247557e-05, 7.203245e-05, 5.234425e-05, 
    3.534233e-05, 2.930656e-05, 3.0206e-05, 4.427705e-05, 2.364902e-05,
  2.378061e-06, 2.673193e-06, 3.002019e-06, 1.638192e-06, 2.247298e-06, 
    2.254749e-06, 3.218192e-06, 3.431445e-06, 5.96317e-06, 7.76991e-06, 
    9.323377e-06, 1.472005e-05, 1.668932e-05, 2.167421e-05, 2.272307e-05,
  3.154639e-06, 2.515334e-06, 2.797486e-06, 2.076653e-06, 2.172384e-06, 
    1.909691e-06, 2.450174e-06, 3.768453e-06, 4.720933e-06, 6.097005e-06, 
    7.468137e-06, 8.108736e-06, 1.294331e-05, 1.43747e-05, 1.693914e-05,
  3.045013e-06, 3.160455e-06, 3.062777e-06, 2.857236e-06, 1.748348e-06, 
    1.578621e-06, 1.201914e-06, 2.235762e-06, 2.194633e-06, 3.433045e-06, 
    4.884779e-06, 5.850113e-06, 5.988333e-06, 9.356698e-06, 9.845727e-06,
  1.943332e-06, 2.128139e-06, 3.932305e-06, 3.031283e-06, 2.987538e-06, 
    1.168219e-06, 4.310571e-07, 8.104162e-07, 1.157969e-06, 1.742003e-06, 
    2.946332e-06, 3.969894e-06, 4.05704e-06, 4.493009e-06, 4.835196e-06,
  2.342789e-06, 9.900069e-07, 1.491324e-06, 2.341126e-06, 4.405728e-06, 
    3.562423e-06, 2.831734e-06, 8.22919e-07, 7.094969e-07, 1.062754e-06, 
    1.736055e-06, 2.397389e-06, 4.016676e-06, 4.951233e-06, 4.670683e-06,
  4.55683e-06, 3.424264e-06, 1.905427e-06, 1.952547e-06, 2.265218e-06, 
    2.449451e-06, 3.968409e-06, 5.185284e-06, 4.60689e-06, 4.668474e-06, 
    1.935204e-06, 1.397641e-06, 2.672131e-06, 3.701941e-06, 5.187532e-06,
  4.231776e-06, 5.672577e-06, 3.185895e-06, 2.816106e-06, 2.926961e-06, 
    2.844018e-06, 2.501941e-06, 2.835802e-06, 2.413392e-06, 2.785572e-06, 
    2.612589e-06, 2.359552e-06, 1.40336e-06, 1.472753e-06, 3.161057e-06,
  3.805998e-06, 3.767303e-06, 5.107127e-06, 3.890226e-06, 2.026438e-06, 
    1.942206e-06, 2.210766e-06, 4.407257e-06, 2.451542e-06, 4.179836e-06, 
    4.686578e-06, 4.60297e-06, 3.611343e-06, 3.22355e-06, 2.736155e-06,
  2.66607e-06, 3.235803e-06, 3.74462e-06, 4.089294e-06, 2.890125e-06, 
    2.518174e-06, 2.347271e-06, 2.976341e-06, 2.512084e-06, 4.184187e-06, 
    2.524334e-06, 2.069793e-06, 3.236561e-06, 3.964709e-06, 4.022559e-06,
  2.841856e-06, 3.35114e-06, 4.092763e-06, 4.496374e-06, 4.372851e-06, 
    3.541004e-06, 4.308387e-06, 4.080333e-06, 2.583856e-06, 3.486701e-06, 
    2.757404e-06, 1.469902e-06, 1.932704e-06, 2.656188e-06, 4.033233e-06,
  8.344462e-06, 5.059575e-06, 3.989569e-06, 3.432788e-06, 2.09968e-06, 
    2.504392e-06, 1.430264e-06, 3.573432e-06, 7.433002e-06, 7.901353e-06, 
    4.277453e-06, 2.018669e-06, 1.400379e-06, 1.42892e-06, 8.600187e-07,
  8.761682e-06, 5.392046e-06, 4.097031e-06, 3.67128e-06, 3.87333e-06, 
    1.798673e-06, 1.107113e-06, 9.832451e-07, 2.498199e-06, 9.586304e-06, 
    7.089587e-06, 3.094893e-06, 2.503219e-06, 1.824726e-06, 1.196221e-06,
  9.510645e-06, 8.752325e-06, 6.879992e-06, 4.309694e-06, 5.037492e-06, 
    5.129126e-06, 2.095173e-06, 1.226155e-06, 7.092507e-07, 2.316785e-06, 
    8.055779e-06, 6.437693e-06, 3.509968e-06, 2.662304e-06, 6.709757e-07,
  9.687411e-06, 1.010102e-05, 7.382589e-06, 6.723035e-06, 5.36674e-06, 
    6.796993e-06, 3.461766e-06, 1.701854e-06, 9.153651e-07, 1.402604e-06, 
    2.455862e-06, 6.214818e-06, 1.264032e-06, 9.593464e-07, 8.702435e-07,
  9.393117e-06, 1.043926e-05, 9.614343e-06, 1.324763e-05, 8.041341e-06, 
    6.171104e-06, 4.838852e-06, 4.101955e-06, 2.389208e-06, 2.376195e-06, 
    1.300335e-06, 1.476221e-06, 2.763383e-06, 2.993568e-06, 7.165463e-07,
  9.747109e-06, 9.124813e-06, 1.27497e-05, 1.320274e-05, 1.288612e-05, 
    1.2984e-05, 7.937134e-06, 1.115394e-05, 5.915562e-06, 6.134341e-06, 
    4.490349e-06, 2.095412e-06, 3.121459e-06, 2.878623e-06, 1.544402e-06,
  9.903228e-06, 1.136356e-05, 1.31003e-05, 1.415477e-05, 1.991659e-05, 
    1.622615e-05, 2.129889e-05, 1.533983e-05, 1.232125e-05, 8.485429e-06, 
    6.361168e-06, 6.178258e-06, 9.095043e-06, 6.696135e-06, 4.079041e-06,
  9.402856e-06, 1.218045e-05, 1.762627e-05, 1.845587e-05, 1.660957e-05, 
    1.893303e-05, 1.520127e-05, 1.393453e-05, 1.34598e-05, 8.404667e-06, 
    8.727116e-06, 6.956335e-06, 7.519318e-06, 1.014385e-05, 1.024727e-05,
  1.027873e-05, 1.165032e-05, 1.311832e-05, 1.669656e-05, 1.788577e-05, 
    1.869342e-05, 1.94104e-05, 2.100314e-05, 1.237397e-05, 1.472972e-05, 
    1.423608e-05, 7.670003e-06, 7.637344e-06, 1.075182e-05, 1.064661e-05,
  1.229412e-05, 1.328633e-05, 1.478178e-05, 1.942212e-05, 1.849971e-05, 
    1.85506e-05, 2.197478e-05, 1.468396e-05, 1.603669e-05, 2.597209e-05, 
    1.873815e-05, 1.406484e-05, 1.629762e-05, 1.130782e-05, 1.109441e-05,
  2.020686e-06, 2.270657e-06, 2.606256e-06, 2.622458e-06, 3.926021e-06, 
    3.855992e-06, 5.252758e-06, 5.407852e-06, 8.949226e-06, 1.548427e-05, 
    1.892385e-05, 1.321915e-05, 1.500603e-05, 1.387641e-05, 7.623028e-06,
  2.507807e-06, 2.52359e-06, 3.336846e-06, 3.241564e-06, 4.376228e-06, 
    5.311682e-06, 4.008402e-06, 3.624843e-06, 7.51593e-06, 1.552622e-05, 
    1.519187e-05, 1.278541e-05, 2.280808e-05, 1.672651e-05, 1.255074e-05,
  3.640853e-06, 3.967291e-06, 5.925738e-06, 3.436078e-06, 3.663908e-06, 
    2.952448e-06, 6.005458e-06, 4.949288e-06, 1.123445e-05, 1.360081e-05, 
    1.376334e-05, 1.950946e-05, 1.964971e-05, 1.915196e-05, 1.446149e-05,
  3.576784e-06, 2.39818e-06, 3.869546e-06, 3.88499e-06, 3.962451e-06, 
    4.198973e-06, 5.457214e-06, 4.29979e-06, 6.841236e-06, 1.064693e-05, 
    1.197643e-05, 1.602746e-05, 1.817112e-05, 1.728957e-05, 1.734134e-05,
  4.33798e-06, 3.845236e-06, 3.516022e-06, 5.988303e-06, 4.486169e-06, 
    4.50051e-06, 3.329756e-06, 5.376656e-06, 8.151665e-06, 1.146165e-05, 
    1.616486e-05, 1.834607e-05, 1.799288e-05, 1.754821e-05, 1.665266e-05,
  2.780968e-06, 4.168866e-06, 6.584487e-06, 3.722525e-06, 3.531237e-06, 
    3.75286e-06, 7.177286e-06, 7.958311e-06, 7.517001e-06, 6.388666e-06, 
    1.306514e-05, 1.793618e-05, 1.833304e-05, 2.007357e-05, 1.535513e-05,
  4.659328e-06, 6.833534e-06, 7.833274e-06, 5.868351e-06, 4.226878e-06, 
    5.020742e-06, 7.402026e-06, 8.112602e-06, 8.077507e-06, 9.595072e-06, 
    1.28644e-05, 1.681027e-05, 2.067369e-05, 1.962643e-05, 1.716004e-05,
  3.312655e-06, 6.617391e-06, 9.762452e-06, 1.191269e-05, 3.073264e-06, 
    3.633549e-06, 4.000909e-06, 4.8091e-06, 1.015482e-05, 9.057113e-06, 
    1.171615e-05, 1.441058e-05, 1.565436e-05, 1.625046e-05, 2.056163e-05,
  3.961905e-06, 6.755708e-06, 1.049469e-05, 9.86722e-06, 3.744011e-06, 
    2.77361e-06, 3.146416e-06, 5.086682e-06, 5.736997e-06, 1.133309e-05, 
    1.337617e-05, 1.109929e-05, 1.496666e-05, 1.64331e-05, 1.752456e-05,
  2.827329e-06, 5.377421e-06, 1.028691e-05, 1.44514e-05, 6.587328e-06, 
    2.864815e-06, 6.086458e-06, 5.899253e-06, 6.862738e-06, 1.286349e-05, 
    1.052357e-05, 1.428401e-05, 1.582042e-05, 1.521113e-05, 1.237475e-05,
  0.000121912, 0.0001466002, 0.0001595332, 0.0001594423, 0.0001652288, 
    0.0001663755, 0.0001655574, 0.000171642, 0.0001754193, 0.0001754171, 
    0.000131184, 8.574746e-05, 6.217247e-05, 5.559692e-05, 3.187181e-05,
  0.0001130236, 0.0001398521, 0.0001526029, 0.0001488601, 0.000140033, 
    0.0001380051, 0.0001341922, 0.000146044, 0.0001413166, 0.0001124335, 
    7.044268e-05, 5.064527e-05, 5.05775e-05, 4.811513e-05, 3.295427e-05,
  0.0001082993, 0.0001335282, 0.0001379374, 0.0001326909, 0.0001183284, 
    0.0001107376, 0.0001176039, 0.0001116116, 8.694396e-05, 5.838163e-05, 
    4.744704e-05, 3.77015e-05, 3.162083e-05, 3.303393e-05, 2.704463e-05,
  0.0001050795, 0.0001094049, 9.237494e-05, 7.906884e-05, 7.690331e-05, 
    7.50482e-05, 6.746346e-05, 5.725715e-05, 3.712934e-05, 2.365934e-05, 
    2.233223e-05, 2.186942e-05, 2.779595e-05, 2.984459e-05, 2.49155e-05,
  9.209304e-05, 7.353193e-05, 6.705736e-05, 6.067187e-05, 5.934385e-05, 
    5.955567e-05, 5.108031e-05, 3.72883e-05, 1.76673e-05, 7.60862e-06, 
    1.228261e-05, 1.607266e-05, 2.494757e-05, 2.726057e-05, 1.890381e-05,
  7.556349e-05, 5.955282e-05, 4.135763e-05, 4.306817e-05, 4.57527e-05, 
    4.040371e-05, 3.054148e-05, 1.550843e-05, 3.754683e-06, 2.849527e-06, 
    5.837053e-06, 1.506588e-05, 2.221532e-05, 2.053523e-05, 1.539995e-05,
  6.185364e-05, 3.150191e-05, 3.565934e-05, 3.746539e-05, 3.546053e-05, 
    2.72812e-05, 7.102456e-06, 2.163815e-06, 9.156264e-07, 5.937215e-06, 
    7.736897e-06, 1.915728e-05, 1.914906e-05, 1.95452e-05, 1.016706e-05,
  4.846287e-05, 3.036917e-05, 4.620574e-05, 3.079876e-05, 2.090375e-05, 
    1.272914e-05, 1.032668e-06, 1.950503e-07, 8.026474e-07, 6.651704e-06, 
    2.271014e-05, 1.413867e-05, 1.252057e-05, 1.101167e-05, 8.995689e-06,
  1.000683e-05, 1.881468e-05, 4.958841e-05, 3.653667e-05, 2.030997e-06, 
    2.692623e-07, 4.029601e-08, 7.698164e-08, 9.367145e-07, 1.081144e-05, 
    2.056225e-05, 2.346156e-05, 1.40579e-05, 1.042549e-05, 7.067585e-06,
  6.290845e-06, 1.304218e-05, 3.252964e-05, 8.185968e-06, 1.351127e-06, 
    8.919659e-08, 1.738275e-09, 3.515161e-09, 1.114196e-06, 8.81011e-06, 
    1.828078e-05, 2.851304e-05, 2.008286e-05, 1.162766e-05, 5.626335e-06,
  5.442744e-06, 3.521841e-06, 2.987632e-06, 7.711348e-07, 2.900455e-06, 
    4.185413e-06, 7.282638e-06, 8.398823e-06, 1.177507e-05, 1.911096e-05, 
    5.768186e-05, 0.0001025509, 0.0001359703, 0.0001550111, 0.0001480694,
  3.650133e-06, 2.762987e-06, 2.319157e-06, 9.069078e-07, 9.412535e-07, 
    1.631848e-06, 3.545101e-06, 6.626048e-06, 1.299277e-05, 3.276586e-05, 
    6.656373e-05, 9.57995e-05, 0.0001170758, 0.0001059881, 0.0001090695,
  3.169155e-06, 2.712674e-06, 2.509676e-06, 1.795215e-06, 8.966252e-07, 
    8.415585e-07, 7.184208e-07, 6.10521e-06, 2.177868e-05, 4.478719e-05, 
    7.489148e-05, 9.530058e-05, 0.0001001864, 9.284366e-05, 8.708471e-05,
  6.131685e-06, 4.425224e-06, 3.340779e-06, 2.588252e-06, 2.112702e-06, 
    1.997323e-06, 5.702207e-06, 1.534677e-05, 3.063486e-05, 4.302193e-05, 
    6.243845e-05, 7.808433e-05, 7.657418e-05, 5.880041e-05, 8.561331e-05,
  2.505294e-06, 4.647349e-06, 3.989372e-06, 5.085006e-06, 6.938861e-06, 
    1.042829e-05, 1.622721e-05, 2.518575e-05, 3.853866e-05, 4.812697e-05, 
    5.830195e-05, 5.420756e-05, 4.154698e-05, 4.205308e-05, 8.395019e-05,
  4.510264e-06, 4.832821e-06, 7.264417e-06, 1.123539e-05, 1.131066e-05, 
    1.413302e-05, 1.725341e-05, 2.384371e-05, 3.581889e-05, 3.784176e-05, 
    3.456102e-05, 2.673722e-05, 2.512915e-05, 4.161288e-05, 0.0001003488,
  5.724633e-06, 7.212546e-06, 9.191846e-06, 1.119352e-05, 1.058744e-05, 
    1.233931e-05, 1.680717e-05, 2.084903e-05, 2.198434e-05, 1.886681e-05, 
    1.937008e-05, 1.522112e-05, 2.895372e-05, 6.808126e-05, 0.0001062757,
  1.294503e-05, 9.864791e-06, 1.191763e-05, 1.450903e-05, 1.340955e-05, 
    1.324771e-05, 1.332532e-05, 9.891753e-06, 1.087828e-05, 7.854231e-06, 
    8.375706e-06, 2.124843e-05, 4.640147e-05, 0.0001252215, 0.0002044319,
  2.218001e-05, 1.889625e-05, 1.602834e-05, 1.518424e-05, 3.205138e-05, 
    2.043537e-05, 1.237295e-05, 8.609095e-06, 4.444919e-06, 4.351859e-06, 
    8.413526e-06, 3.828774e-05, 7.897909e-05, 0.0001353392, 0.0002185391,
  2.68804e-05, 2.884713e-05, 3.126761e-05, 3.693187e-05, 2.692327e-05, 
    1.710881e-05, 9.202136e-06, 6.623524e-06, 7.553658e-06, 7.777929e-06, 
    3.25229e-05, 7.517703e-05, 0.0001071696, 0.000159013, 0.0002263758,
  9.3693e-06, 9.74713e-06, 1.095657e-05, 1.360791e-05, 1.762658e-05, 
    1.905475e-05, 2.079943e-05, 2.38735e-05, 3.744487e-05, 5.029727e-05, 
    3.200828e-05, 2.791206e-05, 2.968137e-05, 4.007472e-05, 3.863552e-05,
  1.004122e-05, 8.114182e-06, 6.967033e-06, 8.972345e-06, 1.132195e-05, 
    1.232734e-05, 1.790241e-05, 2.37532e-05, 3.355985e-05, 4.975684e-05, 
    4.305425e-05, 2.954279e-05, 2.941016e-05, 3.390362e-05, 3.4981e-05,
  8.713138e-06, 6.522811e-06, 7.049341e-06, 7.19117e-06, 7.632845e-06, 
    6.647716e-06, 9.163221e-06, 1.747207e-05, 2.547153e-05, 2.920591e-05, 
    2.877447e-05, 1.884823e-05, 2.347041e-05, 2.594854e-05, 2.682509e-05,
  3.249134e-06, 4.351253e-06, 4.653232e-06, 3.166965e-06, 4.319103e-06, 
    5.089335e-06, 6.406126e-06, 1.303897e-05, 2.172463e-05, 2.007626e-05, 
    1.586588e-05, 1.121062e-05, 1.476509e-05, 1.783379e-05, 1.718929e-05,
  5.489739e-06, 4.10648e-06, 3.080808e-06, 1.773818e-06, 4.488023e-06, 
    4.432487e-06, 3.914669e-06, 7.315173e-06, 8.58887e-06, 1.744885e-05, 
    1.362602e-05, 9.498805e-06, 6.909007e-06, 1.209197e-05, 1.050941e-05,
  7.979223e-06, 7.011717e-06, 4.903353e-06, 4.434714e-06, 4.921626e-06, 
    5.4441e-06, 5.467126e-06, 5.966308e-06, 5.813064e-06, 3.813006e-06, 
    5.824717e-06, 5.96884e-06, 5.02727e-06, 5.617802e-06, 7.608814e-06,
  1.165503e-05, 1.284291e-05, 8.889006e-06, 8.522905e-06, 6.887003e-06, 
    7.298455e-06, 6.965257e-06, 5.525524e-06, 2.934105e-06, 1.613178e-06, 
    8.246994e-07, 1.307377e-06, 1.017728e-06, 2.236613e-06, 3.548573e-06,
  1.543808e-05, 1.527048e-05, 1.682321e-05, 9.691545e-06, 9.03738e-06, 
    7.559211e-06, 7.800029e-06, 6.255456e-06, 2.957803e-06, 6.643578e-07, 
    5.792152e-07, 5.462643e-07, 8.040331e-07, 7.644603e-07, 7.54459e-07,
  1.24584e-05, 1.977056e-05, 2.002306e-05, 1.959896e-05, 1.258411e-05, 
    8.576589e-06, 7.949139e-06, 4.782175e-06, 1.282443e-06, 3.82474e-07, 
    1.42463e-07, 3.953419e-07, 4.995479e-07, 5.938631e-07, 5.318466e-07,
  1.921033e-05, 1.678681e-05, 2.002492e-05, 2.073917e-05, 1.66264e-05, 
    1.178606e-05, 9.028548e-06, 6.617654e-06, 2.776058e-06, 1.103225e-06, 
    5.484692e-07, 7.962277e-07, 6.139663e-07, 6.49293e-08, 1.427798e-06,
  4.351784e-06, 4.586674e-06, 1.023565e-05, 8.763298e-06, 1.302355e-05, 
    1.30731e-05, 1.699282e-05, 1.422887e-05, 2.273725e-05, 1.799975e-05, 
    1.151167e-05, 1.531479e-05, 1.78457e-05, 2.190686e-05, 3.257467e-05,
  1.466521e-06, 5.168611e-06, 9.39549e-06, 1.217797e-05, 1.484966e-05, 
    1.334904e-05, 1.431621e-05, 1.738083e-05, 2.054282e-05, 1.713809e-05, 
    1.208358e-05, 9.770672e-06, 1.32607e-05, 1.377071e-05, 1.81523e-05,
  5.910821e-07, 1.989266e-06, 4.160243e-06, 7.275697e-06, 9.226333e-06, 
    1.578279e-05, 1.349252e-05, 2.455783e-05, 2.751107e-05, 1.110199e-05, 
    1.27877e-05, 8.61968e-06, 9.833253e-06, 1.101496e-05, 1.325674e-05,
  4.690463e-06, 3.163719e-06, 2.368753e-06, 5.686078e-06, 6.099329e-06, 
    1.006293e-05, 1.914635e-05, 1.965003e-05, 2.039706e-05, 2.104144e-05, 
    9.154496e-06, 1.678697e-05, 1.042927e-05, 9.379193e-06, 9.286098e-06,
  4.658373e-06, 3.624398e-06, 3.172202e-06, 5.53428e-06, 7.357229e-06, 
    6.92989e-06, 6.674079e-06, 1.374618e-05, 1.565641e-05, 1.343142e-05, 
    1.690879e-05, 1.480232e-05, 1.775878e-05, 1.500408e-05, 4.198385e-06,
  6.593045e-06, 5.319078e-06, 5.095435e-06, 5.60771e-06, 7.508313e-06, 
    6.593159e-06, 7.581325e-06, 9.185332e-06, 7.337162e-06, 1.233381e-05, 
    1.325196e-05, 1.17123e-05, 1.718185e-05, 1.723258e-05, 9.050667e-06,
  8.27677e-06, 7.032146e-06, 7.500971e-06, 8.866929e-06, 8.295402e-06, 
    7.421936e-06, 7.40938e-06, 7.043272e-06, 7.372473e-06, 7.977581e-06, 
    7.092811e-06, 7.600348e-06, 9.506358e-06, 7.44205e-06, 7.551227e-06,
  8.009977e-06, 8.373087e-06, 1.038798e-05, 9.591636e-06, 9.02008e-06, 
    1.01526e-05, 6.962964e-06, 4.087101e-06, 3.750389e-06, 4.677061e-06, 
    6.428987e-06, 5.707815e-06, 4.856572e-06, 5.943169e-06, 6.459484e-06,
  7.695213e-06, 1.003388e-05, 1.079451e-05, 9.360213e-06, 9.044516e-06, 
    9.224804e-06, 8.772e-06, 6.190964e-06, 5.045386e-06, 4.230862e-06, 
    4.360105e-06, 2.833438e-06, 2.910112e-06, 3.74916e-06, 1.979741e-06,
  7.403721e-06, 8.712792e-06, 8.987777e-06, 9.500223e-06, 8.89745e-06, 
    9.461525e-06, 1.102776e-05, 1.028758e-05, 7.514502e-06, 6.803777e-06, 
    4.216907e-06, 2.324261e-06, 1.568018e-07, 4.393582e-07, 1.232626e-07,
  5.059468e-06, 3.819174e-06, 3.400486e-06, 4.068364e-06, 5.972998e-06, 
    8.367999e-06, 7.054887e-06, 4.242118e-06, 2.469231e-06, 1.665195e-06, 
    2.683004e-06, 4.334496e-06, 9.227368e-06, 1.018527e-05, 9.791031e-06,
  8.301127e-06, 4.476077e-06, 3.396962e-06, 4.441755e-06, 6.054792e-06, 
    5.761125e-06, 5.962218e-06, 5.186091e-06, 3.433298e-06, 1.682909e-06, 
    2.880252e-06, 3.925811e-06, 7.229386e-06, 8.549293e-06, 8.610942e-06,
  8.10134e-06, 6.763463e-06, 4.692852e-06, 4.751638e-06, 5.476424e-06, 
    7.015166e-06, 1.040487e-05, 4.652779e-06, 4.971643e-06, 5.233587e-06, 
    4.048122e-06, 3.481444e-06, 5.586379e-06, 8.791664e-06, 1.095922e-05,
  5.646044e-06, 5.340654e-06, 6.064699e-06, 4.893895e-06, 6.876717e-06, 
    8.088536e-06, 8.877552e-06, 9.186322e-06, 8.846885e-06, 5.46617e-06, 
    6.368658e-06, 4.325788e-06, 6.53584e-06, 1.012176e-05, 1.324235e-05,
  6.372182e-06, 5.459334e-06, 4.806832e-06, 5.927896e-06, 7.225553e-06, 
    7.505746e-06, 7.899564e-06, 9.427403e-06, 6.399372e-06, 5.94663e-06, 
    4.362297e-06, 3.740227e-06, 3.440812e-06, 7.057843e-06, 1.111801e-05,
  7.0349e-06, 7.409901e-06, 4.171991e-06, 5.415327e-06, 5.099995e-06, 
    4.891408e-06, 6.265891e-06, 6.03732e-06, 5.751519e-06, 3.986481e-06, 
    3.192949e-06, 4.789235e-06, 4.332426e-06, 5.929341e-06, 8.004483e-06,
  6.343274e-06, 5.905141e-06, 4.918902e-06, 4.794655e-06, 3.28831e-06, 
    3.92331e-06, 5.149565e-06, 3.940215e-06, 2.625635e-06, 2.013898e-06, 
    3.446819e-06, 3.230535e-06, 3.914988e-06, 4.449802e-06, 5.536489e-06,
  6.949445e-06, 5.942576e-06, 4.218079e-06, 4.529734e-06, 3.541257e-06, 
    2.695435e-06, 2.064143e-06, 1.982201e-06, 3.11956e-06, 3.672319e-06, 
    4.588725e-06, 4.003388e-06, 5.204954e-06, 5.240466e-06, 5.344557e-06,
  6.838418e-06, 6.315137e-06, 7.553814e-06, 5.024525e-06, 3.232339e-06, 
    3.583155e-06, 2.524529e-06, 3.147162e-06, 3.330856e-06, 4.693783e-06, 
    5.291896e-06, 6.526912e-06, 6.92957e-06, 7.454945e-06, 6.158256e-06,
  7.401806e-06, 6.425875e-06, 5.374105e-06, 4.473639e-06, 4.345048e-06, 
    4.202976e-06, 4.248953e-06, 4.134647e-06, 4.055974e-06, 5.585114e-06, 
    6.16326e-06, 6.147766e-06, 8.434467e-06, 7.409402e-06, 7.2117e-06,
  0.0002914674, 0.0002578552, 0.0001686036, 0.0001264693, 5.728534e-05, 
    1.048291e-05, 3.801633e-06, 2.277463e-06, 5.99167e-06, 4.132628e-06, 
    6.808289e-06, 7.407567e-06, 4.575001e-06, 1.546613e-07, 3.804185e-07,
  0.000270632, 0.0002103963, 0.0001428439, 0.0001085007, 7.273279e-05, 
    2.678842e-05, 2.697947e-06, 4.289221e-06, 6.224323e-06, 6.677687e-06, 
    8.729752e-06, 7.293784e-06, 9.204556e-06, 2.413572e-06, 4.170833e-07,
  0.0003154409, 0.0002282035, 0.0001497728, 8.426351e-05, 5.044262e-05, 
    3.305247e-05, 4.740436e-06, 5.409745e-06, 2.010897e-06, 7.942013e-06, 
    8.282432e-06, 8.638495e-06, 6.391149e-06, 1.242975e-06, 1.343937e-06,
  0.0002544865, 0.0002343411, 0.000157522, 8.432843e-05, 3.996933e-05, 
    2.462185e-05, 1.101267e-05, 1.646369e-06, 2.434506e-06, 1.073469e-06, 
    5.746143e-06, 1.03336e-05, 7.183675e-06, 3.929062e-06, 2.493657e-06,
  0.0001782782, 0.0001978513, 0.000144249, 0.00010044, 6.182512e-05, 
    2.808511e-05, 1.416732e-05, 4.8309e-06, 7.317817e-07, 1.782469e-06, 
    4.47397e-06, 6.300442e-06, 7.609548e-06, 2.396944e-06, 2.398843e-06,
  7.898003e-05, 0.0001233081, 8.554929e-05, 6.073539e-05, 5.706597e-05, 
    3.909766e-05, 1.404969e-05, 6.557137e-06, 1.475353e-06, 1.018946e-06, 
    2.595386e-06, 5.768964e-06, 6.797083e-06, 7.361589e-06, 2.31816e-06,
  3.342805e-05, 3.181218e-05, 4.087716e-05, 1.6354e-05, 1.870436e-05, 
    2.117353e-05, 1.324284e-05, 4.858695e-06, 3.274307e-06, 1.211095e-06, 
    1.07741e-06, 2.92555e-06, 9.735202e-06, 8.273741e-06, 9.663658e-06,
  4.683387e-05, 4.96313e-05, 5.818171e-05, 1.801169e-05, 7.49155e-06, 
    9.422512e-06, 7.713788e-06, 5.183577e-06, 2.758669e-06, 1.520979e-06, 
    1.702331e-06, 2.914595e-06, 3.939495e-06, 8.317639e-06, 1.017417e-05,
  5.563948e-05, 4.174306e-05, 3.560602e-05, 1.831052e-05, 9.029836e-06, 
    3.396086e-06, 3.963313e-06, 3.698412e-06, 3.095878e-06, 2.463658e-06, 
    2.515312e-06, 1.44013e-06, 2.139677e-06, 3.67387e-06, 6.098845e-06,
  2.377543e-05, 3.668045e-05, 3.912422e-05, 1.090485e-05, 3.409872e-06, 
    1.684574e-06, 1.975974e-06, 2.823455e-06, 3.503881e-06, 3.772476e-06, 
    3.285076e-06, 2.631894e-06, 1.908797e-06, 2.154861e-06, 2.717879e-06,
  1.068884e-05, 2.265722e-05, 5.286324e-05, 8.70449e-05, 0.0001385926, 
    0.0001724014, 0.0001935086, 0.0002261517, 0.000247177, 0.000243409, 
    0.0002558304, 0.0002615644, 0.0002533496, 0.0002324102, 0.0002056583,
  8.646896e-06, 1.921469e-05, 4.754846e-05, 8.39413e-05, 0.0001205121, 
    0.0001779207, 0.0002267845, 0.0002743898, 0.0003012656, 0.0003097091, 
    0.0003159947, 0.0003374482, 0.0003143053, 0.0002762532, 0.0002433099,
  6.400083e-06, 1.410824e-05, 4.081664e-05, 6.281184e-05, 7.103127e-05, 
    9.939016e-05, 0.0001377357, 0.000160393, 0.0001992667, 0.0002325878, 
    0.0002512364, 0.000231139, 0.0002005263, 0.0002018599, 0.0001579247,
  3.152404e-06, 1.001817e-05, 3.251099e-05, 4.641605e-05, 4.997602e-05, 
    5.489551e-05, 5.790872e-05, 5.59927e-05, 6.626989e-05, 9.043328e-05, 
    9.438536e-05, 7.599044e-05, 6.407068e-05, 5.431009e-05, 4.381288e-05,
  1.525032e-06, 1.048732e-05, 3.141685e-05, 4.13331e-05, 5.003606e-05, 
    4.943923e-05, 2.44635e-05, 2.268572e-05, 1.948276e-05, 2.368004e-05, 
    2.062999e-05, 1.722628e-05, 1.043184e-05, 5.688045e-06, 4.051223e-06,
  4.352335e-07, 7.677276e-06, 3.133554e-05, 5.133832e-05, 7.430304e-05, 
    4.350122e-05, 1.972959e-05, 1.49802e-05, 1.956671e-05, 1.647862e-05, 
    1.298713e-05, 6.693864e-06, 1.818488e-06, 1.963746e-06, 2.583518e-06,
  8.017687e-07, 9.033823e-06, 2.27474e-05, 6.027918e-05, 6.405522e-05, 
    5.449305e-05, 2.693674e-05, 1.906065e-05, 1.562715e-05, 9.39534e-06, 
    1.559924e-06, 9.399683e-07, 3.775089e-06, 5.226801e-06, 3.128775e-06,
  1.760914e-05, 2.522736e-05, 3.56293e-05, 1.757846e-05, 4.9877e-05, 
    3.353676e-05, 4.317386e-05, 3.116348e-05, 9.297882e-06, 1.359577e-06, 
    6.435347e-07, 1.01859e-06, 2.64059e-06, 4.37896e-06, 6.478345e-06,
  4.679347e-05, 5.062448e-05, 4.225939e-05, 5.319759e-05, 3.097688e-05, 
    2.162664e-05, 3.093213e-05, 4.147346e-05, 2.6234e-05, 1.246455e-05, 
    7.340208e-06, 3.029592e-06, 2.345115e-06, 2.781427e-06, 5.098572e-06,
  6.773424e-05, 7.413024e-05, 8.910777e-05, 7.124165e-05, 2.895349e-05, 
    1.034209e-05, 8.325551e-06, 4.527712e-06, 7.610163e-06, 1.014965e-05, 
    7.118762e-06, 6.105676e-06, 4.46483e-06, 4.407099e-06, 2.713783e-06,
  6.568405e-06, 1.173796e-05, 9.303953e-06, 8.155364e-06, 8.677695e-06, 
    1.095072e-05, 8.853057e-06, 1.50682e-05, 8.717828e-06, 1.224306e-05, 
    1.565794e-05, 1.684998e-05, 1.525771e-05, 1.544707e-05, 2.266896e-05,
  5.563554e-06, 7.138818e-06, 8.44827e-06, 1.030084e-05, 6.633029e-06, 
    1.002117e-05, 1.26722e-05, 8.547547e-06, 1.209319e-05, 2.275693e-05, 
    9.666462e-06, 1.239496e-05, 1.602021e-05, 9.638591e-06, 2.004627e-05,
  3.536077e-06, 3.803365e-06, 5.249355e-06, 7.846373e-06, 8.581463e-06, 
    7.436356e-06, 1.113608e-05, 9.824576e-06, 1.729544e-05, 1.207656e-05, 
    9.91402e-06, 8.132252e-06, 9.492225e-06, 1.275076e-05, 1.917449e-05,
  2.465562e-06, 2.3124e-06, 2.931771e-06, 4.354135e-06, 4.349063e-06, 
    6.042683e-06, 6.487291e-06, 7.06372e-06, 5.537217e-06, 7.378685e-06, 
    6.168048e-06, 7.056501e-06, 8.059757e-06, 1.208781e-05, 1.852839e-05,
  1.037015e-06, 4.827288e-07, 9.466338e-07, 8.480281e-07, 1.456446e-06, 
    2.218843e-06, 2.71141e-06, 3.254082e-06, 3.268968e-06, 2.706307e-06, 
    3.088907e-06, 6.30304e-06, 1.137748e-05, 1.546552e-05, 1.567394e-05,
  1.976719e-07, 2.118741e-08, 1.620227e-08, 1.611575e-07, 4.108453e-07, 
    5.958651e-07, 1.582244e-06, 2.710334e-06, 3.022744e-06, 2.407347e-06, 
    3.864397e-06, 1.192277e-05, 1.557242e-05, 1.138235e-05, 1.249848e-05,
  7.670618e-09, 1.049722e-09, 2.305383e-09, 1.261357e-08, 1.663322e-07, 
    3.936525e-07, 2.846009e-07, 3.09455e-07, 1.217712e-06, 4.703292e-06, 
    1.130139e-05, 1.234758e-05, 1.243647e-05, 1.179536e-05, 1.414728e-05,
  3.488259e-09, 9.367953e-10, 1.41108e-07, 8.369661e-09, 1.499126e-07, 
    2.845943e-08, 6.714875e-07, 1.765695e-06, 2.629129e-06, 5.157973e-06, 
    8.059465e-06, 1.018027e-05, 1.043183e-05, 1.159372e-05, 1.504024e-05,
  3.61223e-08, 4.261146e-08, 2.123546e-08, 8.00958e-09, 1.671408e-07, 
    7.992489e-07, 4.267484e-06, 2.631343e-06, 5.215476e-06, 6.668063e-06, 
    6.338203e-06, 6.256477e-06, 9.792937e-06, 1.987479e-05, 3.571629e-05,
  1.684103e-06, 1.117689e-06, 5.477063e-07, 3.736796e-06, 9.295225e-06, 
    5.958822e-06, 4.249495e-06, 3.896376e-06, 6.820255e-06, 6.614423e-06, 
    5.769938e-06, 9.962653e-06, 1.76403e-05, 2.297176e-05, 2.127053e-05,
  1.306359e-07, 1.05926e-07, 1.204182e-07, 8.220771e-08, 3.694567e-07, 
    4.043623e-07, 4.448577e-07, 1.179152e-06, 1.623426e-06, 4.148299e-06, 
    5.789853e-06, 9.319334e-06, 1.983584e-05, 3.030922e-05, 4.301052e-05,
  4.280092e-07, 3.019992e-07, 2.992934e-07, 1.017568e-07, 2.981072e-07, 
    5.389617e-07, 6.180294e-07, 7.784348e-07, 1.587926e-06, 3.595718e-06, 
    1.862657e-05, 2.775234e-05, 3.390746e-05, 3.62039e-05, 3.191951e-05,
  9.339664e-07, 7.965119e-07, 8.074673e-07, 6.796391e-07, 1.023587e-06, 
    1.272435e-06, 1.107123e-06, 1.812981e-06, 3.486557e-06, 1.111949e-05, 
    1.611971e-05, 2.019317e-05, 2.922766e-05, 2.722944e-05, 1.992033e-05,
  1.156947e-06, 1.212031e-06, 1.581442e-06, 1.856419e-06, 2.031124e-06, 
    2.709111e-06, 3.090207e-06, 2.511569e-06, 8.204122e-06, 9.808595e-06, 
    1.07781e-05, 1.142673e-05, 1.142502e-05, 1.336232e-05, 2.117342e-05,
  1.894156e-06, 2.11301e-06, 2.169164e-06, 2.063947e-06, 1.601126e-06, 
    2.688817e-06, 2.830223e-06, 5.698057e-06, 6.838945e-06, 6.572816e-06, 
    6.95681e-06, 8.276739e-06, 8.485386e-06, 9.067009e-06, 8.752783e-06,
  4.719062e-05, 3.527059e-06, 2.975335e-06, 2.265848e-06, 1.796114e-06, 
    2.173055e-06, 2.89592e-06, 4.214199e-06, 4.085523e-06, 4.35629e-06, 
    5.620189e-06, 4.727118e-06, 6.656279e-06, 4.637958e-06, 5.879591e-06,
  0.0001106678, 5.742299e-05, 6.350294e-06, 2.105292e-06, 1.662721e-06, 
    1.475667e-06, 1.622041e-06, 1.18441e-06, 2.178057e-06, 3.362168e-06, 
    2.606422e-06, 3.29663e-06, 3.216749e-06, 3.530722e-06, 4.22916e-06,
  4.040096e-05, 2.375679e-05, 1.804876e-05, 6.700577e-06, 1.975935e-06, 
    1.045379e-06, 1.548488e-06, 1.452431e-06, 1.653106e-06, 1.581433e-06, 
    1.985462e-06, 1.437376e-06, 3.293239e-06, 2.179946e-06, 2.485208e-06,
  1.754256e-05, 1.374084e-05, 8.04409e-06, 5.982245e-06, 1.654243e-06, 
    1.214183e-06, 1.311679e-06, 1.246598e-06, 8.549639e-07, 1.413955e-06, 
    2.073959e-06, 2.17997e-06, 2.256052e-06, 3.313426e-06, 6.891637e-06,
  1.355059e-05, 8.988699e-06, 5.186799e-06, 4.126756e-06, 3.350402e-06, 
    3.405961e-06, 2.200994e-06, 1.61802e-06, 2.744116e-06, 3.05094e-06, 
    4.385759e-06, 4.875084e-06, 1.029069e-05, 1.264374e-05, 1.031106e-05,
  4.092961e-07, 3.33343e-08, 4.921749e-08, 2.589458e-07, 7.910863e-07, 
    1.442634e-06, 2.56813e-06, 5.340601e-06, 6.006884e-06, 4.060938e-06, 
    3.32491e-06, 2.068311e-06, 5.442598e-06, 6.563525e-06, 7.12996e-06,
  1.152989e-06, 1.61241e-07, 2.827043e-07, 2.455906e-07, 1.567049e-07, 
    3.053047e-07, 1.014765e-06, 3.594282e-06, 4.634476e-06, 4.152311e-06, 
    4.406749e-06, 3.212069e-06, 3.93805e-06, 5.020224e-06, 6.105084e-06,
  3.069395e-06, 4.237411e-07, 2.466728e-07, 1.54783e-07, 1.615128e-07, 
    8.882633e-08, 4.269766e-07, 1.013094e-06, 2.761673e-06, 2.804221e-06, 
    2.933849e-06, 2.44006e-06, 2.58574e-06, 3.462028e-06, 5.296492e-06,
  6.730083e-06, 3.118179e-06, 5.005235e-07, 2.922293e-07, 7.250653e-07, 
    3.12323e-07, 3.738084e-07, 5.194362e-07, 1.083391e-06, 8.339131e-07, 
    2.169274e-06, 2.097832e-06, 1.361982e-06, 1.410221e-06, 3.099896e-06,
  5.756541e-06, 8.33461e-06, 1.936648e-06, 3.734215e-07, 3.623185e-07, 
    8.564723e-07, 7.420924e-07, 2.35266e-07, 3.248223e-07, 1.763272e-06, 
    1.47053e-06, 1.525257e-06, 1.435381e-06, 1.679824e-06, 2.367994e-06,
  1.095235e-06, 2.028839e-06, 7.065393e-06, 1.0324e-06, 4.382072e-07, 
    4.710635e-07, 2.822169e-07, 2.859421e-07, 6.035564e-07, 2.081564e-07, 
    2.22188e-07, 6.653428e-07, 1.316975e-06, 1.269493e-06, 1.915481e-06,
  1.836877e-06, 6.37735e-06, 4.63178e-06, 5.918651e-06, 2.554336e-06, 
    1.192717e-06, 1.188443e-06, 9.963138e-07, 7.693906e-07, 7.162583e-07, 
    4.927312e-07, 4.279677e-07, 4.841217e-07, 1.306032e-06, 1.508695e-06,
  7.408271e-06, 7.18843e-06, 5.97048e-06, 1.057049e-05, 9.418348e-06, 
    6.834691e-06, 3.241355e-06, 2.483979e-06, 2.359486e-06, 2.018435e-06, 
    2.295042e-06, 2.680003e-06, 2.872166e-06, 1.724628e-06, 3.233064e-06,
  5.796092e-06, 5.180577e-06, 5.546469e-06, 5.597752e-06, 6.268765e-06, 
    9.363527e-06, 6.446444e-06, 5.630402e-06, 5.009562e-06, 4.040285e-06, 
    3.057136e-06, 3.75326e-06, 2.496936e-06, 3.510936e-06, 3.783438e-06,
  2.550681e-06, 2.588109e-06, 1.978167e-06, 3.656816e-06, 5.675722e-06, 
    8.293449e-06, 1.117363e-05, 1.046346e-05, 1.112628e-05, 5.883077e-06, 
    5.479466e-06, 4.850924e-06, 4.357839e-06, 3.390559e-06, 5.044334e-06,
  6.723724e-06, 7.976554e-06, 8.698486e-06, 7.454117e-06, 1.113006e-05, 
    1.43953e-05, 1.176839e-05, 1.05805e-05, 1.058083e-05, 1.153091e-05, 
    9.549428e-06, 9.967448e-06, 1.017853e-05, 8.99404e-06, 6.675517e-06,
  6.586053e-06, 7.009252e-06, 7.807246e-06, 8.272183e-06, 1.002242e-05, 
    1.150019e-05, 1.106607e-05, 8.707259e-06, 9.810326e-06, 1.000594e-05, 
    1.19726e-05, 1.418193e-05, 1.157224e-05, 1.073358e-05, 9.868085e-06,
  3.788563e-06, 5.696158e-06, 8.419996e-06, 9.289178e-06, 9.269771e-06, 
    8.605218e-06, 9.513431e-06, 8.958461e-06, 9.177379e-06, 1.03552e-05, 
    1.032473e-05, 1.086782e-05, 1.303903e-05, 1.105377e-05, 1.02943e-05,
  5.361e-06, 6.32297e-06, 8.142569e-06, 8.324711e-06, 8.903748e-06, 
    9.943116e-06, 8.36544e-06, 1.04568e-05, 7.562553e-06, 9.493865e-06, 
    7.901815e-06, 7.760676e-06, 8.048585e-06, 1.085518e-05, 8.801088e-06,
  4.450248e-06, 5.895252e-06, 8.447308e-06, 9.072233e-06, 1.005866e-05, 
    7.501912e-06, 7.939952e-06, 6.763358e-06, 6.247602e-06, 7.701748e-06, 
    6.907529e-06, 7.312331e-06, 7.017321e-06, 8.027539e-06, 8.69738e-06,
  2.206216e-06, 4.327546e-06, 8.590149e-06, 8.437278e-06, 9.272342e-06, 
    7.087767e-06, 6.327464e-06, 3.874459e-06, 6.355419e-06, 4.388123e-06, 
    4.603409e-06, 5.381778e-06, 6.791847e-06, 4.761601e-06, 5.373705e-06,
  4.001563e-06, 3.168607e-06, 5.075661e-06, 7.918909e-06, 7.095625e-06, 
    6.617081e-06, 5.045702e-06, 5.900538e-06, 4.004711e-06, 3.830176e-06, 
    4.610293e-06, 4.72205e-06, 5.236033e-06, 6.585296e-06, 4.255272e-06,
  5.635124e-06, 2.438089e-06, 4.439219e-06, 4.523776e-06, 6.710373e-06, 
    6.621326e-06, 7.163027e-06, 6.848336e-06, 5.767561e-06, 4.837313e-06, 
    4.251376e-06, 5.027458e-06, 5.651655e-06, 3.920205e-06, 3.46296e-06,
  3.860503e-06, 1.806891e-06, 1.539639e-06, 3.914945e-06, 6.983526e-06, 
    6.729393e-06, 7.436761e-06, 9.163905e-06, 8.728317e-06, 5.323527e-06, 
    5.403388e-06, 7.20459e-06, 4.399958e-06, 4.390664e-06, 5.698891e-06,
  1.828044e-06, 1.453287e-06, 2.304832e-06, 3.027513e-06, 4.671056e-06, 
    6.354678e-06, 7.802526e-06, 1.193164e-05, 1.140358e-05, 6.505548e-06, 
    7.070893e-06, 6.756344e-06, 6.281226e-06, 6.298544e-06, 5.222653e-06,
  1.280729e-05, 4.656479e-06, 7.437541e-06, 5.955312e-06, 8.076397e-06, 
    5.77936e-06, 7.048874e-06, 5.692387e-06, 7.018056e-06, 5.392909e-06, 
    5.269475e-06, 7.988654e-06, 6.000399e-06, 8.572515e-06, 8.460968e-06,
  8.305074e-08, 3.060016e-08, 2.204991e-07, 8.069681e-07, 5.648874e-08, 
    1.148705e-06, 4.170903e-06, 5.056175e-06, 8.214601e-06, 7.622405e-06, 
    8.766287e-06, 9.592609e-06, 9.347028e-06, 9.606129e-06, 1.087413e-05,
  1.822905e-09, 1.904583e-08, 1.568802e-07, 5.864626e-07, 5.405608e-07, 
    9.336893e-07, 1.528415e-06, 3.587689e-06, 4.842497e-06, 5.838725e-06, 
    6.965499e-06, 7.466304e-06, 8.714064e-06, 8.017244e-06, 8.258206e-06,
  1.217966e-07, 1.896481e-07, 3.39604e-07, 9.138938e-07, 1.887848e-06, 
    2.720818e-06, 2.351922e-06, 3.178801e-06, 3.288053e-06, 3.36224e-06, 
    5.396667e-06, 5.62116e-06, 5.128429e-06, 4.66895e-06, 7.624222e-06,
  7.368254e-07, 1.173164e-06, 1.616665e-06, 3.539482e-06, 5.212628e-06, 
    4.091919e-06, 3.803509e-06, 2.039758e-06, 2.951017e-06, 1.861792e-06, 
    2.714526e-06, 2.156333e-06, 2.741488e-06, 5.188504e-06, 5.942898e-06,
  1.873431e-06, 2.241822e-06, 3.629309e-06, 4.827052e-06, 4.590982e-06, 
    4.021796e-06, 3.469033e-06, 2.524723e-06, 2.860909e-06, 2.209657e-06, 
    3.113162e-06, 2.378469e-06, 3.880757e-06, 2.408539e-06, 3.312185e-06,
  2.903798e-06, 2.788422e-06, 3.812464e-06, 5.01169e-06, 4.675556e-06, 
    3.669186e-06, 5.192468e-06, 4.419695e-06, 3.652569e-06, 3.383429e-06, 
    2.567854e-06, 3.121891e-06, 3.20144e-06, 3.498558e-06, 3.534756e-06,
  4.154317e-06, 4.042458e-06, 3.414911e-06, 4.008422e-06, 4.228785e-06, 
    4.349457e-06, 5.140919e-06, 4.269656e-06, 2.067988e-06, 2.760209e-06, 
    3.129758e-06, 2.655423e-06, 2.422845e-06, 1.918355e-06, 4.162683e-06,
  3.070725e-06, 4.419604e-06, 4.203509e-06, 4.997846e-06, 4.438048e-06, 
    5.962142e-06, 5.595128e-06, 5.383718e-06, 3.83857e-06, 2.291071e-06, 
    2.440804e-06, 2.60848e-06, 2.894044e-06, 2.134606e-06, 4.027778e-06,
  3.13073e-06, 2.700673e-06, 4.560205e-06, 4.520222e-06, 4.655943e-06, 
    5.941451e-06, 5.649164e-06, 5.634368e-06, 5.698383e-06, 4.612773e-06, 
    3.79501e-06, 3.74065e-06, 4.936323e-06, 1.980957e-06, 9.340527e-07,
  2.291355e-06, 2.525171e-06, 1.378538e-06, 3.902971e-06, 5.04941e-06, 
    6.564004e-06, 9.261215e-06, 8.157251e-06, 4.645413e-06, 3.879133e-06, 
    2.415778e-06, 2.962435e-06, 1.433513e-06, 6.840746e-07, 1.032731e-08,
  1.387897e-06, 1.036385e-06, 1.507908e-06, 1.518997e-06, 1.471515e-06, 
    2.766589e-06, 3.990427e-06, 6.962102e-06, 1.137916e-05, 7.22224e-06, 
    5.811185e-06, 3.412696e-06, 1.505886e-06, 1.216569e-06, 4.567588e-07,
  3.289526e-06, 2.103045e-06, 1.97834e-06, 2.043131e-06, 2.331117e-06, 
    2.060944e-06, 2.72739e-06, 3.117523e-06, 6.585014e-06, 1.422924e-05, 
    1.424206e-05, 1.367588e-05, 8.390079e-06, 4.07266e-06, 2.040731e-06,
  4.076866e-06, 4.234065e-06, 3.432669e-06, 4.493284e-06, 3.622461e-06, 
    1.729315e-06, 1.756602e-06, 3.28483e-06, 3.30824e-06, 3.932651e-06, 
    7.350908e-06, 8.770225e-06, 9.532269e-06, 5.202782e-06, 4.749863e-06,
  5.067576e-06, 4.549965e-06, 4.626452e-06, 5.216064e-06, 5.157265e-06, 
    4.015582e-06, 4.119388e-06, 2.496741e-06, 2.109748e-06, 3.07883e-06, 
    3.249624e-06, 3.398529e-06, 4.142978e-06, 5.391712e-06, 8.749035e-06,
  5.935557e-06, 7.205425e-06, 9.223444e-06, 6.392871e-06, 5.36351e-06, 
    6.665704e-06, 6.110109e-06, 5.085875e-06, 3.624047e-06, 2.84498e-06, 
    2.476175e-06, 3.133614e-06, 4.754195e-06, 5.831455e-06, 7.257571e-06,
  6.440592e-06, 7.797682e-06, 6.791531e-06, 8.087456e-06, 4.620395e-06, 
    5.040045e-06, 2.753061e-06, 3.64619e-06, 3.028218e-06, 2.554194e-06, 
    3.869203e-06, 5.159292e-06, 3.943683e-06, 5.22964e-06, 6.297071e-06,
  5.848639e-06, 8.62576e-06, 8.542861e-06, 7.581544e-06, 3.439614e-06, 
    2.009979e-06, 1.790374e-06, 1.18133e-06, 1.527706e-06, 3.927716e-06, 
    4.983256e-06, 1.846543e-06, 1.674956e-06, 3.741553e-06, 5.130901e-06,
  5.537864e-06, 7.36522e-06, 7.490105e-06, 8.481349e-06, 5.654576e-06, 
    1.497481e-06, 5.438124e-07, 8.367707e-07, 1.18004e-06, 1.291356e-06, 
    8.744462e-07, 2.983626e-06, 3.482045e-06, 2.437881e-06, 4.296878e-06,
  6.243548e-06, 7.464965e-06, 7.983506e-06, 7.836358e-06, 9.269041e-06, 
    4.609127e-06, 1.414003e-06, 1.744778e-06, 3.669838e-06, 2.869906e-06, 
    2.854668e-06, 2.360469e-06, 1.890016e-06, 2.996383e-06, 9.850738e-07,
  7.61723e-06, 6.511911e-06, 7.46469e-06, 1.241278e-05, 1.587951e-05, 
    1.603314e-05, 1.40852e-05, 1.967142e-05, 2.313747e-05, 1.214118e-05, 
    1.148418e-05, 9.352565e-06, 4.617554e-06, 2.134597e-06, 2.220193e-06,
  4.318534e-06, 8.240571e-06, 5.268038e-06, 5.479562e-06, 1.015755e-05, 
    1.609503e-05, 1.473914e-05, 1.725874e-05, 1.760131e-05, 1.728895e-05, 
    1.380125e-05, 9.418963e-06, 4.756525e-06, 2.209852e-06, 1.931859e-06,
  4.673951e-06, 2.684106e-06, 5.407977e-06, 8.51969e-06, 4.110774e-06, 
    4.160885e-06, 9.395437e-06, 1.366029e-05, 1.638558e-05, 1.345862e-05, 
    8.051472e-06, 4.178668e-06, 2.546544e-06, 2.982185e-06, 5.319901e-06,
  6.33246e-06, 5.644966e-06, 4.356851e-06, 6.187919e-06, 5.198268e-06, 
    1.007235e-05, 1.0142e-05, 1.451305e-05, 1.644485e-05, 1.217055e-05, 
    7.963797e-06, 4.857662e-06, 1.259565e-06, 4.447342e-06, 4.329248e-06,
  6.961178e-06, 5.372613e-06, 4.819726e-06, 1.179235e-05, 1.043954e-05, 
    1.080617e-05, 1.320698e-05, 1.316543e-05, 1.29538e-05, 6.178506e-06, 
    1.466479e-06, 1.245318e-06, 9.597392e-07, 8.450921e-07, 1.631524e-06,
  6.319323e-06, 6.470892e-06, 5.891779e-06, 7.807224e-06, 1.076914e-05, 
    1.052723e-05, 7.399226e-06, 4.69277e-06, 2.175274e-06, 6.496974e-07, 
    7.06017e-07, 4.729438e-07, 5.322957e-07, 6.089645e-07, 1.050612e-06,
  4.450777e-06, 4.913245e-06, 3.379833e-06, 1.024014e-05, 7.824576e-06, 
    5.835233e-06, 1.987278e-06, 6.024059e-07, 1.110036e-06, 2.626988e-07, 
    4.938547e-07, 8.592637e-07, 2.83965e-07, 4.472147e-07, 6.858269e-07,
  3.366589e-06, 3.484561e-06, 4.386196e-06, 6.218441e-06, 9.765348e-06, 
    5.727791e-06, 1.655743e-06, 5.683436e-07, 1.199189e-07, 1.433503e-07, 
    3.2195e-07, 1.13078e-06, 2.24362e-06, 1.007211e-06, 4.946706e-07,
  1.205285e-05, 8.696868e-06, 4.652456e-06, 2.82717e-06, 3.662342e-06, 
    2.720117e-06, 1.718802e-06, 9.535621e-07, 2.055158e-07, 1.787451e-08, 
    7.730689e-08, 1.586159e-07, 1.159427e-06, 7.955451e-07, 2.021477e-06,
  1.063161e-05, 1.895357e-05, 8.720301e-06, 4.160459e-06, 1.221705e-06, 
    6.716171e-06, 7.819942e-07, 3.729038e-07, 3.51896e-07, 1.915298e-07, 
    7.263585e-07, 1.148314e-06, 6.471888e-07, 3.155264e-07, 4.278541e-07,
  8.932241e-06, 2.076787e-05, 2.410935e-05, 1.41966e-05, 8.21044e-06, 
    1.01045e-05, 7.686404e-06, 8.072626e-06, 8.745675e-06, 9.900353e-06, 
    1.214977e-05, 1.429817e-05, 1.586949e-05, 1.508368e-05, 1.227563e-05,
  7.706491e-06, 2.067583e-05, 2.888958e-05, 2.480663e-05, 2.365338e-05, 
    1.421031e-05, 8.891036e-06, 6.61029e-06, 2.021397e-05, 3.186783e-05, 
    3.991112e-05, 4.825675e-05, 5.188057e-05, 3.122838e-05, 1.936137e-05,
  4.546875e-06, 7.616616e-06, 2.860022e-05, 3.66823e-05, 2.790461e-05, 
    2.585351e-05, 2.728483e-05, 3.549678e-05, 6.429957e-05, 0.0001101914, 
    0.0001536026, 0.000191853, 0.0001927193, 0.0001501396, 8.225112e-05,
  7.233812e-06, 2.232927e-05, 1.113865e-05, 1.573033e-05, 1.380378e-05, 
    1.194832e-05, 1.666604e-05, 2.488783e-05, 4.509641e-05, 8.871222e-05, 
    0.0001407181, 0.0001775744, 0.0001658599, 0.0001111984, 5.409882e-05,
  5.148825e-06, 6.792781e-06, 1.564553e-05, 1.53167e-05, 6.525408e-06, 
    5.892246e-06, 3.14879e-06, 4.474827e-06, 7.919636e-06, 1.118077e-05, 
    6.571461e-06, 3.338725e-06, 1.448147e-06, 4.831688e-07, 8.472186e-07,
  2.878721e-06, 3.578361e-06, 9.676773e-06, 1.624752e-05, 1.311722e-05, 
    9.575904e-06, 4.149055e-06, 3.249352e-06, 2.308505e-06, 2.324827e-06, 
    8.383437e-07, 1.582976e-06, 3.416879e-06, 2.320429e-06, 2.632479e-06,
  2.868241e-06, 1.617424e-06, 2.393476e-06, 8.479342e-06, 1.370762e-05, 
    1.653619e-05, 6.787755e-06, 4.160646e-06, 3.759331e-06, 2.295465e-06, 
    1.382452e-06, 1.438634e-06, 2.029978e-06, 2.363344e-06, 2.444182e-06,
  1.606552e-05, 4.368057e-06, 1.78858e-06, 3.698443e-06, 1.01786e-05, 
    1.244423e-05, 1.008576e-05, 7.732706e-06, 4.268201e-06, 3.278964e-06, 
    2.520392e-06, 1.710842e-06, 1.056001e-05, 2.634973e-05, 2.251342e-05,
  4.240882e-05, 3.366706e-05, 1.409464e-05, 1.623312e-06, 3.707994e-06, 
    9.396766e-06, 1.484988e-05, 9.774542e-06, 6.628328e-06, 1.70765e-05, 
    2.43565e-06, 1.289592e-05, 2.315366e-05, 4.949955e-06, 2.845394e-05,
  6.645545e-05, 3.841435e-05, 3.62381e-05, 1.600596e-05, 3.173165e-06, 
    4.273423e-06, 8.650803e-06, 2.212293e-05, 1.551887e-05, 3.89894e-06, 
    9.90723e-06, 9.662758e-06, 1.018972e-05, 2.602823e-06, 1.123143e-06,
  1.643377e-05, 1.387292e-05, 1.155135e-05, 1.060017e-05, 8.784519e-06, 
    8.192643e-06, 5.957228e-06, 6.300932e-06, 8.278118e-06, 7.953913e-06, 
    8.829464e-06, 1.224913e-05, 1.455221e-05, 1.432816e-05, 1.327884e-05,
  7.223351e-06, 4.671289e-06, 1.752977e-05, 9.508475e-06, 8.707752e-06, 
    6.571787e-06, 6.128745e-06, 6.151858e-06, 6.695098e-06, 8.94511e-06, 
    1.423953e-05, 1.941605e-05, 3.458502e-05, 3.55934e-05, 2.449853e-05,
  1.946151e-05, 1.220498e-05, 7.82704e-06, 1.373182e-05, 1.293154e-05, 
    7.154361e-06, 5.152649e-06, 8.619876e-06, 9.2178e-06, 1.158931e-05, 
    1.908285e-05, 4.736615e-05, 0.0001110801, 0.000174924, 0.0001963802,
  2.267975e-05, 2.273492e-05, 1.876733e-05, 6.029854e-06, 8.092113e-06, 
    4.654352e-06, 3.004803e-06, 7.443442e-06, 5.172023e-06, 3.435536e-06, 
    1.16556e-05, 5.112147e-05, 0.0001388504, 0.0002691007, 0.0003736411,
  2.900136e-06, 5.750888e-06, 1.889767e-05, 2.015694e-05, 1.756961e-05, 
    9.930224e-06, 4.984437e-06, 4.989259e-06, 5.200753e-06, 1.982289e-06, 
    4.533436e-06, 4.285459e-06, 2.41644e-05, 0.0001508411, 0.0003576937,
  1.543696e-06, 2.51222e-06, 9.607751e-06, 1.517109e-05, 2.584853e-05, 
    1.356367e-05, 1.274798e-05, 8.662449e-06, 3.778406e-06, 3.91306e-06, 
    2.623499e-06, 1.057738e-05, 1.24679e-05, 1.594538e-05, 0.0001703737,
  5.487628e-06, 1.494627e-06, 2.125802e-06, 6.309091e-06, 1.873999e-05, 
    2.25282e-05, 1.659344e-05, 9.429436e-06, 7.860461e-06, 8.416135e-06, 
    3.003588e-05, 2.659649e-05, 4.855704e-06, 1.748762e-05, 7.304124e-05,
  1.281145e-05, 3.760563e-06, 1.396762e-06, 3.685131e-06, 7.699389e-06, 
    1.595734e-05, 1.050785e-05, 1.084473e-05, 9.827678e-06, 2.532314e-05, 
    5.197645e-05, 4.026511e-05, 9.31859e-05, 5.233893e-05, 4.403915e-05,
  2.61807e-05, 1.4349e-05, 2.457644e-06, 1.155967e-06, 2.212176e-06, 
    8.676151e-06, 1.450882e-05, 2.124063e-05, 5.899798e-06, 3.913517e-05, 
    6.966564e-05, 6.343498e-05, 2.272446e-05, 4.742866e-05, 4.174905e-05,
  2.125371e-05, 1.730517e-05, 1.308686e-05, 1.065756e-06, 5.277038e-07, 
    2.915706e-06, 3.347613e-06, 2.851861e-05, 0.0001079065, 5.615899e-05, 
    4.76958e-05, 1.313686e-05, 2.980207e-05, 4.987397e-05, 4.59114e-05,
  5.082534e-05, 6.504639e-05, 8.813277e-05, 0.000102737, 0.0001219977, 
    0.000110151, 9.165535e-05, 4.414238e-05, 1.118987e-05, 6.477094e-06, 
    9.483998e-06, 7.772695e-06, 9.708053e-06, 1.321373e-05, 1.820056e-05,
  3.290856e-06, 1.675168e-05, 3.139976e-05, 4.653037e-05, 5.858426e-05, 
    5.186464e-05, 5.807509e-05, 3.679956e-05, 1.083751e-05, 2.460589e-06, 
    6.126209e-06, 8.062705e-06, 7.218882e-06, 1.338322e-05, 2.167641e-05,
  1.800203e-06, 4.757571e-06, 6.697331e-06, 1.133567e-05, 1.719637e-05, 
    2.004186e-05, 1.702004e-05, 1.149054e-05, 5.535397e-06, 5.793809e-07, 
    3.317864e-06, 8.935946e-06, 1.325782e-05, 1.258584e-05, 2.657056e-05,
  1.701636e-07, 6.75062e-07, 1.17739e-06, 2.655839e-06, 6.94357e-06, 
    1.099491e-05, 1.101287e-05, 2.895062e-06, 2.164561e-06, 9.135155e-07, 
    2.059503e-06, 6.249394e-06, 7.795655e-06, 1.083319e-05, 2.704318e-05,
  4.519011e-08, 2.898566e-07, 1.675007e-06, 3.893977e-06, 4.374633e-06, 
    9.327076e-06, 8.902532e-06, 3.624752e-06, 2.463838e-06, 2.202204e-06, 
    1.06462e-06, 2.017593e-06, 3.468396e-06, 4.202413e-06, 3.602367e-05,
  7.588752e-08, 1.608477e-07, 1.153427e-06, 2.428563e-06, 3.977648e-06, 
    9.157427e-06, 7.479746e-06, 3.369252e-06, 9.335807e-07, 5.387078e-06, 
    1.145444e-07, 1.297338e-06, 2.877118e-06, 7.181628e-06, 3.808411e-05,
  1.600657e-06, 1.013937e-06, 4.906519e-07, 9.210439e-07, 2.484479e-06, 
    5.318962e-06, 6.538933e-06, 1.922959e-06, 8.751279e-07, 6.2029e-07, 
    3.45338e-06, 1.164146e-05, 5.982651e-06, 7.254751e-06, 4.558953e-05,
  6.019333e-07, 4.085593e-07, 4.373197e-07, 1.264526e-06, 2.43707e-06, 
    2.294042e-06, 2.969139e-06, 2.602198e-06, 1.044349e-06, 1.233598e-05, 
    4.110789e-06, 3.431474e-06, 2.223407e-05, 1.497338e-05, 3.511242e-05,
  6.823491e-09, 4.883219e-07, 6.485882e-07, 7.941388e-07, 2.910312e-06, 
    1.066475e-06, 4.047949e-06, 1.423309e-06, 1.083004e-05, 1.505733e-05, 
    9.574264e-06, 2.418088e-05, 1.751469e-05, 2.465867e-05, 2.249106e-05,
  1.995209e-07, 4.997669e-07, 4.574616e-07, 5.214613e-07, 1.212249e-06, 
    1.038171e-06, 3.10034e-05, 4.510639e-06, 2.102784e-05, 4.466988e-06, 
    1.782007e-05, 1.393779e-05, 1.381932e-05, 1.651828e-05, 2.416292e-05,
  4.010522e-05, 6.747869e-05, 9.498018e-05, 0.0001381062, 0.0002090683, 
    0.0002982895, 0.000352463, 0.0003771211, 0.0003405609, 0.0002636426, 
    0.0002426287, 0.0002569184, 0.00026969, 0.0002766805, 0.0002901075,
  0.0001534348, 0.0001966763, 0.0002491311, 0.0003100906, 0.0003395541, 
    0.0003535991, 0.0003117237, 0.0002354091, 0.0001668206, 0.0001305895, 
    0.0001552204, 0.0002097036, 0.0002478652, 0.0002655619, 0.0002768275,
  0.0003206905, 0.0003624107, 0.0003855435, 0.000352566, 0.0003066192, 
    0.0002421769, 0.0001728185, 0.0001199476, 0.0001079381, 0.0001118806, 
    0.00013987, 0.0001735387, 0.0002084959, 0.0002219576, 0.0002053673,
  0.0004234968, 0.0004376419, 0.000398614, 0.0003132116, 0.0002420384, 
    0.0001867664, 0.0001494898, 0.0001328982, 0.0001274929, 0.0001439344, 
    0.0001686651, 0.0001759998, 0.0001856204, 0.000172454, 0.0001334779,
  0.0003895306, 0.0003938466, 0.0003288804, 0.0002700081, 0.0002468365, 
    0.0002135029, 0.000187505, 0.0001700812, 0.0001478557, 0.0001396509, 
    0.0001471428, 0.0001539452, 0.0001439189, 0.0001043484, 5.072378e-05,
  0.0002412321, 0.0002482629, 0.0002187831, 0.0002291796, 0.0002328313, 
    0.0002238342, 0.0002097384, 0.0001754943, 0.0001194299, 9.109981e-05, 
    9.877387e-05, 8.504467e-05, 5.485838e-05, 1.493566e-05, 1.45251e-07,
  5.425545e-05, 0.0001020674, 0.0001282494, 0.0001500401, 0.0001769561, 
    0.0001773812, 0.0001747976, 0.0001270737, 5.536267e-05, 4.808075e-05, 
    4.381689e-05, 2.509652e-05, 3.332501e-06, 4.936222e-06, 4.301805e-06,
  8.684045e-06, 3.443335e-05, 6.784687e-05, 8.294514e-05, 0.0001055933, 
    0.0001167457, 0.0001118446, 6.179881e-05, 1.86183e-05, 1.629636e-05, 
    1.040694e-05, 2.058305e-06, 7.141502e-06, 6.246978e-06, 1.014988e-05,
  7.310967e-06, 2.104238e-05, 2.806373e-05, 3.431933e-05, 5.248409e-05, 
    6.777094e-05, 6.108666e-05, 1.940149e-05, 8.897598e-06, 1.936986e-06, 
    1.298892e-06, 3.807995e-06, 6.585239e-06, 1.721327e-05, 2.294436e-05,
  7.878932e-06, 2.366774e-05, 2.288378e-05, 2.589466e-05, 2.823922e-05, 
    3.562742e-05, 2.95891e-05, 6.429926e-06, 1.03193e-05, 4.213872e-07, 
    2.697273e-06, 1.66988e-06, 6.76319e-06, 2.924847e-05, 1.819997e-05,
  7.332537e-06, 3.381754e-06, 1.116365e-06, 9.417548e-07, 7.283386e-07, 
    1.199918e-06, 4.838695e-06, 1.96497e-06, 7.276749e-07, 5.301439e-07, 
    1.473449e-06, 9.144582e-07, 5.930042e-07, 1.480736e-06, 1.08685e-06,
  2.865184e-06, 4.210412e-06, 5.968704e-06, 4.651846e-06, 4.96018e-06, 
    4.667914e-06, 5.472675e-06, 1.946724e-06, 7.596768e-07, 1.674144e-06, 
    2.196238e-06, 2.377035e-06, 2.404824e-06, 3.962788e-06, 8.939614e-06,
  5.875375e-06, 4.702879e-06, 4.638095e-06, 5.231725e-06, 3.673429e-06, 
    5.431873e-06, 4.403049e-06, 2.427276e-06, 1.829228e-06, 3.758473e-06, 
    4.806715e-06, 1.665611e-06, 4.921073e-06, 2.090545e-05, 6.113222e-05,
  8.03396e-06, 5.730383e-06, 8.555763e-06, 3.254155e-06, 2.03404e-06, 
    6.375749e-06, 4.244986e-06, 1.003367e-06, 1.679702e-06, 3.835445e-06, 
    6.220709e-06, 1.972232e-05, 5.626288e-05, 0.0001071572, 0.0001628671,
  6.933529e-06, 5.509893e-06, 7.046007e-06, 3.360114e-06, 3.244546e-06, 
    6.390487e-06, 1.841959e-06, 1.282878e-06, 8.443138e-06, 2.279404e-05, 
    4.754079e-05, 9.293624e-05, 0.0001488326, 0.0002172156, 0.0002720531,
  6.379299e-06, 7.118681e-06, 7.71968e-06, 5.896873e-06, 4.329057e-06, 
    5.503199e-06, 2.243078e-06, 1.455167e-05, 4.599524e-05, 5.337765e-05, 
    8.678518e-05, 0.0001581233, 0.0002304025, 0.0002840781, 0.0002943864,
  1.032038e-05, 5.867842e-06, 6.137132e-06, 7.352511e-06, 6.444891e-06, 
    6.358072e-06, 1.585625e-05, 6.400001e-05, 0.0001129603, 0.0001078019, 
    0.0001430482, 0.0002008893, 0.0002461363, 0.0002411491, 0.0002160274,
  6.476488e-06, 9.725045e-06, 6.903895e-06, 1.051154e-05, 9.453025e-06, 
    1.843847e-05, 4.929798e-05, 0.0001247472, 0.0001397575, 0.0001069811, 
    0.0001150025, 0.0001354327, 9.572837e-05, 6.126447e-05, 8.633077e-05,
  8.846148e-06, 9.085476e-06, 9.827052e-06, 1.788655e-05, 2.328637e-05, 
    3.117424e-05, 5.377003e-05, 9.112433e-05, 6.375977e-05, 8.004049e-05, 
    0.0001128778, 6.057723e-05, 4.787446e-05, 5.135691e-05, 8.039495e-05,
  1.006443e-05, 1.21668e-05, 1.248248e-05, 2.147833e-05, 3.544481e-05, 
    2.819769e-05, 5.029167e-05, 3.489205e-05, 5.506449e-05, 7.671565e-05, 
    3.844669e-05, 2.538146e-05, 3.06076e-05, 5.042434e-05, 2.384544e-05,
  7.333204e-09, 3.137094e-08, 7.129566e-08, 4.125289e-07, 4.330372e-07, 
    3.494424e-07, 1.464047e-08, 3.743689e-07, 6.289166e-07, 1.332951e-06, 
    4.048216e-07, 2.989104e-07, 2.391555e-06, 2.66282e-06, 2.477802e-06,
  9.031012e-07, 5.017882e-08, 3.4103e-08, 2.38041e-08, 6.691973e-08, 
    2.036552e-07, 7.142642e-08, 1.503228e-07, 2.342018e-07, 1.155856e-06, 
    1.502601e-06, 3.013569e-07, 6.587321e-07, 7.842611e-08, 1.009252e-06,
  3.991411e-06, 8.350818e-07, 7.033392e-07, 1.060405e-06, 1.383329e-06, 
    1.584045e-06, 6.779399e-07, 2.520546e-06, 6.164699e-06, 7.502837e-06, 
    4.541105e-06, 7.33175e-07, 3.204298e-07, 7.959353e-07, 2.670003e-06,
  5.547502e-06, 2.865007e-06, 4.743692e-07, 6.513453e-07, 1.146932e-06, 
    1.960992e-06, 2.908228e-06, 6.090511e-06, 7.520131e-06, 6.214144e-06, 
    4.463902e-06, 3.473811e-06, 4.196295e-06, 4.866355e-06, 4.786031e-06,
  2.653007e-06, 1.096293e-06, 7.06157e-07, 4.707524e-07, 6.154388e-07, 
    8.300267e-07, 2.636397e-06, 4.412746e-06, 3.53416e-06, 3.568853e-06, 
    3.827948e-06, 3.514356e-06, 3.746561e-06, 3.849477e-06, 4.117905e-06,
  4.285429e-06, 2.271031e-06, 2.120902e-06, 3.548606e-06, 4.826934e-06, 
    6.568647e-06, 8.350655e-06, 6.507387e-06, 2.827162e-06, 9.058099e-07, 
    1.095084e-06, 1.951553e-06, 3.523357e-06, 3.424092e-06, 5.704922e-06,
  5.78988e-06, 4.758351e-06, 6.991137e-06, 1.105036e-05, 1.25375e-05, 
    1.141966e-05, 1.408858e-05, 5.45073e-06, 4.430846e-06, 2.898886e-06, 
    2.66809e-06, 2.054968e-06, 2.474573e-06, 2.799517e-06, 5.80194e-06,
  8.232882e-06, 8.997887e-06, 1.613671e-05, 2.476754e-05, 2.174352e-05, 
    1.754636e-05, 1.401428e-05, 6.756717e-06, 5.449973e-06, 8.546901e-06, 
    1.027222e-05, 1.206321e-05, 1.286491e-05, 9.872079e-06, 1.654204e-05,
  2.309935e-05, 2.196531e-05, 3.182934e-05, 3.331452e-05, 2.154393e-05, 
    8.870151e-06, 4.761247e-06, 5.763475e-06, 2.601126e-05, 4.643833e-05, 
    3.575579e-05, 2.956898e-05, 2.80836e-05, 2.831097e-05, 2.802254e-05,
  3.736131e-05, 4.347171e-05, 5.163284e-05, 5.784749e-05, 5.92385e-05, 
    2.814467e-05, 1.871651e-05, 2.191805e-05, 4.816262e-05, 5.709744e-05, 
    5.957419e-05, 5.255993e-05, 4.318703e-05, 3.04946e-05, 4.205565e-05,
  2.023477e-06, 1.663702e-06, 2.988052e-06, 2.512289e-06, 1.648297e-06, 
    5.207527e-06, 5.293572e-06, 2.637962e-06, 3.166116e-06, 6.149734e-07, 
    1.802347e-06, 5.232295e-06, 3.666079e-06, 3.382312e-06, 4.205883e-06,
  4.051256e-07, 1.119596e-06, 3.507073e-06, 3.551964e-06, 6.341303e-06, 
    3.9615e-06, 3.495598e-06, 3.781084e-06, 3.600633e-06, 2.529529e-06, 
    2.61068e-06, 1.182727e-06, 1.117494e-06, 2.593914e-06, 3.422001e-06,
  5.067862e-06, 1.464887e-06, 2.811513e-06, 4.277556e-06, 4.497256e-06, 
    5.827972e-06, 5.696992e-06, 5.147689e-06, 5.27175e-06, 4.543854e-06, 
    4.601242e-06, 6.236031e-06, 5.643765e-06, 4.493764e-06, 4.029609e-06,
  8.649656e-06, 4.23997e-06, 3.07687e-06, 2.827707e-06, 1.671924e-06, 
    2.111857e-06, 3.167156e-06, 3.437823e-06, 4.23648e-06, 3.500124e-06, 
    2.364688e-06, 1.532599e-06, 1.141084e-06, 1.325852e-06, 2.134709e-06,
  5.30099e-06, 6.975704e-06, 4.324183e-06, 6.295334e-07, 3.596296e-08, 
    2.351053e-08, 8.308393e-08, 7.891362e-07, 2.070508e-06, 2.190322e-06, 
    2.28506e-06, 1.320304e-06, 1.622063e-06, 2.170877e-06, 2.636031e-06,
  5.577173e-06, 5.580035e-06, 6.540863e-06, 4.534784e-06, 3.977474e-06, 
    1.369569e-06, 2.174707e-06, 1.98082e-06, 1.397359e-06, 1.217091e-06, 
    2.120411e-06, 3.53277e-06, 3.511074e-06, 5.716885e-06, 4.365131e-06,
  6.278049e-06, 7.602992e-06, 8.859498e-06, 6.701965e-06, 2.643021e-06, 
    3.753194e-06, 2.887016e-06, 4.874954e-06, 5.332511e-06, 3.612164e-06, 
    3.875572e-06, 4.591281e-06, 5.932615e-06, 7.64561e-06, 7.836543e-06,
  4.814418e-06, 5.273279e-06, 5.15403e-06, 5.367946e-06, 4.340512e-06, 
    3.157724e-06, 3.660825e-06, 5.454986e-06, 5.877902e-06, 5.313566e-06, 
    3.773177e-06, 4.963969e-06, 5.474982e-06, 5.005862e-06, 6.159996e-06,
  1.10332e-05, 6.777158e-06, 5.384779e-06, 8.715391e-06, 5.896145e-06, 
    1.308079e-06, 1.629421e-06, 7.291703e-06, 9.375954e-06, 7.541954e-06, 
    8.208922e-06, 7.176397e-06, 6.53609e-06, 7.43746e-06, 7.205276e-06,
  1.159177e-05, 9.587729e-06, 5.404992e-06, 7.164157e-06, 7.12154e-06, 
    7.620936e-06, 7.026541e-06, 7.24197e-06, 9.670735e-06, 9.457976e-06, 
    1.015458e-05, 1.277068e-05, 1.651619e-05, 2.19514e-05, 1.393777e-05,
  3.455972e-06, 6.499237e-06, 7.023542e-06, 6.164505e-06, 5.170761e-06, 
    5.582608e-06, 5.0565e-06, 4.872429e-06, 4.665227e-06, 4.029147e-06, 
    3.751022e-06, 3.95841e-06, 5.850091e-06, 7.595479e-06, 6.214302e-06,
  2.717152e-06, 2.753927e-06, 3.830649e-06, 3.893323e-06, 3.256012e-06, 
    3.392867e-06, 2.670811e-06, 2.836765e-06, 2.653931e-06, 3.049655e-06, 
    2.919518e-06, 2.540715e-06, 2.362995e-06, 2.028952e-06, 3.741436e-06,
  2.311796e-06, 1.432961e-08, 2.985409e-08, 6.82744e-07, 6.899654e-07, 
    4.174267e-07, 9.463442e-07, 1.316976e-06, 2.18592e-06, 3.132716e-06, 
    1.838412e-06, 5.132534e-07, 1.515698e-07, 3.294255e-07, 1.237229e-06,
  1.947841e-06, 9.000687e-08, 1.912702e-07, 2.974295e-07, 1.204581e-06, 
    1.716492e-06, 2.745411e-06, 3.865794e-06, 2.671066e-06, 7.30406e-07, 
    9.433023e-08, 8.415895e-08, 4.723389e-07, 2.045163e-07, 9.53863e-08,
  2.446949e-06, 9.583525e-07, 1.887558e-06, 2.226226e-06, 8.037053e-06, 
    9.761231e-06, 7.72871e-06, 6.977901e-06, 5.647087e-06, 7.012831e-06, 
    6.814436e-06, 5.478511e-06, 6.681481e-06, 5.322873e-06, 3.401945e-06,
  3.027899e-06, 6.183413e-06, 5.489127e-06, 7.347819e-06, 1.058799e-05, 
    1.065877e-05, 1.026665e-05, 9.689034e-06, 7.368944e-06, 8.151806e-06, 
    7.478306e-06, 5.92921e-06, 6.154897e-06, 7.058934e-06, 5.932729e-06,
  2.392361e-06, 5.025496e-06, 5.463506e-06, 9.102378e-06, 8.658851e-06, 
    5.452624e-06, 4.812159e-06, 3.929215e-06, 3.625701e-06, 8.227129e-06, 
    8.707442e-06, 7.842174e-06, 8.109069e-06, 9.370951e-06, 9.882268e-06,
  3.43727e-06, 7.685165e-06, 7.648468e-06, 6.712175e-06, 9.81334e-06, 
    1.002484e-05, 3.500234e-06, 2.376378e-06, 4.631581e-06, 1.134672e-05, 
    3.363095e-05, 5.076524e-05, 5.711389e-05, 4.739228e-05, 4.687192e-05,
  6.019503e-06, 7.104388e-06, 5.847008e-06, 6.697711e-06, 5.857439e-06, 
    3.909572e-06, 1.733704e-06, 1.702773e-05, 3.5454e-05, 4.096966e-05, 
    4.242773e-05, 5.570694e-05, 8.327141e-05, 8.279502e-05, 7.631561e-05,
  6.111603e-06, 8.413059e-06, 9.404765e-06, 6.414118e-06, 5.230141e-06, 
    4.545773e-06, 1.038789e-05, 2.844668e-05, 2.784532e-05, 6.529821e-05, 
    7.083771e-05, 8.06256e-05, 0.0001059177, 0.0001208417, 9.247592e-05,
  2.583751e-06, 2.976965e-06, 4.543903e-06, 7.053095e-06, 7.011092e-06, 
    7.55044e-06, 6.376238e-06, 4.123135e-06, 4.180309e-06, 5.450667e-06, 
    5.45223e-06, 5.01621e-06, 9.678258e-06, 7.670542e-06, 8.877389e-06,
  1.621198e-06, 2.073321e-06, 2.28399e-06, 3.201793e-06, 4.296608e-06, 
    4.294636e-06, 5.962943e-06, 5.109148e-06, 4.420328e-06, 4.566923e-06, 
    3.830352e-06, 4.598908e-06, 7.612972e-06, 7.18666e-06, 9.085476e-06,
  1.478079e-06, 1.836906e-06, 1.021442e-06, 3.330532e-06, 1.908452e-06, 
    1.055984e-06, 2.530279e-06, 4.890785e-06, 6.632388e-06, 6.720332e-06, 
    6.839669e-06, 6.165718e-06, 4.576291e-06, 4.795272e-06, 4.026358e-06,
  4.884365e-06, 7.610502e-06, 9.691563e-06, 7.503159e-06, 8.227445e-06, 
    8.831496e-06, 9.618258e-06, 8.323373e-06, 8.896837e-06, 5.300188e-06, 
    4.282315e-06, 3.341942e-06, 3.971264e-06, 2.533446e-06, 1.37503e-07,
  9.580154e-06, 9.375705e-06, 1.080923e-05, 1.285428e-05, 1.085448e-05, 
    8.542863e-06, 8.011191e-06, 5.911495e-06, 5.145023e-06, 4.337797e-06, 
    5.603229e-06, 4.380795e-06, 4.553747e-06, 2.292412e-06, 3.941269e-07,
  1.068792e-05, 1.043928e-05, 1.101552e-05, 1.185269e-05, 1.140973e-05, 
    7.865683e-06, 6.168646e-06, 3.790629e-06, 4.084e-06, 3.967548e-06, 
    3.645777e-06, 4.940337e-06, 5.74898e-06, 4.237946e-06, 4.558518e-06,
  1.036238e-05, 1.268428e-05, 1.185829e-05, 1.202748e-05, 1.148465e-05, 
    5.579554e-06, 1.906001e-06, 2.700618e-06, 4.52852e-06, 1.102996e-05, 
    1.585764e-05, 1.954879e-05, 1.673004e-05, 1.578884e-05, 1.726921e-05,
  1.322319e-05, 1.234783e-05, 1.14485e-05, 8.568855e-06, 6.460053e-06, 
    8.102507e-06, 2.81333e-06, 5.731771e-06, 2.332326e-05, 4.587398e-05, 
    6.974202e-05, 5.38279e-05, 6.374258e-05, 6.028296e-05, 7.316242e-05,
  1.306847e-05, 1.09735e-05, 7.084423e-06, 8.22426e-06, 1.523548e-05, 
    1.827738e-05, 1.943064e-05, 3.669648e-05, 5.773031e-05, 6.821279e-05, 
    7.893142e-05, 6.0372e-05, 6.499292e-05, 5.654784e-05, 6.34025e-05,
  1.833155e-05, 1.285399e-05, 9.344235e-06, 1.044988e-05, 1.816985e-05, 
    1.151104e-05, 5.517213e-05, 6.232603e-05, 0.0001362691, 0.0002021214, 
    0.0001812033, 0.0001227272, 9.885718e-05, 6.379807e-05, 8.313889e-05,
  3.157607e-06, 5.700844e-06, 4.725086e-06, 7.215874e-06, 8.414465e-06, 
    6.691708e-06, 5.192794e-06, 4.365979e-06, 6.074831e-06, 8.72173e-06, 
    4.772482e-06, 8.717792e-06, 6.973685e-06, 3.072653e-06, 2.303431e-06,
  4.2759e-06, 6.052809e-06, 5.295376e-06, 2.463948e-06, 3.89893e-06, 
    3.573184e-06, 4.419326e-06, 4.894222e-06, 7.435851e-06, 6.364716e-06, 
    5.986902e-06, 7.842933e-06, 6.812602e-06, 4.422712e-06, 4.862766e-06,
  7.352158e-06, 8.2088e-06, 6.113616e-06, 6.174455e-06, 5.152474e-06, 
    2.75289e-06, 4.276678e-06, 5.043068e-06, 3.853964e-06, 5.714559e-06, 
    6.835654e-06, 6.413467e-06, 6.359159e-06, 7.260526e-06, 3.376209e-06,
  6.284667e-06, 6.767015e-06, 4.950792e-06, 4.256423e-06, 5.290879e-06, 
    3.4769e-06, 3.233169e-06, 4.612011e-06, 5.724199e-06, 6.078406e-06, 
    7.049123e-06, 9.630575e-06, 7.543908e-06, 5.332477e-06, 4.767456e-06,
  2.62854e-06, 2.620334e-06, 2.433693e-06, 3.03557e-06, 3.640592e-06, 
    3.600391e-06, 4.170066e-06, 3.550839e-06, 3.328779e-06, 1.81457e-06, 
    2.185374e-06, 2.359395e-06, 3.848923e-06, 4.178181e-06, 2.907122e-06,
  2.222966e-06, 2.812919e-06, 1.398345e-06, 2.457284e-06, 2.253018e-06, 
    1.289909e-06, 1.658205e-06, 2.030954e-06, 2.417232e-06, 1.755567e-06, 
    2.850319e-06, 3.597091e-06, 2.039263e-06, 1.689134e-06, 4.27068e-07,
  2.176668e-06, 8.628776e-07, 1.218306e-06, 1.199707e-06, 9.449476e-07, 
    6.952668e-07, 7.333768e-07, 2.817004e-07, 1.010186e-06, 2.268239e-06, 
    3.408286e-06, 3.116467e-06, 6.187828e-06, 6.773614e-06, 6.09196e-06,
  3.000435e-06, 1.506728e-06, 1.341965e-06, 1.472324e-06, 8.013259e-07, 
    1.377094e-06, 1.423788e-06, 2.995745e-06, 4.981954e-06, 7.461275e-06, 
    7.869334e-06, 7.27115e-06, 7.11046e-06, 8.999466e-06, 1.306504e-05,
  4.339995e-06, 2.174601e-06, 1.308569e-06, 1.534457e-06, 1.68284e-06, 
    1.539897e-06, 2.767287e-06, 5.288043e-06, 7.901292e-06, 9.487318e-06, 
    9.114339e-06, 1.064137e-05, 9.357165e-06, 8.469495e-06, 7.076113e-06,
  3.889835e-06, 2.06338e-06, 2.858917e-06, 4.227794e-06, 7.361222e-06, 
    3.373164e-06, 4.126846e-06, 1.132643e-05, 1.014347e-05, 1.187232e-05, 
    1.120715e-05, 1.217079e-05, 1.243138e-05, 1.04105e-05, 7.606576e-06,
  5.439868e-06, 8.855342e-06, 1.126686e-05, 1.458566e-05, 1.92123e-05, 
    1.810398e-05, 1.298357e-05, 1.030779e-05, 7.892441e-06, 8.502158e-06, 
    9.53469e-06, 7.944102e-06, 6.861838e-06, 4.02699e-06, 6.389038e-06,
  1.013966e-05, 9.341235e-06, 1.174858e-05, 1.199087e-05, 9.464099e-06, 
    6.714753e-06, 3.094015e-06, 4.449714e-06, 7.026676e-06, 6.054275e-06, 
    6.8892e-06, 8.078264e-06, 9.712548e-06, 9.621376e-06, 1.047777e-05,
  1.075645e-05, 6.784667e-06, 7.198918e-06, 4.650461e-06, 4.480353e-06, 
    8.543011e-06, 3.800768e-06, 5.436053e-06, 3.595257e-06, 6.240498e-06, 
    1.021717e-05, 2.240102e-05, 3.98432e-05, 5.785693e-05, 6.572685e-05,
  5.51991e-06, 1.368539e-06, 1.585903e-06, 1.904658e-06, 3.476219e-06, 
    6.627662e-06, 5.900545e-06, 5.094648e-06, 1.422721e-05, 2.553683e-05, 
    3.55364e-05, 4.195981e-05, 4.728271e-05, 5.092111e-05, 4.913398e-05,
  2.412451e-06, 1.419003e-06, 6.287715e-07, 1.07811e-06, 1.675965e-06, 
    1.647167e-06, 7.236569e-06, 1.50869e-05, 2.343595e-05, 2.673999e-05, 
    1.764493e-05, 1.253508e-05, 6.050757e-06, 3.379545e-06, 1.809952e-06,
  1.020911e-06, 7.854711e-07, 2.085562e-07, 7.437542e-07, 3.283672e-06, 
    1.10216e-05, 1.889226e-05, 1.783806e-05, 1.554723e-05, 1.336231e-05, 
    9.31893e-06, 4.500979e-06, 8.194273e-07, 2.927264e-07, 2.158742e-07,
  4.626515e-07, 3.004957e-07, 3.411408e-07, 2.45982e-06, 9.407048e-06, 
    1.562132e-05, 1.697494e-05, 1.702585e-05, 1.984866e-05, 2.316078e-05, 
    1.676727e-05, 6.370075e-06, 2.738506e-06, 1.306898e-06, 1.412118e-06,
  1.948422e-07, 7.748939e-07, 2.753833e-06, 7.976183e-06, 1.191705e-05, 
    2.282814e-05, 4.173294e-05, 3.576958e-05, 2.270425e-05, 2.479822e-05, 
    2.456944e-05, 9.375455e-06, 5.610581e-06, 2.09228e-06, 1.090292e-06,
  4.529196e-07, 2.514102e-06, 1.065507e-05, 1.435954e-05, 1.587357e-05, 
    4.452703e-05, 6.355412e-05, 5.271056e-05, 2.802021e-05, 8.624877e-06, 
    1.187226e-05, 1.007037e-05, 2.037077e-05, 1.521971e-05, 3.997815e-06,
  8.055714e-07, 4.336668e-06, 1.99826e-05, 2.613356e-05, 3.012397e-05, 
    4.652132e-05, 6.008018e-05, 5.744547e-05, 6.246613e-05, 6.819041e-05, 
    7.777766e-05, 3.940214e-05, 1.055666e-05, 1.309719e-05, 1.218214e-05,
  2.406912e-06, 1.0965e-06, 1.085247e-06, 1.107416e-06, 1.368297e-06, 
    1.664485e-06, 3.239507e-06, 2.486492e-06, 2.404842e-06, 1.646356e-06, 
    3.157274e-06, 3.604875e-06, 2.918968e-06, 4.343706e-06, 4.964499e-06,
  4.261814e-06, 5.253751e-06, 3.765589e-06, 2.445174e-06, 8.164626e-07, 
    2.071869e-06, 3.897054e-06, 4.043133e-06, 4.537012e-06, 2.672613e-06, 
    2.746205e-06, 1.382975e-06, 1.527345e-06, 1.882865e-06, 2.293591e-06,
  3.594394e-06, 9.599464e-06, 8.10063e-06, 6.246743e-06, 5.412772e-06, 
    3.834096e-06, 3.072325e-06, 1.966595e-06, 1.444285e-06, 1.020123e-06, 
    3.390055e-06, 7.512818e-06, 1.314155e-05, 2.854878e-05, 4.756615e-05,
  4.532838e-06, 4.41353e-06, 4.359783e-06, 5.180115e-06, 5.929477e-06, 
    4.033428e-06, 2.700611e-06, 1.783638e-06, 3.147933e-06, 1.120993e-05, 
    2.745202e-05, 4.304231e-05, 5.828165e-05, 8.488847e-05, 0.0001006932,
  5.202935e-06, 3.60883e-06, 2.990964e-06, 3.167749e-06, 4.994388e-06, 
    2.019408e-06, 2.937263e-06, 5.073132e-06, 1.377301e-05, 2.937425e-05, 
    4.217456e-05, 5.341364e-05, 5.645003e-05, 6.039907e-05, 6.098163e-05,
  4.506553e-06, 4.127325e-06, 2.534031e-06, 4.931804e-06, 3.430478e-06, 
    3.725085e-06, 2.996724e-06, 5.898009e-06, 1.528537e-05, 2.362639e-05, 
    3.553263e-05, 4.112059e-05, 4.204666e-05, 6.108332e-05, 7.784949e-05,
  3.394148e-06, 1.626581e-06, 1.591531e-06, 2.019356e-06, 1.998568e-06, 
    2.31058e-06, 5.922321e-06, 1.052802e-05, 1.262783e-05, 1.607886e-05, 
    1.889163e-05, 8.505624e-06, 5.786737e-06, 9.801833e-06, 3.699675e-05,
  9.243876e-07, 8.11409e-07, 1.716872e-06, 2.573645e-06, 1.824017e-06, 
    3.600013e-06, 5.686548e-06, 8.946773e-06, 2.510657e-05, 7.421825e-05, 
    0.0001203506, 9.180699e-05, 2.517014e-05, 2.095946e-05, 1.907804e-05,
  5.930057e-07, 9.25187e-07, 3.382644e-06, 2.966752e-06, 3.083341e-06, 
    6.852279e-06, 7.098585e-06, 1.141069e-05, 4.356681e-05, 0.0002291588, 
    0.0004694401, 0.0004665305, 0.0002015999, 4.437624e-05, 2.691674e-05,
  3.399654e-08, 1.400832e-06, 5.984601e-06, 6.496148e-06, 1.106365e-05, 
    9.712066e-06, 1.324521e-05, 1.578239e-05, 8.706553e-05, 0.0003387364, 
    0.0007494229, 0.0008615546, 0.0005297232, 0.0001197055, 3.503908e-05,
  1.143784e-05, 1.598652e-05, 1.435012e-05, 1.693886e-05, 1.453603e-05, 
    1.493287e-05, 1.246557e-05, 2.05568e-05, 4.049818e-05, 6.561729e-05, 
    0.0001088985, 0.000174121, 0.0002851328, 0.0004128664, 0.0004958053,
  5.72837e-06, 7.405589e-06, 5.350485e-06, 7.60132e-06, 8.31605e-06, 
    7.666954e-06, 1.702957e-05, 3.25758e-05, 5.152285e-05, 8.631575e-05, 
    0.0001361052, 0.0002086349, 0.0002934667, 0.0003619361, 0.0003976989,
  5.362358e-06, 5.690497e-06, 5.347651e-06, 5.66545e-06, 4.810086e-06, 
    8.827737e-06, 2.21796e-05, 4.771454e-05, 6.740833e-05, 8.90662e-05, 
    0.000124441, 0.0001552075, 0.0001688813, 0.0001787302, 0.0001603059,
  5.645558e-06, 3.909362e-06, 2.774442e-06, 3.928902e-06, 3.863308e-06, 
    9.753382e-06, 2.512378e-05, 4.058318e-05, 5.394593e-05, 6.376519e-05, 
    6.107196e-05, 5.094402e-05, 4.779173e-05, 4.504027e-05, 4.545204e-05,
  6.026294e-06, 3.773258e-06, 3.120807e-06, 5.505493e-06, 5.631812e-06, 
    1.299737e-05, 2.451817e-05, 3.593501e-05, 4.469546e-05, 4.829498e-05, 
    4.776795e-05, 3.656838e-05, 2.429992e-05, 1.405868e-05, 1.525752e-05,
  3.60416e-06, 4.091929e-06, 2.77042e-06, 4.3777e-06, 5.493191e-06, 
    1.472695e-05, 2.562536e-05, 3.925466e-05, 4.436142e-05, 4.57224e-05, 
    4.00821e-05, 2.791742e-05, 1.435368e-05, 8.417415e-06, 1.100972e-05,
  3.063069e-06, 3.919124e-06, 4.186549e-06, 5.823415e-06, 6.930447e-06, 
    1.64772e-05, 3.20534e-05, 4.759285e-05, 4.949493e-05, 4.412626e-05, 
    2.696164e-05, 2.208737e-05, 1.63821e-05, 8.55812e-06, 7.142624e-06,
  3.146907e-06, 4.862762e-06, 8.157665e-06, 6.100464e-06, 8.08656e-06, 
    1.923544e-05, 3.594777e-05, 4.886758e-05, 4.547529e-05, 3.369476e-05, 
    1.913449e-05, 1.069311e-05, 8.983123e-06, 5.958453e-06, 4.249048e-06,
  4.105195e-06, 7.198158e-06, 5.245512e-06, 5.403508e-06, 9.524646e-06, 
    2.333218e-05, 3.706417e-05, 4.305624e-05, 3.508295e-05, 3.130264e-05, 
    1.899457e-05, 9.485692e-06, 4.227507e-06, 1.526687e-06, 2.37847e-06,
  7.128162e-06, 9.429471e-06, 7.005548e-06, 7.198354e-06, 1.50706e-05, 
    3.221184e-05, 4.256994e-05, 3.914119e-05, 3.288988e-05, 3.687212e-05, 
    2.057844e-05, 3.455021e-06, 1.340688e-06, 4.639435e-07, 1.520793e-06,
  6.049765e-07, 1.390937e-06, 1.394888e-06, 2.24173e-06, 3.339808e-06, 
    2.205262e-06, 1.16799e-06, 1.400762e-06, 2.072909e-06, 3.88054e-06, 
    5.336513e-06, 5.346296e-06, 5.623856e-06, 6.302427e-06, 8.519866e-06,
  1.292306e-06, 1.014918e-06, 1.459553e-06, 2.58172e-06, 3.14843e-06, 
    2.497019e-06, 1.842701e-06, 1.163122e-06, 1.623138e-06, 3.213128e-06, 
    3.426168e-06, 5.291515e-06, 4.761137e-06, 6.061996e-06, 8.503741e-06,
  1.004128e-06, 1.795408e-06, 1.335682e-06, 1.441566e-06, 2.022673e-06, 
    2.03362e-06, 1.877462e-06, 1.039102e-06, 1.24325e-06, 2.129621e-06, 
    2.510708e-06, 4.540344e-06, 5.43537e-06, 5.299519e-06, 1.986953e-05,
  9.639909e-07, 1.669068e-06, 8.386971e-07, 1.055065e-06, 1.575249e-06, 
    2.027989e-06, 1.575559e-06, 8.823953e-07, 1.558176e-06, 2.457056e-06, 
    2.034392e-06, 2.930218e-06, 1.19052e-05, 3.128527e-05, 5.164278e-05,
  2.279133e-06, 2.518767e-06, 6.033852e-07, 6.059196e-07, 1.778473e-06, 
    2.962331e-06, 2.90384e-06, 2.083631e-06, 1.638261e-06, 1.645112e-06, 
    3.452547e-06, 1.938923e-05, 4.145661e-05, 6.785737e-05, 7.863541e-05,
  2.333257e-06, 3.201312e-06, 2.882759e-06, 2.185787e-06, 2.901313e-06, 
    3.682017e-06, 3.915437e-06, 2.265466e-06, 1.374992e-06, 2.993376e-06, 
    2.086993e-05, 4.634975e-05, 7.03072e-05, 8.899303e-05, 0.0001091009,
  2.353941e-06, 3.69066e-06, 5.341888e-06, 5.450075e-06, 4.299225e-06, 
    3.825243e-06, 3.673053e-06, 3.327876e-06, 3.941841e-06, 2.122792e-05, 
    4.401699e-05, 6.975332e-05, 9.956209e-05, 0.0001242583, 0.0001402544,
  2.320482e-06, 3.886761e-06, 2.659908e-06, 5.350795e-06, 4.215605e-06, 
    4.213675e-06, 3.75817e-06, 2.990573e-06, 9.78577e-06, 3.267036e-05, 
    6.525064e-05, 9.550957e-05, 0.0001515296, 0.000228799, 0.0002551248,
  3.89301e-06, 6.297395e-06, 5.354314e-06, 5.511091e-06, 3.564896e-06, 
    3.639087e-06, 1.613433e-06, 4.225908e-06, 1.22505e-05, 3.809369e-05, 
    8.442954e-05, 0.0001528897, 0.0002645351, 0.0003471486, 0.0004082465,
  4.509698e-06, 5.47673e-06, 6.679255e-06, 5.695659e-06, 3.352674e-06, 
    2.048678e-06, 2.336194e-06, 5.404255e-06, 1.223414e-05, 4.593422e-05, 
    0.0001341595, 0.0002420138, 0.0003585831, 0.0004387464, 0.0004731717,
  3.072615e-06, 4.676198e-06, 5.269377e-06, 5.898785e-06, 6.845051e-06, 
    6.784549e-06, 6.14047e-06, 4.603755e-06, 5.869223e-06, 7.341692e-06, 
    8.302857e-06, 1.036999e-05, 9.458437e-06, 1.346437e-05, 1.420424e-05,
  2.941059e-06, 4.249031e-06, 3.959595e-06, 4.161119e-06, 2.57492e-06, 
    7.359639e-06, 6.397748e-06, 5.020144e-06, 6.18935e-06, 5.471056e-06, 
    7.59734e-06, 9.415584e-06, 9.706295e-06, 9.717853e-06, 9.186883e-06,
  3.55585e-06, 5.35672e-06, 6.468162e-06, 5.13137e-06, 4.781821e-06, 
    5.205781e-06, 4.709032e-06, 4.59039e-06, 6.644464e-06, 5.670938e-06, 
    6.135886e-06, 7.187745e-06, 9.698248e-06, 8.709967e-06, 7.013601e-06,
  3.430596e-06, 4.348559e-06, 4.826135e-06, 5.218056e-06, 3.314326e-06, 
    5.13179e-06, 3.848696e-06, 4.671788e-06, 6.49533e-06, 5.688044e-06, 
    3.334222e-06, 4.050759e-06, 6.883997e-06, 8.954213e-06, 1.139824e-05,
  3.084512e-06, 3.527292e-06, 4.419001e-06, 4.946641e-06, 3.769441e-06, 
    3.001377e-06, 5.002955e-06, 6.394012e-06, 5.253291e-06, 3.752839e-06, 
    4.009469e-06, 4.55342e-06, 6.175185e-06, 6.077939e-06, 4.797304e-06,
  4.996024e-06, 4.386506e-06, 4.835686e-06, 4.704207e-06, 5.417976e-06, 
    3.557651e-06, 3.153135e-06, 5.907878e-06, 6.563255e-06, 7.277268e-06, 
    5.982267e-06, 5.303364e-06, 5.722529e-06, 3.803161e-06, 3.991856e-06,
  4.518338e-06, 4.2751e-06, 3.173932e-06, 4.563257e-06, 6.067931e-06, 
    6.452603e-06, 5.423707e-06, 4.347241e-06, 4.596322e-06, 5.654962e-06, 
    5.833846e-06, 5.096939e-06, 4.170274e-06, 2.760978e-06, 5.717662e-06,
  7.231341e-06, 7.514349e-06, 6.785072e-06, 5.166136e-06, 6.413695e-06, 
    7.590475e-06, 4.270516e-06, 3.446752e-06, 3.760937e-06, 6.747053e-06, 
    3.689224e-06, 4.192744e-06, 5.511819e-06, 5.640487e-06, 8.661571e-06,
  5.700846e-06, 6.153948e-06, 5.502191e-06, 6.59857e-06, 7.488233e-06, 
    8.404937e-06, 6.896328e-06, 5.156804e-06, 4.332207e-06, 1.969929e-06, 
    1.81881e-06, 1.541979e-06, 6.091349e-06, 6.811957e-06, 5.045621e-06,
  4.179932e-06, 5.579379e-06, 6.165789e-06, 6.71201e-06, 8.168299e-06, 
    5.814492e-06, 5.111498e-06, 7.56027e-06, 3.476979e-06, 3.516213e-06, 
    2.429994e-06, 3.643981e-06, 5.845196e-06, 4.680679e-06, 5.792524e-06,
  5.967236e-06, 6.402415e-06, 8.253473e-06, 8.491908e-06, 8.867265e-06, 
    8.230955e-06, 7.18234e-06, 7.685213e-06, 4.57851e-06, 3.177455e-06, 
    3.482645e-06, 5.748726e-06, 8.909317e-06, 9.001858e-06, 8.389276e-06,
  6.995986e-06, 5.665037e-06, 5.665759e-06, 4.304638e-06, 5.903971e-06, 
    6.168084e-06, 7.26407e-06, 7.269201e-06, 6.068055e-06, 4.958169e-06, 
    2.940284e-06, 3.987955e-06, 3.874903e-06, 3.772791e-06, 8.022564e-06,
  1.093225e-05, 9.738228e-06, 4.014161e-06, 4.758469e-06, 4.760091e-06, 
    7.28827e-06, 7.77236e-06, 4.060428e-06, 4.424202e-06, 5.014933e-06, 
    2.899295e-06, 2.531756e-06, 2.117206e-06, 4.780377e-06, 4.768581e-06,
  8.650034e-06, 8.058464e-06, 8.36479e-06, 5.275992e-06, 3.444528e-06, 
    3.037026e-06, 7.17414e-06, 8.657036e-06, 4.308141e-06, 3.524271e-06, 
    3.250126e-06, 2.891296e-06, 2.518857e-06, 4.149279e-06, 2.771478e-06,
  7.407575e-06, 5.947658e-06, 3.948222e-06, 3.971358e-06, 8.261707e-06, 
    6.377216e-06, 5.289217e-06, 6.385316e-06, 6.492201e-06, 3.580905e-06, 
    3.815014e-06, 4.958819e-06, 3.772513e-06, 2.000728e-06, 2.036209e-06,
  1.026048e-05, 5.926483e-06, 6.77837e-06, 4.92994e-06, 5.621371e-06, 
    6.748419e-06, 7.005809e-06, 4.503592e-06, 6.472852e-06, 4.476813e-06, 
    4.18438e-06, 5.015449e-06, 4.347705e-06, 2.611873e-06, 2.762413e-06,
  8.913586e-06, 5.786379e-06, 6.493459e-06, 9.297435e-06, 4.364334e-06, 
    3.774612e-06, 4.473132e-06, 3.733877e-06, 3.909365e-06, 3.569611e-06, 
    5.378645e-06, 7.678704e-06, 5.651851e-06, 2.176341e-06, 2.740234e-06,
  9.691395e-06, 8.116567e-06, 8.371769e-06, 7.594139e-06, 9.895105e-06, 
    8.915956e-06, 5.930887e-06, 5.299008e-06, 2.85293e-06, 4.465675e-06, 
    3.689495e-06, 5.910227e-06, 3.675175e-06, 2.333578e-06, 2.867476e-06,
  6.531622e-06, 7.951622e-06, 6.976442e-06, 7.859043e-06, 5.484825e-06, 
    3.791517e-06, 5.500928e-06, 3.175041e-06, 3.273403e-06, 5.812366e-06, 
    7.611578e-06, 2.60505e-06, 4.042869e-06, 4.514663e-06, 4.062684e-06,
  6.221539e-06, 7.023457e-06, 5.062619e-06, 6.951003e-06, 6.207313e-06, 
    4.93845e-06, 5.1822e-06, 4.567063e-06, 3.260526e-06, 4.287406e-06, 
    5.588241e-06, 2.122696e-06, 1.818995e-06, 4.086591e-06, 5.344914e-06,
  8.78482e-06, 7.817701e-06, 7.395057e-06, 6.674237e-06, 6.831603e-06, 
    4.666056e-06, 4.315556e-06, 3.44693e-06, 4.044396e-06, 5.110695e-06, 
    8.143575e-06, 1.196527e-05, 9.928032e-06, 8.741563e-06, 7.453452e-06,
  9.881343e-06, 1.02702e-05, 8.791287e-06, 7.286018e-06, 6.617579e-06, 
    1.043326e-05, 8.601308e-06, 6.102122e-06, 4.996383e-06, 3.315896e-06, 
    3.776964e-06, 5.149773e-06, 5.741027e-06, 8.289649e-06, 7.625358e-06,
  7.198835e-06, 1.043437e-05, 8.785251e-06, 7.53961e-06, 8.428705e-06, 
    1.121962e-05, 1.349316e-05, 8.094881e-06, 6.770821e-06, 6.366984e-06, 
    2.710208e-06, 3.257419e-06, 4.205067e-06, 4.318496e-06, 4.204282e-06,
  7.856767e-06, 8.828667e-06, 9.877476e-06, 1.197893e-05, 9.679889e-06, 
    1.112463e-05, 1.320949e-05, 1.26838e-05, 1.101173e-05, 6.818924e-06, 
    2.831151e-06, 2.554941e-06, 4.305621e-06, 3.122391e-06, 3.986181e-06,
  9.665468e-06, 1.04851e-05, 1.123874e-05, 1.229766e-05, 1.046869e-05, 
    1.046383e-05, 7.838918e-06, 8.532439e-06, 6.461687e-06, 7.620931e-06, 
    6.935326e-06, 4.541901e-06, 2.402898e-06, 4.216642e-06, 3.176222e-06,
  1.06778e-05, 1.121307e-05, 1.164687e-05, 1.087145e-05, 1.004368e-05, 
    9.330303e-06, 8.376752e-06, 7.044953e-06, 7.045725e-06, 6.473223e-06, 
    4.622349e-06, 1.941953e-06, 5.02687e-06, 6.049779e-06, 4.241228e-06,
  9.429277e-06, 1.071078e-05, 1.148988e-05, 9.522671e-06, 1.067885e-05, 
    9.446507e-06, 7.508012e-06, 7.625801e-06, 6.072631e-06, 5.107918e-06, 
    4.850919e-06, 4.783091e-06, 5.05267e-06, 4.822761e-06, 5.115382e-06,
  9.860087e-06, 1.019663e-05, 9.146068e-06, 8.160735e-06, 8.74035e-06, 
    7.898581e-06, 8.133836e-06, 6.548226e-06, 5.427695e-06, 6.573414e-06, 
    6.735362e-06, 5.151099e-06, 6.465383e-06, 7.232948e-06, 5.597445e-06,
  8.823084e-06, 6.820356e-06, 7.061764e-06, 6.685079e-06, 7.277341e-06, 
    6.377537e-06, 5.282277e-06, 4.922219e-06, 3.996606e-06, 4.576236e-06, 
    5.623521e-06, 6.371578e-06, 6.176864e-06, 6.063716e-06, 6.343316e-06,
  9.059364e-06, 6.827791e-06, 5.502194e-06, 6.489353e-06, 4.824562e-06, 
    4.067703e-06, 5.147235e-06, 4.935228e-06, 5.54931e-06, 5.797174e-06, 
    6.908917e-06, 5.558373e-06, 5.086318e-06, 4.590405e-06, 4.528877e-06,
  9.249252e-06, 2.140278e-05, 4.002299e-05, 5.98201e-05, 8.639479e-05, 
    9.577999e-05, 8.423688e-05, 6.093322e-05, 6.590183e-05, 6.703581e-05, 
    4.726697e-05, 2.946073e-05, 1.691578e-05, 1.389495e-05, 1.205982e-05,
  4.884336e-06, 7.354794e-06, 1.902396e-05, 4.471792e-05, 6.732965e-05, 
    8.096966e-05, 7.637076e-05, 5.8799e-05, 3.557049e-05, 2.007581e-05, 
    1.089798e-05, 8.344809e-06, 7.901792e-06, 8.362355e-06, 8.051176e-06,
  4.343668e-06, 7.756457e-06, 1.477922e-05, 2.535247e-05, 3.778122e-05, 
    4.536284e-05, 5.178419e-05, 4.059456e-05, 1.910911e-05, 9.676008e-06, 
    7.31391e-06, 5.356631e-06, 5.444624e-06, 5.457858e-06, 4.510242e-06,
  1.268619e-06, 6.35331e-06, 1.301617e-05, 1.354719e-05, 1.682597e-05, 
    2.034045e-05, 2.027529e-05, 1.412241e-05, 1.024423e-05, 1.069302e-05, 
    5.309907e-06, 5.106218e-06, 3.704347e-06, 4.13288e-06, 4.073349e-06,
  1.096797e-06, 1.765197e-06, 4.54134e-06, 4.854121e-06, 5.188463e-06, 
    4.285932e-06, 4.007083e-06, 4.646864e-06, 4.605698e-06, 5.059039e-06, 
    6.1931e-06, 5.96572e-06, 4.214827e-06, 3.237409e-06, 3.13253e-06,
  1.044869e-06, 1.959564e-06, 1.452554e-06, 1.933166e-06, 1.958173e-06, 
    2.751031e-06, 2.352758e-06, 3.590978e-06, 2.837855e-06, 3.265954e-06, 
    4.98968e-06, 7.43741e-06, 5.158049e-06, 4.32011e-06, 3.385899e-06,
  2.105051e-06, 2.213942e-06, 2.419417e-06, 2.665104e-06, 1.933192e-06, 
    2.037194e-06, 2.22019e-06, 3.275902e-06, 6.352367e-06, 7.301044e-06, 
    5.788852e-06, 6.405501e-06, 4.773588e-06, 5.144015e-06, 5.101069e-06,
  2.047618e-06, 2.160996e-06, 2.571166e-06, 3.514205e-06, 3.133638e-06, 
    3.052521e-06, 3.332937e-06, 4.794797e-06, 6.560282e-06, 8.596548e-06, 
    7.189542e-06, 4.26729e-06, 4.664358e-06, 6.304924e-06, 5.977729e-06,
  1.894388e-06, 2.224064e-06, 2.895324e-06, 4.06944e-06, 3.182975e-06, 
    2.35709e-06, 2.241353e-06, 2.262167e-06, 3.508782e-06, 4.706818e-06, 
    3.974686e-06, 3.504803e-06, 5.55091e-06, 8.585379e-06, 7.015477e-06,
  2.729763e-06, 2.92387e-06, 3.490342e-06, 3.340123e-06, 3.171863e-06, 
    4.441476e-06, 3.794715e-06, 3.442075e-06, 3.961017e-06, 3.708303e-06, 
    2.501673e-06, 3.47939e-06, 3.487588e-06, 4.785666e-06, 5.457692e-06,
  1.577288e-11, 1.616381e-17, 3.345161e-11, 5.5774e-10, 1.440884e-07, 
    9.237343e-07, 1.4867e-06, 1.459078e-06, 4.80607e-06, 1.497597e-05, 
    3.18386e-05, 4.896506e-05, 5.823392e-05, 5.58445e-05, 5.371808e-05,
  2.045449e-08, 5.191129e-15, 2.460203e-13, 4.336619e-10, 4.910184e-08, 
    9.331529e-07, 3.364941e-06, 3.947697e-06, 1.322755e-05, 2.856241e-05, 
    4.131398e-05, 5.223641e-05, 5.256426e-05, 4.804186e-05, 4.613253e-05,
  1.935353e-08, 2.375236e-10, 1.186731e-08, 3.851257e-08, 1.842346e-07, 
    1.742606e-06, 4.958403e-06, 1.297469e-05, 2.713477e-05, 3.406264e-05, 
    3.821693e-05, 3.975238e-05, 3.832682e-05, 3.538008e-05, 2.930284e-05,
  1.243473e-06, 9.068119e-07, 1.36459e-06, 2.490661e-06, 4.520884e-06, 
    9.304345e-06, 1.654612e-05, 2.596394e-05, 3.223975e-05, 2.88425e-05, 
    2.488673e-05, 2.409295e-05, 2.505651e-05, 2.63092e-05, 2.638154e-05,
  1.006808e-05, 1.389288e-05, 1.274561e-05, 1.327556e-05, 1.768754e-05, 
    2.323523e-05, 2.868501e-05, 2.860729e-05, 2.184137e-05, 1.509795e-05, 
    1.212166e-05, 1.279265e-05, 1.202843e-05, 1.54158e-05, 2.317026e-05,
  9.651889e-06, 2.100971e-05, 2.374255e-05, 2.151944e-05, 2.18617e-05, 
    2.428943e-05, 2.096524e-05, 1.656421e-05, 1.21351e-05, 8.100255e-06, 
    5.75422e-06, 5.748131e-06, 6.52598e-06, 9.000662e-06, 1.489605e-05,
  2.203066e-06, 5.523527e-06, 6.783935e-06, 7.045807e-06, 8.054407e-06, 
    8.306127e-06, 1.100371e-05, 1.239807e-05, 9.381003e-06, 7.913675e-06, 
    5.946037e-06, 6.010784e-06, 7.285358e-06, 1.082802e-05, 1.284303e-05,
  6.286418e-07, 8.1975e-07, 1.436972e-06, 1.594821e-06, 1.941632e-06, 
    3.478898e-06, 6.110512e-06, 6.405937e-06, 6.501396e-06, 6.758854e-06, 
    6.5197e-06, 6.388513e-06, 4.392565e-06, 5.516167e-06, 4.572964e-06,
  3.900696e-07, 1.463807e-06, 1.247376e-06, 2.284354e-06, 3.588446e-06, 
    3.756928e-06, 3.6507e-06, 2.448532e-06, 2.305203e-06, 3.884552e-06, 
    3.332929e-06, 1.968585e-06, 1.567177e-06, 2.673732e-06, 2.183558e-06,
  1.396351e-07, 3.789571e-07, 1.482343e-06, 3.658464e-06, 3.200387e-06, 
    3.279305e-06, 2.200437e-06, 1.354122e-06, 1.574477e-06, 1.718991e-06, 
    1.835725e-06, 1.437082e-06, 1.107237e-06, 1.570951e-06, 1.269879e-06,
  7.719319e-06, 8.035939e-06, 1.087938e-05, 1.521891e-05, 1.526796e-05, 
    1.640947e-05, 2.016008e-05, 2.793541e-05, 3.321972e-05, 3.924372e-05, 
    3.627831e-05, 2.692841e-05, 1.99071e-05, 8.183061e-06, 1.462509e-06,
  1.130601e-05, 1.681017e-05, 2.482095e-05, 3.133786e-05, 3.067416e-05, 
    2.773074e-05, 3.058838e-05, 3.731162e-05, 4.063337e-05, 4.199349e-05, 
    3.602517e-05, 2.854072e-05, 1.624848e-05, 4.989815e-06, 1.363793e-06,
  1.773566e-05, 3.263922e-05, 4.264836e-05, 5.141925e-05, 5.647429e-05, 
    5.577342e-05, 4.983244e-05, 4.395427e-05, 3.701658e-05, 3.04959e-05, 
    2.351071e-05, 1.682209e-05, 4.027607e-06, 4.29194e-06, 1.590238e-06,
  2.093804e-05, 2.539085e-05, 2.652769e-05, 2.944423e-05, 4.154574e-05, 
    5.422946e-05, 5.348186e-05, 4.181523e-05, 2.959962e-05, 1.756555e-05, 
    1.203531e-05, 7.61378e-06, 3.994837e-06, 1.990204e-06, 3.388384e-06,
  9.574416e-06, 5.202758e-06, 3.861431e-06, 4.419745e-06, 8.838003e-06, 
    1.612722e-05, 2.300164e-05, 2.921917e-05, 3.130229e-05, 2.380354e-05, 
    1.355766e-05, 6.220589e-06, 5.870733e-06, 4.405131e-06, 5.977024e-06,
  2.051697e-06, 1.423795e-06, 1.134025e-06, 1.555391e-06, 1.862554e-06, 
    2.696878e-06, 6.331981e-06, 1.36212e-05, 1.605387e-05, 6.319643e-06, 
    3.53094e-06, 3.643673e-06, 7.209272e-06, 7.861052e-06, 7.891786e-06,
  1.893044e-06, 1.41285e-06, 1.075424e-06, 1.390273e-06, 7.27977e-07, 
    8.036649e-07, 2.045177e-06, 3.313141e-06, 3.173241e-06, 4.192823e-06, 
    5.61778e-06, 8.571369e-06, 8.757744e-06, 1.037128e-05, 8.854178e-06,
  2.311465e-06, 2.179733e-06, 5.064128e-07, 4.657321e-07, 1.514563e-07, 
    3.316404e-07, 8.505868e-07, 1.571872e-06, 2.047801e-06, 1.407709e-06, 
    2.183598e-06, 1.220778e-06, 2.165521e-06, 1.167022e-06, 6.447626e-07,
  2.637076e-06, 8.71679e-07, 5.069138e-07, 2.93875e-07, 3.133237e-07, 
    2.917346e-07, 4.55168e-07, 5.469656e-07, 5.779331e-07, 5.570064e-07, 
    3.029665e-07, 4.518386e-07, 6.484684e-07, 3.901734e-07, 3.544159e-07,
  1.117195e-06, 1.525452e-06, 5.74227e-07, 9.816295e-07, 9.479872e-07, 
    8.616302e-07, 6.998586e-07, 9.418233e-07, 2.348926e-06, 1.975411e-06, 
    2.478801e-06, 2.631252e-06, 2.124831e-06, 3.429081e-06, 8.510276e-07,
  2.315988e-07, 3.262858e-08, 6.240413e-09, 1.410891e-09, 1.695594e-09, 
    3.136766e-10, 2.296242e-10, 1.234176e-10, 2.733868e-11, 5.201499e-08, 
    6.74159e-07, 2.467082e-06, 7.412896e-06, 1.537456e-05, 1.90558e-05,
  1.301931e-06, 4.136305e-07, 1.86264e-07, 2.993352e-08, 5.187299e-08, 
    1.716459e-08, 1.439127e-08, 1.700778e-07, 4.230684e-07, 8.265708e-07, 
    3.82489e-06, 1.060373e-05, 2.061118e-05, 2.803766e-05, 2.722712e-05,
  2.383892e-06, 2.766377e-06, 1.946664e-06, 2.098902e-06, 2.258961e-06, 
    1.489872e-06, 2.902172e-06, 2.831992e-06, 5.610254e-06, 8.589384e-06, 
    1.484911e-05, 2.352988e-05, 3.13898e-05, 3.045123e-05, 2.844769e-05,
  7.825126e-06, 1.967631e-05, 2.004897e-05, 1.642674e-05, 1.778446e-05, 
    1.840377e-05, 1.720069e-05, 1.797272e-05, 2.09395e-05, 2.481633e-05, 
    3.063561e-05, 3.69865e-05, 3.626548e-05, 3.471068e-05, 2.529002e-05,
  2.216328e-05, 3.747301e-05, 2.544027e-05, 1.516227e-05, 1.421067e-05, 
    1.991573e-05, 1.897224e-05, 2.259613e-05, 2.931912e-05, 4.503141e-05, 
    5.64783e-05, 5.758473e-05, 5.100225e-05, 4.218052e-05, 3.368465e-05,
  1.909512e-05, 2.210411e-05, 1.658859e-05, 1.020519e-05, 8.602418e-06, 
    4.951719e-06, 5.446861e-06, 6.692523e-06, 2.374607e-05, 4.880337e-05, 
    6.33694e-05, 6.617226e-05, 6.593574e-05, 6.152556e-05, 4.544113e-05,
  9.074434e-06, 8.263506e-06, 7.509676e-06, 6.658911e-06, 5.354848e-06, 
    4.555565e-06, 4.283216e-06, 5.448996e-06, 1.017708e-05, 1.577463e-05, 
    1.816439e-05, 1.598463e-05, 1.603547e-05, 2.033896e-05, 2.289311e-05,
  4.558878e-06, 2.921595e-06, 2.880362e-06, 2.777594e-06, 1.955753e-06, 
    3.550543e-06, 3.265543e-06, 3.338585e-06, 4.626449e-06, 4.919275e-06, 
    4.291408e-06, 4.336408e-06, 4.552997e-06, 7.160379e-06, 7.736147e-06,
  4.247264e-06, 4.612834e-06, 3.973811e-06, 1.945828e-06, 1.807723e-06, 
    1.688078e-06, 1.730861e-06, 1.60083e-06, 1.098958e-06, 6.738545e-07, 
    1.242468e-06, 1.835613e-06, 1.786371e-06, 1.689209e-06, 2.144117e-06,
  4.530777e-06, 4.573455e-06, 3.724252e-06, 2.025614e-06, 2.227653e-06, 
    3.647214e-06, 2.810889e-06, 2.232623e-06, 5.45011e-06, 5.245411e-06, 
    4.219221e-06, 4.462225e-06, 4.87291e-06, 4.886921e-06, 5.055829e-06,
  2.197836e-06, 2.727645e-06, 2.990058e-06, 2.899031e-06, 4.894326e-06, 
    4.626699e-06, 5.102249e-06, 5.941128e-06, 6.211058e-06, 8.695588e-06, 
    1.046729e-05, 1.240258e-05, 1.235521e-05, 1.432633e-05, 1.338429e-05,
  3.649478e-06, 2.936166e-06, 2.383958e-06, 1.222421e-06, 7.875148e-07, 
    7.042044e-07, 2.124834e-06, 3.141617e-06, 3.458296e-06, 4.213732e-06, 
    5.243875e-06, 4.346344e-06, 5.610529e-06, 5.969206e-06, 4.734985e-06,
  6.973091e-06, 5.501315e-06, 4.085283e-06, 3.20075e-06, 2.371911e-06, 
    1.525369e-06, 5.726225e-07, 2.506432e-07, 1.716127e-07, 2.290446e-07, 
    3.843149e-07, 1.592185e-06, 1.588027e-06, 1.431272e-06, 2.140292e-06,
  1.22325e-05, 1.412115e-05, 1.004563e-05, 6.629087e-06, 4.997667e-06, 
    4.157219e-06, 2.97271e-06, 8.402229e-07, 3.415135e-07, 6.712184e-08, 
    7.664354e-09, 1.962621e-07, 1.417669e-07, 1.052054e-07, 1.28256e-07,
  2.001988e-05, 2.056364e-05, 1.958311e-05, 1.260314e-05, 6.773606e-06, 
    6.07123e-06, 6.024037e-06, 3.889873e-06, 2.612843e-06, 5.478443e-07, 
    2.479553e-07, 8.688901e-08, 9.519078e-08, 3.904857e-07, 3.432547e-07,
  2.003326e-05, 1.883472e-05, 1.58758e-05, 1.449171e-05, 9.068541e-06, 
    1.02345e-05, 1.02045e-05, 1.157596e-05, 1.044638e-05, 1.04087e-05, 
    8.470399e-06, 6.690799e-06, 8.436062e-06, 7.764246e-06, 7.259303e-06,
  7.416671e-06, 6.124601e-06, 9.508426e-06, 9.035468e-06, 8.5201e-06, 
    8.392877e-06, 8.955595e-06, 1.20447e-05, 1.242743e-05, 1.534488e-05, 
    1.613983e-05, 1.522429e-05, 1.545358e-05, 1.072411e-05, 1.355949e-05,
  1.464611e-06, 1.257382e-06, 1.512359e-06, 2.255758e-06, 3.540528e-06, 
    3.928209e-06, 5.294001e-06, 6.270303e-06, 7.38335e-06, 8.962117e-06, 
    9.634648e-06, 9.683712e-06, 1.123356e-05, 9.886765e-06, 7.935891e-06,
  2.625779e-06, 1.598226e-06, 1.365768e-06, 2.541075e-06, 2.721296e-06, 
    2.286067e-06, 2.143223e-06, 2.374729e-06, 1.808181e-06, 2.222439e-06, 
    2.943317e-06, 2.007017e-06, 1.666667e-06, 2.329828e-06, 2.015791e-06,
  4.240406e-06, 3.264233e-06, 2.605347e-06, 3.325883e-06, 3.143383e-06, 
    5.252565e-06, 4.418019e-06, 2.153319e-05, 1.147117e-05, 2.024154e-05, 
    1.3696e-05, 1.677763e-05, 2.327062e-06, 2.070297e-06, 8.326291e-06,
  3.097191e-06, 3.482806e-06, 2.083007e-06, 1.632037e-06, 2.96109e-06, 
    2.854252e-06, 2.93359e-06, 3.292479e-06, 3.92842e-06, 4.022329e-06, 
    5.658404e-06, 8.112139e-06, 9.351963e-06, 9.01685e-06, 1.036014e-05,
  3.122875e-06, 2.55403e-06, 1.49351e-06, 1.418371e-06, 6.063298e-07, 
    1.110238e-06, 2.107053e-06, 2.475988e-06, 2.550308e-06, 4.059566e-06, 
    5.547538e-06, 6.698618e-06, 9.903601e-06, 8.902313e-06, 1.125311e-05,
  2.884476e-06, 5.348581e-06, 3.895325e-06, 1.649237e-06, 1.672011e-06, 
    1.301479e-06, 8.34013e-07, 7.978594e-07, 1.525727e-06, 3.304994e-06, 
    3.026295e-06, 4.237251e-06, 5.119882e-06, 6.850772e-06, 7.506113e-06,
  4.612829e-06, 3.77332e-06, 3.652272e-06, 3.701089e-06, 3.11844e-06, 
    1.544774e-06, 6.126074e-07, 3.137002e-07, 1.057038e-06, 5.008914e-07, 
    1.430706e-06, 2.166222e-06, 2.420984e-06, 3.776712e-06, 4.74651e-06,
  5.267196e-06, 6.200731e-06, 4.486277e-06, 4.685915e-06, 3.532057e-06, 
    4.408472e-06, 1.609828e-06, 1.740536e-06, 5.656297e-07, 3.859239e-07, 
    9.103634e-07, 1.387468e-06, 1.499193e-06, 1.520274e-06, 2.855708e-06,
  1.057854e-05, 7.48412e-06, 6.955193e-06, 5.09109e-06, 3.411956e-06, 
    4.359979e-06, 5.095704e-06, 4.194612e-06, 1.636258e-06, 3.715972e-07, 
    7.921482e-07, 1.662067e-06, 1.016421e-06, 8.838129e-07, 1.785607e-06,
  1.150504e-05, 1.359969e-05, 6.394365e-06, 5.691603e-06, 3.182337e-06, 
    5.279271e-06, 3.887234e-06, 5.408671e-06, 5.649059e-06, 5.219353e-06, 
    2.750571e-06, 3.524063e-06, 3.809164e-06, 2.84274e-06, 2.588381e-06,
  1.174506e-05, 1.072384e-05, 1.023009e-05, 8.388858e-06, 6.5272e-06, 
    6.505397e-06, 7.288035e-06, 2.169096e-05, 7.491664e-06, 7.806611e-06, 
    7.473852e-06, 6.781954e-06, 5.05786e-06, 7.151235e-06, 4.834718e-06,
  9.508534e-06, 9.993444e-06, 8.895248e-06, 9.827759e-06, 8.804101e-06, 
    6.764905e-06, 7.514412e-06, 8.227096e-06, 8.270846e-06, 6.993173e-06, 
    5.36793e-06, 6.492961e-06, 5.133123e-06, 4.792723e-06, 5.664927e-06,
  6.582819e-06, 6.748028e-06, 6.577448e-06, 1.024481e-05, 1.047691e-05, 
    1.003283e-05, 1.031228e-05, 1.236112e-05, 9.821163e-06, 9.766622e-06, 
    1.096993e-05, 8.175264e-06, 8.425159e-06, 6.329103e-06, 5.477356e-06,
  7.087785e-06, 1.138744e-05, 1.033472e-05, 7.063024e-06, 7.497066e-06, 
    8.382247e-06, 5.972911e-06, 3.481118e-06, 3.638801e-06, 4.150898e-06, 
    4.086115e-06, 3.355145e-06, 4.089159e-06, 3.436737e-06, 3.263837e-06,
  5.922785e-06, 7.012094e-06, 1.014661e-05, 7.603629e-06, 8.215219e-06, 
    7.704172e-06, 6.111828e-06, 5.262131e-06, 3.248031e-06, 3.928845e-06, 
    3.429721e-06, 4.372201e-06, 3.659389e-06, 3.699244e-06, 4.644332e-06,
  3.401492e-06, 5.119941e-06, 3.406851e-06, 5.618608e-06, 5.965358e-06, 
    6.900053e-06, 4.557015e-06, 3.049899e-06, 3.496132e-06, 5.379238e-06, 
    5.449556e-06, 3.461244e-06, 4.395292e-06, 3.807581e-06, 5.813334e-06,
  7.660503e-06, 2.388087e-06, 4.357825e-06, 4.970391e-06, 4.288864e-06, 
    4.138186e-06, 3.929656e-06, 3.813958e-06, 6.044209e-06, 4.138082e-06, 
    5.654985e-06, 3.889908e-06, 2.383153e-06, 3.43899e-06, 3.932284e-06,
  1.140135e-05, 1.009517e-05, 7.561957e-06, 5.37366e-06, 4.913981e-06, 
    5.575412e-06, 5.047209e-06, 3.940335e-06, 3.994873e-06, 3.842605e-06, 
    3.405485e-06, 3.825672e-06, 3.130709e-06, 2.475993e-06, 1.585408e-06,
  8.953251e-06, 1.073839e-05, 9.928141e-06, 1.53152e-06, 3.872773e-06, 
    4.60164e-06, 4.857457e-06, 4.782795e-06, 4.733197e-06, 3.698987e-06, 
    5.257891e-06, 2.13093e-06, 2.149648e-06, 3.212704e-06, 2.807438e-06,
  5.228728e-06, 9.680228e-06, 5.841698e-06, 4.147586e-06, 2.351957e-06, 
    1.464312e-06, 3.126535e-06, 5.42254e-06, 6.105127e-06, 7.884732e-06, 
    5.46262e-06, 5.331662e-06, 3.860097e-06, 3.905046e-06, 3.726125e-06,
  6.624392e-06, 6.16684e-06, 5.019197e-06, 3.077381e-06, 4.425305e-06, 
    6.045812e-06, 3.782702e-06, 6.732188e-06, 1.093707e-05, 8.434784e-06, 
    9.113544e-06, 7.858506e-06, 4.268962e-06, 4.088553e-06, 5.884962e-06,
  1.908887e-05, 1.854806e-05, 1.014451e-05, 4.589132e-06, 4.494185e-06, 
    3.462089e-06, 4.399491e-06, 5.303609e-06, 2.155376e-06, 4.410623e-06, 
    6.701189e-06, 9.795564e-06, 9.8511e-06, 8.345504e-06, 5.892348e-06,
  3.831912e-05, 3.076769e-05, 3.242242e-05, 2.142326e-05, 1.185841e-05, 
    5.578388e-06, 5.767047e-06, 4.055303e-06, 3.779894e-06, 2.176867e-06, 
    5.257003e-06, 7.674736e-06, 8.036413e-06, 9.822471e-06, 9.666634e-06,
  4.340084e-06, 4.663944e-06, 8.401474e-06, 5.981748e-06, 3.614671e-06, 
    4.006959e-06, 2.76564e-06, 3.136345e-06, 3.857428e-06, 5.991305e-06, 
    8.477737e-06, 5.080852e-06, 4.138415e-06, 3.444164e-06, 5.443213e-06,
  2.993701e-06, 4.709858e-06, 6.118228e-06, 5.686183e-06, 4.002502e-06, 
    3.490416e-06, 3.519944e-06, 3.281202e-06, 2.436898e-06, 5.514965e-06, 
    5.517499e-06, 6.407242e-06, 3.870562e-06, 4.597867e-06, 4.583969e-06,
  2.892725e-06, 2.734723e-06, 4.593973e-06, 5.612127e-06, 4.501736e-06, 
    4.023644e-06, 4.370248e-06, 3.543064e-06, 1.518924e-06, 6.240665e-06, 
    5.461023e-06, 5.259782e-06, 2.309726e-06, 3.615854e-06, 5.07252e-06,
  1.771023e-06, 2.55372e-06, 3.441626e-06, 3.981205e-06, 4.764836e-06, 
    4.431218e-06, 5.528449e-06, 3.708547e-06, 5.339281e-06, 6.877111e-06, 
    6.276323e-06, 6.027374e-06, 4.834621e-06, 5.033703e-06, 3.81863e-06,
  2.091398e-06, 2.880375e-06, 3.645986e-06, 7.484413e-06, 1.140301e-05, 
    1.543303e-05, 1.758788e-05, 2.891094e-05, 3.439888e-05, 2.262804e-05, 
    1.863186e-05, 1.425523e-05, 5.826474e-06, 4.475492e-06, 3.778218e-06,
  6.048602e-06, 9.648562e-06, 1.460577e-05, 2.18257e-05, 3.222041e-05, 
    5.606999e-05, 0.0001221327, 0.0001317113, 0.0001078777, 5.485241e-05, 
    2.199146e-05, 1.110634e-05, 2.379555e-06, 2.969411e-06, 4.542609e-06,
  9.818279e-06, 1.684922e-05, 1.995342e-05, 1.831158e-05, 3.558309e-05, 
    0.0001474098, 0.0002945441, 0.0003117271, 0.0002614121, 0.0001509417, 
    5.210676e-05, 1.217647e-05, 5.25364e-06, 5.787649e-06, 4.089976e-06,
  1.871952e-05, 3.448057e-05, 3.628814e-05, 2.652568e-05, 9.110675e-05, 
    0.0003978808, 0.0005052621, 0.0005753009, 0.0003959097, 0.0002046065, 
    5.904925e-05, 2.559282e-05, 1.300521e-05, 6.533378e-06, 2.018149e-05,
  3.626078e-05, 3.375909e-05, 2.451041e-05, 5.399081e-05, 0.0003110843, 
    0.0006610663, 0.0006820547, 0.0007510724, 0.0006392548, 0.0002570532, 
    8.876514e-05, 2.905266e-05, 2.328575e-05, 2.23121e-05, 2.347809e-05,
  3.474733e-05, 2.99184e-05, 3.056309e-05, 0.0001659174, 0.0008616444, 
    0.001039778, 0.0009715434, 0.001063524, 0.0007901517, 0.0002927332, 
    5.325529e-05, 3.107946e-05, 3.062266e-05, 3.954682e-05, 2.920542e-05,
  1.693606e-06, 2.111185e-06, 2.247477e-06, 4.297322e-06, 4.666275e-06, 
    2.316341e-06, 1.94304e-06, 3.59091e-06, 4.814976e-06, 5.886801e-06, 
    7.665264e-06, 7.084954e-06, 3.361343e-06, 1.431882e-06, 9.216451e-07,
  2.752796e-06, 2.417984e-06, 1.053669e-05, 2.49978e-05, 1.085462e-05, 
    3.736199e-06, 2.371986e-06, 2.562186e-06, 3.477651e-06, 4.258212e-06, 
    7.108695e-06, 1.231315e-05, 1.461776e-05, 1.311011e-05, 1.032243e-05,
  5.04757e-06, 1.910261e-05, 0.0001690149, 0.0002299702, 6.014444e-05, 
    1.033928e-05, 5.978222e-06, 6.188823e-06, 7.269392e-06, 9.688686e-06, 
    1.206405e-05, 1.656973e-05, 1.856714e-05, 1.972891e-05, 2.064917e-05,
  1.121616e-05, 6.885947e-05, 0.0004674848, 0.0006017194, 0.0003083155, 
    5.559115e-05, 5.082042e-05, 4.747187e-05, 4.028036e-05, 4.511463e-05, 
    5.416694e-05, 5.991135e-05, 5.758826e-05, 4.918254e-05, 3.684344e-05,
  2.760632e-05, 0.0001306214, 0.0006593093, 0.0008967063, 0.0006591682, 
    0.0001634441, 0.0001324111, 0.0001518372, 0.0001351388, 9.678305e-05, 
    7.343143e-05, 5.996106e-05, 6.194396e-05, 6.239676e-05, 6.157508e-05,
  4.332804e-05, 0.0001431768, 0.0005258175, 0.001022784, 0.0009032522, 
    0.000325022, 0.000192964, 0.0002306927, 0.0001963323, 0.0001185594, 
    6.299746e-05, 2.395218e-05, 1.749401e-05, 2.415703e-05, 2.068561e-05,
  4.569723e-05, 0.0001530371, 0.0003770829, 0.0008989031, 0.001097369, 
    0.0005419724, 0.0002037731, 0.0001704852, 0.0001142876, 7.94073e-05, 
    6.746606e-05, 3.045389e-05, 2.794275e-05, 2.458964e-05, 1.405232e-05,
  3.009222e-05, 0.00011644, 0.0002824413, 0.0006693635, 0.001201596, 
    0.0007255671, 0.0001507644, 3.180527e-05, 3.322434e-05, 1.994556e-05, 
    9.744901e-06, 1.431788e-05, 4.33083e-06, 7.154039e-06, 5.629074e-06,
  3.636277e-05, 8.132162e-05, 0.0002193485, 0.0005211092, 0.001167388, 
    0.0008106727, 7.622373e-05, 1.793862e-06, 4.012037e-07, 1.704505e-05, 
    9.486419e-06, 8.376472e-06, 7.353849e-08, 5.973213e-08, 7.59336e-06,
  1.449174e-05, 5.192357e-05, 0.0001370861, 0.0003862258, 0.001149374, 
    0.0006797341, 1.332236e-05, 4.577596e-07, 2.959778e-07, 2.592673e-06, 
    4.135428e-06, 4.7186e-08, 8.027292e-06, 1.497174e-05, 1.891617e-05,
  1.221802e-05, 0.0004634882, 0.0005616456, 0.0004184764, 0.0001847454, 
    0.0001582461, 0.0001175678, 5.511994e-05, 1.738957e-05, 8.630734e-06, 
    1.169519e-05, 1.121847e-05, 1.099673e-05, 8.776261e-06, 1.090597e-05,
  1.025394e-05, 0.0003106802, 0.0006332406, 0.0004704455, 0.0001172775, 
    3.157423e-05, 2.787227e-05, 2.116103e-05, 1.306122e-05, 6.955765e-06, 
    8.553657e-06, 9.212036e-06, 9.63051e-06, 9.314929e-06, 9.607232e-06,
  6.007008e-06, 6.338418e-05, 0.0005353628, 0.0004447298, 0.0002273667, 
    3.93749e-05, 2.073776e-05, 1.488935e-05, 7.567202e-06, 6.539659e-06, 
    7.912719e-06, 6.811884e-06, 1.026648e-05, 9.85977e-06, 8.685118e-06,
  6.172329e-06, 1.518857e-05, 0.0002386399, 0.0002184913, 0.000151813, 
    4.290567e-05, 1.426495e-05, 7.663834e-06, 2.995862e-06, 3.665446e-06, 
    5.077211e-06, 5.39057e-06, 1.073268e-05, 1.011506e-05, 7.948093e-06,
  5.095744e-06, 3.119578e-06, 3.812329e-06, 2.879818e-05, 5.687464e-05, 
    3.092906e-05, 8.521443e-06, 2.4771e-06, 1.232039e-06, 8.591977e-07, 
    1.576764e-06, 2.194528e-06, 8.554057e-06, 1.067578e-05, 8.874741e-06,
  2.939377e-06, 4.124892e-06, 5.828733e-06, 1.675524e-05, 4.421482e-05, 
    2.66302e-05, 3.462407e-06, 2.688318e-07, 4.818237e-07, 2.664485e-07, 
    1.896986e-07, 6.234437e-07, 5.02171e-06, 9.716216e-06, 1.228371e-05,
  1.657779e-06, 8.682101e-06, 1.452303e-05, 3.060559e-05, 4.868672e-05, 
    1.952295e-05, 7.235511e-07, 1.351207e-07, 3.385054e-07, 1.786223e-07, 
    2.843851e-08, 1.003553e-06, 2.114334e-06, 5.395516e-06, 7.158808e-06,
  2.170165e-06, 8.898312e-06, 3.259356e-05, 5.912934e-05, 3.911995e-05, 
    4.168799e-06, 4.236124e-07, 2.475313e-08, 9.632535e-08, 2.093223e-07, 
    1.191783e-07, 1.40768e-06, 1.02594e-06, 6.604951e-07, 6.759489e-07,
  3.438722e-06, 5.01487e-06, 1.08529e-05, 1.870695e-05, 1.585374e-05, 
    9.727229e-07, 6.55177e-07, 3.188625e-07, 5.207936e-08, 8.517798e-07, 
    3.348127e-07, 1.168336e-06, 7.859875e-08, 1.300648e-08, 4.63612e-08,
  1.14714e-06, 3.30292e-06, 4.244152e-06, 5.392801e-06, 3.793199e-06, 
    1.793732e-06, 1.926188e-06, 1.822436e-07, 2.972887e-08, 1.893327e-06, 
    1.001092e-05, 3.262054e-07, 2.562741e-08, 4.481873e-06, 8.993179e-07,
  1.028003e-05, 6.669845e-06, 6.432196e-06, 7.463802e-06, 6.192057e-06, 
    6.155477e-06, 1.072242e-05, 3.733312e-05, 4.421288e-05, 3.57557e-05, 
    2.894118e-05, 2.406485e-05, 2.437094e-05, 2.129844e-05, 1.903593e-05,
  1.138534e-05, 1.315617e-05, 1.125697e-05, 1.11616e-05, 9.364636e-06, 
    8.40076e-06, 1.238346e-05, 2.045493e-05, 2.031347e-05, 1.898414e-05, 
    1.827547e-05, 2.033978e-05, 1.811397e-05, 1.888169e-05, 2.053761e-05,
  1.637832e-05, 2.456474e-05, 3.095911e-05, 2.982032e-05, 2.80247e-05, 
    2.894334e-05, 2.92469e-05, 2.979707e-05, 2.77649e-05, 2.754661e-05, 
    2.350794e-05, 1.693229e-05, 1.774073e-05, 1.728321e-05, 1.708612e-05,
  3.192089e-05, 5.403098e-05, 5.447862e-05, 5.055885e-05, 4.420181e-05, 
    4.021874e-05, 3.331478e-05, 2.896243e-05, 2.527815e-05, 2.209754e-05, 
    1.453516e-05, 1.439998e-05, 1.382849e-05, 1.495727e-05, 1.661199e-05,
  1.905286e-05, 1.688583e-05, 1.024164e-05, 2.285528e-06, 1.664882e-06, 
    2.279809e-06, 4.530746e-06, 5.41664e-06, 6.740297e-06, 9.632978e-06, 
    9.612753e-06, 1.105643e-05, 1.413338e-05, 1.196382e-05, 1.393875e-05,
  5.286812e-06, 1.766616e-07, 1.215327e-07, 6.29777e-08, 7.421825e-08, 
    1.697985e-07, 7.347693e-07, 1.561771e-06, 5.532125e-06, 4.21601e-06, 
    3.35132e-06, 6.133751e-06, 1.075256e-05, 7.399155e-06, 1.281488e-05,
  7.872701e-08, 2.718288e-08, 4.43619e-08, 2.491645e-08, 4.76885e-08, 
    8.909364e-09, 7.411431e-09, 3.07289e-07, 9.561272e-07, 9.016413e-07, 
    7.341679e-07, 1.872248e-06, 5.516875e-06, 9.179364e-06, 9.703963e-06,
  2.96496e-07, 7.848803e-09, 6.01339e-09, 6.085928e-09, 1.194151e-07, 
    2.43288e-08, 7.153371e-09, 5.692649e-09, 7.356345e-09, 6.63199e-07, 
    3.248055e-06, 4.981679e-06, 1.509283e-05, 1.386101e-05, 3.420453e-05,
  2.531825e-07, 2.831119e-07, 1.849828e-08, 3.316681e-07, 1.254172e-07, 
    3.89213e-09, 3.035797e-09, 1.900121e-07, 3.710495e-07, 3.064778e-06, 
    4.672409e-05, 8.140792e-05, 0.000107162, 9.445662e-05, 3.453446e-05,
  5.667939e-07, 4.277994e-07, 1.572416e-07, 4.319906e-07, 5.424349e-07, 
    5.01949e-07, 1.898667e-06, 1.058301e-05, 3.339662e-05, 2.68644e-05, 
    8.354508e-05, 3.97761e-05, 1.129196e-05, 1.421339e-05, 4.219254e-06,
  0.0001601688, 0.0001755777, 0.0001131424, 4.354495e-05, 5.229798e-06, 
    1.502661e-06, 9.503738e-07, 1.068959e-06, 8.762721e-07, 1.011296e-06, 
    1.030941e-06, 1.331311e-06, 1.221136e-06, 1.507707e-06, 1.298529e-06,
  7.108047e-05, 0.0001080434, 0.0001370279, 0.0001409067, 8.361754e-05, 
    2.894411e-05, 3.598803e-06, 1.041308e-06, 9.650724e-07, 1.506829e-06, 
    2.239215e-06, 2.380749e-06, 2.549554e-06, 1.985473e-06, 1.733795e-06,
  1.433416e-05, 1.35232e-05, 1.969676e-05, 3.269269e-05, 5.409099e-05, 
    4.727821e-05, 2.496082e-05, 1.394308e-05, 2.92118e-06, 7.052016e-07, 
    3.204031e-06, 2.405022e-06, 3.239652e-06, 3.944762e-06, 6.573334e-06,
  2.586264e-05, 3.419125e-05, 4.063936e-05, 4.35121e-05, 4.185173e-05, 
    5.431349e-05, 6.838412e-05, 5.00096e-05, 3.349724e-05, 1.586451e-05, 
    1.406086e-05, 1.175352e-05, 7.540873e-06, 9.83762e-06, 9.095622e-06,
  1.538133e-05, 1.265532e-05, 1.163894e-05, 9.68578e-06, 1.598771e-05, 
    3.049662e-05, 5.286103e-05, 8.051693e-05, 0.0001077507, 0.0001194807, 
    8.469157e-05, 3.081649e-05, 8.246254e-06, 8.77414e-06, 6.490593e-06,
  1.287907e-05, 7.275095e-06, 1.793043e-06, 2.339475e-06, 1.966519e-06, 
    1.836821e-06, 1.673192e-06, 2.660089e-06, 8.780356e-06, 3.756952e-05, 
    7.39317e-05, 7.261898e-05, 5.253377e-05, 2.222763e-05, 8.081878e-06,
  5.627547e-06, 3.622194e-06, 2.297647e-06, 9.845398e-07, 1.259342e-06, 
    5.723756e-07, 2.717825e-07, 6.860095e-08, 2.659992e-07, 2.275747e-06, 
    5.398459e-06, 7.863169e-06, 6.991029e-06, 9.931355e-06, 6.335132e-06,
  2.914193e-06, 1.83077e-06, 1.22474e-06, 1.008303e-06, 1.572845e-06, 
    6.888338e-07, 2.239316e-06, 3.955013e-06, 4.438583e-06, 1.690458e-06, 
    1.303136e-06, 3.162606e-06, 4.425331e-06, 6.173404e-06, 1.339893e-05,
  3.804852e-06, 1.822983e-06, 3.208879e-06, 2.41179e-06, 8.917241e-06, 
    5.373499e-06, 7.553139e-06, 7.453586e-06, 8.780115e-06, 1.181201e-05, 
    1.064921e-05, 2.589562e-05, 2.238953e-05, 3.082589e-05, 2.426925e-05,
  1.23489e-06, 2.30837e-06, 1.148527e-06, 2.165874e-06, 6.496362e-06, 
    1.175577e-05, 1.131227e-05, 2.397486e-05, 2.624089e-05, 3.54579e-05, 
    8.061837e-06, 3.419714e-06, 4.785058e-06, 9.323111e-06, 9.082616e-06,
  7.65209e-05, 0.0001108784, 0.0001245431, 5.852987e-05, 1.593767e-05, 
    4.285243e-06, 3.522659e-06, 1.623961e-06, 1.619823e-06, 2.226919e-07, 
    3.345632e-07, 2.257612e-08, 5.89186e-09, 4.633746e-09, 3.494155e-09,
  8.289177e-06, 1.521189e-05, 7.645819e-05, 0.000144737, 0.0001902676, 
    0.0001309291, 2.93441e-05, 6.423093e-06, 4.521497e-06, 1.609443e-06, 
    6.31566e-07, 1.233313e-07, 4.670165e-08, 2.228774e-08, 6.834421e-09,
  5.114137e-06, 1.388967e-06, 4.649134e-06, 2.326616e-05, 0.0001036802, 
    0.0001725309, 0.0001849989, 0.0001475621, 8.255794e-05, 2.694928e-05, 
    1.082253e-05, 9.284207e-07, 1.561718e-07, 1.885962e-08, 1.411634e-08,
  4.186794e-06, 5.201894e-07, 7.292393e-07, 1.540124e-06, 7.36296e-06, 
    2.889384e-05, 6.861563e-05, 0.0001423027, 0.0001759609, 0.0001620752, 
    8.953873e-05, 3.48791e-05, 1.529523e-05, 1.0497e-07, 2.013339e-08,
  3.491159e-06, 2.880377e-06, 1.104906e-06, 1.50986e-06, 1.296149e-06, 
    4.316553e-06, 9.116641e-06, 2.150539e-05, 4.771367e-05, 0.0001309133, 
    0.0001968354, 0.0001581989, 7.438339e-05, 1.37238e-05, 1.343872e-07,
  1.359098e-06, 2.337028e-06, 1.025581e-06, 1.828686e-06, 1.51699e-06, 
    2.958421e-06, 4.184281e-06, 1.823374e-06, 6.280937e-06, 3.696425e-05, 
    7.40976e-05, 0.000159791, 0.0002027338, 0.0001080383, 1.410764e-05,
  1.954952e-06, 8.841894e-07, 2.753062e-06, 5.922105e-06, 1.50302e-06, 
    2.173482e-06, 2.821165e-06, 6.270775e-06, 2.036049e-06, 5.151075e-06, 
    1.108336e-05, 2.174231e-05, 5.885774e-05, 0.0001200587, 9.455652e-05,
  2.694468e-06, 4.395058e-06, 5.751243e-06, 3.789493e-06, 8.26733e-07, 
    1.126059e-06, 1.954091e-06, 4.985611e-06, 4.473361e-06, 4.346699e-06, 
    8.932533e-06, 1.521523e-05, 1.641359e-05, 1.656796e-05, 1.555398e-05,
  4.128327e-06, 5.222944e-06, 3.746438e-06, 3.753268e-06, 3.776298e-06, 
    7.053188e-06, 8.307709e-06, 1.225957e-05, 1.290053e-05, 7.58811e-06, 
    1.644601e-05, 1.148217e-05, 2.996391e-05, 2.044052e-05, 1.244997e-05,
  4.775311e-06, 2.170409e-06, 2.459673e-06, 4.343645e-06, 4.293641e-06, 
    9.348357e-06, 9.120653e-06, 7.46429e-06, 3.170239e-06, 7.366065e-06, 
    5.796844e-06, 5.08368e-06, 1.005432e-05, 1.789943e-05, 1.65337e-05,
  6.652132e-06, 5.539979e-06, 6.143173e-06, 5.908185e-06, 4.96449e-06, 
    4.348108e-06, 8.359387e-06, 7.22032e-06, 9.442915e-06, 1.044097e-05, 
    9.047963e-06, 8.402753e-06, 3.516473e-06, 1.648582e-06, 4.32071e-07,
  6.210425e-06, 6.898389e-06, 6.576967e-06, 6.304623e-06, 1.82007e-06, 
    1.607099e-06, 5.874487e-06, 4.637944e-06, 6.632536e-06, 1.119974e-05, 
    1.18842e-05, 1.137399e-05, 6.373358e-06, 3.25062e-06, 5.791568e-07,
  3.84662e-06, 5.052567e-06, 4.566007e-06, 5.573136e-06, 2.832867e-06, 
    1.770975e-06, 6.227991e-06, 1.871374e-06, 2.923537e-06, 5.84904e-06, 
    1.024333e-05, 2.771194e-05, 2.626004e-05, 8.65738e-06, 3.138081e-06,
  6.283389e-07, 2.225226e-06, 2.932356e-06, 3.742939e-06, 2.884541e-06, 
    2.87509e-06, 1.527987e-06, 5.681016e-07, 9.516149e-07, 1.876219e-06, 
    8.450871e-06, 2.912178e-05, 3.923208e-05, 1.619605e-05, 4.245937e-06,
  2.305112e-07, 1.993665e-07, 5.296004e-07, 2.025614e-06, 2.752581e-06, 
    2.527451e-06, 4.510852e-07, 1.919887e-07, 2.410466e-07, 5.799772e-07, 
    1.607985e-07, 9.382088e-06, 2.700828e-05, 1.473237e-05, 6.305874e-07,
  1.173303e-07, 5.243995e-07, 6.171744e-07, 2.214473e-06, 3.090878e-06, 
    4.345536e-06, 2.289865e-06, 1.536746e-06, 9.426689e-07, 1.732121e-06, 
    1.17754e-07, 1.269948e-05, 1.19633e-05, 5.539551e-06, 1.590624e-06,
  1.308453e-06, 1.307918e-06, 3.740887e-06, 3.462278e-06, 9.657782e-07, 
    5.365895e-07, 5.983431e-06, 4.167965e-06, 9.838846e-06, 6.144535e-06, 
    7.204542e-06, 1.418332e-05, 1.198269e-05, 5.102538e-06, 5.100733e-07,
  1.711677e-06, 1.806912e-06, 2.220744e-06, 2.266237e-06, 1.917443e-06, 
    5.103082e-06, 1.345192e-06, 4.359347e-06, 3.154801e-06, 5.325276e-06, 
    9.114272e-06, 1.294466e-05, 1.575718e-05, 7.282471e-06, 2.815009e-06,
  2.582857e-06, 1.959647e-06, 1.585486e-06, 2.23729e-06, 2.648299e-06, 
    5.249697e-06, 9.716696e-06, 4.795562e-06, 3.516726e-06, 5.463209e-06, 
    1.144292e-05, 2.316818e-05, 6.804907e-06, 6.456211e-06, 3.931981e-06,
  1.528152e-06, 1.121948e-06, 8.227614e-07, 8.075177e-07, 1.699284e-06, 
    4.723147e-06, 5.066122e-06, 1.268384e-05, 1.693663e-05, 1.073548e-05, 
    2.111056e-05, 2.241257e-05, 1.657685e-05, 8.093106e-06, 7.840137e-06,
  1.890645e-05, 3.668168e-05, 5.215517e-05, 7.074989e-05, 8.268495e-05, 
    7.512107e-05, 4.875311e-05, 2.735366e-05, 1.396458e-05, 1.21394e-05, 
    1.064067e-05, 6.694628e-06, 2.301006e-06, 9.14698e-07, 3.163594e-07,
  1.455229e-05, 3.610433e-05, 5.05509e-05, 6.559307e-05, 6.311572e-05, 
    3.878661e-05, 2.101404e-05, 1.054845e-05, 1.115918e-05, 1.064703e-05, 
    7.195706e-06, 3.380982e-06, 4.769212e-07, 3.405259e-08, 2.701604e-08,
  1.664188e-05, 3.340694e-05, 4.667644e-05, 4.781174e-05, 2.995575e-05, 
    1.23623e-05, 6.851392e-06, 3.515786e-06, 7.415e-06, 6.681113e-06, 
    2.392878e-06, 3.716403e-07, 2.614477e-08, 5.989657e-10, 6.44404e-09,
  1.897207e-05, 3.338019e-05, 3.185281e-05, 1.880538e-05, 3.825613e-06, 
    9.002593e-07, 9.650545e-07, 2.686843e-07, 9.083109e-07, 1.138434e-06, 
    2.346449e-07, 4.413794e-08, 1.178425e-09, 1.441689e-10, 8.932609e-10,
  2.286346e-05, 2.95531e-05, 1.59696e-05, 1.219454e-06, 2.503282e-07, 
    1.257339e-07, 2.413463e-08, 3.83826e-08, 6.402188e-08, 1.268276e-07, 
    2.546061e-08, 4.521148e-09, 1.67212e-10, 1.209027e-10, 1.32584e-08,
  2.681748e-05, 2.306181e-05, 2.19894e-06, 1.870854e-07, 3.894844e-07, 
    1.51865e-08, 1.903693e-08, 8.170429e-09, 9.884911e-07, 3.939727e-06, 
    5.123962e-09, 3.541905e-09, 1.397102e-10, 1.386485e-08, 1.245042e-07,
  2.458005e-05, 1.336447e-06, 5.552031e-07, 1.414474e-07, 1.479926e-07, 
    9.453224e-07, 1.609303e-06, 3.645349e-06, 7.038929e-06, 9.786776e-06, 
    8.074795e-06, 4.130784e-06, 1.323889e-06, 6.061186e-07, 3.752173e-07,
  2.220692e-06, 5.106053e-07, 8.541392e-07, 4.063098e-07, 1.311986e-08, 
    1.06615e-06, 3.394205e-07, 1.482221e-06, 3.716738e-06, 8.819623e-06, 
    6.773176e-06, 5.472426e-06, 5.104531e-06, 3.482113e-06, 2.037545e-06,
  8.397643e-07, 1.605522e-06, 2.384128e-06, 1.633171e-06, 9.127946e-07, 
    3.895337e-07, 7.213219e-07, 1.066817e-06, 2.324806e-06, 5.157274e-06, 
    6.367107e-06, 9.579377e-06, 8.276417e-06, 8.278385e-06, 8.818974e-06,
  1.542192e-06, 1.787088e-06, 1.848823e-06, 2.929986e-06, 4.894287e-07, 
    4.030296e-07, 8.040331e-07, 1.266104e-06, 1.532261e-06, 2.429345e-06, 
    4.945054e-06, 6.970575e-06, 7.669137e-06, 1.596451e-05, 1.96518e-05,
  3.310872e-06, 4.289731e-06, 3.046187e-06, 1.123918e-06, 3.010484e-06, 
    2.5396e-05, 5.546094e-05, 7.863113e-05, 9.023723e-05, 9.317307e-05, 
    8.797398e-05, 7.279225e-05, 5.280274e-05, 3.739006e-05, 2.960691e-05,
  6.345555e-06, 4.320331e-06, 2.389559e-06, 2.055643e-06, 1.764987e-05, 
    4.880857e-05, 7.192348e-05, 7.477662e-05, 6.865779e-05, 5.459857e-05, 
    3.29967e-05, 2.037009e-05, 1.535018e-05, 1.47595e-05, 1.300724e-05,
  5.092949e-06, 4.152397e-06, 2.910681e-06, 1.932667e-05, 4.684604e-05, 
    6.226944e-05, 6.65143e-05, 5.841802e-05, 3.905021e-05, 2.540898e-05, 
    1.920306e-05, 2.062871e-05, 2.295597e-05, 2.405923e-05, 2.26856e-05,
  2.779442e-06, 5.657728e-06, 1.916721e-05, 4.302821e-05, 6.110936e-05, 
    6.093884e-05, 4.460654e-05, 2.875426e-05, 2.616866e-05, 2.943375e-05, 
    2.883718e-05, 2.393338e-05, 2.644436e-05, 2.579413e-05, 2.201875e-05,
  9.303905e-06, 2.503975e-05, 4.179744e-05, 5.422758e-05, 4.197382e-05, 
    3.162636e-05, 2.804388e-05, 3.741862e-05, 3.599516e-05, 2.041872e-05, 
    1.982737e-05, 1.909703e-05, 1.351108e-05, 1.133884e-05, 8.675433e-06,
  2.552259e-05, 3.8535e-05, 3.956875e-05, 3.39798e-05, 2.675428e-05, 
    2.872979e-05, 1.705031e-05, 1.328309e-05, 1.830263e-05, 2.794541e-05, 
    3.997365e-05, 3.595096e-05, 6.899454e-05, 6.415255e-05, 1.011392e-05,
  5.037066e-05, 3.929594e-05, 2.385625e-05, 1.821965e-05, 1.738362e-05, 
    1.657466e-05, 1.519964e-05, 1.450749e-05, 2.826025e-05, 2.849742e-05, 
    4.365123e-05, 4.209855e-05, 4.647986e-05, 2.247037e-05, 1.809227e-05,
  3.24922e-05, 2.428639e-05, 2.120099e-05, 1.729384e-05, 1.313383e-05, 
    8.320113e-06, 6.587133e-06, 4.682806e-06, 5.988134e-06, 1.743101e-05, 
    1.642576e-05, 1.568424e-05, 2.189213e-05, 1.948955e-05, 2.269901e-05,
  3.084668e-05, 1.834551e-05, 1.425965e-05, 9.485936e-06, 5.540295e-06, 
    4.290516e-06, 3.121321e-06, 2.84321e-06, 5.130199e-06, 5.696561e-06, 
    6.659827e-06, 7.444035e-06, 1.2614e-05, 1.834222e-05, 2.661255e-05,
  1.897618e-05, 1.205407e-05, 1.514618e-05, 7.348968e-06, 2.98894e-06, 
    1.898424e-06, 2.276151e-06, 2.506238e-06, 3.489053e-06, 4.8992e-06, 
    4.202141e-06, 7.442584e-06, 5.947399e-06, 1.390641e-05, 1.046871e-05,
  9.65213e-06, 8.056083e-06, 5.121851e-06, 4.724712e-06, 4.099713e-06, 
    3.84551e-06, 3.135707e-06, 2.684045e-06, 1.449803e-06, 1.478244e-06, 
    1.426188e-06, 7.611801e-07, 3.217614e-06, 2.710687e-06, 2.659576e-06,
  4.986345e-06, 3.250686e-06, 4.910422e-06, 5.776835e-06, 3.463054e-06, 
    2.382713e-06, 1.400498e-06, 1.850136e-06, 1.533211e-06, 6.205539e-07, 
    7.514138e-07, 1.64299e-06, 1.581355e-06, 4.313075e-07, 1.599769e-06,
  7.90655e-06, 2.482868e-06, 2.257478e-06, 1.991631e-06, 5.760457e-07, 
    6.572139e-07, 8.440651e-07, 9.042e-07, 7.474075e-07, 9.372952e-07, 
    6.006256e-07, 6.099664e-07, 7.243113e-07, 2.843444e-06, 1.041633e-06,
  1.170646e-05, 5.703973e-06, 1.443887e-06, 1.001165e-06, 5.262091e-07, 
    2.457011e-06, 1.203627e-06, 1.945972e-06, 2.642651e-06, 5.077731e-06, 
    4.857735e-06, 3.133218e-06, 2.896553e-06, 6.39284e-06, 8.831118e-06,
  2.054156e-05, 1.621023e-05, 1.011176e-05, 9.583333e-06, 8.354409e-06, 
    7.198144e-06, 4.618973e-06, 5.573823e-06, 7.501479e-06, 8.374451e-06, 
    7.714693e-06, 9.364507e-06, 8.241826e-06, 9.003918e-06, 1.052905e-05,
  1.71401e-05, 1.973532e-05, 1.910232e-05, 1.913865e-05, 1.423121e-05, 
    1.402567e-05, 1.357534e-05, 1.514037e-05, 1.515701e-05, 1.832648e-05, 
    1.601673e-05, 3.471108e-05, 4.737867e-05, 6.410154e-05, 6.460799e-05,
  3.430608e-05, 3.516275e-05, 2.254455e-05, 1.631326e-05, 1.593585e-05, 
    1.487158e-05, 1.191055e-05, 1.150571e-05, 2.450681e-05, 4.233652e-05, 
    7.668735e-05, 7.103247e-05, 7.570304e-05, 0.0001320958, 0.000165369,
  3.244328e-05, 3.077049e-05, 1.998878e-05, 1.234616e-05, 1.034154e-05, 
    8.419945e-06, 1.300659e-05, 1.996834e-05, 4.055158e-05, 7.778249e-05, 
    7.64595e-05, 0.0001128969, 0.0001373266, 6.302629e-05, 5.513187e-05,
  3.127293e-05, 1.797176e-05, 9.617536e-06, 7.388487e-06, 7.413516e-06, 
    7.178578e-06, 1.407758e-05, 1.851443e-05, 2.193741e-05, 4.53853e-05, 
    4.766816e-05, 3.846846e-05, 4.918875e-05, 3.190935e-05, 4.315607e-05,
  1.671283e-05, 8.953015e-06, 4.930921e-06, 5.776454e-06, 1.004253e-05, 
    1.905827e-05, 1.235521e-05, 1.455366e-05, 1.094095e-05, 8.377646e-06, 
    1.421548e-05, 1.290158e-05, 2.375691e-05, 2.048236e-05, 1.572746e-05,
  9.135288e-06, 7.605125e-06, 6.543282e-06, 5.052831e-06, 4.935327e-06, 
    3.012351e-06, 2.62197e-06, 2.151447e-06, 5.10192e-06, 5.804181e-06, 
    6.596293e-06, 8.094788e-06, 1.078934e-05, 1.127378e-05, 9.513725e-06,
  5.769432e-06, 7.088756e-06, 7.337896e-06, 6.162573e-06, 4.062126e-06, 
    4.92311e-06, 4.865622e-06, 3.347988e-06, 2.723711e-06, 3.522173e-06, 
    4.001166e-06, 6.903516e-06, 6.031499e-06, 7.56224e-06, 8.010244e-06,
  6.537644e-06, 3.723585e-06, 3.2489e-06, 4.594034e-06, 4.262301e-06, 
    4.527613e-06, 5.542713e-06, 5.825723e-06, 6.245515e-06, 3.982542e-06, 
    6.905008e-06, 4.946588e-06, 7.830786e-06, 9.144809e-06, 5.890073e-06,
  9.683069e-06, 3.202398e-06, 4.513509e-06, 3.919265e-06, 5.241509e-06, 
    5.245582e-06, 1.62051e-06, 3.700279e-06, 4.723562e-06, 7.025314e-06, 
    6.657803e-06, 6.735659e-06, 5.802306e-06, 7.784447e-06, 5.307815e-06,
  1.81597e-05, 9.479885e-06, 4.054947e-06, 1.329356e-06, 1.584702e-06, 
    2.123759e-06, 2.584489e-06, 3.593775e-06, 3.904576e-06, 4.860238e-06, 
    1.474541e-06, 2.45144e-06, 2.982508e-06, 2.71422e-06, 1.440124e-06,
  2.971508e-05, 2.627203e-05, 1.073654e-05, 7.89398e-06, 7.869886e-06, 
    5.492306e-06, 2.989553e-06, 3.21197e-06, 2.078645e-06, 5.284483e-06, 
    6.748019e-06, 5.840046e-06, 3.814277e-06, 4.113042e-06, 1.787226e-06,
  2.775377e-05, 2.164084e-05, 1.383047e-05, 7.414896e-06, 7.6112e-06, 
    1.543588e-05, 9.538773e-06, 1.069333e-05, 1.110205e-05, 1.996305e-05, 
    1.307542e-05, 1.210039e-05, 1.193641e-05, 1.033521e-05, 7.732589e-06,
  1.446125e-05, 1.686573e-05, 1.656272e-05, 2.130035e-05, 1.466992e-05, 
    1.60955e-05, 1.903363e-05, 2.271968e-05, 2.413395e-05, 2.862093e-05, 
    2.944057e-05, 3.308229e-05, 5.680903e-05, 2.816015e-05, 2.654953e-05,
  5.798336e-06, 8.28612e-06, 8.132191e-06, 1.504747e-05, 2.043284e-05, 
    1.74531e-05, 2.113965e-05, 1.753885e-05, 2.182633e-05, 2.720956e-05, 
    2.925029e-05, 3.460481e-05, 2.343336e-05, 3.175944e-05, 4.44277e-05,
  4.70796e-06, 6.533995e-06, 6.693053e-06, 9.04819e-06, 8.748184e-06, 
    8.081834e-06, 1.043715e-05, 7.148278e-06, 8.665193e-06, 6.142331e-06, 
    6.032099e-06, 6.998765e-06, 1.583513e-05, 1.520076e-05, 1.552425e-05,
  8.163816e-06, 8.789309e-06, 7.132399e-06, 1.183744e-05, 1.316665e-05, 
    1.022129e-05, 7.868143e-06, 7.344829e-06, 1.084384e-05, 7.014162e-06, 
    4.992073e-06, 8.769885e-06, 6.756668e-06, 8.774476e-06, 1.299089e-05,
  1.585199e-05, 6.667534e-06, 8.965643e-06, 4.868745e-06, 6.858604e-06, 
    9.437881e-06, 8.988928e-06, 6.269751e-06, 3.838694e-06, 6.096349e-06, 
    6.644304e-06, 6.487294e-06, 6.920272e-06, 9.397989e-06, 8.54634e-06,
  4.752824e-05, 5.980784e-06, 8.464898e-06, 8.262206e-06, 5.695832e-06, 
    5.232086e-06, 6.386502e-06, 5.673484e-06, 6.692935e-06, 5.228646e-06, 
    6.216469e-06, 7.602435e-06, 7.303121e-06, 7.146224e-06, 6.829417e-06,
  0.0001721582, 2.494496e-05, 6.275931e-06, 6.63345e-06, 6.630645e-06, 
    5.726164e-06, 1.815415e-06, 4.668064e-06, 5.986836e-06, 3.611808e-06, 
    2.533362e-06, 7.186812e-06, 9.252727e-06, 5.832027e-06, 4.608117e-06,
  0.0001733298, 9.0074e-05, 3.011952e-05, 6.895221e-06, 9.736899e-07, 
    1.217632e-06, 4.163385e-06, 5.057184e-06, 4.210037e-06, 4.830174e-06, 
    5.754533e-06, 3.316253e-06, 6.065013e-06, 4.193015e-06, 4.903839e-06,
  0.0001160647, 0.0001212285, 3.900238e-05, 3.777473e-05, 1.769965e-05, 
    2.574061e-06, 9.251809e-07, 7.349866e-06, 2.05884e-06, 2.6019e-06, 
    2.21351e-06, 3.833199e-06, 7.50465e-06, 2.188062e-06, 5.619987e-06,
  0.00015235, 0.0001277087, 0.0001025812, 9.099794e-05, 5.317368e-05, 
    1.687958e-05, 1.174684e-05, 5.877142e-06, 3.508065e-06, 4.28159e-06, 
    7.711182e-06, 6.647605e-06, 6.470036e-06, 5.312568e-06, 5.572291e-06,
  6.56932e-05, 9.536783e-05, 4.774562e-05, 4.799681e-05, 3.699777e-05, 
    2.750451e-05, 2.037612e-05, 2.920845e-05, 1.471946e-05, 1.253778e-05, 
    5.447072e-06, 4.875756e-06, 5.286637e-06, 4.681739e-06, 4.973343e-06,
  2.840994e-05, 2.078685e-05, 2.631602e-05, 3.331785e-05, 3.14838e-05, 
    4.103404e-05, 4.385837e-05, 4.542675e-05, 4.461973e-05, 2.960033e-05, 
    1.797159e-05, 1.41614e-05, 7.97623e-06, 5.918103e-06, 5.770767e-06,
  2.516707e-05, 3.80879e-05, 3.313364e-05, 2.370829e-05, 1.851352e-05, 
    1.172839e-05, 1.322255e-05, 1.07204e-05, 1.463769e-05, 2.917337e-05, 
    3.358732e-05, 2.474631e-05, 1.95496e-05, 1.835624e-05, 1.084197e-05,
  1.695591e-05, 3.94038e-06, 4.442432e-06, 5.663073e-06, 5.519389e-06, 
    6.694278e-06, 8.930101e-06, 9.189102e-06, 7.037156e-06, 6.156177e-06, 
    5.833049e-06, 6.303393e-06, 5.743208e-06, 8.551804e-06, 6.578404e-06,
  2.23035e-05, 7.191928e-06, 5.306798e-06, 6.09045e-06, 4.734272e-06, 
    4.44626e-06, 7.568043e-06, 1.01762e-05, 9.568394e-06, 6.105816e-06, 
    5.245567e-06, 5.235413e-06, 8.559919e-06, 5.680836e-06, 6.805855e-06,
  5.22775e-05, 6.71347e-06, 6.452536e-06, 5.404418e-06, 3.189732e-06, 
    1.090958e-05, 5.553576e-06, 3.765067e-06, 6.108186e-06, 6.92912e-06, 
    7.239257e-06, 6.598822e-06, 6.140074e-06, 5.738485e-06, 4.666159e-06,
  0.0001430667, 3.650703e-05, 6.926122e-06, 4.57707e-06, 1.58578e-06, 
    2.456727e-06, 2.220014e-06, 4.954807e-06, 5.034612e-06, 7.680633e-06, 
    7.888032e-06, 6.787045e-06, 7.150231e-06, 4.963226e-06, 4.717778e-06,
  0.000200104, 0.0001373908, 6.159655e-05, 2.110353e-05, 4.623045e-06, 
    1.0637e-06, 2.253996e-06, 1.907438e-06, 3.195116e-06, 6.718743e-06, 
    7.086775e-06, 6.012963e-06, 5.343868e-06, 6.255437e-06, 4.20584e-06,
  0.0003760408, 0.000234233, 0.0002113229, 9.020374e-05, 6.76163e-05, 
    8.758387e-06, 1.357018e-06, 1.59345e-06, 5.311268e-06, 2.769841e-06, 
    4.264167e-06, 4.214256e-06, 6.940134e-06, 7.01226e-06, 6.388908e-06,
  0.0003464631, 0.0002842579, 0.0001949891, 0.0001378297, 0.0001181197, 
    6.492962e-05, 2.232886e-05, 1.013056e-05, 3.03875e-06, 2.178906e-06, 
    2.886163e-06, 4.292504e-06, 6.491751e-06, 8.505519e-06, 1.050975e-05,
  0.0002532709, 0.000222274, 0.0002917169, 0.0001769177, 0.0001534281, 
    5.330671e-05, 7.167919e-05, 4.991295e-05, 4.152595e-06, 3.708522e-06, 
    2.026156e-06, 2.396358e-06, 3.534437e-06, 5.617376e-06, 7.565449e-06,
  0.0001468381, 0.0002043002, 0.0002190217, 0.000203249, 0.0002303965, 
    0.0001220011, 7.395227e-05, 0.0001068314, 2.767662e-05, 1.416983e-05, 
    5.517325e-06, 2.359964e-06, 1.937565e-06, 2.502334e-06, 3.034803e-06,
  8.909549e-05, 0.0001128875, 0.0001729436, 0.0001967696, 0.0001968034, 
    0.0002338122, 0.0001336715, 7.912547e-05, 0.0001065187, 4.593771e-05, 
    2.538453e-05, 1.200647e-05, 3.436264e-06, 7.758977e-06, 1.217413e-06,
  3.156681e-06, 3.89448e-06, 3.434752e-06, 4.657759e-06, 3.661667e-06, 
    4.017673e-06, 2.318858e-06, 2.019116e-06, 1.343763e-06, 1.431573e-06, 
    1.88356e-06, 2.454024e-06, 2.922656e-06, 3.092645e-06, 3.162532e-06,
  6.852437e-06, 4.826996e-06, 3.450295e-06, 4.660085e-06, 5.214377e-06, 
    6.170201e-06, 4.40645e-06, 2.578426e-06, 1.849504e-06, 2.118796e-06, 
    2.623116e-06, 2.693621e-06, 2.94343e-06, 2.286135e-06, 3.083979e-06,
  1.337094e-05, 9.235017e-06, 5.980099e-06, 4.819781e-06, 2.963933e-06, 
    4.855761e-06, 4.049634e-06, 4.466388e-06, 5.354153e-06, 2.530256e-06, 
    2.690749e-06, 3.972456e-06, 3.624875e-06, 3.276062e-06, 2.574062e-06,
  1.577487e-05, 1.078483e-05, 8.00157e-06, 5.545643e-06, 3.121176e-06, 
    2.920019e-06, 2.831817e-06, 2.169224e-06, 3.888463e-06, 3.293841e-06, 
    2.909227e-06, 4.378752e-06, 4.174974e-06, 4.403753e-06, 5.360104e-06,
  5.561279e-05, 3.763562e-05, 1.663073e-05, 3.160375e-06, 3.043133e-06, 
    4.135046e-06, 4.453763e-06, 3.162382e-06, 3.766105e-06, 3.427808e-06, 
    3.380143e-06, 3.069385e-06, 4.296386e-06, 4.487122e-06, 6.125583e-06,
  0.0004684302, 0.0005690593, 0.0003677317, 0.0001248675, 4.701028e-06, 
    3.81884e-06, 4.399841e-06, 3.63849e-06, 4.994288e-06, 5.16499e-06, 
    3.765277e-06, 4.790762e-06, 4.230892e-06, 4.683407e-06, 5.36793e-06,
  0.0007232654, 0.001040588, 0.0009350845, 0.0004906895, 0.0001449584, 
    8.390509e-06, 3.398844e-06, 3.745402e-06, 5.115505e-06, 7.719904e-06, 
    8.000885e-06, 9.081928e-06, 8.787232e-06, 7.87828e-06, 8.374992e-06,
  0.0003653914, 0.0006545925, 0.0009588298, 0.0007602573, 0.0003070402, 
    0.000102499, 1.734002e-05, 4.269118e-06, 2.971413e-06, 4.596993e-06, 
    5.804908e-06, 5.951509e-06, 8.593775e-06, 1.045115e-05, 1.204414e-05,
  0.0001534629, 0.0003541888, 0.0006700752, 0.0007793299, 0.0005695385, 
    0.0002229447, 8.737162e-05, 2.262476e-05, 6.206008e-06, 1.833701e-06, 
    2.469819e-06, 2.876878e-06, 3.579979e-06, 3.68274e-06, 4.124959e-06,
  7.371179e-05, 0.0001309485, 0.0002674962, 0.0005274014, 0.0007550413, 
    0.0004981961, 0.0001335841, 7.477666e-05, 4.430356e-05, 1.043018e-05, 
    4.588951e-06, 6.063964e-06, 5.680427e-06, 6.085869e-06, 5.844972e-06,
  5.892673e-06, 6.148328e-06, 4.654662e-06, 2.716604e-06, 1.327753e-06, 
    7.743178e-07, 1.32791e-07, 3.149012e-07, 8.749903e-07, 3.075671e-06, 
    4.718071e-06, 6.365807e-06, 5.985994e-06, 7.417835e-06, 6.196037e-06,
  5.320592e-06, 5.038215e-06, 4.432648e-06, 4.500441e-06, 3.249404e-06, 
    1.929644e-06, 1.425393e-06, 1.880272e-06, 9.601596e-07, 5.640122e-07, 
    8.953901e-07, 1.959126e-06, 1.908829e-06, 2.706196e-06, 3.434847e-06,
  5.399469e-06, 4.998431e-06, 3.888825e-06, 4.565872e-06, 4.191228e-06, 
    3.449827e-06, 2.946002e-06, 3.006058e-06, 1.615596e-06, 2.34246e-06, 
    1.063929e-06, 9.391722e-07, 5.316954e-07, 9.293801e-07, 8.741064e-07,
  9.771634e-06, 8.211304e-06, 5.604368e-06, 3.374192e-06, 3.870822e-06, 
    2.794926e-06, 2.735174e-06, 3.489132e-06, 3.112833e-06, 2.887945e-06, 
    2.511424e-06, 1.903263e-06, 1.443372e-06, 6.559798e-07, 4.399044e-07,
  1.48229e-05, 1.456325e-05, 1.333938e-05, 8.734341e-06, 4.700431e-06, 
    4.097471e-06, 3.031642e-06, 4.324316e-06, 4.875898e-06, 6.860842e-06, 
    7.074128e-06, 6.01722e-06, 5.727825e-06, 6.344801e-06, 4.946101e-06,
  2.335498e-05, 2.044745e-05, 1.983115e-05, 2.094564e-05, 1.755166e-05, 
    1.562596e-05, 1.015873e-05, 7.577331e-06, 6.972597e-06, 7.368486e-06, 
    6.692045e-06, 7.589652e-06, 8.296704e-06, 8.916884e-06, 8.412747e-06,
  0.0001177258, 0.000152352, 0.0001381513, 0.0001146462, 6.436647e-05, 
    6.003055e-06, 5.138652e-06, 3.998452e-06, 4.202109e-06, 3.706051e-06, 
    3.528978e-06, 3.246543e-06, 4.239506e-06, 4.638435e-06, 4.954088e-06,
  0.0002161762, 0.0002813465, 0.0003172267, 0.0003882408, 0.0003285899, 
    0.0001663056, 5.441052e-05, 4.95788e-05, 4.775635e-05, 3.795419e-05, 
    1.916087e-05, 5.491237e-06, 8.72936e-07, 9.451273e-07, 3.406344e-06,
  0.0001666099, 0.0002543538, 0.000419308, 0.0005752806, 0.0005258533, 
    0.000387483, 0.0002504091, 0.0002105855, 0.0002472261, 0.0002181489, 
    0.0001576283, 8.428661e-05, 2.547014e-05, 1.404812e-05, 1.493216e-05,
  7.635788e-05, 0.000174441, 0.0002125331, 0.0005544024, 0.0006254196, 
    0.0004796289, 0.0004262322, 0.0004276591, 0.0004474007, 0.0003964306, 
    0.0003288107, 0.0001746243, 6.049339e-05, 3.984318e-05, 3.531334e-05,
  4.184482e-06, 5.471285e-06, 6.53405e-06, 6.805675e-06, 8.407721e-06, 
    7.478641e-06, 7.787214e-06, 6.060422e-06, 7.420142e-06, 5.796667e-06, 
    6.628224e-06, 4.793498e-06, 4.898287e-06, 1.229352e-06, 1.069299e-06,
  1.928152e-06, 2.671952e-06, 3.179757e-06, 3.277353e-06, 3.894417e-06, 
    4.778048e-06, 2.5314e-06, 6.069113e-07, 5.407351e-07, 1.93372e-07, 
    9.515944e-08, 1.510144e-07, 2.972447e-07, 2.271893e-07, 3.259449e-07,
  2.262288e-06, 2.767314e-06, 1.645183e-06, 1.240386e-06, 8.948062e-07, 
    9.047257e-07, 7.162612e-07, 1.590125e-06, 1.620116e-07, 6.698287e-07, 
    9.57289e-08, 2.192073e-07, 1.996587e-07, 1.577668e-08, 2.601176e-07,
  2.467308e-06, 2.615684e-06, 2.402501e-06, 2.448789e-06, 1.822047e-06, 
    1.627834e-06, 1.488679e-06, 1.895659e-06, 2.292061e-06, 1.801191e-07, 
    8.118931e-07, 1.181442e-06, 2.424171e-06, 3.871972e-06, 5.70777e-06,
  3.18525e-06, 3.168902e-06, 2.93638e-06, 3.964349e-06, 3.166936e-06, 
    3.375062e-06, 2.654399e-06, 3.040844e-06, 3.672642e-06, 3.642543e-06, 
    4.933515e-06, 9.896272e-06, 1.128958e-05, 1.519568e-05, 1.676285e-05,
  3.092845e-06, 2.442818e-06, 1.999538e-06, 3.729487e-06, 3.35723e-06, 
    3.678394e-06, 4.105835e-06, 6.532499e-06, 1.044363e-05, 1.582711e-05, 
    2.35427e-05, 2.253314e-05, 2.239009e-05, 1.683696e-05, 1.084753e-05,
  2.178742e-06, 1.598046e-06, 1.826589e-06, 3.377018e-06, 5.512422e-06, 
    5.142716e-06, 4.296386e-06, 4.964204e-06, 8.347038e-06, 1.232191e-05, 
    1.797459e-05, 2.133078e-05, 2.419527e-05, 4.683681e-05, 0.0001076165,
  2.196909e-06, 6.594103e-07, 1.229223e-06, 2.248279e-06, 3.108758e-06, 
    2.210679e-06, 3.881074e-06, 6.402554e-06, 2.220807e-05, 0.00010605, 
    0.0002412865, 0.0003000528, 0.0003200639, 0.0003374417, 0.0003277522,
  1.218547e-06, 8.943338e-07, 3.653549e-07, 8.953822e-07, 1.996225e-06, 
    4.727083e-06, 1.332508e-05, 3.361881e-05, 9.298372e-05, 0.0002517153, 
    0.000387514, 0.0004708272, 0.0004881706, 0.00039308, 0.0002592375,
  1.25925e-06, 1.979774e-06, 3.780577e-06, 5.262173e-06, 6.161575e-06, 
    2.119424e-05, 5.432891e-05, 9.769489e-05, 0.0001420653, 0.0002233314, 
    0.0002846761, 0.0003179094, 0.0003117953, 0.0002274107, 0.0002524942,
  9.561025e-06, 1.370326e-05, 1.492922e-05, 1.853264e-05, 1.981107e-05, 
    2.03773e-05, 2.065093e-05, 2.270159e-05, 2.768018e-05, 3.099297e-05, 
    3.77855e-05, 4.543856e-05, 5.221091e-05, 5.529227e-05, 5.790044e-05,
  7.130974e-06, 1.035748e-05, 1.605672e-05, 1.854696e-05, 2.221405e-05, 
    2.074265e-05, 2.247856e-05, 2.490169e-05, 2.839362e-05, 2.99555e-05, 
    3.620908e-05, 3.615489e-05, 4.697836e-05, 5.309013e-05, 6.276881e-05,
  5.138531e-06, 6.601655e-06, 9.348772e-06, 1.435926e-05, 1.766048e-05, 
    1.971312e-05, 1.634449e-05, 1.995925e-05, 2.402659e-05, 2.711482e-05, 
    2.956292e-05, 3.350294e-05, 3.37841e-05, 4.043416e-05, 5.188325e-05,
  5.787143e-06, 6.242503e-06, 6.484499e-06, 7.386135e-06, 1.071667e-05, 
    1.388692e-05, 1.27603e-05, 1.570075e-05, 1.803723e-05, 1.950716e-05, 
    2.005717e-05, 2.209949e-05, 2.698957e-05, 3.367435e-05, 3.358986e-05,
  4.17604e-06, 3.774576e-06, 5.360489e-06, 6.962161e-06, 8.516046e-06, 
    8.315359e-06, 1.087649e-05, 1.381172e-05, 1.406417e-05, 1.4802e-05, 
    1.540975e-05, 1.74216e-05, 1.782225e-05, 2.093483e-05, 2.585674e-05,
  3.238966e-06, 3.150709e-06, 3.927486e-06, 4.427857e-06, 5.532835e-06, 
    7.306136e-06, 9.722479e-06, 1.048417e-05, 1.112716e-05, 1.203934e-05, 
    1.250077e-05, 1.334179e-05, 1.633997e-05, 1.798469e-05, 1.826615e-05,
  2.291883e-06, 3.224774e-06, 3.599246e-06, 4.694567e-06, 5.225983e-06, 
    5.596859e-06, 7.305183e-06, 7.61173e-06, 1.01834e-05, 1.074573e-05, 
    1.039197e-05, 1.197006e-05, 1.290457e-05, 1.430836e-05, 1.627017e-05,
  1.527738e-06, 2.885499e-06, 2.822414e-06, 3.580208e-06, 4.011867e-06, 
    5.158241e-06, 6.57684e-06, 6.875163e-06, 7.316059e-06, 8.178352e-06, 
    9.510253e-06, 1.138292e-05, 1.513474e-05, 1.607687e-05, 1.730492e-05,
  1.259221e-06, 1.215467e-06, 1.481944e-06, 2.277623e-06, 3.177459e-06, 
    4.486028e-06, 5.917255e-06, 6.09117e-06, 6.781879e-06, 1.135667e-05, 
    9.879634e-06, 1.173367e-05, 1.363445e-05, 1.516887e-05, 1.688313e-05,
  3.481542e-07, 8.12876e-08, 1.492214e-06, 1.755472e-06, 2.536015e-06, 
    2.633954e-06, 3.267387e-06, 3.679542e-06, 4.882394e-06, 6.872624e-06, 
    8.927566e-06, 9.87332e-06, 1.029433e-05, 1.145842e-05, 1.465064e-05,
  9.003653e-06, 7.298934e-06, 5.114901e-06, 5.223135e-06, 2.323199e-06, 
    1.670943e-06, 1.426943e-06, 2.155789e-06, 2.267869e-06, 2.817476e-06, 
    2.085641e-06, 2.018956e-06, 3.496252e-06, 5.784575e-06, 8.951868e-06,
  9.253459e-06, 6.142076e-06, 7.370259e-06, 6.230282e-06, 4.534062e-06, 
    1.316698e-06, 1.410348e-06, 1.506759e-06, 2.212186e-06, 1.951994e-06, 
    2.4642e-06, 1.425596e-06, 3.218166e-06, 3.886678e-06, 4.137068e-06,
  8.4327e-06, 1.086682e-05, 9.875439e-06, 9.918562e-06, 7.54396e-06, 
    3.536395e-06, 1.911929e-06, 1.541336e-06, 2.148028e-06, 1.23214e-06, 
    2.069035e-06, 1.508508e-06, 1.733806e-06, 2.383117e-06, 3.189574e-06,
  5.142315e-06, 3.718145e-06, 7.222764e-06, 1.17017e-05, 1.117238e-05, 
    3.323695e-06, 1.560788e-06, 1.665885e-06, 1.897552e-06, 2.091344e-06, 
    1.497981e-06, 1.233625e-06, 1.505636e-06, 1.120461e-06, 1.233135e-06,
  2.957648e-06, 3.184857e-06, 3.979439e-06, 5.915198e-06, 1.243185e-05, 
    4.525577e-06, 1.60185e-06, 2.38646e-06, 2.692949e-06, 1.856557e-06, 
    1.971116e-06, 1.282954e-06, 1.158323e-06, 1.548045e-06, 1.495557e-06,
  2.072564e-06, 1.208385e-06, 4.645323e-06, 6.398368e-06, 4.072157e-06, 
    2.204865e-06, 2.933454e-06, 5.43673e-06, 6.466189e-06, 3.808035e-06, 
    2.088577e-06, 6.704903e-07, 1.368718e-06, 1.780961e-06, 6.40532e-07,
  2.108186e-06, 1.834638e-06, 1.090613e-06, 1.779755e-06, 3.372614e-06, 
    3.67096e-06, 2.630368e-06, 9.79778e-06, 1.013775e-05, 9.270118e-06, 
    3.566246e-06, 4.300128e-06, 1.750389e-06, 1.204668e-06, 6.995936e-07,
  6.022365e-06, 3.522631e-06, 3.293749e-06, 3.122405e-06, 2.063004e-06, 
    4.292103e-06, 3.616863e-06, 4.198567e-06, 1.098852e-05, 9.449953e-06, 
    9.198087e-06, 5.427328e-06, 4.917074e-06, 5.812473e-07, 4.650212e-07,
  3.6631e-06, 3.883116e-06, 4.227872e-06, 4.956762e-06, 5.197697e-06, 
    5.240336e-06, 6.578962e-06, 5.486706e-06, 5.005538e-06, 5.799805e-06, 
    7.693329e-06, 1.058236e-05, 7.725894e-06, 2.581356e-06, 1.75471e-06,
  2.463393e-06, 1.940779e-06, 2.516478e-06, 3.683887e-06, 5.242854e-06, 
    6.068099e-06, 6.437543e-06, 4.850102e-06, 4.632333e-06, 3.650765e-06, 
    5.04112e-06, 8.502883e-06, 1.028829e-05, 6.120513e-06, 5.53382e-06,
  1.291362e-06, 2.15337e-06, 5.603521e-06, 6.423205e-06, 7.925988e-06, 
    9.017048e-06, 9.713191e-06, 9.967129e-06, 1.009843e-05, 1.026972e-05, 
    9.517409e-06, 7.626213e-06, 7.491215e-06, 1.140543e-05, 7.411514e-06,
  6.74275e-07, 1.462725e-06, 2.933996e-06, 4.971691e-06, 6.278889e-06, 
    6.566224e-06, 7.135347e-06, 8.397022e-06, 7.000695e-06, 8.323644e-06, 
    7.782327e-06, 8.655238e-06, 7.137254e-06, 5.145012e-06, 7.166968e-06,
  4.916542e-07, 1.188556e-06, 2.338395e-06, 3.649447e-06, 4.746269e-06, 
    5.635336e-06, 7.39423e-06, 6.176499e-06, 7.379636e-06, 8.69423e-06, 
    6.381067e-06, 8.158614e-06, 6.749924e-06, 4.537679e-06, 4.593421e-06,
  3.19787e-07, 1.16409e-06, 2.010046e-06, 2.500017e-06, 3.009308e-06, 
    5.77747e-06, 4.172816e-06, 4.865051e-06, 7.307616e-06, 7.383449e-06, 
    6.380402e-06, 5.345771e-06, 4.461801e-06, 3.292659e-06, 3.182746e-06,
  5.306578e-07, 1.190511e-06, 3.522882e-06, 3.671987e-06, 1.841599e-06, 
    4.302321e-06, 3.534501e-06, 3.276482e-06, 5.374071e-06, 6.473598e-06, 
    6.713451e-06, 4.881641e-06, 4.61482e-06, 3.56953e-06, 3.04055e-06,
  3.406777e-07, 7.905201e-07, 3.528005e-06, 1.853665e-06, 1.915163e-06, 
    2.120054e-06, 2.833403e-06, 4.157444e-06, 5.125685e-06, 5.470844e-06, 
    8.196331e-06, 7.21448e-06, 6.779283e-06, 4.890845e-06, 4.898666e-06,
  4.592238e-07, 1.214022e-06, 2.445817e-06, 2.895627e-06, 2.597848e-06, 
    2.659995e-06, 5.553317e-06, 4.762088e-06, 3.137513e-06, 4.868895e-06, 
    6.74596e-06, 1.007785e-05, 8.829345e-06, 6.856162e-06, 7.721854e-06,
  5.682252e-07, 6.945867e-07, 1.964327e-06, 4.680002e-06, 4.492507e-06, 
    4.509945e-06, 3.912123e-06, 3.223764e-06, 5.456369e-06, 4.108182e-06, 
    4.610884e-06, 5.800508e-06, 7.702019e-06, 8.144761e-06, 9.563974e-06,
  5.873629e-07, 7.11829e-07, 1.694208e-06, 4.902774e-06, 6.807102e-06, 
    8.431051e-06, 8.365843e-06, 6.414752e-06, 4.593321e-06, 2.694047e-06, 
    2.871489e-06, 4.777489e-06, 7.34332e-06, 8.24717e-06, 8.397333e-06,
  2.419919e-07, 9.662834e-07, 2.520262e-06, 6.892333e-06, 1.034999e-05, 
    1.154612e-05, 1.328507e-05, 1.270331e-05, 1.008133e-05, 3.447505e-06, 
    5.06283e-06, 3.094493e-06, 4.179364e-06, 7.501875e-06, 9.102766e-06,
  6.370728e-05, 9.751691e-05, 9.788597e-05, 8.276263e-05, 5.864146e-05, 
    3.164494e-05, 1.265838e-05, 5.984091e-06, 5.006466e-06, 6.927368e-06, 
    1.269129e-05, 1.165468e-05, 4.426198e-06, 1.083103e-06, 5.262122e-07,
  6.383405e-05, 8.672443e-05, 7.205042e-05, 4.764858e-05, 2.546189e-05, 
    8.853607e-06, 4.407746e-06, 5.180131e-06, 7.070259e-06, 9.022899e-06, 
    8.222042e-06, 6.207075e-06, 2.563029e-06, 6.295732e-07, 6.945318e-07,
  4.63324e-05, 4.709474e-05, 3.984802e-05, 2.182379e-05, 5.843879e-06, 
    4.521685e-06, 3.679549e-06, 6.025859e-06, 8.374607e-06, 7.126496e-06, 
    5.720956e-06, 3.138263e-06, 2.728024e-06, 1.068443e-06, 6.599078e-07,
  1.564065e-05, 2.2932e-05, 1.647404e-05, 3.669622e-06, 4.141963e-06, 
    6.35886e-06, 8.19154e-06, 6.931256e-06, 4.937502e-06, 2.652868e-06, 
    2.661931e-06, 3.417915e-06, 2.985545e-06, 1.216519e-06, 4.653719e-07,
  1.835464e-05, 2.467037e-05, 4.683922e-07, 2.392485e-06, 4.963882e-06, 
    6.909482e-06, 5.859406e-06, 5.104939e-06, 1.812267e-06, 9.637457e-07, 
    2.733547e-06, 5.820786e-06, 9.214871e-06, 5.607717e-06, 5.826726e-07,
  9.163412e-06, 6.299398e-06, 1.681547e-06, 2.885171e-06, 4.189777e-06, 
    5.231855e-06, 3.11189e-06, 2.813516e-06, 1.635163e-06, 1.139745e-06, 
    4.224887e-06, 1.502557e-05, 2.972069e-05, 3.808501e-05, 1.417524e-05,
  6.890323e-08, 7.232052e-08, 1.355692e-06, 1.939124e-06, 3.757e-06, 
    2.542034e-06, 2.306849e-06, 3.96427e-06, 2.71813e-06, 1.536494e-06, 
    6.81498e-06, 3.107928e-05, 6.639554e-05, 7.479641e-05, 4.18616e-05,
  8.839951e-09, 1.773385e-07, 2.744723e-07, 8.651974e-07, 1.12844e-06, 
    1.634412e-06, 2.910733e-06, 3.580503e-06, 6.061336e-06, 1.333803e-06, 
    1.312383e-05, 4.22368e-05, 7.054881e-05, 5.854556e-05, 2.382327e-05,
  1.628529e-07, 1.030545e-07, 7.22498e-07, 1.976576e-06, 6.717303e-06, 
    1.059893e-05, 1.926409e-05, 2.572769e-05, 1.838567e-05, 6.750422e-06, 
    1.697888e-05, 4.600007e-05, 4.995646e-05, 1.909716e-05, 2.545671e-06,
  1.672528e-08, 1.061075e-07, 9.263969e-07, 2.769575e-06, 1.239008e-05, 
    1.612739e-05, 2.597943e-05, 3.898968e-05, 5.330367e-05, 5.239952e-06, 
    2.857504e-05, 2.139906e-05, 2.124097e-05, 8.164004e-06, 1.589198e-06,
  1.101411e-05, 2.439098e-05, 5.44494e-05, 0.0001069729, 0.0001572553, 
    0.0001847234, 0.0001941165, 0.0001950409, 0.0001605843, 0.0001446704, 
    0.000126839, 0.0001167543, 0.0001082232, 8.900635e-05, 7.038622e-05,
  2.111503e-05, 4.526348e-05, 8.05399e-05, 0.0001273863, 0.0001627885, 
    0.0001707057, 0.0001229248, 9.54956e-05, 8.122833e-05, 7.37855e-05, 
    7.631258e-05, 7.002562e-05, 7.668285e-05, 7.520452e-05, 6.964197e-05,
  3.787775e-05, 5.279732e-05, 7.964679e-05, 8.899195e-05, 9.760738e-05, 
    7.954628e-05, 5.749486e-05, 4.316719e-05, 4.369966e-05, 4.540967e-05, 
    4.46018e-05, 4.979724e-05, 5.592057e-05, 6.181915e-05, 6.981371e-05,
  3.539836e-05, 3.341023e-05, 4.009901e-05, 5.109411e-05, 4.632072e-05, 
    3.840612e-05, 2.412683e-05, 2.31443e-05, 2.730739e-05, 3.19269e-05, 
    3.539272e-05, 4.521406e-05, 5.821693e-05, 7.273439e-05, 8.258816e-05,
  4.266883e-05, 3.963411e-05, 5.683e-05, 3.692419e-05, 2.60821e-05, 
    2.498475e-05, 2.596766e-05, 2.23584e-05, 2.567963e-05, 2.205308e-05, 
    3.208597e-05, 4.24967e-05, 5.828224e-05, 8.308461e-05, 0.0001150533,
  8.733012e-05, 9.353019e-05, 7.515257e-05, 5.96391e-05, 4.701033e-05, 
    3.698617e-05, 2.851448e-05, 2.047016e-05, 2.127784e-05, 1.696684e-05, 
    2.183161e-05, 2.940842e-05, 4.367317e-05, 7.23921e-05, 0.0001194291,
  0.0001567957, 0.000147296, 0.0001135113, 7.800095e-05, 5.064883e-05, 
    3.469301e-05, 3.034768e-05, 2.512606e-05, 2.696206e-05, 2.856496e-05, 
    2.458223e-05, 2.401212e-05, 3.608354e-05, 5.73139e-05, 8.202882e-05,
  0.0002184907, 0.0001857212, 0.0001430196, 0.0001056961, 6.936065e-05, 
    4.725145e-05, 3.915844e-05, 2.545718e-05, 2.341894e-05, 1.877705e-05, 
    2.003856e-05, 2.931642e-05, 3.90231e-05, 5.871472e-05, 7.689346e-05,
  0.0002274607, 0.0001975481, 0.0001582891, 0.0001237995, 9.630107e-05, 
    8.106932e-05, 5.367785e-05, 3.181896e-05, 3.222233e-05, 1.503508e-05, 
    2.375386e-05, 4.0464e-05, 8.075115e-05, 0.0001021246, 0.0001187849,
  0.0001821527, 0.0001560661, 0.0001140956, 8.487488e-05, 5.727509e-05, 
    5.182076e-05, 4.64556e-05, 4.649936e-05, 3.96315e-05, 3.742247e-05, 
    3.926723e-05, 6.919921e-05, 0.000104967, 0.0001228177, 0.0001185254,
  8.586982e-06, 9.544436e-06, 1.022456e-05, 1.117244e-05, 9.658002e-06, 
    1.084821e-05, 1.008278e-05, 1.106655e-05, 7.73998e-06, 1.132686e-05, 
    9.777877e-06, 1.262296e-05, 1.174981e-05, 1.334055e-05, 1.935897e-05,
  1.06924e-05, 1.118259e-05, 1.135652e-05, 1.093188e-05, 1.056456e-05, 
    9.762082e-06, 7.647534e-06, 7.090479e-06, 9.930885e-06, 1.265592e-05, 
    1.105309e-05, 1.310674e-05, 9.9993e-06, 1.286808e-05, 1.323982e-05,
  1.295378e-05, 9.765704e-06, 1.004889e-05, 9.228415e-06, 8.094924e-06, 
    8.15368e-06, 6.198778e-06, 7.13949e-06, 8.283912e-06, 1.191659e-05, 
    9.396065e-06, 1.363432e-05, 1.210503e-05, 1.233845e-05, 1.366269e-05,
  1.758499e-05, 1.399182e-05, 1.219828e-05, 9.753145e-06, 8.018128e-06, 
    7.44828e-06, 5.884905e-06, 7.735652e-06, 1.140195e-05, 3.728108e-06, 
    1.304081e-05, 1.622281e-05, 1.312618e-05, 1.763651e-05, 1.51083e-05,
  1.211679e-05, 1.307079e-05, 1.374393e-05, 1.550321e-05, 1.303971e-05, 
    1.084003e-05, 1.209331e-05, 1.213105e-05, 8.644061e-06, 6.762854e-06, 
    1.493155e-05, 1.686643e-05, 1.879215e-05, 1.763815e-05, 1.657034e-05,
  1.868557e-05, 1.70982e-05, 1.175762e-05, 1.101382e-05, 8.42883e-06, 
    1.261471e-05, 1.60937e-05, 1.614305e-05, 1.164715e-05, 8.968623e-06, 
    1.671875e-05, 1.570224e-05, 1.67347e-05, 1.279472e-05, 1.136638e-05,
  1.932785e-05, 1.925276e-05, 1.764411e-05, 9.433551e-06, 8.610838e-06, 
    1.187539e-05, 1.337073e-05, 1.540948e-05, 1.36918e-05, 1.680482e-05, 
    1.91238e-05, 2.004155e-05, 1.679549e-05, 1.621811e-05, 1.103165e-05,
  1.358479e-05, 1.22255e-05, 1.292936e-05, 1.965211e-05, 1.716069e-05, 
    1.569394e-05, 1.400648e-05, 1.116798e-05, 1.283166e-05, 1.60539e-05, 
    1.625295e-05, 1.908532e-05, 1.661156e-05, 1.608875e-05, 1.625223e-05,
  1.339662e-05, 1.400681e-05, 1.400217e-05, 1.78217e-05, 1.60509e-05, 
    1.41583e-05, 1.249163e-05, 1.199727e-05, 1.213606e-05, 1.24405e-05, 
    1.158114e-05, 1.248674e-05, 1.431746e-05, 1.495095e-05, 1.764262e-05,
  5.580951e-05, 4.124554e-05, 3.603341e-05, 3.607012e-05, 3.521331e-05, 
    3.639677e-05, 2.892597e-05, 1.932251e-05, 1.530305e-05, 1.192354e-05, 
    1.449048e-05, 1.367693e-05, 1.251428e-05, 1.11347e-05, 1.251382e-05,
  1.184971e-05, 1.274373e-05, 7.270464e-06, 8.690876e-06, 7.579975e-06, 
    7.592957e-06, 6.304977e-06, 7.562132e-06, 7.225029e-06, 5.872868e-06, 
    5.667035e-06, 8.053386e-06, 6.799691e-06, 9.905965e-06, 8.55167e-06,
  1.627544e-05, 1.228847e-05, 1.212021e-05, 8.936846e-06, 6.968224e-06, 
    6.28377e-06, 5.028192e-06, 5.509766e-06, 5.449913e-06, 6.013322e-06, 
    5.438761e-06, 5.652374e-06, 5.920432e-06, 6.531416e-06, 5.730139e-06,
  1.958062e-05, 1.574152e-05, 1.441456e-05, 1.039645e-05, 5.65993e-06, 
    5.38072e-06, 6.195755e-06, 4.290624e-06, 5.70425e-06, 3.598574e-06, 
    5.773978e-06, 5.959628e-06, 6.862216e-06, 7.015632e-06, 5.67904e-06,
  2.202426e-05, 2.0416e-05, 1.58437e-05, 1.087561e-05, 6.070339e-06, 
    5.128588e-06, 4.796556e-06, 5.531608e-06, 3.957994e-06, 4.078388e-06, 
    3.619844e-06, 4.720594e-06, 5.428908e-06, 6.241474e-06, 5.988437e-06,
  4.702294e-05, 2.709275e-05, 1.751145e-05, 1.388209e-05, 1.413707e-05, 
    7.551334e-06, 6.659696e-06, 6.070557e-06, 5.383133e-06, 4.204808e-06, 
    3.504509e-06, 3.182159e-06, 4.750721e-06, 4.780803e-06, 6.11744e-06,
  0.000119176, 7.611216e-05, 3.896025e-05, 2.316718e-05, 1.046227e-05, 
    9.528075e-06, 8.563179e-06, 8.286567e-06, 9.406797e-06, 6.28881e-06, 
    6.196945e-06, 5.676067e-06, 5.370076e-06, 4.807806e-06, 5.243327e-06,
  0.0002610221, 0.0001858833, 0.0001244854, 7.642622e-05, 2.626537e-05, 
    6.132234e-06, 7.460113e-06, 9.611682e-06, 7.048261e-06, 8.984282e-06, 
    8.832853e-06, 7.100002e-06, 7.878031e-06, 6.061493e-06, 6.201362e-06,
  0.0004392596, 0.0003603477, 0.0002575581, 0.0001701942, 7.43803e-05, 
    8.294459e-06, 6.666173e-06, 8.887626e-06, 8.334357e-06, 1.155391e-05, 
    9.701921e-06, 8.007748e-06, 6.511362e-06, 6.194479e-06, 1.023922e-05,
  0.0005568559, 0.0005035065, 0.0004166913, 0.0002881976, 0.0001520524, 
    2.765381e-05, 1.318489e-05, 5.7547e-06, 6.654866e-06, 7.661451e-06, 
    8.668941e-06, 8.552089e-06, 8.580386e-06, 9.188985e-06, 1.110937e-05,
  0.0005857096, 0.0004995597, 0.0003929026, 0.0003132043, 0.0001907011, 
    8.388363e-05, 3.637219e-05, 9.978434e-06, 4.876888e-06, 7.640783e-06, 
    7.255834e-06, 7.798973e-06, 8.062526e-06, 7.827696e-06, 1.059966e-05,
  2.291283e-05, 1.40414e-05, 1.237733e-05, 1.119189e-05, 1.744195e-05, 
    1.802239e-05, 1.696363e-05, 1.200479e-05, 7.005523e-06, 8.274265e-06, 
    7.364354e-06, 8.624918e-06, 9.342642e-06, 1.062889e-05, 7.088105e-06,
  0.0001018353, 0.0001335266, 0.0001069658, 3.872826e-05, 1.395568e-05, 
    1.52497e-05, 1.763469e-05, 1.05281e-05, 5.826621e-06, 3.884306e-06, 
    5.633626e-06, 6.918642e-06, 6.239807e-06, 6.866899e-06, 5.158176e-06,
  0.0001762916, 0.0002173554, 0.0001953591, 9.473271e-05, 2.514107e-05, 
    1.298795e-05, 1.557338e-05, 8.217681e-06, 5.054062e-06, 2.99845e-06, 
    4.024358e-06, 5.255908e-06, 7.524822e-06, 6.047242e-06, 4.07297e-06,
  0.0001656131, 0.0001959932, 0.0001719855, 9.610662e-05, 3.211234e-05, 
    8.643852e-06, 1.367389e-05, 6.664514e-06, 3.322801e-06, 2.072666e-06, 
    2.342445e-06, 4.764255e-06, 5.033214e-06, 5.265459e-06, 4.014236e-06,
  0.0001122779, 0.0001009886, 7.025994e-05, 3.758437e-05, 1.158278e-05, 
    1.012975e-05, 8.985176e-06, 8.538354e-06, 5.497507e-06, 2.090819e-06, 
    1.889561e-06, 3.150888e-06, 3.402221e-06, 5.802925e-06, 5.074588e-06,
  0.0001063974, 7.093202e-05, 4.550876e-05, 2.241138e-05, 1.249127e-05, 
    8.553258e-06, 8.259465e-06, 9.226609e-06, 7.276701e-06, 5.954998e-06, 
    2.962579e-06, 2.313895e-06, 3.424039e-06, 4.839723e-06, 6.319961e-06,
  0.0001337031, 9.577506e-05, 8.151502e-05, 5.369472e-05, 2.754008e-05, 
    1.073454e-05, 7.823368e-06, 9.201258e-06, 1.196998e-05, 1.08175e-05, 
    5.994163e-06, 2.52107e-06, 2.400158e-06, 5.54227e-06, 5.584654e-06,
  0.0001145733, 0.0001007422, 9.51304e-05, 9.310854e-05, 6.750586e-05, 
    3.091881e-05, 1.293338e-05, 1.149616e-05, 1.12694e-05, 1.164121e-05, 
    9.458166e-06, 6.20551e-06, 3.648013e-06, 4.819019e-06, 5.007353e-06,
  6.707499e-05, 7.734045e-05, 7.733747e-05, 8.046569e-05, 7.90443e-05, 
    5.835e-05, 2.946188e-05, 1.450362e-05, 1.076494e-05, 1.081664e-05, 
    9.143363e-06, 7.736447e-06, 5.706941e-06, 3.625678e-06, 3.45674e-06,
  6.615506e-05, 6.716915e-05, 7.045164e-05, 6.72653e-05, 8.876721e-05, 
    7.59481e-05, 4.967533e-05, 2.507897e-05, 1.418982e-05, 8.375491e-06, 
    9.485923e-06, 8.682713e-06, 6.845498e-06, 4.644774e-06, 3.780385e-06,
  1.187517e-05, 3.491503e-05, 5.069329e-05, 0.0001011555, 0.0001837955, 
    0.0002560671, 0.0002762411, 0.0002771313, 0.0002383582, 0.0001918245, 
    0.000137427, 0.0001066686, 7.498121e-05, 7.005001e-05, 6.118572e-05,
  1.784116e-05, 6.057534e-05, 0.0001444183, 0.0002845925, 0.0003538094, 
    0.0003574485, 0.0003268275, 0.0003127699, 0.000282361, 0.0002327486, 
    0.0001783989, 0.0001352507, 0.0001028012, 7.099504e-05, 4.723177e-05,
  1.923197e-05, 7.943637e-05, 0.0001959249, 0.0003624749, 0.0004698085, 
    0.0004654013, 0.0004110329, 0.0003981635, 0.0003712937, 0.0003290341, 
    0.0002702022, 0.0002110861, 0.0001544552, 9.578017e-05, 3.914843e-05,
  2.490269e-05, 7.439785e-05, 0.0001782582, 0.0003099464, 0.0004174206, 
    0.0004524063, 0.0004253205, 0.0003996127, 0.0004012385, 0.0003627279, 
    0.0003233383, 0.0002614208, 0.0001796964, 9.666062e-05, 3.561364e-05,
  4.213256e-05, 4.927349e-05, 0.0001040379, 0.0001606065, 0.0002061774, 
    0.0002208783, 0.000222992, 0.0002413446, 0.0002745169, 0.0002870843, 
    0.000282689, 0.0002378359, 0.0001383349, 5.884399e-05, 1.931774e-05,
  4.264821e-05, 1.441407e-05, 3.616609e-05, 5.923638e-05, 7.740694e-05, 
    8.084847e-05, 7.967647e-05, 0.0001031904, 0.0001430556, 0.0001929698, 
    0.0002185899, 0.0002118054, 0.0001216664, 3.324483e-05, 7.118279e-06,
  2.674719e-05, 1.40962e-05, 2.185156e-05, 4.305748e-05, 5.291466e-05, 
    5.512673e-05, 6.451272e-05, 7.785783e-05, 9.8734e-05, 0.0001258333, 
    0.0001603621, 0.0001577886, 9.176244e-05, 3.564892e-05, 8.455049e-06,
  3.174676e-05, 5.432738e-05, 3.512618e-05, 4.301816e-05, 4.221862e-05, 
    4.744229e-05, 7.001297e-05, 7.828921e-05, 7.020515e-05, 5.980525e-05, 
    5.522467e-05, 4.721902e-05, 4.212203e-05, 2.340603e-05, 8.291352e-06,
  2.87962e-05, 4.590791e-05, 5.590317e-05, 3.669347e-05, 3.960029e-05, 
    4.012823e-05, 4.031173e-05, 3.228235e-05, 2.625316e-05, 2.612604e-05, 
    1.465232e-05, 1.209806e-05, 1.196495e-05, 9.415709e-06, 6.063535e-06,
  6.554562e-05, 6.67585e-05, 6.581484e-05, 7.940053e-05, 0.0001056484, 
    0.0001603313, 0.0001917656, 0.0001888308, 0.0001333178, 3.547371e-05, 
    4.902942e-06, 5.177993e-06, 4.183961e-06, 3.983613e-06, 2.204616e-06,
  4.776273e-05, 7.422396e-05, 7.787698e-05, 8.476614e-05, 3.842167e-05, 
    1.453327e-05, 7.956128e-06, 5.686859e-06, 5.603637e-06, 5.391659e-06, 
    3.886788e-06, 3.168688e-06, 4.578207e-06, 1.081283e-05, 2.047089e-05,
  1.653485e-05, 2.034812e-05, 2.622299e-05, 3.692439e-05, 1.112831e-05, 
    2.904488e-06, 4.464634e-06, 6.699365e-06, 5.043045e-06, 5.405393e-06, 
    4.07977e-06, 1.21767e-06, 3.231355e-06, 1.100222e-05, 3.613024e-05,
  3.558499e-06, 3.033854e-06, 1.725154e-06, 1.643223e-06, 1.659495e-06, 
    3.155988e-06, 3.961849e-06, 5.435103e-06, 5.547909e-06, 3.929038e-06, 
    6.52961e-07, 3.582713e-07, 1.783396e-06, 1.399307e-05, 8.905678e-05,
  3.365303e-07, 2.880077e-09, 7.306815e-08, 1.664022e-06, 2.749489e-06, 
    1.958766e-06, 7.381028e-07, 3.987691e-07, 1.046772e-06, 3.710934e-07, 
    1.978332e-07, 3.563966e-07, 4.456415e-06, 6.338402e-05, 0.0001180685,
  6.775335e-10, 1.562892e-08, 3.605916e-08, 1.512138e-07, 5.799345e-08, 
    3.392183e-08, 1.268545e-07, 2.179521e-07, 6.861701e-08, 1.108918e-08, 
    3.122173e-08, 7.226574e-07, 3.553474e-05, 0.0001015185, 0.0001173336,
  1.345695e-10, 1.079174e-09, 3.273274e-09, 5.710938e-08, 1.492649e-10, 
    1.671647e-10, 1.34357e-09, 1.367644e-07, 4.406219e-07, 1.182222e-08, 
    1.324455e-07, 1.398084e-05, 8.274502e-05, 0.0003291691, 0.0005386513,
  9.197261e-11, 1.040326e-10, 9.377602e-11, 3.690549e-09, 2.9776e-12, 
    4.682445e-11, 5.02943e-10, 9.147732e-09, 1.409254e-08, 1.307896e-06, 
    4.207818e-05, 0.0002064305, 0.0004289112, 0.0006101966, 0.0007012509,
  1.066148e-09, 1.459788e-09, 2.824142e-08, 1.081505e-08, 6.656231e-09, 
    3.556401e-09, 5.405876e-09, 7.859771e-07, 4.262805e-06, 3.328531e-05, 
    0.0001301224, 0.0002191835, 0.000228348, 0.0001794163, 0.0002023486,
  2.990779e-07, 9.004848e-08, 7.054899e-08, 1.766793e-07, 5.509765e-08, 
    3.914049e-08, 6.151577e-07, 2.43537e-06, 1.043081e-05, 3.683076e-05, 
    5.680942e-05, 2.027736e-05, 7.645875e-06, 3.779411e-05, 0.0001356486,
  3.507799e-05, 4.834542e-05, 4.259078e-05, 3.369301e-05, 3.379694e-05, 
    3.703685e-05, 1.313669e-05, 4.120518e-06, 9.247256e-06, 3.3856e-05, 
    7.800579e-06, 1.042829e-05, 3.095476e-05, 0.0001245296, 0.0003276905,
  1.418285e-05, 7.48439e-06, 1.288765e-05, 2.714554e-05, 6.5464e-05, 
    9.888784e-05, 0.0001165972, 0.0001224409, 0.0001166289, 0.000103117, 
    9.583192e-05, 7.861492e-05, 5.033156e-05, 2.756605e-05, 1.223132e-05,
  6.340056e-05, 4.13501e-05, 3.892534e-05, 4.180737e-05, 5.882316e-05, 
    9.009815e-05, 8.081368e-05, 6.452369e-05, 6.582629e-05, 5.995171e-05, 
    4.853394e-05, 3.949819e-05, 2.849073e-05, 1.834354e-05, 2.062856e-05,
  6.585568e-05, 6.992694e-05, 7.240674e-05, 5.031033e-05, 6.791105e-05, 
    4.652894e-05, 4.421023e-05, 3.62872e-05, 2.410659e-05, 3.229992e-05, 
    1.981638e-05, 2.011586e-05, 1.066075e-05, 1.239775e-05, 3.288297e-05,
  2.206434e-05, 2.473001e-05, 5.400482e-05, 4.917333e-05, 4.057092e-05, 
    3.319168e-05, 2.503179e-05, 1.59758e-05, 8.346561e-06, 1.306766e-05, 
    1.188422e-05, 1.09738e-05, 5.991659e-06, 1.027439e-05, 6.706244e-05,
  4.372064e-06, 1.04834e-05, 2.589292e-05, 2.996458e-05, 3.483255e-05, 
    3.222323e-05, 2.954579e-05, 1.948761e-05, 1.723628e-05, 1.436746e-05, 
    1.338595e-05, 1.133549e-05, 8.926117e-06, 2.720039e-05, 7.108242e-05,
  1.791329e-06, 1.898012e-06, 6.739641e-06, 1.615732e-05, 2.48486e-05, 
    4.664248e-05, 3.439824e-05, 4.105764e-05, 3.914874e-05, 3.010414e-05, 
    2.571598e-05, 2.055379e-05, 2.174735e-05, 3.533679e-05, 6.467881e-05,
  6.110882e-07, 1.431419e-06, 3.310431e-06, 6.675089e-06, 1.584383e-05, 
    2.422158e-05, 3.204534e-05, 4.523033e-05, 3.503878e-05, 3.982215e-05, 
    4.601187e-05, 5.506414e-05, 6.693287e-05, 5.317962e-05, 4.400339e-05,
  7.066314e-07, 1.612557e-06, 2.284721e-06, 7.063245e-06, 8.625519e-06, 
    1.381656e-05, 2.15756e-05, 2.706749e-05, 4.408835e-05, 4.703366e-05, 
    4.480048e-05, 5.270778e-05, 4.314552e-05, 1.93489e-05, 4.505449e-05,
  1.53141e-06, 1.364777e-06, 1.469257e-06, 2.407313e-06, 3.565872e-06, 
    5.721536e-06, 1.107783e-05, 1.706029e-05, 2.425907e-05, 2.991702e-05, 
    2.648622e-05, 4.969082e-05, 9.890126e-05, 0.0001262884, 0.0001617728,
  5.525999e-06, 3.333079e-06, 1.007827e-05, 1.602273e-05, 2.446957e-05, 
    6.903309e-05, 0.0001124307, 0.0001190239, 0.0001557242, 0.000211602, 
    0.0002343091, 0.0002697346, 0.0002822572, 0.0003007329, 0.0003039509,
  1.945852e-06, 1.720121e-06, 1.423826e-06, 2.738166e-06, 3.362356e-06, 
    7.03362e-06, 8.985104e-06, 9.005253e-06, 1.512872e-05, 2.385807e-05, 
    4.636545e-05, 8.909004e-05, 8.489739e-05, 8.432007e-05, 7.99073e-05,
  1.62217e-06, 1.568534e-06, 1.396393e-06, 2.401428e-06, 4.188869e-06, 
    6.093426e-06, 8.102988e-06, 8.425802e-06, 1.75823e-05, 2.113399e-05, 
    2.973475e-05, 6.837464e-05, 7.924209e-05, 6.441728e-05, 7.100019e-05,
  1.261234e-06, 8.758952e-07, 1.559303e-06, 2.666616e-06, 2.560759e-06, 
    4.31291e-06, 7.359862e-06, 1.097468e-05, 1.433475e-05, 1.47291e-05, 
    1.552857e-05, 2.222306e-05, 3.010974e-05, 3.441446e-05, 4.022269e-05,
  1.151846e-06, 1.529422e-06, 1.602931e-06, 2.058705e-06, 2.327763e-06, 
    4.154846e-06, 5.802168e-06, 6.501859e-06, 8.213025e-06, 8.826234e-06, 
    1.125931e-05, 1.628573e-05, 1.729593e-05, 1.543589e-05, 2.242939e-05,
  1.476883e-06, 1.302875e-06, 1.849828e-06, 1.886005e-06, 2.282052e-06, 
    2.706798e-06, 3.350765e-06, 4.293934e-06, 4.788532e-06, 6.6505e-06, 
    6.329603e-06, 1.081323e-05, 1.375027e-05, 1.201897e-05, 1.360928e-05,
  1.212491e-06, 1.196859e-06, 1.315598e-06, 1.731374e-06, 1.833806e-06, 
    1.923652e-06, 2.562615e-06, 2.786797e-06, 3.576898e-06, 3.530173e-06, 
    5.190216e-06, 6.987691e-06, 1.010234e-05, 1.363553e-05, 1.33082e-05,
  8.875867e-07, 8.148301e-07, 1.361969e-06, 1.061483e-06, 1.903971e-06, 
    1.538944e-06, 1.302981e-06, 1.612351e-06, 2.09886e-06, 3.15937e-06, 
    4.463596e-06, 8.173018e-06, 1.649358e-05, 3.636638e-05, 4.890269e-05,
  7.002509e-07, 1.272131e-06, 1.68384e-06, 1.093819e-06, 7.985192e-07, 
    6.853531e-07, 7.986555e-07, 1.001495e-06, 1.662554e-06, 3.89803e-06, 
    7.779883e-06, 1.411552e-05, 3.424529e-05, 5.293912e-05, 4.470215e-05,
  5.796035e-07, 9.918751e-07, 8.481955e-07, 7.585328e-07, 6.170158e-07, 
    9.330441e-07, 1.457914e-06, 2.14814e-06, 4.040416e-06, 5.315459e-06, 
    1.666673e-05, 1.554463e-05, 3.804309e-05, 2.625482e-05, 2.162041e-05,
  4.004174e-07, 3.785426e-07, 4.73071e-07, 5.49702e-07, 3.138301e-07, 
    2.419266e-07, 8.264735e-07, 1.439653e-06, 4.56904e-06, 8.379066e-06, 
    1.085213e-05, 1.889773e-05, 1.667023e-05, 2.083583e-05, 2.060566e-05,
  2.456222e-08, 5.158745e-08, 8.970134e-09, 2.010985e-07, 9.278795e-07, 
    2.091625e-06, 3.31519e-06, 2.371022e-06, 2.276314e-06, 3.71399e-06, 
    5.023006e-06, 9.333505e-06, 1.327632e-05, 1.579466e-05, 1.286531e-05,
  1.164401e-07, 1.237997e-07, 9.672201e-09, 9.611903e-09, 6.87478e-07, 
    6.271292e-07, 5.92207e-07, 1.242863e-06, 5.81076e-07, 1.45371e-06, 
    3.68273e-06, 7.44019e-06, 1.047459e-05, 9.25438e-06, 1.174586e-05,
  3.678724e-07, 2.860521e-07, 1.944546e-07, 5.557972e-08, 1.188583e-07, 
    5.188549e-07, 1.800668e-06, 1.602314e-06, 1.093692e-06, 7.546781e-07, 
    1.964906e-06, 4.866416e-06, 8.471232e-06, 1.025928e-05, 1.046837e-05,
  6.928408e-07, 4.872108e-07, 2.358594e-07, 5.279633e-07, 2.184965e-07, 
    5.804471e-07, 1.075901e-06, 2.033051e-06, 2.777073e-06, 2.192308e-06, 
    1.870057e-06, 4.323326e-06, 5.07074e-06, 5.998225e-06, 9.289468e-06,
  1.050845e-06, 7.642628e-07, 2.289306e-09, 3.132133e-09, 7.674882e-08, 
    3.080272e-07, 7.052159e-07, 1.115252e-06, 1.365377e-06, 2.022259e-06, 
    2.811565e-06, 2.531597e-06, 3.326744e-06, 3.001324e-06, 3.306161e-06,
  2.83553e-06, 6.039471e-07, 7.266995e-08, 6.943388e-08, 2.092949e-07, 
    2.780354e-07, 7.091681e-07, 9.877622e-07, 1.583658e-06, 1.627119e-06, 
    2.187552e-06, 1.825315e-06, 2.185074e-06, 1.969881e-06, 1.421934e-06,
  5.363382e-06, 3.636455e-06, 1.407727e-06, 5.170662e-07, 5.12698e-07, 
    9.817139e-07, 1.512238e-06, 1.715149e-06, 2.003075e-06, 2.027981e-06, 
    2.449022e-06, 3.678424e-06, 2.045765e-06, 1.319931e-06, 2.035692e-06,
  5.427738e-06, 4.975652e-06, 2.873535e-06, 3.799787e-06, 3.078435e-06, 
    4.182014e-06, 4.10766e-06, 3.570556e-06, 2.737415e-06, 3.782661e-06, 
    4.585906e-06, 4.276465e-06, 2.805072e-06, 3.151292e-06, 2.213086e-06,
  9.81647e-06, 4.248735e-06, 2.778829e-06, 5.024886e-06, 5.239295e-06, 
    8.109996e-06, 9.825511e-06, 8.131933e-06, 6.104543e-06, 5.966043e-06, 
    6.452204e-06, 5.895794e-06, 3.947679e-06, 3.11983e-06, 2.165285e-06,
  7.689887e-06, 9.887138e-06, 5.485047e-06, 6.449134e-06, 6.574752e-06, 
    7.971323e-06, 1.129513e-05, 1.165282e-05, 8.246317e-06, 5.607343e-06, 
    5.190043e-06, 3.283491e-06, 2.469892e-06, 2.164267e-06, 1.959954e-06,
  1.067746e-05, 7.459919e-06, 8.958992e-06, 5.033468e-06, 6.102918e-06, 
    6.069983e-06, 6.319807e-06, 5.90055e-06, 6.301206e-06, 3.692276e-06, 
    3.27807e-06, 3.125364e-06, 4.593565e-06, 5.439693e-06, 3.54488e-06,
  1.404304e-05, 1.222474e-05, 1.006463e-05, 6.410124e-06, 6.839068e-06, 
    5.933189e-06, 5.533515e-06, 4.595987e-06, 4.89681e-06, 4.420011e-06, 
    4.165738e-06, 6.035982e-06, 3.823777e-06, 4.659027e-06, 3.106447e-06,
  7.719641e-06, 8.325746e-06, 5.69165e-06, 4.620868e-06, 5.899129e-06, 
    5.404986e-06, 3.85499e-06, 5.342095e-06, 5.119472e-06, 4.884488e-06, 
    3.660856e-06, 5.545285e-06, 6.962181e-06, 5.061087e-06, 1.869072e-06,
  2.652444e-06, 1.43542e-06, 1.826143e-06, 4.355799e-06, 4.275501e-06, 
    5.526638e-06, 6.175063e-06, 8.523854e-06, 8.626476e-06, 6.434262e-06, 
    6.335643e-06, 5.503725e-06, 7.159609e-06, 7.736257e-06, 3.667546e-06,
  2.927015e-06, 3.481327e-06, 1.79496e-06, 1.628903e-06, 3.516264e-06, 
    5.681624e-06, 7.144095e-06, 8.679571e-06, 7.536527e-06, 8.798738e-06, 
    8.591511e-06, 5.286173e-06, 5.01317e-06, 5.093213e-06, 5.155093e-06,
  3.482756e-06, 3.590507e-06, 2.99551e-06, 1.853151e-06, 2.804388e-06, 
    4.312399e-06, 4.624938e-06, 6.984135e-06, 8.618687e-06, 6.646358e-06, 
    1.050874e-05, 8.978443e-06, 7.350885e-06, 5.624306e-06, 7.245552e-06,
  4.002183e-06, 3.367219e-06, 3.271193e-06, 3.108956e-06, 3.777592e-06, 
    3.517673e-06, 5.542311e-06, 7.958241e-06, 1.137902e-05, 1.113865e-05, 
    1.236412e-05, 1.167667e-05, 1.073719e-05, 7.038319e-06, 4.810609e-06,
  4.911101e-06, 4.458972e-06, 4.778416e-06, 4.392878e-06, 4.737036e-06, 
    5.721287e-06, 8.317167e-06, 8.475065e-06, 1.021537e-05, 8.844534e-06, 
    1.022541e-05, 1.591369e-05, 1.237387e-05, 1.190366e-05, 9.942734e-06,
  3.9549e-06, 4.638305e-06, 4.868406e-06, 6.042435e-06, 5.125533e-06, 
    9.693504e-06, 1.761768e-06, 2.287113e-06, 5.876988e-06, 7.587421e-06, 
    1.13333e-05, 7.44905e-06, 7.072166e-06, 1.038313e-05, 1.122675e-05,
  3.552615e-06, 4.819904e-06, 5.454453e-06, 6.81514e-06, 7.784204e-06, 
    5.862111e-06, 4.981103e-06, 7.605267e-06, 6.028902e-06, 4.964695e-06, 
    6.440219e-06, 6.135889e-06, 5.537167e-06, 4.595455e-06, 6.679847e-06,
  2.084931e-05, 1.109706e-05, 9.362981e-06, 9.12405e-06, 5.790308e-06, 
    7.24583e-06, 7.756018e-06, 5.898828e-06, 7.640499e-06, 9.49765e-06, 
    1.151933e-05, 9.329933e-06, 1.074913e-05, 8.911872e-06, 7.459123e-06,
  9.66097e-06, 4.613987e-06, 5.321811e-06, 4.282399e-06, 4.165033e-06, 
    4.310082e-06, 6.568991e-06, 9.094073e-06, 8.901161e-06, 9.256049e-06, 
    1.311589e-05, 1.186716e-05, 1.439066e-05, 1.267173e-05, 7.795945e-06,
  6.006022e-06, 6.225525e-06, 2.269051e-06, 2.719197e-06, 2.469549e-06, 
    4.654801e-06, 9.208889e-06, 9.641808e-06, 1.221013e-05, 1.145862e-05, 
    1.181984e-05, 1.250872e-05, 1.225973e-05, 1.16078e-05, 8.437579e-06,
  6.365426e-06, 5.550436e-06, 2.674767e-06, 1.962118e-06, 2.197337e-06, 
    4.224384e-06, 1.076442e-05, 1.196636e-05, 1.169754e-05, 1.4333e-05, 
    1.337306e-05, 1.539213e-05, 1.318936e-05, 1.213124e-05, 9.020017e-06,
  7.283835e-06, 4.538294e-06, 2.778541e-06, 1.38102e-06, 1.348805e-06, 
    4.989367e-06, 1.06147e-05, 9.778058e-06, 9.379279e-06, 9.371494e-06, 
    1.162694e-05, 1.076667e-05, 1.035624e-05, 1.224173e-05, 9.475479e-06,
  6.73482e-06, 4.20463e-06, 1.672812e-06, 6.472729e-07, 1.861174e-06, 
    3.135612e-06, 5.789352e-06, 7.116876e-06, 1.066482e-05, 9.683164e-06, 
    9.462188e-06, 1.132298e-05, 9.292025e-06, 5.817918e-06, 4.777729e-06,
  6.615433e-06, 2.436356e-06, 1.135546e-06, 1.104854e-06, 2.099342e-06, 
    2.008895e-06, 5.927191e-06, 1.004661e-05, 1.185223e-05, 9.108786e-06, 
    1.273702e-05, 1.110129e-05, 8.417169e-06, 6.087379e-06, 6.609549e-06,
  5.130772e-06, 2.271701e-06, 2.145522e-06, 2.101928e-06, 2.993589e-06, 
    4.039365e-06, 5.74569e-06, 1.08227e-05, 1.118679e-05, 8.938367e-06, 
    1.015363e-05, 9.683283e-06, 5.60443e-06, 7.268566e-06, 3.01661e-06,
  5.645639e-06, 1.526619e-06, 2.22654e-06, 3.008689e-06, 3.281933e-06, 
    4.926168e-06, 8.085782e-06, 7.807005e-06, 6.859273e-06, 8.977531e-06, 
    8.302434e-06, 6.245166e-06, 6.488936e-06, 7.181021e-06, 6.753804e-06,
  5.478186e-06, 5.52557e-06, 4.632824e-06, 4.336665e-06, 4.825606e-06, 
    4.765167e-06, 5.905594e-06, 6.724582e-06, 6.038969e-06, 5.927191e-06, 
    6.668153e-06, 6.73261e-06, 6.605409e-06, 7.745057e-06, 7.383596e-06,
  0.000251099, 6.953382e-05, 4.857077e-05, 2.300535e-05, 1.583185e-05, 
    1.138703e-05, 5.40429e-06, 4.351928e-06, 2.456119e-06, 4.41192e-06, 
    4.161025e-06, 5.257442e-06, 6.241385e-06, 6.938417e-06, 4.734095e-06,
  7.488246e-05, 3.757076e-05, 1.283685e-05, 4.705627e-06, 4.716886e-06, 
    5.368309e-06, 5.604707e-06, 2.412492e-06, 2.591512e-06, 2.378908e-06, 
    1.891944e-06, 2.161171e-06, 3.230085e-06, 4.127777e-06, 5.020361e-06,
  5.594401e-05, 5.130296e-05, 2.7282e-05, 1.025242e-05, 6.870237e-06, 
    6.631009e-06, 3.938121e-06, 3.734444e-06, 2.116841e-06, 2.704555e-06, 
    2.06157e-06, 4.128795e-06, 4.366173e-06, 5.036119e-06, 4.83721e-06,
  6.802752e-05, 4.703004e-05, 2.046248e-05, 7.393257e-06, 7.90059e-06, 
    6.839787e-06, 8.233967e-06, 3.931178e-06, 3.880337e-06, 3.893571e-06, 
    6.524165e-06, 5.104238e-06, 5.283544e-06, 4.737841e-06, 4.194546e-06,
  8.146268e-05, 2.295805e-05, 6.94526e-06, 5.440621e-06, 7.593227e-06, 
    8.34087e-06, 5.613756e-06, 4.480481e-06, 7.70654e-07, 3.475872e-06, 
    5.870825e-06, 5.693213e-06, 6.413929e-06, 4.437923e-06, 2.874123e-06,
  3.251643e-05, 2.493384e-05, 8.423754e-06, 1.034101e-05, 6.632236e-06, 
    5.904067e-06, 5.437269e-06, 6.35036e-06, 8.24784e-06, 7.345493e-06, 
    7.61414e-06, 7.610273e-06, 6.174555e-06, 3.273947e-06, 2.282794e-06,
  7.177036e-06, 3.710464e-06, 5.409401e-06, 5.898474e-06, 7.127788e-06, 
    6.23732e-06, 6.417773e-06, 9.034232e-06, 8.59831e-06, 6.212176e-06, 
    6.239105e-06, 4.178833e-06, 5.245208e-06, 4.566425e-06, 3.69149e-06,
  3.351268e-06, 3.264932e-06, 3.421369e-06, 5.430049e-06, 7.218114e-06, 
    7.042868e-06, 1.010099e-05, 7.840691e-06, 5.415785e-06, 6.08237e-06, 
    5.184132e-06, 3.98466e-06, 5.171041e-06, 6.054324e-06, 5.167647e-06,
  9.080069e-07, 2.136966e-06, 3.442233e-06, 5.853847e-06, 8.867766e-06, 
    9.682137e-06, 8.843103e-06, 6.829342e-06, 3.805243e-06, 6.832272e-06, 
    6.023845e-06, 5.37536e-06, 6.394665e-06, 5.942381e-06, 5.64295e-06,
  1.483272e-06, 2.119706e-06, 3.194329e-06, 3.680087e-06, 5.206812e-06, 
    7.758894e-06, 7.220546e-06, 7.690057e-06, 6.770005e-06, 5.628163e-06, 
    6.705004e-06, 7.403146e-06, 7.467629e-06, 6.871908e-06, 7.822709e-06,
  2.426331e-05, 5.680633e-05, 8.474536e-05, 8.73844e-05, 9.753156e-05, 
    8.675428e-05, 6.698117e-05, 5.576375e-05, 9.886714e-05, 0.0001388886, 
    3.716547e-05, 5.964488e-06, 6.134937e-06, 6.178705e-06, 4.910966e-06,
  2.635297e-05, 0.0001364836, 0.0001242902, 0.0001391202, 0.0001393303, 
    0.0001381822, 0.0001274896, 0.0001115514, 0.000196192, 0.0001718019, 
    0.000101761, 1.834018e-05, 1.044132e-05, 7.048357e-06, 4.890675e-06,
  1.590488e-05, 0.0001600913, 0.0001711346, 0.000158166, 0.0001197801, 
    0.0001140721, 0.0001245917, 8.874913e-05, 7.264435e-05, 0.0001221405, 
    0.000152057, 4.274002e-05, 8.520647e-06, 5.49107e-06, 6.152972e-06,
  1.047894e-05, 0.0001998384, 0.0002061106, 0.0001599979, 0.000110452, 
    0.0001061645, 0.0001048105, 7.884201e-05, 6.14905e-05, 0.0001607059, 
    0.0002124121, 7.013523e-05, 6.654697e-06, 6.136113e-06, 6.99761e-06,
  1.967587e-05, 0.0001024985, 0.0001867591, 0.000132227, 8.047438e-05, 
    6.568256e-05, 6.066411e-05, 7.618716e-05, 8.831577e-05, 0.0001794495, 
    0.0001615385, 6.478091e-05, 7.3018e-06, 6.469123e-06, 4.532953e-06,
  3.782513e-05, 7.844333e-05, 8.588121e-05, 7.887935e-05, 7.1043e-05, 
    6.434447e-05, 5.950117e-05, 7.817381e-05, 0.0001312524, 0.0001459282, 
    0.0002270398, 7.953523e-05, 7.427789e-06, 6.328818e-06, 5.458118e-06,
  9.670361e-05, 6.581173e-05, 0.0001160901, 5.309956e-05, 5.453561e-05, 
    6.401506e-05, 6.810707e-05, 0.0001025273, 8.341132e-05, 0.0001186754, 
    0.0001879956, 6.940015e-05, 7.969989e-06, 4.856733e-06, 5.010058e-06,
  7.356487e-05, 4.645884e-05, 5.093309e-05, 4.624094e-05, 4.357141e-05, 
    4.390867e-05, 4.5759e-05, 5.153033e-05, 7.01338e-05, 7.200761e-05, 
    0.0001278487, 4.261898e-05, 6.67734e-06, 4.206966e-06, 4.110501e-06,
  4.649553e-05, 3.031245e-05, 4.47731e-05, 3.915329e-05, 3.416257e-05, 
    3.204285e-05, 4.214287e-05, 3.782762e-05, 6.251802e-05, 6.440782e-05, 
    6.666876e-05, 2.519854e-05, 5.551195e-06, 3.964445e-06, 3.284237e-06,
  2.36529e-05, 2.198144e-05, 2.502268e-05, 3.096717e-05, 1.678558e-05, 
    3.525343e-05, 3.982446e-05, 3.722108e-05, 8.513275e-05, 7.046633e-05, 
    4.009808e-05, 1.42793e-05, 3.733938e-06, 2.900631e-06, 3.385919e-06,
  1.880472e-05, 2.237259e-05, 3.957346e-05, 4.492444e-05, 4.154323e-05, 
    3.538207e-05, 1.903587e-05, 3.104773e-05, 8.053752e-05, 0.0001896665, 
    0.0002385901, 0.0001376845, 7.809624e-05, 7.306322e-05, 6.672535e-05,
  4.686271e-06, 1.283147e-05, 2.531686e-05, 3.503511e-05, 4.332837e-05, 
    4.677378e-05, 1.839365e-05, 3.488733e-05, 3.766434e-05, 0.0001199309, 
    0.0002985322, 0.0002524108, 0.0001368824, 8.730119e-05, 7.160826e-05,
  2.095136e-06, 4.43792e-06, 1.160122e-05, 2.088095e-05, 4.396514e-05, 
    4.232585e-05, 2.016499e-05, 3.784816e-05, 9.406896e-06, 9.345768e-05, 
    0.000194009, 0.0003432767, 0.0002580128, 0.0001249254, 7.622514e-05,
  1.591663e-06, 1.207347e-06, 3.678296e-06, 1.050097e-05, 1.710812e-05, 
    2.261937e-05, 4.678948e-05, 3.006916e-05, 2.573917e-05, 3.397543e-05, 
    9.068768e-05, 0.0003362945, 0.0002854931, 0.0001966642, 0.0001121838,
  1.994645e-06, 1.242983e-06, 1.708822e-06, 4.042304e-06, 4.844019e-06, 
    2.183462e-05, 3.260023e-05, 3.992111e-05, 3.677898e-05, 3.690842e-05, 
    5.948525e-05, 0.0001657505, 0.0002535399, 0.0002334585, 0.0001829406,
  1.641737e-06, 8.915236e-07, 1.350214e-06, 1.276909e-06, 2.489619e-06, 
    6.743327e-06, 1.268268e-05, 2.705402e-05, 4.046155e-05, 4.300637e-05, 
    5.705476e-05, 0.0001271105, 0.0001903501, 0.0001861854, 0.0001742851,
  1.385874e-05, 4.508564e-06, 6.199891e-07, 1.296181e-06, 1.649808e-06, 
    2.642615e-06, 6.736174e-06, 1.072282e-05, 1.71387e-05, 2.522324e-05, 
    3.368251e-05, 8.823761e-05, 0.0001520854, 0.0001324476, 0.000131558,
  2.439552e-05, 1.426343e-05, 6.055257e-06, 2.566515e-06, 1.448995e-06, 
    1.867983e-06, 2.264548e-06, 5.135271e-06, 8.230827e-06, 8.38123e-06, 
    1.115802e-05, 0.0001024691, 0.0001037282, 0.0001136864, 0.0001091243,
  1.27064e-05, 6.781931e-06, 4.296772e-06, 2.3234e-06, 1.726263e-06, 
    1.864934e-06, 1.93395e-06, 1.963308e-06, 1.382981e-06, 2.886117e-06, 
    1.96184e-05, 6.308281e-05, 0.0001135221, 0.000113511, 0.0001046665,
  1.352235e-06, 2.167836e-06, 1.622145e-06, 9.033502e-07, 9.4725e-07, 
    1.627741e-06, 1.482729e-06, 1.939153e-06, 1.86567e-06, 7.373794e-06, 
    7.712984e-05, 0.0001014477, 0.0001159715, 0.0001105252, 0.0001086152,
  3.289884e-05, 6.560543e-05, 3.30093e-05, 3.175849e-05, 2.022849e-05, 
    1.856237e-05, 2.975388e-05, 1.657157e-05, 2.195486e-05, 2.903385e-05, 
    3.701239e-05, 6.520212e-05, 6.136307e-05, 9.154937e-05, 0.000107176,
  1.148423e-05, 5.302716e-05, 3.286233e-05, 3.695397e-05, 3.003049e-05, 
    1.670846e-05, 1.585526e-05, 1.676678e-05, 2.264519e-05, 2.057151e-05, 
    4.124988e-05, 5.433768e-05, 6.680247e-05, 6.83423e-05, 9.295688e-05,
  8.947571e-06, 1.558352e-05, 4.954867e-05, 4.545278e-05, 2.889629e-05, 
    8.832907e-06, 7.080244e-06, 9.340908e-06, 1.284095e-05, 1.932834e-05, 
    3.619647e-05, 0.0001123331, 7.835041e-05, 0.0001058568, 0.000119643,
  1.611591e-06, 5.203663e-06, 1.356477e-05, 2.241881e-05, 2.831696e-05, 
    8.399225e-06, 7.283496e-06, 4.832033e-06, 4.369421e-06, 3.794676e-06, 
    1.254548e-05, 7.788909e-05, 0.0001499893, 0.0002167144, 0.0001239987,
  5.718224e-08, 2.166994e-07, 3.702033e-06, 7.945639e-06, 1.741413e-05, 
    1.788797e-05, 1.961113e-05, 1.235868e-05, 8.724085e-06, 7.050009e-06, 
    6.226137e-06, 1.394448e-05, 0.000108197, 0.0001536945, 0.0001301457,
  1.381942e-07, 2.296545e-08, 6.28212e-07, 3.122007e-07, 7.602777e-06, 
    9.659203e-06, 1.586763e-05, 2.684308e-05, 2.299035e-05, 2.073428e-05, 
    2.073426e-05, 3.68735e-05, 5.716279e-05, 0.0001436589, 0.0001171029,
  4.439888e-06, 3.484309e-07, 6.110068e-08, 2.903955e-07, 2.720899e-07, 
    2.189598e-06, 1.263948e-05, 1.597539e-05, 2.839227e-05, 3.577048e-05, 
    4.100046e-05, 5.994174e-05, 6.828134e-05, 8.945482e-05, 7.681271e-05,
  3.011991e-05, 4.798991e-06, 1.660654e-06, 9.513404e-07, 1.26287e-06, 
    2.46269e-06, 4.794207e-06, 6.018772e-06, 1.056757e-05, 1.249517e-05, 
    1.647064e-05, 2.107935e-05, 2.230575e-05, 1.845494e-05, 1.37148e-05,
  0.0001151305, 6.143977e-05, 1.491945e-05, 2.518462e-06, 2.21179e-06, 
    4.390437e-06, 3.719933e-06, 4.436881e-06, 5.524682e-06, 5.528901e-06, 
    7.685263e-06, 8.567325e-06, 6.97042e-06, 6.5236e-06, 6.582932e-06,
  0.000137451, 0.0001119203, 9.231903e-05, 3.523881e-05, 3.136597e-06, 
    2.022735e-06, 3.693064e-06, 5.658238e-06, 7.983499e-06, 5.681963e-06, 
    7.085569e-06, 6.540567e-06, 4.60695e-06, 4.113779e-06, 4.506011e-06,
  1.003381e-05, 1.752023e-05, 2.797956e-05, 3.144775e-05, 2.603819e-05, 
    1.165598e-05, 1.163647e-05, 1.242113e-05, 1.430626e-05, 1.247288e-05, 
    1.684994e-05, 2.564882e-05, 2.180662e-05, 1.463624e-05, 1.025999e-05,
  3.493676e-06, 3.265674e-06, 1.39605e-05, 1.322951e-05, 2.427453e-05, 
    1.700869e-05, 2.414615e-05, 1.681109e-05, 2.646633e-05, 2.092464e-05, 
    1.954773e-05, 2.893295e-05, 3.116106e-05, 3.514431e-05, 1.292338e-05,
  3.082496e-06, 2.715031e-06, 6.741472e-06, 5.837914e-06, 9.528847e-06, 
    9.343713e-06, 2.400096e-05, 3.194264e-05, 3.92555e-05, 3.871049e-05, 
    4.538924e-05, 5.371207e-05, 5.475015e-05, 4.906906e-05, 4.787028e-05,
  2.468629e-06, 3.758809e-06, 4.000017e-06, 1.306549e-06, 2.38922e-06, 
    3.519826e-06, 3.606594e-06, 9.954537e-06, 2.443377e-05, 7.814609e-05, 
    8.536095e-05, 6.985181e-05, 0.0001222657, 0.0001346221, 8.455393e-05,
  8.340995e-07, 4.171658e-06, 2.456738e-06, 3.572096e-06, 3.587714e-06, 
    5.951561e-06, 5.89867e-06, 3.983668e-06, 3.866915e-06, 6.499122e-06, 
    1.705484e-05, 8.648919e-05, 0.0001461879, 0.0001269504, 0.0001289581,
  9.455248e-09, 1.570853e-07, 1.617953e-06, 4.431637e-06, 3.872236e-06, 
    6.436574e-06, 9.336639e-06, 1.281258e-05, 5.253924e-06, 5.354603e-06, 
    6.682326e-06, 2.382261e-05, 7.048655e-05, 0.0001137841, 0.0001239388,
  3.573214e-10, 6.292739e-10, 5.298736e-08, 1.488441e-06, 1.453919e-06, 
    4.048778e-06, 6.992163e-06, 9.549618e-06, 2.005474e-05, 1.536828e-05, 
    1.342811e-05, 2.110267e-05, 6.557559e-05, 9.592596e-05, 6.647999e-05,
  1.22629e-06, 9.34938e-08, 5.633473e-09, 2.002492e-08, 7.388603e-08, 
    1.008791e-06, 3.886139e-06, 9.269051e-06, 1.123013e-05, 1.216554e-05, 
    3.194139e-05, 3.557258e-05, 5.516199e-05, 5.167274e-05, 3.228613e-05,
  1.121129e-05, 1.135083e-05, 5.238049e-06, 3.740181e-08, 1.885016e-09, 
    1.082942e-07, 9.452658e-07, 3.516959e-06, 6.460351e-06, 7.215766e-06, 
    1.137191e-05, 1.571536e-05, 2.678795e-05, 2.368901e-05, 1.155253e-05,
  8.883637e-05, 0.0001016295, 4.61745e-05, 1.556567e-05, 4.140554e-07, 
    1.002789e-06, 3.676366e-07, 1.385397e-06, 2.381899e-06, 3.915712e-06, 
    5.031528e-06, 6.126119e-06, 8.073982e-06, 6.678429e-06, 6.052337e-06,
  9.402152e-07, 4.583524e-06, 5.303866e-06, 3.630315e-06, 1.153472e-05, 
    1.01973e-05, 1.545975e-05, 1.465492e-05, 1.203851e-05, 4.923634e-06, 
    5.738583e-06, 8.630269e-06, 1.43126e-05, 2.103039e-05, 4.355612e-05,
  2.249476e-06, 2.11699e-06, 3.281169e-06, 3.390388e-06, 6.588368e-06, 
    1.143815e-05, 1.666786e-05, 1.198062e-05, 1.414649e-05, 7.696714e-06, 
    5.725982e-06, 6.412349e-06, 1.118424e-05, 1.848301e-05, 3.446613e-05,
  9.483787e-07, 1.687965e-06, 1.305097e-06, 2.064218e-06, 3.078327e-06, 
    4.794807e-06, 1.845066e-05, 2.964008e-05, 1.843829e-05, 1.068622e-05, 
    1.046006e-05, 1.373971e-05, 1.049829e-05, 1.604181e-05, 3.034348e-05,
  9.660214e-07, 2.424518e-06, 3.707917e-06, 2.565633e-06, 2.161358e-06, 
    2.335793e-06, 8.45867e-06, 2.086381e-05, 2.866533e-05, 1.871256e-05, 
    2.78265e-05, 2.086877e-05, 2.980797e-05, 9.440717e-06, 1.529121e-05,
  1.951288e-07, 1.460828e-06, 5.036752e-06, 6.183801e-06, 2.31278e-06, 
    2.239326e-06, 2.282388e-06, 1.701883e-06, 4.846523e-06, 2.692089e-05, 
    2.574592e-05, 3.321473e-05, 3.688635e-05, 7.490671e-05, 2.154667e-05,
  6.231589e-07, 1.948344e-07, 9.131762e-07, 4.80867e-06, 2.236214e-06, 
    2.40039e-06, 1.492895e-06, 1.787837e-06, 4.575777e-06, 4.87687e-06, 
    1.135614e-05, 3.404787e-05, 4.968562e-05, 4.251651e-05, 3.70125e-05,
  1.265587e-09, 1.236783e-10, 3.897249e-07, 9.981669e-07, 5.879556e-07, 
    1.397889e-06, 2.243135e-06, 2.634511e-06, 2.447223e-06, 3.626124e-06, 
    6.681679e-06, 2.063448e-05, 3.408716e-05, 2.859342e-05, 3.842651e-05,
  1.021986e-08, 6.060056e-09, 1.681e-09, 1.54817e-08, 9.185804e-08, 
    4.830703e-07, 2.291151e-06, 3.356837e-06, 3.119314e-06, 3.624632e-06, 
    4.495069e-06, 1.164034e-05, 3.234003e-05, 3.759948e-05, 3.502341e-05,
  2.690317e-06, 1.150226e-06, 6.01026e-07, 1.948452e-08, 2.782262e-08, 
    2.748615e-07, 3.89274e-07, 1.598876e-06, 3.257341e-06, 3.323359e-06, 
    4.148715e-06, 5.985205e-06, 1.768974e-05, 2.170669e-05, 3.373752e-05,
  3.526424e-06, 1.698325e-06, 3.01847e-06, 3.235058e-07, 3.005741e-08, 
    1.989576e-08, 3.228519e-08, 2.421878e-07, 1.80601e-06, 3.093374e-06, 
    3.29051e-06, 7.87375e-06, 2.239577e-05, 2.385415e-05, 1.294866e-05,
  0.0001140329, 0.0001422838, 0.0001735898, 0.0001949739, 0.0001471621, 
    6.758943e-05, 2.096209e-05, 8.448732e-06, 1.64792e-06, 7.623107e-07, 
    4.612677e-06, 1.02218e-05, 6.859019e-06, 8.899283e-06, 1.579672e-05,
  9.5925e-05, 0.0001301117, 0.0001703687, 0.000208682, 0.0001819216, 
    9.328809e-05, 3.368422e-05, 1.238981e-05, 2.956089e-06, 1.497134e-07, 
    2.015111e-06, 5.883233e-06, 1.430107e-05, 1.019281e-05, 8.554954e-06,
  7.710601e-05, 0.0001089346, 0.0001471998, 0.0002045227, 0.0001967754, 
    0.0001242487, 5.139532e-05, 1.841118e-05, 1.012885e-05, 2.977797e-07, 
    6.914087e-07, 3.149468e-06, 1.083979e-05, 1.450124e-05, 8.305958e-06,
  5.922973e-05, 8.094103e-05, 0.0001180495, 0.0001712423, 0.0002074711, 
    0.0001720262, 7.385974e-05, 2.212908e-05, 1.275015e-05, 4.657721e-06, 
    2.494383e-07, 1.343778e-06, 6.341181e-06, 1.021628e-05, 1.323207e-05,
  4.532824e-05, 5.422412e-05, 8.161565e-05, 0.0001201117, 0.0001813134, 
    0.0001992939, 0.0001197689, 3.516101e-05, 1.098789e-05, 8.370995e-06, 
    6.732605e-07, 3.783555e-07, 2.352408e-06, 7.278033e-06, 1.485395e-05,
  3.379029e-05, 3.501051e-05, 4.340339e-05, 6.557316e-05, 0.0001296094, 
    0.0001806952, 0.0001447576, 4.419377e-05, 8.452977e-06, 1.02821e-05, 
    6.273803e-06, 1.197992e-06, 2.164596e-06, 3.666169e-06, 8.610634e-06,
  1.891139e-05, 2.691471e-05, 2.629841e-05, 3.104471e-05, 6.214003e-05, 
    0.0001178725, 0.0001058254, 3.016948e-05, 2.835838e-06, 4.111781e-06, 
    7.43976e-06, 3.888182e-06, 3.288288e-06, 3.100685e-06, 7.570679e-06,
  1.14683e-05, 1.84908e-05, 1.673047e-05, 1.71811e-05, 5.352988e-05, 
    3.22858e-05, 4.126839e-05, 9.2935e-06, 3.696563e-07, 9.309094e-07, 
    3.807944e-06, 4.155878e-06, 2.386325e-06, 3.169425e-06, 5.663815e-06,
  5.449318e-06, 2.469908e-05, 2.151101e-05, 2.202261e-05, 1.704976e-05, 
    1.332032e-05, 6.490088e-06, 1.929528e-06, 1.119606e-07, 2.753017e-07, 
    6.02308e-07, 1.839549e-06, 3.120477e-06, 5.312771e-06, 2.841839e-06,
  5.693984e-06, 2.39491e-05, 7.76575e-06, 5.72772e-06, 2.401368e-06, 
    1.028943e-06, 1.669459e-06, 1.414023e-07, 9.543948e-09, 1.40193e-08, 
    3.596629e-07, 1.054121e-06, 2.672922e-06, 3.737545e-06, 7.205684e-06,
  4.244851e-06, 3.013394e-06, 3.195894e-06, 4.335314e-06, 1.110412e-05, 
    2.177762e-05, 3.509447e-05, 3.931922e-05, 5.622058e-05, 6.62197e-05, 
    8.171864e-05, 9.785406e-05, 0.0001098564, 0.0001038992, 8.060217e-05,
  4.040597e-06, 3.734089e-06, 3.052374e-06, 6.098643e-06, 2.063987e-05, 
    3.772865e-05, 3.472879e-05, 3.786231e-05, 4.823305e-05, 7.381745e-05, 
    7.165578e-05, 7.839346e-05, 9.716301e-05, 9.253799e-05, 6.700352e-05,
  3.810808e-06, 4.620144e-06, 4.348314e-06, 8.842213e-06, 3.568751e-05, 
    4.48021e-05, 3.914992e-05, 4.397531e-05, 4.470639e-05, 6.087999e-05, 
    5.866641e-05, 6.299772e-05, 9.105833e-05, 9.931598e-05, 0.0001025681,
  1.092376e-05, 1.263494e-05, 1.106168e-05, 1.270918e-05, 3.329608e-05, 
    4.970667e-05, 5.465054e-05, 6.120752e-05, 4.680876e-05, 4.014249e-05, 
    4.983629e-05, 5.662327e-05, 0.0001163177, 0.000121116, 0.000111204,
  2.478708e-05, 3.176926e-05, 2.389246e-05, 1.676838e-05, 4.05823e-05, 
    4.32187e-05, 7.257692e-05, 9.440976e-05, 8.495234e-05, 9.054617e-05, 
    0.0001110431, 0.0001226049, 0.0001317447, 0.0001291793, 7.682362e-05,
  1.741661e-05, 2.187089e-05, 2.382775e-05, 2.650562e-05, 2.680048e-05, 
    3.45097e-05, 9.066502e-05, 0.0001415275, 0.0001987226, 0.0001943231, 
    0.000174698, 0.0001450149, 0.0001673642, 0.0001092406, 5.107481e-05,
  7.976355e-06, 9.580242e-06, 1.333558e-05, 1.138426e-05, 2.39514e-05, 
    8.699296e-05, 0.000222219, 0.0002743377, 0.000274366, 0.0002662238, 
    0.0001913335, 0.0001348609, 8.564894e-05, 6.475923e-05, 3.043059e-05,
  4.692352e-06, 1.137306e-05, 1.554891e-05, 2.28135e-05, 3.257531e-05, 
    8.09749e-05, 0.0002465326, 0.0003642635, 0.0003254596, 0.0003157673, 
    0.0002605717, 0.0001302097, 5.9331e-05, 3.287672e-05, 3.520418e-05,
  8.305591e-06, 1.369772e-05, 2.150517e-05, 3.750554e-05, 5.908189e-05, 
    7.777498e-05, 0.0001387902, 0.0002495696, 0.0002937438, 0.0003236362, 
    0.0003176101, 0.0002029861, 7.517796e-05, 2.974792e-05, 1.806565e-05,
  1.451417e-05, 2.496182e-05, 3.553753e-05, 6.316558e-05, 5.799944e-05, 
    5.754284e-05, 5.790951e-05, 9.490726e-05, 0.0001329709, 0.0002037996, 
    0.000292282, 0.0002685146, 0.0001663658, 7.488339e-05, 2.603763e-05,
  1.845708e-06, 1.967244e-06, 2.704272e-06, 4.063709e-06, 4.60209e-06, 
    3.940583e-06, 2.688779e-06, 2.895314e-06, 2.871271e-06, 3.634729e-06, 
    4.434869e-06, 5.930939e-06, 9.662319e-06, 8.821491e-06, 1.021778e-05,
  1.267828e-06, 2.227687e-06, 2.470532e-06, 3.166267e-06, 4.076562e-06, 
    3.780369e-06, 4.13471e-06, 3.492205e-06, 3.580496e-06, 4.368502e-06, 
    4.327886e-06, 4.666223e-06, 9.318449e-06, 9.124927e-06, 9.997494e-06,
  2.250867e-06, 2.277701e-06, 4.109354e-06, 4.317851e-06, 4.468837e-06, 
    3.973403e-06, 4.156979e-06, 3.872847e-06, 4.247388e-06, 5.319972e-06, 
    6.350646e-06, 6.412881e-06, 6.716823e-06, 4.942508e-06, 1.584016e-05,
  2.40618e-06, 3.009679e-06, 3.847814e-06, 4.761379e-06, 4.956041e-06, 
    4.758012e-06, 4.832849e-06, 4.822111e-06, 4.529245e-06, 6.437131e-06, 
    8.321637e-06, 7.272245e-06, 3.234445e-06, 5.779213e-06, 2.141445e-05,
  3.379575e-06, 5.165739e-06, 4.232394e-06, 4.166049e-06, 4.757429e-06, 
    5.537442e-06, 4.849425e-06, 5.951532e-06, 5.703591e-06, 5.48131e-06, 
    8.065746e-06, 9.123089e-06, 2.891452e-06, 9.67145e-06, 3.25628e-05,
  3.353739e-06, 4.709354e-06, 4.269024e-06, 4.585115e-06, 5.409245e-06, 
    5.659577e-06, 5.633537e-06, 6.915491e-06, 5.555683e-06, 5.480543e-06, 
    6.794095e-06, 8.558663e-06, 4.348556e-06, 1.381851e-05, 4.336505e-05,
  4.855033e-06, 5.099074e-06, 5.477169e-06, 5.209173e-06, 4.838882e-06, 
    5.469906e-06, 5.63346e-06, 8.250012e-06, 7.640115e-06, 5.919556e-06, 
    7.412834e-06, 7.781282e-06, 5.099012e-06, 2.02502e-05, 5.521112e-05,
  6.649606e-06, 5.712337e-06, 5.6926e-06, 5.364182e-06, 4.326626e-06, 
    5.25196e-06, 7.273584e-06, 7.943004e-06, 7.900304e-06, 7.713633e-06, 
    7.575982e-06, 4.843895e-06, 5.551439e-06, 2.710481e-05, 7.080367e-05,
  7.194784e-06, 4.697946e-06, 6.07719e-06, 4.96615e-06, 4.262466e-06, 
    5.190331e-06, 7.627811e-06, 9.04801e-06, 7.685238e-06, 6.839653e-06, 
    4.921993e-06, 4.915e-06, 1.601387e-05, 3.049897e-05, 4.964535e-05,
  6.689362e-06, 6.377599e-06, 5.742656e-06, 5.735355e-06, 4.78494e-06, 
    5.196401e-06, 8.008874e-06, 9.796627e-06, 7.954166e-06, 5.52394e-06, 
    6.977563e-06, 1.310386e-05, 1.583478e-05, 2.379412e-05, 3.271428e-05,
  3.414912e-06, 2.556568e-06, 3.630229e-06, 8.279221e-06, 9.059581e-06, 
    1.146456e-05, 1.396439e-05, 1.454209e-05, 1.112813e-05, 9.720836e-06, 
    8.6004e-06, 8.161485e-06, 1.008944e-05, 1.670304e-05, 1.63761e-05,
  3.516176e-06, 3.915914e-06, 4.437152e-06, 5.053355e-06, 9.188188e-06, 
    1.079025e-05, 1.02399e-05, 1.28339e-05, 9.20552e-06, 6.474717e-06, 
    5.384055e-06, 6.102543e-06, 7.3304e-06, 1.13897e-05, 1.124335e-05,
  2.466572e-06, 2.69282e-06, 5.517226e-06, 5.497168e-06, 7.422779e-06, 
    8.444312e-06, 7.978309e-06, 6.19324e-06, 5.410534e-06, 4.980673e-06, 
    6.341307e-06, 9.298839e-06, 1.174249e-05, 9.886929e-06, 4.890588e-06,
  7.595041e-07, 3.234201e-06, 4.883496e-06, 6.375522e-06, 5.745391e-06, 
    7.011659e-06, 7.79448e-06, 5.333143e-06, 6.599449e-06, 6.253985e-06, 
    7.562056e-06, 9.360729e-06, 6.912731e-06, 6.809468e-06, 2.608742e-06,
  1.488531e-07, 3.004342e-06, 4.640361e-06, 5.867334e-06, 5.123093e-06, 
    5.373593e-06, 5.756372e-06, 3.144362e-06, 7.035607e-06, 7.701649e-06, 
    7.250283e-06, 4.788087e-06, 3.084828e-06, 2.471432e-06, 1.453857e-06,
  1.305914e-06, 7.778066e-07, 3.409611e-06, 4.483965e-06, 4.900692e-06, 
    3.648415e-06, 3.435581e-06, 2.51979e-06, 7.362003e-06, 8.436353e-06, 
    7.926382e-06, 7.106764e-06, 3.543064e-06, 2.336957e-06, 1.516567e-06,
  1.329131e-06, 1.135632e-06, 1.66596e-06, 3.482791e-06, 4.560444e-06, 
    5.044711e-06, 5.094445e-06, 3.559962e-06, 6.211204e-06, 6.972096e-06, 
    6.144354e-06, 4.928007e-06, 3.732976e-06, 4.886474e-06, 1.101551e-05,
  9.891342e-07, 9.880343e-07, 1.766997e-06, 2.916098e-06, 3.886563e-06, 
    5.923428e-06, 5.573098e-06, 4.338478e-06, 4.458735e-06, 6.188916e-06, 
    5.627351e-06, 2.571292e-06, 4.657057e-06, 9.14611e-06, 2.697197e-05,
  9.057546e-07, 9.873318e-07, 1.947966e-06, 2.774219e-06, 3.809979e-06, 
    5.739626e-06, 6.193813e-06, 5.341034e-06, 3.591452e-06, 3.826337e-06, 
    4.619144e-06, 1.874104e-06, 3.034637e-06, 1.488983e-05, 2.793332e-05,
  1.645212e-06, 1.219528e-06, 1.253676e-06, 2.309785e-06, 3.434334e-06, 
    5.577509e-06, 6.472811e-06, 5.506621e-06, 3.499306e-06, 2.826967e-06, 
    1.390413e-06, 2.312516e-06, 3.748451e-06, 1.185078e-05, 2.089519e-05,
  2.708501e-05, 4.25116e-05, 3.934801e-05, 5.310045e-05, 5.817959e-05, 
    6.939764e-05, 7.804616e-05, 8.4498e-05, 0.0001129327, 0.0001172098, 
    0.0001386542, 0.000120479, 9.154844e-05, 7.740351e-05, 4.845811e-05,
  1.987645e-05, 2.591354e-05, 3.089588e-05, 3.891035e-05, 3.605354e-05, 
    4.24578e-05, 6.182449e-05, 5.807278e-05, 7.636873e-05, 0.0001081519, 
    8.488288e-05, 8.962203e-05, 4.837894e-05, 4.52934e-05, 1.597055e-05,
  1.094725e-05, 1.890655e-05, 1.645595e-05, 2.259061e-05, 3.77019e-05, 
    4.077061e-05, 3.974891e-05, 4.118148e-05, 3.843029e-05, 3.196085e-05, 
    4.618498e-05, 4.60929e-05, 3.583304e-05, 1.987976e-05, 4.874623e-06,
  1.776887e-05, 1.879601e-05, 1.814372e-05, 7.960246e-06, 3.327931e-05, 
    3.09948e-05, 3.531068e-05, 3.45519e-05, 3.25504e-05, 1.888724e-05, 
    1.912894e-05, 1.97571e-05, 1.785531e-05, 1.024581e-05, 5.550707e-06,
  4.32167e-06, 4.942352e-06, 7.839427e-06, 1.340132e-05, 1.771182e-05, 
    1.201181e-05, 1.303652e-05, 2.372461e-05, 2.120717e-05, 2.410425e-05, 
    1.414141e-05, 1.085924e-05, 8.767863e-06, 4.163407e-06, 3.441891e-06,
  1.180945e-05, 1.184069e-05, 1.028348e-05, 1.321268e-05, 1.509686e-05, 
    1.043746e-05, 1.923703e-05, 1.342015e-05, 1.335042e-05, 1.109606e-05, 
    9.694979e-06, 5.908473e-06, 5.377458e-06, 4.151563e-06, 2.632671e-06,
  7.411822e-06, 9.81736e-06, 1.321592e-05, 2.042025e-05, 1.940288e-05, 
    1.59577e-05, 1.344448e-05, 1.406776e-05, 1.155443e-05, 8.847676e-06, 
    4.737793e-06, 4.095147e-06, 4.4678e-06, 3.406021e-06, 6.136856e-06,
  1.227369e-05, 7.642696e-06, 1.404289e-05, 1.38099e-05, 1.241941e-05, 
    1.176095e-05, 1.027993e-05, 1.052929e-05, 7.676317e-06, 5.021094e-06, 
    4.402087e-06, 6.34243e-06, 2.857615e-06, 7.175424e-06, 1.288678e-05,
  8.227901e-06, 7.976539e-06, 4.351833e-06, 2.8168e-06, 3.812071e-06, 
    3.691869e-06, 8.145317e-06, 8.948236e-06, 7.294213e-06, 3.945962e-06, 
    2.66355e-06, 2.248824e-06, 3.607504e-06, 7.608748e-06, 2.668009e-05,
  2.698279e-06, 2.302057e-06, 1.673478e-06, 7.429203e-07, 1.016668e-06, 
    1.716821e-06, 3.923933e-06, 5.712235e-06, 3.95076e-06, 3.919648e-06, 
    2.725921e-06, 1.812209e-06, 1.824866e-06, 1.054554e-05, 2.399464e-05,
  3.104097e-05, 4.26198e-05, 6.098855e-05, 6.704778e-05, 8.070622e-05, 
    8.503967e-05, 7.757158e-05, 7.637741e-05, 7.235199e-05, 6.327691e-05, 
    6.920209e-05, 6.859584e-05, 7.409404e-05, 0.0001226102, 0.0001595949,
  9.847248e-06, 1.462597e-05, 3.700037e-05, 5.968481e-05, 6.311864e-05, 
    6.428445e-05, 7.913243e-05, 0.0001000488, 8.949627e-05, 0.0001067789, 
    8.945075e-05, 0.0001149981, 0.0001519886, 0.0001142933, 0.000121629,
  3.667738e-06, 8.831123e-06, 1.578429e-05, 2.790194e-05, 4.757717e-05, 
    6.045153e-05, 6.833218e-05, 9.058495e-05, 9.838428e-05, 0.0001095721, 
    0.0001274438, 0.0001418865, 0.0001329334, 0.0001458678, 0.000116365,
  4.210281e-07, 2.76604e-06, 1.262642e-05, 1.244441e-05, 3.816885e-05, 
    4.834896e-05, 4.441557e-05, 8.02902e-05, 7.777193e-05, 7.379502e-05, 
    0.0001067322, 0.000115333, 0.0001284358, 0.0001555622, 0.0001242501,
  6.18232e-06, 5.10167e-06, 4.114002e-06, 8.379117e-06, 1.63429e-05, 
    2.395679e-05, 3.126092e-05, 6.051021e-05, 9.180701e-05, 0.0001135708, 
    9.344565e-05, 0.000112799, 7.897476e-05, 0.0001060146, 0.0001435391,
  2.383898e-05, 2.076421e-05, 2.937174e-05, 1.74915e-05, 1.515278e-05, 
    1.700819e-05, 3.174947e-05, 4.251591e-05, 6.835604e-05, 5.009286e-05, 
    8.492094e-05, 0.0001092982, 0.0001171115, 9.465638e-05, 0.0001297598,
  8.062827e-06, 4.792452e-05, 6.06819e-05, 3.548605e-05, 1.961039e-05, 
    3.711659e-05, 3.966093e-05, 3.866599e-05, 4.188781e-05, 5.091182e-05, 
    8.135771e-05, 8.921321e-05, 0.0001232839, 0.0001106273, 8.867398e-05,
  1.952222e-06, 2.213445e-05, 2.202363e-05, 3.041391e-05, 3.838282e-05, 
    2.524394e-05, 2.640729e-05, 4.548625e-05, 5.765277e-05, 8.203503e-05, 
    7.267476e-05, 6.236321e-05, 7.477737e-05, 7.307263e-05, 7.100408e-05,
  3.870919e-08, 1.464912e-06, 1.4731e-05, 2.493126e-05, 3.266076e-05, 
    2.393948e-05, 2.17004e-05, 4.867023e-05, 5.098069e-05, 4.202716e-05, 
    6.137622e-05, 5.92535e-05, 5.348938e-05, 5.395756e-05, 5.133621e-05,
  3.839933e-06, 2.60229e-06, 5.743005e-06, 7.596465e-06, 7.114294e-06, 
    1.131179e-05, 9.457613e-06, 1.131009e-05, 1.974043e-05, 2.659553e-05, 
    4.021222e-05, 3.900493e-05, 3.622805e-05, 3.738197e-05, 3.36843e-05,
  8.330503e-06, 1.656871e-05, 2.472667e-05, 3.288631e-05, 2.191927e-05, 
    6.510473e-05, 7.247803e-05, 2.5671e-05, 7.370562e-05, 7.138222e-05, 
    9.311439e-05, 5.483063e-05, 8.081747e-05, 6.259923e-05, 0.0001159902,
  1.123075e-06, 1.238105e-06, 6.127742e-06, 1.493421e-05, 1.653913e-05, 
    2.693495e-05, 4.51608e-05, 4.959887e-05, 2.814245e-05, 5.274444e-05, 
    7.422922e-05, 8.851473e-05, 3.086502e-05, 4.577793e-05, 7.07289e-05,
  1.520855e-06, 5.697936e-07, 2.672837e-06, 2.898428e-06, 3.281397e-06, 
    4.647966e-06, 5.527622e-06, 1.293454e-05, 1.134525e-05, 1.545578e-05, 
    2.045338e-05, 5.202444e-05, 3.172694e-05, 2.628392e-05, 3.432717e-05,
  7.180782e-07, 5.398275e-07, 1.265527e-06, 4.287598e-06, 2.487964e-06, 
    5.101909e-06, 9.469953e-06, 1.085647e-05, 7.078629e-06, 1.13649e-05, 
    1.181325e-05, 3.275867e-05, 4.457064e-05, 1.58387e-05, 1.697861e-05,
  7.766442e-07, 7.955653e-07, 3.702135e-06, 3.935024e-06, 6.509777e-06, 
    2.41561e-06, 2.767224e-06, 1.04154e-05, 3.068991e-06, 1.495894e-05, 
    1.718132e-05, 2.126162e-06, 8.239108e-06, 1.099445e-05, 1.842852e-05,
  9.587709e-08, 1.155605e-06, 6.256148e-06, 2.13953e-06, 7.806366e-06, 
    9.488721e-06, 4.594018e-06, 1.248964e-05, 4.34327e-05, 3.481664e-05, 
    3.743335e-05, 4.794345e-05, 5.216848e-05, 1.295012e-05, 8.902295e-06,
  6.254796e-08, 7.853147e-07, 1.366021e-06, 5.050086e-06, 8.342486e-06, 
    1.208294e-05, 3.222959e-05, 4.561675e-05, 6.158204e-05, 5.484075e-05, 
    4.469865e-05, 5.623653e-05, 4.376648e-05, 2.01937e-05, 5.561138e-05,
  1.047873e-07, 2.141222e-07, 4.043187e-06, 3.904649e-06, 1.017459e-05, 
    2.166397e-05, 4.425522e-05, 6.506847e-05, 5.384099e-05, 7.154298e-05, 
    4.108567e-05, 3.445909e-05, 8.355866e-05, 9.240009e-05, 4.453736e-05,
  3.586932e-07, 2.633178e-06, 9.901713e-06, 1.494764e-05, 3.782021e-05, 
    3.426114e-05, 3.462939e-05, 2.5797e-05, 3.422059e-05, 5.706716e-05, 
    5.947996e-05, 4.569552e-05, 6.146096e-05, 6.251479e-05, 2.20763e-05,
  9.613888e-07, 1.151573e-06, 6.282606e-06, 9.429423e-06, 1.597125e-05, 
    1.541413e-05, 2.140336e-05, 2.054359e-05, 1.984196e-05, 2.306807e-05, 
    2.893424e-05, 3.157425e-05, 3.148587e-05, 4.289965e-05, 3.768271e-05,
  7.450545e-07, 1.26252e-06, 1.829668e-06, 1.95132e-06, 2.374625e-06, 
    3.498145e-06, 5.190871e-06, 6.914933e-06, 1.043604e-05, 1.448754e-05, 
    1.868689e-05, 2.286379e-05, 2.560982e-05, 2.939212e-05, 3.431274e-05,
  1.644826e-07, 4.298834e-07, 6.620697e-07, 8.478355e-07, 1.553699e-06, 
    1.55263e-06, 2.629482e-06, 2.984499e-06, 4.386543e-06, 7.73309e-06, 
    1.014725e-05, 1.291285e-05, 1.46575e-05, 2.160566e-05, 2.827779e-05,
  3.370466e-08, 4.388602e-07, 6.072548e-07, 1.05345e-06, 1.21564e-06, 
    1.307189e-06, 1.796124e-06, 3.124266e-06, 2.9314e-06, 5.730004e-06, 
    8.828517e-06, 1.034221e-05, 1.304261e-05, 1.290769e-05, 1.535706e-05,
  5.58919e-08, 1.538099e-07, 6.068836e-07, 4.383963e-07, 4.165331e-07, 
    5.759957e-07, 8.895001e-07, 1.372938e-06, 1.673672e-06, 2.475386e-06, 
    3.511707e-06, 4.429285e-06, 6.909333e-06, 7.645282e-06, 1.062468e-05,
  2.366662e-07, 1.770088e-07, 4.877489e-08, 6.825928e-08, 3.899749e-07, 
    3.901177e-07, 4.763974e-07, 8.87957e-07, 1.196284e-06, 1.053642e-06, 
    1.626456e-06, 2.048449e-06, 2.509896e-06, 3.194853e-06, 5.494316e-06,
  3.558834e-07, 5.810207e-07, 3.58437e-07, 5.173633e-07, 5.480389e-07, 
    5.287679e-07, 3.897631e-07, 5.206647e-07, 4.341306e-07, 6.020529e-07, 
    6.150829e-07, 1.07016e-06, 1.070381e-06, 1.764885e-06, 2.30932e-06,
  9.629596e-08, 2.73726e-07, 7.23293e-07, 1.077336e-06, 1.367336e-06, 
    1.210465e-06, 9.216154e-07, 1.037161e-06, 1.041748e-06, 5.28052e-07, 
    4.115097e-07, 1.244561e-07, 1.116051e-06, 5.811121e-07, 1.273945e-06,
  8.85422e-09, 2.89404e-07, 5.175208e-07, 7.692801e-07, 8.699656e-07, 
    1.236424e-06, 1.313364e-06, 1.229992e-06, 1.653297e-06, 2.031554e-06, 
    1.101719e-06, 1.254196e-06, 3.386454e-07, 3.717784e-07, 8.47765e-07,
  1.033089e-08, 2.754212e-08, 3.652225e-07, 6.141648e-07, 1.54843e-06, 
    1.501955e-06, 2.334636e-06, 1.807262e-06, 1.988047e-06, 3.321959e-06, 
    4.289398e-06, 6.228365e-06, 5.678132e-06, 7.178453e-06, 1.235345e-05,
  8.278213e-07, 8.996069e-07, 1.260385e-06, 1.368616e-06, 1.863297e-06, 
    3.316259e-06, 5.692831e-06, 5.892972e-06, 7.96921e-06, 7.759383e-06, 
    8.482514e-06, 1.722683e-05, 2.037881e-05, 1.684932e-05, 1.843899e-05,
  3.376265e-06, 2.779108e-06, 4.550954e-06, 4.556149e-06, 4.943236e-06, 
    4.779778e-06, 6.391303e-06, 7.181699e-06, 8.518846e-06, 9.644308e-06, 
    1.10786e-05, 1.227888e-05, 1.746525e-05, 3.063213e-05, 5.222414e-05,
  1.153113e-06, 1.057887e-06, 1.469473e-06, 1.664276e-06, 2.955653e-06, 
    3.383689e-06, 3.605863e-06, 4.374368e-06, 5.859452e-06, 8.260956e-06, 
    1.029575e-05, 9.150074e-06, 7.882909e-06, 9.791062e-06, 1.333081e-05,
  2.687373e-08, 2.289076e-07, 8.2283e-07, 1.211812e-06, 8.954304e-07, 
    1.385849e-06, 1.457661e-06, 2.785141e-06, 3.707522e-06, 4.945624e-06, 
    7.241605e-06, 8.921918e-06, 8.588902e-06, 9.020881e-06, 9.6771e-06,
  1.122193e-06, 1.901873e-07, 7.922711e-08, 5.608596e-08, 4.019766e-08, 
    1.058228e-06, 1.296072e-06, 7.21867e-07, 1.626861e-06, 2.656232e-06, 
    3.637996e-06, 5.702411e-06, 5.905419e-06, 7.520106e-06, 8.24302e-06,
  7.435063e-07, 4.782172e-07, 5.953006e-08, 3.574263e-09, 6.939219e-08, 
    3.681137e-08, 1.777388e-07, 3.292827e-07, 8.1514e-07, 9.691556e-07, 
    1.869205e-06, 2.806255e-06, 4.044828e-06, 5.145308e-06, 6.316669e-06,
  1.085577e-06, 5.963783e-08, 5.17947e-09, 5.878696e-08, 1.117572e-08, 
    1.775923e-07, 1.450122e-07, 1.794767e-07, 3.56802e-07, 4.755108e-07, 
    1.15735e-06, 1.875469e-06, 2.643303e-06, 3.066036e-06, 4.971349e-06,
  1.009367e-06, 1.437546e-07, 4.96639e-09, 6.013999e-09, 3.846063e-09, 
    1.333263e-08, 2.422329e-07, 4.272724e-07, 3.514463e-07, 7.516775e-08, 
    1.085126e-06, 9.676082e-07, 1.304438e-06, 1.761475e-06, 2.81749e-06,
  2.003873e-06, 1.484789e-07, 1.388105e-08, 6.269157e-09, 4.253253e-09, 
    1.408567e-08, 7.041537e-08, 6.694961e-08, 6.108225e-08, 6.900264e-07, 
    7.190554e-07, 1.108241e-06, 1.015353e-06, 9.829071e-07, 1.429263e-06,
  1.61137e-06, 1.061501e-07, 1.029718e-07, 1.57997e-07, 8.962725e-09, 
    8.315262e-09, 3.615878e-08, 2.604835e-08, 2.510407e-07, 1.072599e-06, 
    1.148609e-06, 9.689635e-07, 2.68061e-07, 1.637322e-07, 3.33625e-07,
  1.331198e-06, 6.131825e-07, 7.950285e-08, 2.690642e-08, 4.009383e-08, 
    3.348777e-08, 9.986059e-09, 1.731156e-07, 5.639549e-07, 7.116764e-07, 
    1.311645e-06, 6.136774e-07, 1.404566e-06, 1.364599e-06, 4.354885e-07,
  8.267315e-06, 7.701768e-06, 7.161652e-06, 7.058109e-06, 5.477201e-06, 
    4.827159e-06, 4.464733e-06, 5.679007e-06, 2.360226e-05, 6.180966e-05, 
    8.632152e-05, 6.374807e-05, 4.117642e-05, 4.021322e-05, 4.109626e-05,
  6.3602e-06, 5.122121e-06, 4.53748e-06, 5.377411e-06, 5.543899e-06, 
    4.66833e-06, 4.300243e-06, 5.736338e-06, 7.574396e-06, 1.080513e-05, 
    3.373413e-05, 5.406334e-05, 6.252274e-05, 4.47041e-05, 4.031728e-05,
  1.680716e-06, 7.752333e-07, 9.634637e-07, 1.423308e-06, 2.241934e-06, 
    4.550198e-06, 4.141722e-06, 2.644329e-06, 2.965033e-06, 3.515537e-06, 
    8.536453e-06, 2.189269e-05, 2.265778e-05, 3.984728e-05, 3.791937e-05,
  1.806471e-07, 2.506831e-07, 4.523269e-09, 1.284548e-07, 2.768705e-07, 
    1.794599e-06, 2.132329e-06, 1.872555e-06, 7.703829e-07, 3.785644e-07, 
    9.683285e-07, 2.879564e-06, 8.021215e-06, 1.190002e-05, 1.95221e-05,
  4.662024e-07, 4.426541e-07, 5.429275e-08, 4.475737e-08, 5.862748e-07, 
    3.773837e-07, 2.224437e-07, 3.335003e-07, 6.362836e-07, 1.773807e-06, 
    6.624179e-07, 7.841662e-07, 1.187397e-06, 2.382518e-06, 1.086193e-05,
  1.864524e-06, 2.258764e-06, 1.473024e-06, 8.026037e-08, 2.950928e-07, 
    8.067225e-08, 3.112857e-09, 1.297094e-07, 8.675028e-08, 1.165727e-06, 
    2.018824e-06, 1.262963e-06, 1.037785e-06, 2.036008e-06, 2.438173e-06,
  3.858995e-06, 2.361008e-06, 4.617663e-07, 1.270815e-07, 5.971484e-07, 
    8.682113e-08, 4.716584e-09, 4.0231e-07, 1.002666e-06, 3.460203e-07, 
    9.183373e-07, 1.643435e-06, 2.577474e-06, 1.887439e-06, 1.09855e-06,
  1.378342e-06, 1.978398e-06, 8.971527e-07, 4.72749e-08, 1.678407e-07, 
    3.345934e-08, 1.008748e-07, 1.629667e-07, 9.410781e-08, 5.749735e-07, 
    1.032871e-06, 2.24067e-06, 3.159097e-06, 2.658166e-06, 4.126586e-06,
  1.072464e-06, 1.867161e-06, 5.172988e-07, 3.563653e-08, 7.418265e-09, 
    6.573418e-08, 5.035337e-08, 3.469983e-08, 2.989956e-07, 8.543077e-07, 
    6.223701e-07, 1.024266e-06, 1.688943e-06, 2.525099e-06, 4.515919e-06,
  1.216364e-06, 5.608832e-07, 4.43227e-08, 1.043692e-07, 1.620383e-07, 
    2.872411e-07, 1.493291e-07, 1.653682e-07, 2.126274e-07, 6.196586e-07, 
    1.389419e-06, 4.955766e-07, 8.235658e-07, 1.165766e-06, 2.523809e-06,
  9.224987e-06, 8.668006e-06, 6.480285e-06, 6.674068e-06, 7.705243e-06, 
    8.776914e-06, 9.873798e-06, 1.639749e-05, 1.890823e-05, 2.229516e-05, 
    2.948392e-05, 4.422188e-05, 4.975811e-05, 3.966461e-05, 3.148388e-05,
  6.073215e-06, 7.129613e-06, 4.072397e-06, 3.722719e-06, 4.576628e-06, 
    4.436138e-06, 6.731012e-06, 7.937525e-06, 8.121197e-06, 8.259635e-06, 
    8.18897e-06, 1.056948e-05, 1.74178e-05, 2.518262e-05, 2.686665e-05,
  1.515388e-06, 8.816095e-07, 2.999017e-07, 4.106911e-07, 2.057433e-06, 
    3.980204e-06, 5.05247e-06, 7.122068e-06, 7.056055e-06, 7.381152e-06, 
    7.476707e-06, 4.829079e-06, 5.966979e-06, 1.121161e-05, 1.294795e-05,
  1.105889e-07, 1.125193e-07, 8.563738e-09, 1.890676e-07, 1.239689e-06, 
    2.831486e-06, 2.128786e-06, 3.175097e-06, 5.084575e-06, 5.895176e-06, 
    7.568126e-06, 5.766331e-06, 4.728112e-06, 1.838684e-06, 3.209947e-06,
  2.212347e-09, 2.70695e-12, 3.07895e-10, 1.641474e-07, 4.398537e-07, 
    7.4026e-07, 1.581803e-06, 4.302486e-07, 1.627771e-07, 9.02493e-07, 
    3.551019e-06, 1.649582e-06, 1.334639e-06, 3.525549e-07, 1.35655e-07,
  3.30496e-11, 1.869457e-12, 2.101205e-08, 2.690178e-08, 1.258058e-06, 
    2.319902e-06, 8.751232e-07, 2.142992e-07, 1.349581e-07, 5.830074e-07, 
    8.085279e-07, 8.452482e-07, 1.125129e-06, 8.803402e-07, 1.057629e-06,
  2.539298e-08, 2.881495e-10, 2.795508e-07, 9.141916e-07, 3.96504e-06, 
    3.388169e-06, 3.911095e-06, 2.855314e-06, 5.619455e-06, 5.221526e-06, 
    3.064142e-06, 3.400289e-06, 3.151374e-06, 5.301416e-06, 3.175753e-06,
  6.674574e-08, 9.816637e-08, 1.95705e-07, 2.85606e-06, 2.308483e-06, 
    4.939244e-06, 7.937981e-06, 3.8289e-06, 7.193068e-06, 6.384129e-06, 
    3.245263e-06, 5.439499e-06, 7.799344e-06, 6.653023e-06, 4.234903e-06,
  9.674417e-09, 2.469867e-08, 1.929163e-07, 4.505784e-06, 2.794225e-06, 
    3.250781e-06, 5.164388e-06, 2.833131e-06, 2.758616e-06, 5.563669e-06, 
    5.689536e-06, 5.429104e-06, 8.852253e-06, 7.361995e-06, 3.833634e-06,
  6.997375e-08, 9.899972e-09, 1.603184e-07, 4.973145e-06, 2.613137e-06, 
    2.734893e-06, 4.699412e-06, 4.977302e-06, 4.088261e-06, 2.586666e-06, 
    1.000124e-05, 8.66516e-06, 1.065124e-05, 3.351794e-06, 5.92521e-06,
  6.073172e-05, 6.444775e-05, 6.356581e-05, 5.718559e-05, 5.304979e-05, 
    5.026342e-05, 5.086121e-05, 4.49323e-05, 4.223522e-05, 3.524303e-05, 
    4.452358e-05, 5.458144e-05, 7.183099e-05, 0.0001022637, 0.0001564363,
  1.263714e-05, 1.987561e-05, 3.215062e-05, 3.791258e-05, 3.7799e-05, 
    3.961542e-05, 4.593231e-05, 3.689881e-05, 3.248457e-05, 2.854582e-05, 
    2.604524e-05, 2.450954e-05, 2.640362e-05, 3.235403e-05, 4.459972e-05,
  2.004795e-05, 2.53228e-05, 3.171648e-05, 3.203041e-05, 2.933501e-05, 
    2.894579e-05, 3.363572e-05, 3.52403e-05, 3.084008e-05, 2.99943e-05, 
    2.942326e-05, 2.628022e-05, 2.788136e-05, 3.305867e-05, 4.116981e-05,
  1.820565e-05, 2.53885e-05, 2.831603e-05, 2.268572e-05, 1.78764e-05, 
    1.687009e-05, 1.355606e-05, 1.764018e-05, 1.855813e-05, 2.38051e-05, 
    2.390649e-05, 2.439578e-05, 2.414024e-05, 2.758036e-05, 3.285263e-05,
  1.997169e-05, 2.638324e-05, 1.996282e-05, 1.227621e-05, 1.011359e-05, 
    8.368785e-06, 8.655885e-06, 1.105262e-05, 1.584385e-05, 1.884948e-05, 
    2.493226e-05, 2.416457e-05, 2.868697e-05, 2.445254e-05, 2.753699e-05,
  1.483652e-05, 1.800803e-05, 1.66333e-05, 1.019334e-05, 5.509818e-06, 
    5.42831e-06, 5.864833e-06, 8.907174e-06, 1.065609e-05, 1.179936e-05, 
    1.273572e-05, 1.320007e-05, 1.991026e-05, 2.289284e-05, 3.25698e-05,
  5.64324e-06, 1.55012e-05, 1.628889e-05, 1.293707e-05, 1.087427e-05, 
    8.653552e-06, 8.35394e-06, 1.205404e-05, 1.416581e-05, 1.139117e-05, 
    1.637241e-05, 2.077603e-05, 2.621366e-05, 3.240733e-05, 3.986865e-05,
  6.711061e-06, 1.384041e-05, 1.123097e-05, 9.976267e-06, 7.846758e-06, 
    1.17957e-05, 8.531303e-06, 1.570853e-05, 1.252972e-05, 6.736524e-06, 
    8.91017e-06, 1.60539e-05, 1.86108e-05, 2.429895e-05, 3.656134e-05,
  6.198733e-06, 1.500381e-05, 5.125774e-06, 4.671347e-06, 4.453737e-06, 
    9.646103e-06, 1.188543e-05, 7.633957e-06, 3.698949e-06, 4.854818e-06, 
    7.025142e-06, 9.907983e-06, 1.000211e-05, 1.613753e-05, 1.617459e-05,
  6.140398e-06, 9.753579e-06, 7.450267e-06, 5.21892e-06, 5.801578e-06, 
    6.737899e-06, 9.276325e-06, 7.091953e-06, 1.130994e-05, 1.009147e-05, 
    9.298441e-06, 7.457997e-06, 4.923001e-06, 5.491373e-06, 4.524084e-06,
  1.914215e-05, 2.007647e-05, 1.95278e-05, 1.819617e-05, 1.137767e-05, 
    1.750825e-05, 1.456177e-05, 1.392891e-05, 1.078466e-05, 1.127557e-05, 
    7.529422e-06, 4.579188e-06, 1.528728e-06, 7.534591e-07, 2.728986e-07,
  1.235814e-05, 1.952863e-05, 2.472527e-05, 2.871095e-05, 1.514574e-05, 
    1.136483e-05, 1.038934e-05, 1.326927e-05, 1.15609e-05, 1.38378e-05, 
    1.124777e-05, 6.047957e-06, 2.564424e-06, 2.09556e-06, 1.542747e-06,
  4.3531e-06, 1.307298e-05, 1.658881e-05, 1.793732e-05, 2.258963e-05, 
    1.507371e-05, 1.383664e-05, 2.041268e-05, 1.09714e-05, 1.4412e-05, 
    1.547216e-05, 1.022751e-05, 4.357595e-06, 3.584015e-06, 2.010545e-06,
  2.913492e-06, 6.383622e-06, 1.197909e-05, 1.254869e-05, 1.608349e-05, 
    2.157765e-05, 2.050157e-05, 1.31379e-05, 1.430565e-05, 1.727574e-05, 
    1.985655e-05, 1.368358e-05, 9.220731e-06, 4.766588e-06, 4.079658e-06,
  1.071161e-06, 3.898455e-06, 6.926697e-06, 1.426946e-05, 1.734936e-05, 
    1.716411e-05, 1.957788e-05, 1.777515e-05, 1.638301e-05, 1.693497e-05, 
    1.751712e-05, 2.171516e-05, 1.423561e-05, 9.316019e-06, 8.424168e-06,
  5.839518e-07, 1.172109e-06, 3.494393e-06, 9.440651e-06, 1.210113e-05, 
    1.486184e-05, 1.977282e-05, 2.238503e-05, 2.015142e-05, 1.687563e-05, 
    1.779242e-05, 1.394421e-05, 1.439119e-05, 1.943937e-05, 8.557577e-06,
  5.250736e-07, 6.178959e-07, 1.211042e-06, 4.104502e-06, 8.216217e-06, 
    1.258695e-05, 1.617473e-05, 1.936725e-05, 2.022461e-05, 1.528478e-05, 
    1.593632e-05, 1.340417e-05, 1.666821e-05, 2.291081e-05, 2.278048e-05,
  3.354406e-08, 3.612564e-08, 2.70735e-08, 1.83851e-06, 5.538931e-06, 
    8.387517e-06, 1.586538e-05, 1.601033e-05, 1.471172e-05, 1.461596e-05, 
    1.436388e-05, 1.747331e-05, 2.726026e-05, 3.623744e-05, 4.014263e-05,
  8.299638e-07, 5.744812e-07, 5.238926e-07, 1.230013e-06, 2.96524e-06, 
    1.077608e-05, 2.072503e-05, 2.035948e-05, 2.268995e-05, 3.499311e-05, 
    3.337256e-05, 4.203046e-05, 5.28792e-05, 5.173276e-05, 4.194514e-05,
  8.806574e-06, 1.250302e-05, 1.006468e-05, 8.044645e-06, 1.283265e-05, 
    2.440188e-05, 3.174607e-05, 4.050054e-05, 5.561695e-05, 6.572699e-05, 
    5.519811e-05, 6.722871e-05, 8.897133e-05, 9.201842e-05, 7.325839e-05,
  2.845408e-05, 1.104808e-05, 2.015988e-06, 3.990204e-06, 7.531118e-06, 
    1.083501e-05, 1.313486e-05, 1.231787e-05, 1.498731e-05, 1.234738e-05, 
    9.969959e-06, 1.045647e-05, 1.081676e-05, 1.137109e-05, 7.664971e-06,
  4.674221e-05, 6.359212e-06, 2.648771e-06, 1.481821e-06, 4.181762e-06, 
    7.489163e-06, 9.052096e-06, 1.397219e-05, 1.305126e-05, 1.286348e-05, 
    1.36468e-05, 9.114457e-06, 9.433241e-06, 1.143534e-05, 1.136192e-05,
  3.650467e-05, 1.225871e-05, 3.86266e-06, 1.249808e-06, 2.64023e-06, 
    5.177491e-06, 8.770811e-06, 1.154674e-05, 1.156494e-05, 1.312403e-05, 
    1.678432e-05, 1.178383e-05, 1.030647e-05, 1.057956e-05, 1.426699e-05,
  1.764203e-05, 1.530203e-05, 5.997228e-06, 2.425423e-06, 7.659475e-07, 
    3.306677e-06, 5.648442e-06, 8.250998e-06, 1.093916e-05, 1.03889e-05, 
    1.135987e-05, 1.181719e-05, 1.28308e-05, 1.29312e-05, 9.29606e-06,
  2.80447e-05, 2.166366e-05, 6.636244e-06, 7.977417e-06, 5.154914e-07, 
    1.909954e-08, 3.091831e-06, 6.641572e-06, 9.373037e-06, 8.374403e-06, 
    1.145617e-05, 1.29305e-05, 1.381618e-05, 9.568949e-06, 1.331141e-05,
  1.430535e-05, 1.081883e-05, 1.263005e-05, 4.883649e-06, 3.560782e-06, 
    1.628556e-08, 1.78916e-06, 3.469911e-06, 6.714701e-06, 7.371382e-06, 
    8.788619e-06, 1.242283e-05, 1.366184e-05, 1.387008e-05, 1.3812e-05,
  1.884568e-05, 8.850413e-06, 1.002291e-05, 8.832301e-06, 5.753448e-06, 
    4.69962e-06, 1.141171e-06, 2.930651e-06, 5.253009e-06, 6.608641e-06, 
    7.976787e-06, 8.41783e-06, 1.24533e-05, 1.857606e-05, 1.682516e-05,
  1.196337e-05, 1.169619e-05, 9.444044e-06, 1.374558e-05, 1.146957e-05, 
    5.383577e-06, 3.398084e-06, 1.142578e-06, 4.13144e-06, 4.474758e-06, 
    7.557356e-06, 8.949268e-06, 9.053007e-06, 8.935574e-06, 1.106683e-05,
  4.909595e-06, 1.169577e-05, 1.121969e-05, 1.704312e-05, 1.694517e-05, 
    1.47274e-05, 5.813543e-06, 2.661012e-06, 7.005655e-07, 3.355802e-06, 
    3.136333e-06, 8.693813e-06, 9.234546e-06, 8.968881e-06, 8.277667e-06,
  5.376975e-06, 6.102874e-06, 9.954566e-06, 2.040289e-05, 2.872506e-05, 
    3.459223e-05, 2.711669e-05, 9.171073e-06, 2.352852e-06, 2.181109e-06, 
    6.176131e-07, 3.413455e-06, 5.517819e-06, 8.017986e-06, 9.410774e-06,
  0.0008204607, 0.0007410458, 0.0007007229, 0.000686562, 0.0006639893, 
    0.0006545869, 0.0005197831, 0.0003528311, 0.000213122, 0.0001182258, 
    4.562347e-05, 1.64405e-05, 9.940379e-06, 9.519269e-06, 1.047541e-05,
  0.0005974846, 0.0005976605, 0.0005717739, 0.0005648016, 0.0005770598, 
    0.0005389, 0.0004524497, 0.0003231522, 0.0002208742, 0.0001260501, 
    6.047108e-05, 2.001673e-05, 7.612842e-06, 7.954701e-06, 8.753642e-06,
  0.0003267088, 0.0003860499, 0.0003811633, 0.0003654301, 0.0003657583, 
    0.0003531261, 0.0002925849, 0.0001994513, 0.0001516004, 8.381508e-05, 
    4.271055e-05, 1.814053e-05, 7.250979e-06, 5.966661e-06, 7.404468e-06,
  6.86486e-05, 0.0001491766, 0.000168308, 0.0001801795, 0.0001960505, 
    0.0001697096, 0.0001200588, 7.686342e-05, 6.031808e-05, 3.52327e-05, 
    1.441473e-05, 9.764288e-06, 7.482035e-06, 5.008998e-06, 5.17076e-06,
  1.564767e-05, 2.348179e-05, 3.227219e-05, 2.616465e-05, 4.429732e-05, 
    3.810759e-05, 2.947731e-05, 2.420909e-05, 2.36591e-05, 2.028595e-05, 
    1.485557e-05, 1.176374e-05, 6.698167e-06, 5.928183e-06, 6.783448e-06,
  3.305603e-05, 1.806329e-05, 1.575431e-05, 1.195949e-05, 3.773593e-06, 
    3.935728e-06, 1.328427e-05, 1.356764e-05, 1.865508e-05, 1.311041e-05, 
    9.803902e-06, 9.391852e-06, 9.888109e-06, 7.593379e-06, 6.698571e-06,
  3.473722e-05, 2.321853e-05, 1.45977e-05, 6.821869e-06, 4.615136e-06, 
    2.948344e-06, 3.401416e-05, 2.104272e-05, 3.041778e-05, 8.264813e-06, 
    8.589982e-06, 1.203243e-05, 1.312126e-05, 9.841738e-06, 8.753125e-06,
  2.364105e-05, 3.090771e-05, 4.149597e-05, 1.240313e-05, 3.993681e-05, 
    0.0001308023, 9.006645e-05, 2.203233e-05, 6.665418e-06, 3.581295e-06, 
    8.481859e-06, 1.119445e-05, 1.250484e-05, 1.144202e-05, 1.03113e-05,
  2.61168e-05, 2.042255e-05, 3.972127e-05, 4.016761e-05, 9.810267e-05, 
    0.0001933418, 8.998939e-05, 1.391483e-05, 3.443405e-06, 1.993593e-06, 
    5.032242e-06, 1.074322e-05, 1.331633e-05, 1.132442e-05, 1.03854e-05,
  2.127456e-05, 2.341238e-05, 1.593402e-05, 1.964457e-05, 7.404312e-05, 
    0.0001207629, 5.218324e-05, 1.320767e-05, 1.394107e-06, 6.385411e-07, 
    2.329172e-06, 9.165855e-06, 1.170938e-05, 1.030172e-05, 1.006852e-05,
  7.214716e-06, 1.178537e-05, 1.53835e-05, 1.986461e-05, 2.571124e-05, 
    7.848105e-05, 0.0001569123, 0.0002426697, 0.0003623621, 0.0004273512, 
    0.000374291, 0.0002630326, 0.0001655286, 9.797537e-05, 7.175935e-05,
  5.086972e-06, 1.097164e-05, 1.219783e-05, 2.159659e-05, 2.956322e-05, 
    5.833014e-05, 0.0001032629, 0.0001860861, 0.0002842626, 0.0003269723, 
    0.0003210596, 0.0002354321, 0.0001226918, 5.466751e-05, 3.737788e-05,
  4.976023e-06, 5.472884e-06, 1.343279e-05, 1.673106e-05, 1.573355e-05, 
    3.315053e-05, 6.868517e-05, 0.0001205016, 0.0001774381, 0.0002195915, 
    0.0002052288, 0.0001478298, 8.608549e-05, 3.960045e-05, 2.640082e-05,
  3.784225e-06, 6.13335e-06, 5.351743e-06, 7.738902e-06, 1.448078e-05, 
    2.163682e-05, 4.881238e-05, 6.81129e-05, 9.140313e-05, 0.0001269861, 
    0.0001388556, 0.0001003184, 7.535877e-05, 4.61511e-05, 2.913697e-05,
  3.178269e-06, 3.898067e-06, 3.479273e-06, 6.947523e-06, 1.122995e-05, 
    1.838968e-05, 3.857285e-05, 5.2582e-05, 6.019484e-05, 9.451127e-05, 
    0.0001091853, 8.965265e-05, 6.968775e-05, 7.59822e-05, 6.764221e-05,
  1.33261e-06, 2.277814e-06, 2.253755e-06, 4.755569e-06, 4.643876e-06, 
    8.590059e-06, 2.407973e-05, 4.102357e-05, 4.456543e-05, 6.351358e-05, 
    7.032973e-05, 5.74817e-05, 6.555126e-05, 0.0001258967, 0.0001453269,
  8.045149e-07, 1.562257e-06, 2.550429e-06, 3.014546e-06, 1.055367e-05, 
    1.912047e-05, 1.090689e-05, 4.631539e-05, 9.658313e-05, 0.0001139968, 
    3.119513e-05, 3.393973e-05, 7.19861e-05, 0.0001775576, 0.000233478,
  7.170172e-07, 1.682319e-06, 2.073002e-06, 2.238248e-05, 2.445374e-05, 
    6.3859e-05, 2.971745e-05, 7.348586e-05, 0.000105307, 6.874493e-05, 
    1.973978e-05, 3.079042e-05, 9.915001e-05, 0.0002076391, 0.0002432093,
  1.03978e-06, 1.658394e-06, 8.25203e-06, 2.217091e-05, 3.35716e-05, 
    5.220336e-05, 8.325917e-05, 6.490628e-05, 7.361598e-05, 6.863442e-05, 
    2.574887e-05, 4.578634e-05, 0.0001142929, 0.0001839335, 0.000156567,
  2.139742e-06, 5.106665e-06, 1.33484e-05, 2.018244e-05, 3.673744e-05, 
    3.30332e-05, 6.954254e-05, 8.89865e-05, 5.515123e-05, 4.906498e-05, 
    6.460202e-05, 9.800616e-05, 0.0001832766, 0.0001138547, 7.854751e-05,
  3.994264e-06, 5.824789e-06, 1.022568e-05, 1.304002e-05, 1.675199e-05, 
    1.494405e-05, 2.481672e-05, 3.4262e-05, 4.165321e-05, 4.91631e-05, 
    4.780122e-05, 4.011026e-05, 5.728119e-05, 7.002206e-05, 6.546885e-05,
  4.982195e-06, 5.233675e-06, 6.824959e-06, 1.103418e-05, 1.221665e-05, 
    1.542476e-05, 1.741035e-05, 2.258007e-05, 3.412249e-05, 4.487481e-05, 
    4.595328e-05, 4.503758e-05, 6.163921e-05, 6.129121e-05, 5.984274e-05,
  8.739678e-06, 1.120212e-05, 8.014908e-06, 7.722972e-06, 8.880438e-06, 
    1.142866e-05, 1.366467e-05, 1.832275e-05, 2.251093e-05, 3.427533e-05, 
    3.494084e-05, 3.707394e-05, 4.74525e-05, 4.802869e-05, 4.372939e-05,
  1.178663e-05, 9.415688e-06, 9.442957e-06, 8.369992e-06, 8.725839e-06, 
    8.466026e-06, 1.077273e-05, 1.131132e-05, 1.22994e-05, 2.048761e-05, 
    2.82918e-05, 3.104231e-05, 3.38983e-05, 4.392702e-05, 6.684411e-05,
  1.307013e-05, 1.371875e-05, 1.444312e-05, 9.943323e-06, 1.388036e-05, 
    1.026864e-05, 8.805713e-06, 1.074681e-05, 1.188435e-05, 1.165714e-05, 
    1.639437e-05, 1.72612e-05, 2.314375e-05, 4.338684e-05, 0.0001040801,
  1.092232e-05, 1.296524e-05, 1.243534e-05, 1.307627e-05, 1.025601e-05, 
    1.09782e-05, 1.049917e-05, 9.694559e-06, 1.179992e-05, 1.048668e-05, 
    1.005524e-05, 1.513289e-05, 2.042332e-05, 3.621698e-05, 0.0001235709,
  9.035328e-06, 1.342563e-05, 1.698703e-05, 6.70467e-06, 1.100014e-05, 
    1.155262e-05, 1.076925e-05, 1.271944e-05, 1.218419e-05, 1.140543e-05, 
    1.39144e-05, 1.227208e-05, 1.559182e-05, 2.382397e-05, 0.0001052357,
  5.84884e-06, 1.217253e-05, 1.434527e-05, 1.223051e-05, 1.604338e-05, 
    1.232495e-05, 1.244846e-05, 1.365792e-05, 1.199878e-05, 1.261917e-05, 
    1.242398e-05, 1.135894e-05, 1.256722e-05, 3.153424e-05, 6.640373e-05,
  3.720097e-06, 8.546734e-06, 1.452783e-05, 1.658081e-05, 1.575295e-05, 
    1.603794e-05, 1.609579e-05, 1.289259e-05, 1.171564e-05, 1.307039e-05, 
    1.367201e-05, 1.087572e-05, 1.676181e-05, 3.735106e-05, 9.308934e-05,
  4.215235e-06, 9.240734e-06, 1.39121e-05, 1.400118e-05, 1.764588e-05, 
    2.083777e-05, 2.037154e-05, 1.574127e-05, 1.195512e-05, 1.208013e-05, 
    1.215807e-05, 1.155895e-05, 2.319197e-05, 5.861229e-05, 8.389397e-05,
  3.82076e-06, 4.474318e-06, 1.036096e-05, 1.79645e-05, 2.828164e-05, 
    3.449094e-05, 5.255722e-05, 6.306714e-05, 5.687066e-05, 5.625783e-05, 
    7.01667e-05, 0.0001026193, 0.0001609503, 0.0002355105, 0.0002749732,
  2.070845e-06, 4.61522e-06, 8.671157e-06, 1.411257e-05, 2.399534e-05, 
    3.974116e-05, 4.499775e-05, 6.013877e-05, 6.648929e-05, 7.477555e-05, 
    8.3974e-05, 0.0001115289, 0.0001900132, 0.0002569746, 0.0002597793,
  8.432791e-07, 1.964107e-06, 5.092164e-06, 8.318e-06, 1.511808e-05, 
    3.149096e-05, 4.137901e-05, 5.640407e-05, 6.83947e-05, 8.905068e-05, 
    9.647452e-05, 0.0001490264, 0.0001972124, 0.0002339937, 0.0001814438,
  5.232151e-07, 1.620427e-06, 3.004869e-06, 7.147463e-06, 1.342003e-05, 
    2.419157e-05, 3.90217e-05, 4.949889e-05, 6.983768e-05, 6.856443e-05, 
    7.602727e-05, 0.0001331446, 0.0001653794, 0.0001683465, 0.0001463551,
  9.462807e-07, 1.181296e-06, 2.503193e-06, 5.469696e-06, 8.89966e-06, 
    1.627223e-05, 3.31863e-05, 4.646285e-05, 6.90216e-05, 7.727162e-05, 
    0.0001078632, 0.0001234349, 0.0001547057, 0.0001401231, 0.0001020598,
  1.424599e-06, 1.058487e-06, 1.728887e-06, 4.116138e-06, 7.397684e-06, 
    1.289844e-05, 2.604523e-05, 4.344742e-05, 5.58003e-05, 9.258775e-05, 
    0.0001012413, 0.0001125105, 0.0001313457, 0.0001242231, 0.0001025427,
  2.868657e-06, 2.470001e-06, 2.359106e-06, 8.188046e-06, 5.785021e-06, 
    1.09563e-05, 2.079033e-05, 3.969284e-05, 6.055645e-05, 7.768709e-05, 
    7.536806e-05, 9.822231e-05, 0.0001080177, 0.0001108194, 8.755588e-05,
  3.648615e-06, 1.675842e-06, 2.965433e-06, 4.38015e-06, 8.941526e-06, 
    1.263174e-05, 1.895137e-05, 2.716849e-05, 4.76752e-05, 6.563612e-05, 
    7.154077e-05, 0.0001060246, 0.0001239278, 0.0001073938, 7.801025e-05,
  1.708904e-06, 1.584309e-06, 2.832145e-06, 3.82882e-06, 6.613388e-06, 
    1.113145e-05, 1.208929e-05, 1.867453e-05, 3.046378e-05, 4.778187e-05, 
    7.151591e-05, 8.502689e-05, 0.0001107743, 0.0001260761, 0.0001086853,
  1.215488e-06, 1.650227e-06, 2.805361e-06, 3.773196e-06, 5.058037e-06, 
    7.451119e-06, 1.177254e-05, 1.721067e-05, 2.160566e-05, 3.09495e-05, 
    4.841161e-05, 6.041423e-05, 7.126544e-05, 0.0001012881, 7.456292e-05,
  1.730386e-07, 1.669008e-07, 1.966887e-07, 6.147354e-07, 2.174851e-06, 
    4.72901e-06, 8.582772e-06, 1.723476e-05, 2.792964e-05, 5.105032e-05, 
    5.939473e-05, 8.519828e-05, 9.251457e-05, 6.288842e-05, 4.87787e-05,
  4.235843e-08, 3.707517e-08, 1.820469e-07, 8.119224e-07, 2.799594e-06, 
    3.828831e-06, 7.761112e-06, 1.944971e-05, 2.624543e-05, 3.914832e-05, 
    6.039668e-05, 8.522592e-05, 0.0001082901, 8.069335e-05, 5.881304e-05,
  2.25992e-09, 5.118351e-08, 1.440139e-07, 3.430449e-07, 1.396712e-06, 
    3.183237e-06, 6.95842e-06, 1.342446e-05, 1.986733e-05, 3.457621e-05, 
    4.959922e-05, 8.540091e-05, 0.0001149849, 0.0001078952, 7.986058e-05,
  8.511628e-09, 9.220843e-09, 7.898046e-08, 2.452133e-07, 9.440829e-07, 
    3.081225e-06, 6.84634e-06, 1.071873e-05, 1.727591e-05, 2.458772e-05, 
    4.093396e-05, 6.803381e-05, 6.58284e-05, 0.0001251352, 8.065722e-05,
  2.764048e-08, 1.025766e-09, 8.234421e-08, 1.915443e-07, 8.685211e-07, 
    1.727386e-06, 5.642759e-06, 9.771657e-06, 1.417771e-05, 1.847488e-05, 
    3.328422e-05, 3.760158e-05, 9.084848e-05, 9.851769e-05, 8.335165e-05,
  5.833035e-08, 9.509498e-09, 3.800818e-08, 1.554144e-07, 8.42586e-07, 
    1.918228e-06, 4.782753e-06, 7.55426e-06, 1.029158e-05, 1.776049e-05, 
    2.216065e-05, 5.393289e-05, 7.274599e-05, 6.410289e-05, 8.42514e-05,
  5.340906e-08, 7.107403e-09, 3.753469e-08, 1.25633e-07, 3.68931e-07, 
    1.787141e-06, 3.00631e-06, 7.43157e-06, 1.241067e-05, 1.622846e-05, 
    1.825617e-05, 3.429345e-05, 5.013915e-05, 5.872558e-05, 6.680582e-05,
  7.884668e-08, 1.335074e-08, 1.499995e-08, 2.97873e-07, 5.110317e-07, 
    1.301079e-06, 3.110566e-06, 5.036034e-06, 8.023171e-06, 1.415682e-05, 
    1.824901e-05, 1.853841e-05, 3.46386e-05, 4.281734e-05, 5.149652e-05,
  1.423505e-07, 2.003013e-08, 1.214846e-07, 1.32722e-07, 3.422664e-07, 
    7.48423e-07, 2.039354e-06, 4.688352e-06, 6.3477e-06, 1.240089e-05, 
    1.840674e-05, 2.21382e-05, 2.236144e-05, 2.942751e-05, 3.688573e-05,
  2.190269e-08, 5.321121e-09, 1.133443e-07, 3.837997e-07, 2.558874e-07, 
    9.913856e-07, 1.563968e-06, 3.46244e-06, 5.117183e-06, 1.020253e-05, 
    1.593507e-05, 2.586294e-05, 3.164598e-05, 3.60817e-05, 7.275441e-05,
  4.481505e-06, 6.330572e-06, 9.774267e-06, 1.073294e-05, 1.043654e-05, 
    9.311239e-06, 7.316958e-06, 7.806281e-06, 1.307548e-05, 4.341733e-05, 
    0.0001033421, 0.0001094412, 7.323e-05, 3.74701e-05, 2.014808e-05,
  5.229269e-06, 7.551164e-06, 1.136487e-05, 1.218442e-05, 1.397369e-05, 
    1.324058e-05, 9.120202e-06, 4.656316e-06, 7.303333e-06, 1.516995e-05, 
    3.680065e-05, 7.143188e-05, 8.872725e-05, 7.233366e-05, 3.989539e-05,
  4.232915e-07, 2.854063e-06, 1.009377e-05, 1.489276e-05, 1.240921e-05, 
    1.339379e-05, 1.169573e-05, 7.140955e-06, 5.925905e-06, 7.642214e-06, 
    1.418991e-05, 2.748797e-05, 5.223817e-05, 6.990208e-05, 6.365393e-05,
  6.385429e-07, 2.388747e-07, 1.276182e-06, 3.646917e-06, 5.024137e-06, 
    5.273983e-06, 7.744997e-06, 7.145373e-06, 5.177896e-06, 4.604806e-06, 
    5.62634e-06, 9.22289e-06, 1.737388e-05, 2.94985e-05, 4.589944e-05,
  4.068415e-07, 3.212757e-07, 2.032787e-07, 3.074162e-07, 3.074491e-07, 
    4.571583e-07, 7.207737e-07, 1.816465e-06, 9.696931e-07, 7.641951e-07, 
    6.960367e-07, 4.254093e-06, 7.090587e-06, 1.174207e-05, 1.722003e-05,
  4.618249e-07, 1.472367e-07, 4.301332e-08, 1.68392e-07, 1.091052e-08, 
    5.315885e-08, 8.502301e-08, 5.919659e-07, 1.886407e-07, 3.097117e-07, 
    1.186602e-06, 2.621066e-06, 5.140144e-06, 6.786192e-06, 1.113832e-05,
  3.05583e-07, 9.644904e-08, 3.274705e-06, 1.294292e-06, 1.39862e-06, 
    4.568811e-08, 1.370126e-07, 3.894574e-07, 7.972783e-08, 3.538226e-07, 
    1.322207e-06, 1.82572e-06, 5.444116e-06, 4.604514e-06, 8.307111e-06,
  1.474089e-06, 3.237604e-07, 2.906263e-06, 5.064799e-07, 1.434213e-08, 
    1.141916e-07, 3.931561e-07, 1.86247e-07, 1.689311e-07, 7.836464e-08, 
    9.921727e-07, 1.699598e-06, 4.420601e-06, 3.712354e-06, 7.067552e-06,
  3.537309e-06, 2.234635e-06, 2.239519e-06, 1.361275e-07, 1.591706e-08, 
    3.398215e-07, 3.966614e-08, 7.746873e-08, 4.160071e-09, 2.796397e-07, 
    6.75586e-07, 1.671531e-06, 3.061298e-06, 4.532313e-06, 6.695492e-06,
  3.294403e-06, 3.194794e-06, 4.828933e-07, 1.400406e-08, 1.496162e-11, 
    4.404621e-10, 6.421256e-13, 5.440368e-12, 1.817397e-10, 3.49408e-07, 
    6.403914e-07, 5.40887e-07, 2.925555e-06, 2.415841e-06, 6.65429e-06,
  9.311419e-07, 2.924308e-06, 8.02862e-06, 1.552642e-05, 1.880233e-05, 
    2.544066e-05, 2.424475e-05, 1.536043e-05, 6.016575e-06, 2.148595e-06, 
    1.437037e-06, 2.861878e-06, 9.657235e-07, 1.1894e-07, 1.170476e-06,
  2.38971e-05, 1.253188e-05, 8.973798e-06, 1.672566e-05, 2.356938e-05, 
    2.740662e-05, 2.193687e-05, 1.164178e-05, 6.318553e-06, 4.405612e-06, 
    2.462107e-06, 4.203687e-06, 3.443724e-06, 5.394298e-07, 5.413822e-07,
  4.704974e-06, 3.038137e-06, 6.308551e-06, 1.317695e-05, 2.000746e-05, 
    1.60795e-05, 9.603856e-06, 6.335952e-06, 5.484142e-06, 6.519974e-06, 
    4.853785e-06, 5.311022e-06, 3.857821e-06, 3.497063e-06, 2.170383e-06,
  2.910085e-05, 1.454778e-05, 8.340826e-06, 6.570349e-06, 5.282136e-06, 
    1.171916e-05, 1.512849e-05, 1.52278e-05, 1.54211e-05, 1.270685e-05, 
    1.199109e-05, 1.114018e-05, 8.918469e-06, 8.324588e-06, 5.636372e-06,
  1.102519e-05, 8.805984e-06, 1.0119e-07, 1.246266e-06, 6.296613e-07, 
    4.605811e-07, 4.792402e-06, 6.909314e-06, 1.744056e-05, 2.303915e-05, 
    2.07912e-05, 1.248142e-05, 1.254846e-05, 1.346472e-05, 1.143807e-05,
  1.261502e-08, 1.047087e-08, 7.206482e-09, 2.884532e-09, 1.667598e-09, 
    3.927497e-08, 9.004529e-07, 3.386946e-06, 5.694025e-06, 3.391589e-06, 
    6.637834e-06, 5.580751e-06, 2.065208e-05, 1.51712e-05, 1.753724e-05,
  3.54882e-09, 1.193765e-09, 7.53254e-10, 6.035086e-08, 1.879725e-06, 
    5.159216e-07, 5.914881e-07, 5.001516e-07, 1.408102e-06, 2.558992e-06, 
    3.020325e-06, 4.604205e-06, 9.418695e-06, 9.448227e-06, 1.336746e-05,
  3.231576e-10, 4.417997e-08, 5.507306e-07, 3.183148e-06, 2.664392e-06, 
    1.742703e-06, 2.566178e-06, 3.289156e-06, 1.104244e-06, 2.63228e-06, 
    6.035453e-06, 5.174502e-06, 5.496911e-06, 5.980643e-06, 1.282575e-05,
  1.934153e-08, 9.854894e-07, 3.145685e-06, 3.662261e-06, 4.515007e-06, 
    4.446753e-06, 3.876621e-06, 3.754745e-06, 2.006311e-06, 3.346805e-06, 
    3.905912e-06, 2.3491e-06, 2.307991e-06, 1.950552e-06, 2.48973e-06,
  2.064427e-07, 2.33601e-06, 1.88847e-06, 1.244497e-06, 1.713852e-06, 
    3.535708e-06, 3.917281e-06, 3.361447e-06, 3.252769e-06, 4.854112e-07, 
    2.5839e-08, 5.554608e-07, 2.762513e-07, 1.219044e-06, 3.783199e-06,
  7.797783e-06, 8.523811e-06, 9.632059e-06, 1.057171e-05, 9.853402e-06, 
    1.02619e-05, 2.454893e-05, 4.863057e-05, 8.324584e-05, 0.0001129697, 
    0.0001552395, 0.0002091004, 0.0002612806, 0.0002834701, 0.000291088,
  2.878791e-06, 2.013661e-06, 2.067368e-06, 1.900825e-06, 5.920389e-06, 
    1.705959e-05, 4.742697e-05, 9.364507e-05, 0.0001415933, 0.0001847015, 
    0.0002326901, 0.0002622083, 0.0002745768, 0.000233946, 0.0002420217,
  1.437167e-05, 1.090676e-05, 7.086573e-06, 1.269964e-05, 2.17355e-05, 
    4.781238e-05, 9.970277e-05, 0.0001650026, 0.0002129537, 0.0002504203, 
    0.000269522, 0.0002637309, 0.0002264857, 0.0002033224, 0.0001418684,
  6.250555e-05, 5.625932e-05, 8.760727e-05, 0.0001083176, 0.0001263424, 
    0.00016824, 0.0002200116, 0.0002719828, 0.0002841573, 0.000306885, 
    0.0002787477, 0.0002266515, 0.000186058, 0.0001116548, 0.0001291759,
  7.515227e-05, 0.0001335328, 0.0002561722, 0.0001919228, 0.0002742756, 
    0.0003350443, 0.0003765031, 0.0003586767, 0.0003342216, 0.0002623343, 
    0.0002250373, 0.0001742517, 0.0001230976, 0.0001086258, 0.0001016915,
  7.004105e-05, 0.0001903022, 0.0002041122, 0.000295959, 0.00028545, 
    0.0003211613, 0.0003355978, 0.0003201989, 0.0002862581, 0.000236595, 
    0.0002042662, 0.0001659353, 0.0001073209, 6.709845e-05, 0.0001131936,
  3.671687e-05, 0.0001004444, 0.0001646378, 0.0002149089, 0.0002494048, 
    0.0002939046, 0.0002829316, 0.0002686603, 0.0002687783, 0.0002243954, 
    0.000186113, 0.0001489449, 0.000115756, 8.81169e-05, 7.162958e-05,
  1.7333e-05, 0.0001067622, 0.0001133944, 0.0001641175, 0.0002037325, 
    0.0002230991, 0.0002405022, 0.0002372156, 0.0002303201, 0.0002009134, 
    0.0001582387, 0.0001305814, 7.877938e-05, 7.459192e-05, 5.960676e-05,
  8.631002e-06, 7.969823e-05, 8.899141e-05, 0.0001173962, 0.000140711, 
    0.0001664013, 0.0001919472, 0.0001976104, 0.0002020009, 0.0001736195, 
    0.0001262284, 8.413978e-05, 5.789306e-05, 5.883647e-05, 7.700299e-05,
  5.431502e-06, 7.657176e-05, 6.371586e-05, 7.479246e-05, 9.498589e-05, 
    0.0001088673, 0.0001345887, 0.0001598136, 0.0001422314, 0.0001178126, 
    7.635283e-05, 4.376696e-05, 3.54875e-05, 5.571117e-05, 6.805811e-05,
  8.214858e-06, 8.390267e-06, 9.544552e-06, 1.156824e-05, 2.154913e-05, 
    2.854382e-05, 3.499598e-05, 3.280686e-05, 4.483225e-05, 5.741269e-05, 
    5.224955e-05, 9.66681e-05, 0.0001369464, 0.0001024532, 7.961981e-05,
  5.523585e-06, 7.174314e-06, 6.958786e-06, 9.123302e-06, 1.085324e-05, 
    1.07358e-05, 9.313048e-06, 3.163774e-05, 4.058642e-05, 4.330766e-05, 
    5.336357e-05, 4.98488e-05, 7.34324e-05, 4.123759e-05, 0.0001182753,
  4.836471e-06, 4.29757e-06, 5.85133e-06, 5.104926e-06, 5.297207e-06, 
    5.270474e-06, 1.225541e-05, 1.296371e-05, 2.899474e-05, 3.22857e-05, 
    2.763691e-05, 4.855119e-05, 5.86759e-05, 3.564095e-05, 2.410994e-05,
  5.600629e-06, 3.673646e-06, 6.459374e-06, 3.045818e-06, 4.984458e-06, 
    5.001558e-06, 6.540233e-06, 1.181539e-05, 9.162221e-06, 1.232095e-05, 
    3.016374e-05, 3.09023e-05, 1.597862e-05, 1.36269e-05, 3.665156e-06,
  4.52553e-06, 4.336317e-06, 4.674559e-06, 5.065384e-06, 3.02609e-06, 
    6.275081e-06, 4.51112e-06, 7.508983e-06, 9.402236e-06, 8.749088e-06, 
    9.693788e-06, 8.721076e-06, 3.236852e-06, 3.190318e-06, 2.661409e-06,
  5.421217e-06, 4.032439e-06, 5.639925e-06, 5.195911e-06, 2.776871e-06, 
    3.940445e-06, 3.410283e-06, 4.763212e-06, 2.477389e-06, 2.939272e-06, 
    2.925901e-06, 1.823357e-06, 1.903641e-06, 2.694998e-06, 2.642e-06,
  3.573864e-06, 4.700591e-06, 5.035818e-06, 3.113604e-06, 2.330932e-06, 
    2.146667e-06, 1.958137e-06, 1.78582e-06, 2.501486e-06, 1.213716e-06, 
    2.498195e-06, 1.66407e-06, 2.323921e-06, 2.690519e-06, 2.917372e-06,
  2.965107e-06, 2.808981e-06, 1.486275e-06, 7.702386e-07, 6.526959e-07, 
    1.358112e-06, 1.3722e-06, 1.676796e-06, 2.084153e-06, 2.970472e-06, 
    1.973041e-06, 1.818299e-06, 2.931147e-06, 4.812758e-06, 5.217233e-06,
  2.142094e-06, 9.65023e-07, 4.12022e-07, 1.892139e-08, 3.521146e-07, 
    1.210094e-06, 2.091347e-06, 2.468134e-06, 1.563336e-06, 1.2303e-06, 
    1.65592e-06, 2.022061e-06, 3.31192e-06, 6.060437e-06, 5.971427e-06,
  5.844653e-07, 3.840737e-10, 8.740169e-09, 2.071917e-08, 5.173332e-07, 
    1.603201e-06, 2.515684e-06, 2.272038e-06, 1.547396e-06, 7.515845e-07, 
    6.475552e-07, 7.843497e-07, 2.55436e-06, 2.285585e-06, 3.895197e-06,
  3.075785e-06, 2.600854e-06, 2.332834e-06, 8.104328e-07, 1.509799e-06, 
    1.09427e-06, 1.721701e-06, 3.085777e-06, 3.715438e-06, 3.79294e-06, 
    4.990526e-06, 5.816888e-06, 1.172875e-05, 1.348731e-05, 9.133474e-06,
  1.607155e-06, 9.618007e-07, 9.421838e-07, 1.445019e-06, 1.841171e-06, 
    1.243104e-06, 1.084366e-06, 1.092054e-06, 1.776471e-06, 2.223783e-06, 
    2.59338e-06, 3.276158e-06, 4.678811e-06, 6.123951e-06, 9.155787e-06,
  1.880775e-06, 8.55124e-07, 1.237759e-06, 1.096991e-06, 1.74514e-06, 
    1.672809e-06, 1.418419e-06, 1.965091e-06, 1.719324e-06, 1.162796e-06, 
    1.255085e-06, 1.467488e-06, 3.044992e-06, 1.065972e-05, 1.909404e-05,
  2.296287e-06, 1.302551e-06, 1.048283e-06, 1.06191e-06, 1.205988e-06, 
    1.694999e-06, 1.324296e-06, 1.360165e-06, 1.037038e-06, 1.330184e-06, 
    2.011427e-06, 2.875208e-06, 1.13714e-05, 1.923616e-05, 2.95045e-05,
  2.107504e-06, 1.649959e-06, 1.34691e-06, 1.178289e-06, 1.032715e-06, 
    9.00887e-07, 1.143581e-06, 1.656884e-06, 2.244901e-06, 2.878844e-06, 
    4.043717e-06, 8.797892e-06, 1.542496e-05, 1.603655e-05, 2.571791e-05,
  1.27435e-06, 1.282485e-06, 1.651105e-06, 1.646959e-06, 1.937599e-06, 
    2.199048e-06, 2.672271e-06, 2.560158e-06, 4.635434e-06, 4.730044e-06, 
    5.851783e-06, 8.669124e-06, 8.035541e-06, 5.070303e-06, 1.533629e-05,
  6.692846e-07, 2.017462e-06, 3.019616e-06, 3.232022e-06, 2.930898e-06, 
    3.520391e-06, 5.369831e-06, 5.572488e-06, 5.058351e-06, 4.734826e-06, 
    4.702213e-06, 4.260044e-06, 4.772141e-06, 4.35391e-06, 6.963547e-06,
  1.288657e-06, 2.806481e-06, 3.913622e-06, 4.589348e-06, 4.66599e-06, 
    5.321777e-06, 5.184055e-06, 5.61846e-06, 4.137079e-06, 3.866529e-06, 
    2.991662e-06, 3.07634e-06, 3.886979e-06, 3.346159e-06, 4.239349e-06,
  2.37637e-06, 4.552565e-06, 4.758449e-06, 4.80635e-06, 5.662797e-06, 
    5.891676e-06, 5.614451e-06, 3.216858e-06, 3.362123e-06, 4.591514e-06, 
    4.08126e-06, 3.668337e-06, 3.394939e-06, 3.30169e-06, 4.64296e-06,
  3.512651e-06, 6.552311e-06, 6.817424e-06, 5.434939e-06, 4.891544e-06, 
    5.646976e-06, 5.81623e-06, 5.340803e-06, 4.466174e-06, 3.17053e-06, 
    3.321942e-06, 4.478035e-06, 3.38678e-06, 3.387491e-06, 4.243263e-06,
  6.659183e-05, 6.011483e-05, 5.235149e-05, 6.659905e-05, 6.696936e-05, 
    7.499553e-05, 9.790781e-05, 9.15639e-05, 7.317279e-05, 4.345334e-05, 
    1.706071e-05, 1.186371e-05, 1.092933e-05, 1.316302e-05, 1.261152e-05,
  0.0001060262, 0.0001091285, 8.385265e-05, 7.358113e-05, 6.703822e-05, 
    8.866273e-05, 7.976013e-05, 7.402878e-05, 6.093626e-05, 3.320701e-05, 
    1.271078e-05, 1.071381e-05, 8.304651e-06, 8.588543e-06, 9.403279e-06,
  0.0001142396, 0.0001110745, 0.0001301591, 9.920587e-05, 0.0001003124, 
    0.0001064, 8.494386e-05, 7.026042e-05, 4.866942e-05, 3.058396e-05, 
    1.433945e-05, 9.494767e-06, 8.648227e-06, 7.117828e-06, 7.243675e-06,
  5.572151e-05, 7.810258e-05, 9.394612e-05, 6.183111e-05, 5.199981e-05, 
    3.855631e-05, 2.636115e-05, 1.546491e-05, 1.832573e-05, 1.513946e-05, 
    1.032027e-05, 1.0821e-05, 1.094641e-05, 1.024708e-05, 5.928271e-06,
  6.267962e-05, 6.769258e-05, 4.792576e-05, 4.497609e-05, 1.74936e-05, 
    4.769436e-06, 6.632464e-06, 9.293812e-06, 1.028229e-05, 8.960492e-06, 
    1.071006e-05, 1.098515e-05, 1.063803e-05, 9.845417e-06, 5.793925e-06,
  1.328818e-05, 9.343126e-06, 8.959044e-06, 2.983782e-06, 3.334301e-06, 
    5.168675e-06, 5.909411e-06, 8.122004e-06, 9.347308e-06, 7.799455e-06, 
    8.972987e-06, 9.024712e-06, 1.165327e-05, 9.143385e-06, 5.40743e-06,
  1.026433e-05, 6.440599e-06, 1.506325e-05, 7.207438e-06, 6.083375e-06, 
    5.761533e-06, 8.023758e-06, 9.29486e-06, 1.059893e-05, 9.95963e-06, 
    7.73371e-06, 8.208379e-06, 1.197843e-05, 7.523374e-06, 6.849463e-06,
  5.082532e-06, 8.077413e-06, 3.912158e-06, 6.596446e-06, 5.990314e-06, 
    7.15615e-06, 9.805712e-06, 1.305796e-05, 1.465269e-05, 1.048033e-05, 
    8.379241e-06, 1.096852e-05, 1.184992e-05, 1.085839e-05, 7.740082e-06,
  2.326373e-06, 3.033892e-06, 3.82903e-06, 5.336981e-06, 7.739225e-06, 
    8.938315e-06, 9.612302e-06, 1.181172e-05, 1.364245e-05, 1.120711e-05, 
    6.821807e-06, 1.021843e-05, 1.130236e-05, 1.11588e-05, 1.1803e-05,
  1.942981e-06, 3.185188e-06, 3.886507e-06, 4.520127e-06, 5.665623e-06, 
    8.449102e-06, 1.084176e-05, 1.303469e-05, 1.391008e-05, 7.468572e-06, 
    6.218726e-06, 7.119905e-06, 1.007079e-05, 1.04987e-05, 9.680723e-06,
  3.088333e-05, 3.554019e-05, 1.936392e-05, 1.018108e-05, 9.313045e-06, 
    7.245832e-06, 9.253274e-06, 2.090832e-05, 3.376552e-05, 6.986693e-05, 
    8.303566e-05, 8.665877e-05, 9.65552e-05, 9.793406e-05, 0.0001145696,
  1.137703e-05, 1.25028e-05, 9.756185e-06, 4.889481e-06, 5.597328e-06, 
    5.661552e-06, 8.661766e-06, 1.967883e-05, 5.010523e-05, 9.01442e-05, 
    8.596885e-05, 0.0001092936, 0.0001151123, 0.0001336684, 0.0001574963,
  1.881476e-05, 1.604664e-05, 1.199041e-05, 8.257574e-06, 5.66855e-06, 
    6.463983e-06, 2.012069e-05, 6.5623e-05, 7.975216e-05, 8.381446e-05, 
    0.0001265524, 0.0001480268, 0.0001610332, 0.00019318, 0.0001972918,
  4.638133e-05, 5.766079e-05, 4.08738e-05, 1.13974e-05, 1.025191e-05, 
    3.805603e-05, 3.897069e-05, 6.891461e-05, 5.601017e-05, 8.281494e-05, 
    0.0001129396, 0.0001906224, 0.0001624433, 0.0001899284, 0.0001823597,
  3.659126e-05, 3.119301e-05, 2.932058e-05, 3.488435e-05, 5.6853e-05, 
    5.449604e-05, 6.199862e-05, 7.287991e-05, 5.198568e-05, 7.41526e-05, 
    7.524608e-05, 9.245108e-05, 0.0001067044, 0.0001260129, 0.0001223176,
  4.954507e-05, 4.579557e-05, 4.741402e-05, 7.215232e-05, 6.441559e-05, 
    4.260816e-05, 4.541224e-05, 8.108108e-05, 4.570607e-05, 4.934649e-05, 
    5.053437e-05, 6.214527e-05, 7.219805e-05, 6.68261e-05, 7.187438e-05,
  9.009875e-05, 0.0001270631, 0.0001277812, 0.0001472246, 0.0001172653, 
    0.0001243948, 0.0001403063, 0.0001677642, 0.000168001, 0.0001763911, 
    0.0001640822, 0.0002104906, 0.0002027157, 0.0001514365, 0.0001584558,
  0.0001870835, 0.000244637, 0.0002544875, 0.0002336223, 0.0002197161, 
    0.0001917849, 0.0001830546, 0.0002082327, 0.0002249261, 0.0002273699, 
    0.0002323459, 0.0002207562, 0.0002142737, 0.0001899626, 0.0001446233,
  0.0002131319, 0.0002140177, 0.000211258, 0.000156361, 0.0001067804, 
    0.0001051222, 8.301043e-05, 0.0001144635, 0.0001185382, 0.0001430837, 
    0.0001357508, 0.0001290517, 0.0001099347, 7.488586e-05, 9.765877e-05,
  0.0001026807, 0.0001062383, 0.0001156799, 9.65587e-05, 8.601666e-05, 
    6.281489e-05, 7.413916e-05, 9.806669e-05, 9.893424e-05, 9.94121e-05, 
    8.165444e-05, 7.268443e-05, 5.893649e-05, 8.207203e-05, 0.0001052061,
  2.137465e-05, 7.85568e-05, 9.235831e-05, 6.825117e-05, 1.389816e-05, 
    6.970904e-06, 3.977975e-06, 8.141375e-06, 6.684371e-06, 7.533398e-06, 
    1.045878e-05, 1.810357e-05, 2.800159e-05, 3.968721e-05, 4.176222e-05,
  1.811987e-05, 3.178258e-05, 0.000133891, 9.441273e-05, 5.480815e-05, 
    1.991441e-05, 8.094861e-06, 6.565547e-06, 7.184404e-06, 6.933755e-06, 
    7.980219e-06, 9.819239e-06, 1.575337e-05, 2.188474e-05, 2.356685e-05,
  2.494455e-05, 1.891387e-05, 5.674197e-05, 0.0001548245, 7.686945e-05, 
    3.198955e-05, 8.572247e-06, 7.110199e-06, 6.541144e-06, 8.177592e-06, 
    7.850223e-06, 1.010253e-05, 9.762431e-06, 1.072672e-05, 1.25378e-05,
  2.197175e-05, 3.738637e-05, 6.786826e-05, 7.450287e-05, 0.0001027645, 
    2.993065e-05, 8.631404e-06, 3.048679e-06, 5.751582e-06, 5.769359e-06, 
    7.359745e-06, 7.38599e-06, 6.770167e-06, 5.319735e-06, 6.317785e-06,
  3.495298e-05, 5.312202e-05, 6.373123e-05, 5.796154e-05, 9.271782e-05, 
    4.970645e-05, 1.775723e-05, 3.283845e-06, 2.263811e-06, 3.014851e-06, 
    3.294612e-06, 2.586347e-06, 3.817627e-06, 4.684085e-06, 5.912877e-06,
  3.557124e-05, 3.683309e-05, 4.037514e-05, 4.653529e-05, 0.0001111732, 
    8.262315e-05, 4.006559e-05, 1.413149e-05, 3.985363e-06, 7.333757e-07, 
    6.560005e-07, 9.39889e-07, 1.478834e-06, 1.126081e-06, 1.173019e-06,
  1.547811e-05, 2.602217e-05, 7.669673e-05, 5.743091e-05, 7.132001e-05, 
    6.750407e-05, 3.748393e-05, 2.091628e-05, 2.447604e-06, 2.446838e-07, 
    4.276734e-09, 4.131939e-09, 5.828744e-08, 1.64427e-07, 2.472833e-07,
  1.119502e-05, 1.130913e-05, 3.548439e-05, 1.444805e-05, 4.824452e-05, 
    3.739087e-05, 4.839001e-05, 2.332643e-05, 9.814024e-06, 5.362953e-06, 
    2.352228e-06, 5.345907e-06, 6.297459e-06, 9.315e-06, 8.060999e-06,
  2.026614e-05, 3.448551e-06, 2.218852e-05, 1.774359e-05, 3.895651e-05, 
    6.433474e-05, 7.905288e-05, 9.064632e-05, 5.0018e-05, 3.488359e-05, 
    4.758753e-05, 4.48049e-05, 5.136342e-05, 3.384416e-05, 2.114015e-05,
  2.590752e-05, 8.053997e-06, 1.649775e-05, 4.150902e-05, 7.854131e-05, 
    0.0001472315, 0.0001281323, 0.0001363192, 8.645462e-05, 9.476531e-05, 
    8.365398e-05, 6.079124e-05, 9.375188e-05, 4.213172e-05, 2.659485e-05,
  6.698273e-06, 6.283563e-06, 5.674419e-06, 5.447232e-06, 7.267131e-06, 
    9.018167e-06, 6.315658e-06, 4.408649e-06, 5.55765e-06, 6.823097e-06, 
    7.449421e-06, 6.487678e-06, 6.605544e-06, 3.131361e-06, 3.017047e-06,
  7.827451e-06, 7.793034e-06, 5.922749e-06, 5.610739e-06, 6.995286e-06, 
    1.203616e-05, 1.109154e-05, 1.640361e-05, 2.010951e-05, 1.670261e-05, 
    5.587804e-06, 3.742952e-07, 3.757485e-09, 9.312352e-08, 3.000625e-07,
  9.578896e-06, 8.267627e-06, 6.632103e-06, 5.105623e-06, 7.612827e-06, 
    7.958967e-06, 9.660512e-06, 1.604595e-05, 1.894816e-05, 1.68999e-05, 
    3.751098e-06, 3.675801e-10, 1.584651e-08, 6.942249e-10, 1.7866e-09,
  6.39572e-06, 8.37001e-06, 7.146662e-06, 5.21616e-06, 5.44158e-06, 
    3.490543e-06, 5.160473e-06, 8.158784e-06, 1.030256e-05, 8.772237e-06, 
    2.435591e-06, 1.778254e-07, 2.112124e-09, 1.035469e-07, 4.800861e-07,
  2.944522e-06, 7.25029e-06, 7.254199e-06, 7.261584e-06, 9.071163e-06, 
    1.047851e-05, 5.845529e-06, 4.421052e-06, 6.23965e-06, 3.878262e-06, 
    2.670964e-06, 1.038738e-06, 4.635853e-07, 1.783588e-06, 7.574015e-06,
  2.26838e-06, 3.458706e-06, 6.581774e-06, 1.015572e-05, 1.307471e-05, 
    1.909287e-05, 4.622192e-06, 3.209464e-06, 2.541551e-06, 2.346996e-06, 
    1.576003e-06, 1.440019e-06, 3.221376e-06, 8.726168e-06, 1.11591e-05,
  8.611506e-07, 2.115705e-06, 5.421416e-06, 1.502855e-05, 1.306843e-05, 
    2.457915e-05, 8.305838e-06, 3.476821e-06, 3.50266e-06, 2.251683e-06, 
    1.880304e-06, 2.785256e-06, 9.809684e-06, 1.102333e-05, 1.115221e-05,
  6.655694e-06, 9.385722e-07, 4.521055e-06, 8.170913e-06, 2.329713e-05, 
    2.482772e-05, 1.376089e-05, 3.141118e-06, 3.229888e-06, 3.399112e-06, 
    4.630135e-06, 1.002583e-05, 1.065377e-05, 1.035341e-05, 3.988264e-06,
  1.201291e-05, 1.155681e-06, 2.967677e-06, 7.607418e-06, 1.882903e-05, 
    1.127859e-05, 2.565762e-06, 3.847952e-06, 9.481407e-06, 5.314771e-06, 
    6.633669e-06, 6.002223e-06, 3.954009e-06, 4.724499e-06, 1.708218e-05,
  2.472844e-05, 8.906916e-07, 1.759634e-06, 5.81864e-06, 1.20566e-05, 
    1.370387e-05, 2.654541e-05, 4.852388e-05, 1.381564e-05, 3.606094e-06, 
    1.010819e-05, 2.613042e-06, 1.349792e-05, 6.110051e-05, 0.0001760343,
  2.965886e-05, 1.658307e-05, 5.507584e-06, 1.998494e-06, 1.21548e-06, 
    1.446204e-06, 6.305599e-07, 2.529531e-07, 9.162923e-07, 8.434773e-07, 
    1.091979e-06, 1.962201e-06, 1.134228e-05, 1.654613e-05, 1.616905e-05,
  2.474439e-05, 1.272329e-05, 2.061489e-06, 3.694257e-09, 6.885137e-07, 
    8.121689e-07, 1.58889e-06, 2.822173e-06, 3.078698e-06, 2.450131e-06, 
    1.481862e-06, 8.62755e-07, 2.482559e-06, 5.866631e-06, 7.030964e-06,
  2.58192e-05, 1.302875e-05, 4.056723e-06, 2.232678e-07, 2.681884e-07, 
    8.440118e-07, 1.44284e-06, 3.237361e-06, 5.67776e-06, 2.343145e-06, 
    2.967752e-07, 2.330106e-08, 1.914565e-06, 5.939822e-06, 5.42338e-06,
  2.435162e-05, 1.709233e-05, 6.462812e-06, 1.404492e-06, 1.614299e-06, 
    1.195612e-06, 1.450372e-06, 2.280283e-06, 1.641773e-06, 9.891817e-07, 
    4.701615e-07, 1.627211e-06, 3.006809e-06, 5.248116e-06, 2.907443e-06,
  1.936839e-05, 1.088594e-05, 7.410723e-06, 3.871745e-06, 8.667683e-07, 
    4.354457e-07, 4.935595e-07, 1.152445e-06, 8.290651e-07, 5.471197e-07, 
    6.002219e-07, 1.746387e-06, 3.221023e-06, 2.759816e-06, 1.607015e-06,
  0.0001030714, 4.033485e-05, 1.398864e-05, 3.054073e-06, 1.711261e-06, 
    9.784493e-07, 9.998882e-07, 5.255243e-07, 5.080333e-07, 6.584413e-07, 
    1.033695e-06, 1.457009e-06, 1.988986e-06, 3.467798e-06, 6.529466e-06,
  0.0005398506, 0.0003342339, 0.0001355509, 3.724404e-05, 6.681892e-06, 
    1.13193e-06, 1.286115e-06, 7.402447e-07, 9.309907e-07, 9.074722e-07, 
    9.381159e-07, 1.258079e-06, 2.792148e-06, 7.158426e-06, 7.407015e-06,
  0.0006087104, 0.0004892935, 0.0002884184, 0.0001187346, 4.37198e-05, 
    8.081742e-06, 1.299264e-06, 2.156544e-06, 1.002354e-06, 1.220752e-06, 
    1.15506e-06, 1.280814e-06, 5.03239e-06, 8.83419e-06, 5.403468e-06,
  0.0005723115, 0.0005048311, 0.0003632208, 0.0001954178, 6.699219e-05, 
    1.373671e-05, 5.467352e-06, 1.146766e-06, 8.945318e-07, 2.880495e-06, 
    2.588865e-06, 3.246016e-06, 6.619649e-06, 4.767478e-06, 6.930603e-06,
  0.000456376, 0.0004924556, 0.0004955758, 0.0003967294, 0.0001919862, 
    4.641209e-05, 1.335775e-05, 1.51728e-05, 1.631524e-05, 1.16347e-06, 
    8.276441e-07, 3.245241e-06, 6.699768e-06, 7.415264e-06, 2.850002e-05,
  3.24814e-05, 1.033542e-05, 4.364882e-06, 5.822862e-07, 3.332524e-08, 
    1.006914e-07, 4.313979e-07, 1.754882e-06, 1.635414e-06, 1.539581e-06, 
    2.050286e-06, 2.623568e-06, 2.000735e-06, 3.734385e-06, 7.9581e-06,
  1.065208e-05, 2.817828e-06, 1.220103e-06, 7.599219e-08, 4.629144e-08, 
    1.197301e-06, 1.594066e-06, 2.023962e-06, 2.181615e-06, 1.305771e-06, 
    6.904488e-07, 2.085644e-07, 4.429457e-07, 2.664463e-06, 2.374228e-06,
  5.970086e-06, 1.470873e-06, 9.228962e-07, 4.677362e-07, 9.159567e-07, 
    2.025088e-06, 2.509498e-06, 2.184597e-06, 2.779663e-06, 1.765242e-06, 
    1.513461e-06, 5.262989e-07, 1.478544e-07, 2.052877e-09, 5.843467e-08,
  3.26309e-06, 5.627379e-07, 8.654767e-07, 8.351841e-07, 1.46479e-06, 
    1.786859e-06, 2.19016e-06, 1.824056e-06, 2.18085e-06, 1.422028e-06, 
    2.244515e-06, 9.104093e-07, 2.463061e-07, 6.225788e-10, 2.642358e-07,
  4.625902e-07, 1.214503e-07, 9.084303e-07, 1.212904e-06, 1.78321e-06, 
    1.691508e-06, 1.935714e-06, 2.06811e-06, 2.717748e-06, 5.002283e-06, 
    3.162614e-06, 1.724791e-06, 2.190524e-09, 1.889435e-08, 4.203265e-07,
  1.822316e-06, 2.209517e-06, 1.41527e-06, 1.868335e-06, 3.243417e-06, 
    2.683625e-06, 1.991488e-06, 3.681364e-06, 4.337665e-06, 4.737421e-06, 
    5.059393e-06, 3.750519e-06, 2.521423e-06, 1.276824e-06, 4.514244e-07,
  7.973469e-05, 8.697424e-05, 2.53239e-05, 1.387007e-05, 1.225971e-05, 
    4.80784e-06, 3.345914e-06, 4.078292e-06, 4.513434e-06, 5.063189e-06, 
    4.766199e-06, 4.877484e-06, 4.667434e-06, 3.755043e-06, 2.886508e-06,
  0.0003371749, 0.0003481358, 0.0001040661, 5.870085e-05, 5.251056e-05, 
    3.478437e-05, 1.107065e-05, 4.747397e-06, 6.96985e-06, 6.479426e-06, 
    6.307345e-06, 6.881199e-06, 6.681154e-06, 4.513245e-06, 5.589397e-06,
  0.0004853968, 0.0003732705, 0.0001308207, 9.239437e-05, 8.158083e-05, 
    7.551e-05, 3.521176e-05, 1.734672e-05, 9.499296e-06, 1.201531e-05, 
    1.133987e-05, 1.176503e-05, 9.128333e-06, 8.409655e-06, 5.576256e-06,
  9.376687e-05, 0.0001128201, 9.982645e-05, 7.855675e-05, 9.171964e-05, 
    0.0001434715, 9.27275e-05, 4.270571e-05, 2.1651e-05, 2.097473e-05, 
    3.001699e-05, 3.249825e-05, 2.491148e-05, 1.854316e-05, 1.448664e-05,
  1.954186e-05, 1.834901e-05, 2.99949e-05, 3.234451e-05, 2.716881e-05, 
    2.965134e-05, 2.917601e-05, 3.277076e-05, 3.074312e-05, 3.839635e-05, 
    4.793592e-05, 4.821784e-05, 6.793118e-05, 6.774255e-05, 3.144603e-05,
  1.248734e-05, 2.091141e-05, 2.647971e-05, 2.116414e-05, 2.653836e-05, 
    3.45315e-05, 4.152818e-05, 2.807992e-05, 3.660083e-05, 4.122091e-05, 
    4.210621e-05, 4.155013e-05, 2.961134e-05, 1.85055e-05, 1.115645e-05,
  5.923421e-06, 1.598019e-05, 1.574308e-05, 1.337891e-05, 1.602521e-05, 
    2.043668e-05, 2.471398e-05, 2.311208e-05, 2.735777e-05, 2.356545e-05, 
    3.162142e-05, 1.777051e-05, 7.671365e-06, 1.170524e-06, 3.742098e-07,
  4.282082e-06, 6.566622e-06, 4.753058e-06, 4.890526e-06, 6.058688e-06, 
    6.603192e-06, 1.024091e-05, 8.954164e-06, 1.204021e-05, 1.413854e-05, 
    9.071006e-06, 6.691543e-06, 3.318298e-06, 1.119989e-06, 2.366265e-07,
  3.241695e-06, 1.39404e-06, 1.093479e-06, 1.218848e-06, 1.131687e-06, 
    2.377499e-06, 3.147973e-06, 4.060002e-06, 5.869929e-06, 6.032039e-06, 
    4.323106e-06, 3.578578e-06, 2.146462e-06, 7.945061e-07, 5.221336e-07,
  3.244847e-07, 3.800506e-07, 4.525303e-07, 5.013521e-07, 8.039983e-07, 
    1.411681e-06, 1.818752e-06, 3.693896e-06, 5.441271e-06, 4.307298e-06, 
    3.304076e-06, 3.399284e-06, 2.09837e-06, 1.039491e-06, 9.541342e-07,
  2.026872e-07, 3.666855e-07, 9.308635e-07, 1.676358e-06, 3.435571e-06, 
    3.424721e-06, 1.206095e-06, 3.061206e-06, 3.833491e-06, 3.448901e-06, 
    2.865337e-06, 1.674764e-06, 8.560013e-07, 1.09333e-06, 2.030267e-06,
  7.113459e-07, 1.049249e-06, 2.958367e-06, 6.821117e-06, 2.324643e-05, 
    9.055897e-06, 3.30403e-06, 2.204463e-06, 4.52333e-06, 4.974173e-06, 
    1.769675e-06, 1.152167e-06, 1.320393e-06, 1.474713e-06, 5.471192e-07,
  1.073906e-06, 2.268065e-06, 4.24861e-06, 1.349082e-05, 2.798331e-05, 
    7.528567e-06, 2.677544e-06, 9.553862e-07, 3.79935e-06, 4.608416e-06, 
    5.866933e-06, 3.929316e-06, 4.106501e-06, 6.376084e-06, 5.645509e-06,
  1.524417e-06, 2.901688e-06, 7.640181e-06, 1.834289e-05, 4.508361e-05, 
    3.519808e-05, 3.414826e-06, 2.724558e-06, 8.55387e-06, 5.524125e-06, 
    9.236785e-06, 7.208151e-06, 8.956253e-06, 1.529959e-05, 2.134021e-05,
  2.991935e-05, 7.414336e-06, 4.485414e-07, 1.395743e-08, 1.670763e-07, 
    2.177807e-06, 5.807944e-06, 5.877347e-06, 6.58501e-06, 8.343545e-06, 
    1.480263e-05, 1.464879e-05, 1.102464e-05, 8.38172e-06, 1.160351e-05,
  5.294867e-05, 2.223527e-05, 7.625946e-06, 4.172334e-06, 1.553862e-06, 
    1.710777e-07, 5.400028e-07, 2.830975e-06, 3.479564e-06, 3.788054e-06, 
    5.315234e-06, 7.534822e-06, 8.568896e-06, 1.84039e-05, 2.383276e-05,
  3.921182e-05, 3.109684e-05, 3.200148e-05, 1.720572e-05, 9.47492e-06, 
    7.623982e-06, 2.486683e-06, 1.881264e-06, 3.587873e-06, 3.768465e-06, 
    7.503238e-06, 1.14437e-05, 1.560881e-05, 1.920669e-05, 1.673703e-05,
  5.300552e-06, 2.12534e-05, 3.359548e-05, 3.867676e-05, 2.843827e-05, 
    2.051178e-05, 1.456314e-05, 9.84194e-06, 9.106479e-06, 8.056086e-06, 
    1.121704e-05, 1.207873e-05, 8.876087e-06, 7.777987e-06, 6.923186e-06,
  6.770136e-08, 9.691456e-07, 6.862544e-06, 2.159698e-05, 2.830181e-05, 
    3.339976e-05, 2.054637e-05, 1.9751e-05, 1.419735e-05, 1.121645e-05, 
    9.081115e-06, 6.29162e-06, 6.755165e-06, 4.941613e-06, 5.822611e-06,
  2.04052e-07, 6.554701e-08, 1.556996e-07, 7.956538e-07, 5.292849e-06, 
    1.714105e-05, 1.782052e-05, 2.438186e-05, 2.280315e-05, 1.362462e-05, 
    1.123524e-05, 8.63467e-06, 9.715242e-06, 7.215516e-06, 7.188013e-06,
  2.153211e-07, 1.974192e-08, 2.10549e-07, 3.756573e-07, 4.330217e-07, 
    5.143449e-07, 5.851457e-06, 1.23323e-05, 1.730206e-05, 2.267085e-05, 
    1.986801e-05, 1.244824e-05, 1.098506e-05, 1.00793e-05, 1.056623e-05,
  6.119105e-07, 5.175596e-07, 2.329743e-06, 6.50352e-07, 6.42125e-07, 
    1.282493e-07, 9.779715e-08, 1.116425e-06, 3.075585e-06, 7.319473e-06, 
    9.440535e-06, 1.055522e-05, 9.100391e-06, 9.217341e-06, 1.24071e-05,
  1.328422e-06, 1.471314e-06, 6.889185e-06, 1.009911e-05, 8.857472e-06, 
    2.493682e-06, 1.478298e-06, 1.451129e-06, 1.204583e-06, 1.513849e-06, 
    2.8215e-06, 3.292231e-06, 5.295531e-06, 3.643608e-06, 4.484171e-06,
  1.568052e-06, 6.312911e-07, 7.697474e-06, 4.359708e-05, 5.435276e-05, 
    2.517954e-05, 6.96753e-06, 1.722675e-06, 1.440957e-06, 3.686703e-06, 
    2.031776e-06, 2.640136e-06, 2.514335e-06, 1.897064e-06, 3.637115e-06,
  1.054004e-05, 1.417565e-06, 2.67174e-09, 4.934028e-08, 1.351304e-06, 
    4.174198e-06, 4.74765e-06, 4.282361e-06, 8.18994e-06, 9.927552e-06, 
    1.435555e-05, 1.72672e-05, 2.873934e-05, 4.32683e-05, 5.114546e-05,
  1.888759e-05, 6.215172e-06, 3.570022e-08, 2.558827e-08, 3.632077e-07, 
    4.046367e-07, 4.036314e-06, 4.549471e-06, 5.501495e-06, 8.363375e-06, 
    1.087514e-05, 1.296241e-05, 1.647648e-05, 2.257646e-05, 2.86092e-05,
  3.06246e-05, 1.114616e-05, 7.048861e-06, 1.691516e-07, 1.766717e-07, 
    2.897859e-07, 1.100433e-06, 2.964425e-06, 3.377143e-06, 5.23921e-06, 
    6.694929e-06, 9.745858e-06, 1.004763e-05, 1.326539e-05, 1.590509e-05,
  1.96962e-05, 1.826579e-05, 1.254793e-05, 5.275933e-06, 5.133581e-08, 
    2.672548e-09, 5.414701e-08, 9.406107e-07, 2.412161e-06, 3.377869e-06, 
    5.433008e-06, 6.918085e-06, 9.605363e-06, 1.051387e-05, 1.134952e-05,
  5.127618e-06, 1.317568e-05, 2.091388e-05, 8.231321e-06, 4.000869e-06, 
    6.409696e-07, 1.070854e-07, 8.313903e-07, 1.393333e-06, 1.930438e-06, 
    2.02527e-06, 4.403451e-06, 6.629975e-06, 8.658372e-06, 9.675062e-06,
  1.570483e-05, 4.467636e-06, 7.499579e-06, 1.573501e-05, 8.350755e-06, 
    5.41437e-06, 3.712662e-06, 1.807878e-06, 3.902348e-06, 3.679946e-06, 
    2.144756e-06, 2.189803e-06, 4.641588e-06, 5.428982e-06, 7.845319e-06,
  3.083428e-05, 1.830565e-05, 1.059929e-05, 6.680546e-06, 5.764346e-06, 
    9.133277e-06, 8.320717e-06, 1.201391e-05, 1.538485e-05, 1.224159e-05, 
    5.981294e-06, 2.22305e-06, 5.058217e-06, 4.602888e-06, 5.202459e-06,
  5.708419e-05, 4.939236e-05, 2.412242e-05, 7.018932e-06, 3.561452e-06, 
    6.733578e-06, 8.995579e-06, 1.449176e-05, 2.333004e-05, 2.579047e-05, 
    2.475942e-05, 2.011201e-05, 1.409978e-05, 5.312988e-06, 4.021127e-06,
  2.610576e-05, 3.594915e-05, 5.719729e-05, 8.64531e-05, 7.3947e-05, 
    1.06881e-05, 8.211849e-06, 9.979506e-06, 1.208803e-05, 1.623018e-05, 
    2.106855e-05, 2.912759e-05, 3.12154e-05, 2.958953e-05, 2.117619e-05,
  7.108491e-06, 2.243699e-05, 6.278018e-05, 0.0003880153, 0.0005016229, 
    0.0001608155, 6.393111e-06, 5.627716e-06, 6.988566e-06, 8.650931e-06, 
    1.094185e-05, 1.931501e-05, 2.924294e-05, 3.856039e-05, 3.99692e-05,
  3.051194e-08, 2.695596e-08, 4.625428e-08, 7.387631e-07, 1.68291e-06, 
    2.644701e-06, 2.913171e-06, 1.368266e-06, 4.864709e-06, 6.836744e-06, 
    1.021961e-05, 1.371472e-05, 2.09361e-05, 3.695006e-05, 4.533499e-05,
  1.344878e-06, 9.732204e-08, 3.422407e-07, 4.750494e-07, 9.945808e-07, 
    2.117696e-06, 1.74199e-06, 9.118607e-07, 3.329113e-06, 6.523623e-06, 
    8.08775e-06, 1.351423e-05, 1.912867e-05, 3.12025e-05, 5.274967e-05,
  9.786351e-07, 2.050635e-06, 3.314892e-07, 1.362009e-06, 1.32305e-06, 
    1.899611e-06, 1.866679e-06, 8.76439e-07, 1.813055e-06, 3.113455e-06, 
    5.852222e-06, 8.302795e-06, 1.466939e-05, 2.537192e-05, 4.464974e-05,
  7.496201e-07, 1.569136e-06, 5.320276e-07, 2.02716e-06, 1.054981e-06, 
    2.200493e-06, 2.597729e-06, 2.281098e-06, 2.36291e-06, 3.056294e-06, 
    4.167414e-06, 6.94954e-06, 1.263717e-05, 2.063601e-05, 2.703337e-05,
  2.113294e-06, 6.484954e-07, 6.012842e-07, 2.785593e-06, 3.092145e-06, 
    1.722702e-06, 3.233186e-06, 2.047905e-06, 4.258897e-06, 3.244767e-06, 
    3.772961e-06, 6.521562e-06, 1.012036e-05, 1.49257e-05, 1.631907e-05,
  4.396346e-06, 3.468102e-06, 1.892458e-06, 5.377831e-06, 4.596816e-06, 
    5.23957e-06, 2.973446e-06, 3.278521e-06, 2.342832e-06, 3.64012e-06, 
    3.698868e-06, 5.080466e-06, 8.255346e-06, 1.069513e-05, 1.16426e-05,
  2.2476e-05, 8.5457e-06, 4.716991e-06, 2.672178e-06, 5.142072e-06, 
    9.904274e-06, 5.728591e-06, 3.298262e-06, 2.938283e-06, 2.457364e-06, 
    3.247648e-06, 4.203082e-06, 7.505673e-06, 7.793621e-06, 8.612617e-06,
  2.470344e-05, 1.580509e-05, 1.133925e-05, 7.566635e-06, 6.50868e-06, 
    9.38945e-06, 7.028391e-06, 4.166237e-06, 2.411693e-06, 1.822158e-06, 
    2.025212e-06, 3.269048e-06, 3.695873e-06, 5.865123e-06, 6.738929e-06,
  3.874613e-05, 2.137231e-05, 1.194264e-05, 1.046302e-05, 1.07416e-05, 
    1.026753e-05, 1.013859e-05, 1.348736e-05, 7.672755e-06, 2.9152e-06, 
    1.527271e-06, 1.062124e-06, 1.666828e-06, 1.928635e-06, 2.569945e-06,
  4.598429e-05, 3.924613e-05, 8.157807e-05, 4.438254e-05, 2.131319e-05, 
    1.851302e-05, 1.295246e-05, 1.442676e-05, 1.170289e-05, 4.10431e-06, 
    2.634666e-06, 3.6888e-06, 1.758487e-06, 1.125966e-06, 2.207196e-06,
  8.178121e-06, 6.455141e-06, 6.686637e-06, 1.124394e-05, 6.557499e-06, 
    4.24083e-06, 4.951817e-06, 3.57131e-06, 2.311023e-06, 2.538515e-06, 
    2.899235e-06, 4.283655e-06, 3.923144e-06, 9.228997e-07, 1.112644e-06,
  1.043087e-05, 9.596091e-06, 1.044947e-05, 7.099688e-06, 4.694173e-06, 
    5.315256e-06, 4.637796e-06, 1.568211e-06, 2.452812e-06, 2.396121e-06, 
    2.341778e-06, 2.251459e-06, 2.695884e-06, 1.996416e-06, 2.555093e-06,
  1.323528e-05, 1.048064e-05, 6.815631e-06, 5.247196e-06, 5.762406e-06, 
    3.841487e-06, 2.549394e-06, 2.342575e-06, 2.216758e-06, 2.611951e-06, 
    2.941389e-06, 4.786838e-06, 4.741065e-06, 6.732766e-06, 6.264432e-06,
  1.072583e-05, 7.758483e-06, 6.250024e-06, 6.437091e-06, 3.94148e-06, 
    3.214299e-06, 2.091906e-06, 3.27057e-06, 3.064161e-06, 3.491654e-06, 
    5.104421e-06, 7.243615e-06, 8.418971e-06, 7.001256e-06, 5.887707e-06,
  7.84472e-06, 7.394515e-06, 6.600851e-06, 5.680014e-06, 3.252513e-06, 
    4.051918e-06, 2.808133e-06, 3.619555e-06, 5.392071e-06, 5.141806e-06, 
    6.612883e-06, 8.206085e-06, 8.821543e-06, 7.010224e-06, 7.549142e-06,
  7.857302e-06, 6.227634e-06, 5.968677e-06, 6.907082e-06, 5.112277e-06, 
    3.014618e-06, 3.601464e-06, 3.906805e-06, 4.943885e-06, 6.234752e-06, 
    7.275079e-06, 7.138618e-06, 7.163136e-06, 5.350834e-06, 4.947392e-06,
  8.313465e-06, 6.73512e-06, 6.460135e-06, 8.438837e-06, 5.130812e-06, 
    4.564139e-06, 3.29726e-06, 3.858494e-06, 4.085196e-06, 5.703986e-06, 
    7.361747e-06, 6.864772e-06, 6.339654e-06, 5.064443e-06, 5.770765e-06,
  7.440652e-06, 8.086419e-06, 6.804261e-06, 7.315402e-06, 7.412516e-06, 
    4.913576e-06, 3.248696e-06, 3.008227e-06, 3.486583e-06, 4.008712e-06, 
    4.758999e-06, 5.427553e-06, 5.196772e-06, 4.983113e-06, 6.657369e-06,
  6.774902e-06, 9.501057e-06, 8.815102e-06, 7.467812e-06, 8.81819e-06, 
    6.122448e-06, 3.359958e-06, 2.155186e-06, 2.58125e-06, 3.097248e-06, 
    3.458348e-06, 3.492014e-06, 4.348447e-06, 5.940541e-06, 1.011766e-05,
  6.17098e-06, 7.428315e-06, 1.002498e-05, 1.092861e-05, 9.466563e-06, 
    9.384807e-06, 4.706022e-06, 2.823069e-06, 1.842608e-06, 2.431313e-06, 
    2.75265e-06, 2.548127e-06, 3.323707e-06, 6.61469e-06, 1.262604e-05,
  1.225746e-05, 1.224344e-05, 8.578392e-06, 5.745578e-06, 5.867439e-06, 
    6.678303e-06, 5.019398e-06, 2.826939e-06, 1.201135e-06, 4.448511e-07, 
    4.467922e-09, 1.245204e-07, 1.466801e-07, 3.001481e-06, 1.851724e-06,
  1.432234e-05, 1.137734e-05, 8.675157e-06, 6.792817e-06, 4.650453e-06, 
    1.822897e-06, 2.816016e-06, 3.443138e-06, 3.906623e-06, 3.9587e-08, 
    4.120859e-08, 1.250248e-07, 7.070205e-08, 4.408857e-07, 3.805746e-06,
  1.388013e-05, 8.689321e-06, 6.08178e-06, 5.412814e-06, 2.741915e-06, 
    1.700214e-06, 2.168436e-06, 2.438912e-06, 1.251534e-06, 2.83133e-08, 
    3.715362e-08, 1.280353e-07, 7.112986e-08, 2.386046e-08, 1.198564e-06,
  1.033115e-05, 6.509872e-06, 2.980042e-06, 3.480548e-06, 2.429831e-06, 
    2.409223e-06, 1.30542e-06, 1.021214e-06, 7.917058e-07, 5.768827e-08, 
    8.516528e-08, 3.010939e-07, 8.645585e-08, 3.203015e-07, 2.408579e-06,
  6.839801e-06, 3.886089e-06, 1.983249e-06, 2.882971e-06, 2.949027e-06, 
    1.877892e-06, 1.394952e-06, 1.737736e-06, 4.607077e-06, 1.855985e-06, 
    1.576185e-07, 2.011569e-07, 6.877478e-07, 1.755511e-06, 2.029971e-06,
  4.435944e-06, 2.693536e-06, 2.172755e-06, 1.837469e-06, 1.893482e-06, 
    2.215388e-06, 2.003855e-06, 2.499522e-06, 3.03778e-06, 1.602445e-06, 
    2.037768e-07, 7.958181e-07, 8.673916e-07, 1.383875e-06, 1.822987e-06,
  4.00527e-06, 3.393484e-06, 2.697539e-06, 1.469621e-06, 2.175486e-06, 
    2.628148e-06, 3.290255e-06, 2.581507e-06, 3.363253e-06, 1.362148e-07, 
    1.99991e-06, 1.044935e-06, 1.252725e-06, 1.736557e-06, 3.878421e-06,
  3.943464e-06, 5.671856e-06, 3.340263e-06, 1.99592e-06, 1.716625e-06, 
    3.651758e-06, 5.223916e-06, 3.114426e-06, 2.03304e-06, 3.220074e-06, 
    2.60221e-06, 3.338659e-06, 2.342293e-06, 3.98254e-06, 1.301038e-05,
  2.884764e-06, 5.021619e-06, 4.350677e-06, 3.043034e-06, 2.732055e-06, 
    3.818432e-06, 3.640712e-06, 3.718401e-06, 1.593632e-06, 2.111225e-06, 
    2.365509e-06, 3.19259e-06, 3.502796e-06, 5.751296e-06, 1.440523e-05,
  2.684993e-06, 5.918906e-06, 6.523328e-06, 5.514333e-06, 3.363099e-06, 
    3.408031e-06, 3.675192e-06, 3.332208e-06, 2.882713e-06, 2.732236e-06, 
    2.193281e-06, 3.00668e-06, 3.766294e-06, 7.238814e-06, 1.222728e-05,
  1.565615e-05, 8.103431e-06, 1.543501e-06, 1.863775e-08, 3.948541e-07, 
    3.683999e-06, 2.107791e-06, 3.28046e-07, 4.04992e-06, 4.368209e-06, 
    6.451497e-06, 7.358624e-06, 4.13577e-06, 4.599531e-06, 1.135943e-05,
  5.753457e-06, 3.961604e-06, 1.566657e-07, 1.521668e-08, 6.458521e-07, 
    1.357037e-06, 1.333395e-06, 4.581963e-07, 2.226506e-06, 4.597898e-06, 
    5.037174e-06, 6.317924e-06, 4.497274e-06, 3.91362e-06, 6.154298e-06,
  3.928898e-06, 1.519588e-06, 2.378646e-08, 3.296239e-08, 2.270131e-07, 
    5.025069e-07, 1.002367e-06, 9.789611e-07, 3.23593e-06, 5.949596e-06, 
    6.294368e-06, 6.061328e-06, 5.967404e-06, 2.738539e-06, 4.074177e-06,
  5.662464e-06, 1.60025e-06, 4.582807e-10, 8.721547e-09, 8.410265e-08, 
    4.210437e-07, 3.737185e-07, 2.624894e-06, 4.924285e-06, 3.40478e-06, 
    5.209629e-06, 8.463164e-06, 7.823975e-06, 6.155003e-06, 3.555907e-06,
  3.473243e-06, 5.551429e-07, 7.834496e-10, 1.480176e-09, 5.362556e-07, 
    4.97674e-07, 8.501591e-08, 1.572831e-06, 4.176588e-06, 4.901743e-06, 
    4.434737e-06, 4.797544e-06, 5.604431e-06, 6.014142e-06, 6.787197e-06,
  9.24447e-07, 5.636701e-07, 7.688874e-10, 7.349603e-10, 9.344685e-07, 
    5.393631e-07, 3.633842e-07, 2.093688e-06, 4.443627e-06, 2.962051e-06, 
    4.136275e-06, 5.699557e-06, 6.017831e-06, 5.724308e-06, 6.459923e-06,
  2.245734e-06, 7.716155e-07, 4.904479e-09, 8.860081e-08, 9.876735e-07, 
    1.419362e-06, 9.087865e-07, 1.85075e-06, 5.47635e-06, 4.482551e-06, 
    3.384495e-06, 4.019209e-06, 5.588779e-06, 5.562736e-06, 6.796767e-06,
  4.958643e-06, 1.454524e-06, 8.145684e-08, 3.65376e-07, 2.211804e-07, 
    7.4361e-07, 1.995721e-07, 2.282265e-06, 2.225641e-06, 3.782466e-06, 
    3.135436e-06, 3.761562e-06, 5.420997e-06, 7.438263e-06, 8.667898e-06,
  3.325131e-06, 2.530759e-06, 9.524989e-07, 6.03409e-07, 6.470488e-07, 
    1.127903e-06, 1.417316e-06, 1.773214e-06, 1.750421e-06, 2.115487e-06, 
    2.837461e-06, 5.157038e-06, 5.412861e-06, 1.106596e-05, 1.242896e-05,
  2.077065e-06, 3.097573e-06, 2.594124e-06, 7.266827e-07, 8.901803e-07, 
    2.330575e-06, 1.322095e-06, 1.920256e-06, 3.174985e-06, 4.081983e-06, 
    4.351883e-06, 6.005451e-06, 1.183992e-05, 1.618911e-05, 1.77566e-05,
  8.033833e-05, 9.56374e-05, 0.0001196529, 0.000131407, 0.0002132076, 
    0.0002950355, 0.0003068079, 0.0001782471, 0.0001645228, 0.0001413691, 
    0.0001023765, 6.351052e-05, 1.745658e-05, 4.25047e-06, 9.202375e-06,
  5.254405e-05, 5.886894e-05, 4.948619e-05, 0.0001064727, 9.536115e-05, 
    0.000114664, 0.000305422, 9.317943e-05, 0.0002318255, 0.0001579389, 
    6.924842e-05, 3.664771e-05, 7.080682e-06, 6.994077e-06, 7.602677e-06,
  3.932441e-05, 4.147461e-05, 5.779669e-05, 5.644633e-05, 0.0001007351, 
    6.8464e-05, 0.0001304928, 0.0001439036, 7.622151e-05, 4.199177e-05, 
    2.169817e-05, 5.299187e-06, 5.001313e-06, 6.351719e-06, 4.38186e-06,
  1.274403e-05, 3.930456e-05, 2.737573e-05, 3.050718e-05, 6.766121e-05, 
    2.785556e-05, 8.946892e-05, 5.079324e-05, 1.052979e-05, 6.793422e-06, 
    4.90412e-06, 4.377182e-06, 4.674598e-06, 6.587342e-06, 4.660979e-06,
  8.223248e-06, 2.597613e-05, 2.440601e-05, 2.135048e-05, 1.729204e-05, 
    1.970762e-05, 2.510776e-05, 2.561501e-05, 7.893078e-06, 2.80341e-06, 
    5.012247e-06, 6.898157e-06, 6.875542e-06, 7.116658e-06, 5.817444e-06,
  4.815063e-06, 1.656843e-05, 1.609228e-05, 3.030555e-05, 1.749587e-05, 
    9.016537e-06, 2.066049e-05, 1.544235e-05, 3.00326e-06, 3.308876e-06, 
    6.08436e-06, 7.631076e-06, 7.575745e-06, 5.398313e-06, 4.869624e-06,
  4.125135e-06, 8.807367e-06, 1.627593e-05, 1.347692e-05, 1.548883e-05, 
    2.061913e-05, 1.1665e-05, 2.41817e-06, 2.843178e-06, 2.423653e-06, 
    4.88848e-06, 4.907625e-06, 5.280895e-06, 4.916096e-06, 4.588157e-06,
  4.264177e-06, 5.413212e-06, 1.140179e-05, 5.560724e-06, 6.516184e-06, 
    2.991579e-06, 2.584587e-06, 5.137176e-06, 3.610429e-06, 1.936007e-06, 
    3.182764e-06, 5.359572e-06, 2.914456e-06, 2.477906e-06, 4.62625e-06,
  8.402439e-06, 7.241718e-06, 5.739892e-06, 3.220545e-06, 2.069777e-06, 
    2.442603e-06, 4.728059e-07, 4.684792e-06, 3.904989e-06, 2.439845e-06, 
    2.364707e-06, 3.226782e-06, 1.366257e-06, 2.107212e-06, 5.211596e-06,
  1.298577e-05, 1.020813e-05, 4.763418e-06, 1.943669e-06, 1.970419e-06, 
    4.428238e-07, 7.36893e-07, 5.961633e-06, 2.635937e-06, 3.175041e-06, 
    1.081807e-06, 2.633721e-06, 2.594267e-06, 3.266945e-06, 5.402482e-06,
  8.089763e-06, 3.054408e-05, 1.513902e-05, 3.852674e-05, 4.0193e-05, 
    2.641949e-05, 2.314521e-05, 1.728534e-05, 1.819902e-05, 1.690689e-05, 
    7.56925e-05, 8.138735e-05, 0.0001248784, 0.0001263181, 0.000106314,
  8.484631e-06, 1.518904e-05, 2.434048e-05, 1.62659e-05, 3.30369e-05, 
    3.363437e-05, 2.483101e-05, 1.62809e-05, 1.564667e-05, 3.090213e-05, 
    7.273803e-05, 0.0001352322, 0.0001669004, 0.0001165879, 0.0001068817,
  1.529277e-06, 5.195569e-06, 1.310254e-05, 1.592976e-05, 1.597642e-05, 
    2.947604e-05, 4.687754e-05, 3.612145e-05, 4.20819e-05, 0.0001100013, 
    0.0001474437, 0.0001475373, 0.0001298221, 0.0001694942, 8.014531e-05,
  1.050774e-05, 9.054171e-06, 1.721568e-05, 6.677684e-06, 1.614517e-05, 
    3.2837e-05, 2.133395e-05, 4.478149e-05, 3.343136e-05, 5.060532e-05, 
    4.226698e-05, 5.898873e-05, 0.0001402447, 0.0001255631, 0.0001669573,
  1.200371e-05, 7.570042e-06, 1.396773e-05, 1.183588e-05, 5.9346e-05, 
    4.399737e-05, 4.659108e-05, 6.346731e-05, 5.472391e-05, 5.574762e-05, 
    6.213222e-05, 3.800975e-05, 0.0001327578, 0.0001478118, 0.0001214135,
  4.753813e-06, 2.032723e-05, 1.849447e-05, 1.594804e-05, 2.99003e-05, 
    5.164603e-05, 5.235123e-05, 8.776333e-05, 8.260876e-05, 7.392492e-05, 
    5.957923e-05, 8.941202e-05, 8.253135e-05, 0.0001202476, 0.0001364567,
  4.195344e-06, 1.334521e-05, 3.650442e-05, 3.542451e-05, 4.345751e-05, 
    4.647571e-05, 7.205638e-05, 6.408219e-05, 7.186909e-05, 7.039292e-05, 
    5.549291e-05, 4.553326e-05, 0.0001030117, 9.106101e-05, 0.0001437389,
  1.769049e-05, 1.997743e-05, 4.700093e-05, 4.980569e-05, 4.758843e-05, 
    4.856255e-05, 5.657701e-05, 7.037872e-05, 6.070484e-05, 7.252247e-05, 
    8.066971e-05, 7.036529e-05, 6.64123e-05, 7.494951e-05, 7.664986e-05,
  1.562504e-05, 1.888323e-05, 2.796341e-05, 3.758099e-05, 5.041071e-05, 
    5.806354e-05, 4.709406e-05, 6.820667e-05, 8.185613e-05, 6.654819e-05, 
    7.660051e-05, 6.301275e-05, 7.715073e-05, 5.666975e-05, 8.586507e-05,
  3.431606e-06, 1.954339e-05, 2.921253e-05, 5.684984e-05, 6.753771e-05, 
    4.170705e-05, 0.0001024459, 9.790708e-05, 7.393851e-05, 9.196825e-05, 
    8.87796e-05, 9.565872e-05, 5.790201e-05, 6.3491e-05, 6.298738e-05,
  4.896127e-06, 1.523951e-05, 1.562947e-05, 2.33239e-05, 3.662488e-05, 
    4.662043e-05, 5.024555e-05, 6.221029e-05, 9.541935e-05, 0.0001509944, 
    0.0001393841, 0.0001357743, 0.0001865682, 0.000195104, 0.00020458,
  1.869244e-06, 9.070917e-06, 9.508432e-06, 1.510391e-05, 2.03031e-05, 
    3.540405e-05, 4.898285e-05, 4.840364e-05, 6.394964e-05, 7.405031e-05, 
    8.624131e-05, 8.603297e-05, 9.921425e-05, 9.745279e-05, 0.0001072955,
  1.28698e-07, 1.835388e-06, 5.777504e-06, 9.738926e-06, 1.400859e-05, 
    2.019487e-05, 3.047119e-05, 4.07677e-05, 5.727879e-05, 6.515766e-05, 
    7.053341e-05, 7.045939e-05, 8.634608e-05, 7.346013e-05, 6.90103e-05,
  8.795428e-08, 1.020276e-07, 5.883632e-07, 2.674195e-06, 7.66181e-06, 
    9.3862e-06, 1.373734e-05, 2.306349e-05, 3.503534e-05, 4.456178e-05, 
    5.431947e-05, 5.722659e-05, 6.040143e-05, 5.391142e-05, 4.136371e-05,
  4.804874e-08, 7.113886e-07, 8.901829e-08, 4.137715e-07, 5.606793e-07, 
    2.324754e-06, 8.860679e-06, 8.570752e-06, 1.248179e-05, 2.012547e-05, 
    2.064807e-05, 2.422703e-05, 2.285586e-05, 1.953632e-05, 1.736032e-05,
  6.797502e-07, 3.447889e-07, 1.582229e-07, 1.300048e-07, 1.408869e-07, 
    3.88774e-07, 7.339892e-07, 1.756898e-06, 6.655075e-06, 6.406351e-06, 
    7.331755e-06, 8.626362e-06, 7.771616e-06, 6.632612e-06, 8.368836e-06,
  1.861476e-06, 3.187091e-07, 2.270623e-07, 7.208702e-07, 1.565631e-06, 
    1.115308e-06, 9.215465e-07, 2.438899e-06, 2.189251e-06, 2.944625e-06, 
    4.515231e-06, 6.617687e-06, 6.448789e-06, 6.254083e-06, 7.565731e-06,
  1.967065e-05, 3.135459e-06, 7.156927e-08, 1.41075e-07, 5.751888e-07, 
    8.509833e-07, 2.4224e-06, 2.248993e-06, 1.230046e-06, 1.51489e-06, 
    3.680479e-06, 3.928439e-06, 5.059576e-06, 4.087286e-06, 4.521809e-06,
  4.407235e-05, 2.116885e-05, 8.205041e-07, 7.709413e-08, 4.145409e-07, 
    6.509667e-07, 1.775243e-06, 2.176493e-06, 1.626273e-06, 9.339489e-07, 
    1.154893e-06, 1.812325e-06, 1.592241e-06, 2.885113e-06, 1.614247e-06,
  4.343315e-05, 4.91485e-05, 5.690157e-06, 1.694477e-06, 6.415189e-07, 
    1.957475e-06, 6.956795e-07, 7.439342e-07, 1.632917e-06, 1.810645e-06, 
    1.197262e-06, 1.546079e-06, 2.502529e-06, 2.627486e-06, 3.131436e-06,
  9.829049e-06, 7.173458e-06, 1.02725e-05, 4.302713e-06, 4.463039e-06, 
    5.859009e-06, 7.658352e-06, 8.597473e-06, 1.233013e-05, 2.81197e-05, 
    3.983542e-05, 6.920304e-05, 8.691116e-05, 0.0001123235, 9.891562e-05,
  1.278707e-05, 9.598552e-06, 6.520321e-06, 9.364585e-06, 5.55638e-06, 
    5.0016e-06, 4.913967e-06, 4.227562e-06, 4.306838e-06, 5.868634e-06, 
    1.139746e-05, 2.86595e-05, 3.842387e-05, 4.553243e-05, 4.770657e-05,
  1.789723e-05, 1.035531e-05, 6.693243e-06, 4.005273e-06, 2.655585e-06, 
    3.43034e-06, 3.46143e-06, 3.662098e-06, 3.055916e-06, 4.540711e-06, 
    5.856116e-06, 1.147463e-05, 1.538103e-05, 2.156868e-05, 2.840569e-05,
  1.277554e-05, 1.391763e-05, 1.083232e-05, 1.002819e-05, 7.078054e-07, 
    3.072907e-06, 4.791488e-06, 6.512503e-06, 5.333856e-06, 4.307195e-06, 
    5.299956e-06, 6.864732e-06, 1.04909e-05, 1.722495e-05, 2.940175e-05,
  1.64712e-05, 1.818127e-05, 1.863749e-05, 1.296112e-05, 4.387606e-06, 
    1.668814e-06, 3.148683e-06, 4.31645e-06, 5.117359e-06, 7.332972e-06, 
    6.307757e-06, 9.359284e-06, 1.299988e-05, 1.939317e-05, 2.760578e-05,
  2.517099e-05, 2.112907e-05, 1.718418e-05, 1.785405e-05, 6.840308e-06, 
    9.392252e-07, 8.447761e-07, 2.211658e-06, 2.944252e-06, 4.137236e-06, 
    6.393259e-06, 9.845746e-06, 1.236466e-05, 1.348885e-05, 1.72078e-05,
  3.824101e-05, 2.985055e-05, 3.674016e-05, 3.063183e-05, 1.17733e-05, 
    2.167721e-06, 1.169018e-06, 1.379588e-06, 2.102641e-06, 2.493588e-06, 
    4.750897e-06, 5.027266e-06, 5.373232e-06, 9.860028e-06, 1.227086e-05,
  2.928329e-05, 4.296169e-05, 5.009872e-05, 6.236912e-05, 2.574732e-05, 
    1.635802e-05, 2.64511e-06, 2.466596e-06, 1.59104e-06, 1.562491e-06, 
    1.596318e-06, 2.503038e-06, 4.313461e-06, 4.559351e-06, 4.657531e-06,
  3.398126e-05, 5.051132e-05, 6.790014e-05, 4.315145e-05, 2.863222e-05, 
    1.44485e-05, 2.874161e-06, 8.668423e-07, 9.567123e-07, 7.150939e-07, 
    8.972069e-07, 6.880736e-07, 2.789319e-06, 4.38357e-06, 2.417846e-06,
  1.278764e-05, 2.912837e-05, 4.448681e-05, 6.195992e-05, 6.433563e-05, 
    2.641222e-05, 1.204826e-05, 4.517831e-06, 3.165655e-06, 1.55909e-06, 
    1.402626e-06, 1.795018e-06, 2.216546e-06, 2.762123e-06, 2.916152e-06,
  2.185269e-05, 3.012425e-05, 3.899757e-05, 3.244408e-05, 7.405132e-05, 
    8.673834e-05, 0.0001112113, 8.551678e-05, 0.0001303446, 0.0001042686, 
    7.625662e-05, 3.901605e-05, 3.703705e-05, 7.327892e-05, 0.0001255573,
  2.245494e-05, 1.396504e-05, 2.811683e-05, 3.849005e-05, 6.340277e-05, 
    9.327864e-05, 7.842821e-05, 8.708845e-05, 7.522028e-05, 6.686485e-05, 
    4.720683e-05, 2.612391e-05, 2.044991e-05, 3.139854e-05, 3.31611e-05,
  9.449717e-06, 1.199233e-05, 1.478225e-05, 1.492874e-05, 3.31947e-05, 
    4.478849e-05, 1.506225e-05, 5.321269e-05, 4.81517e-05, 6.195383e-05, 
    8.453651e-06, 2.177422e-05, 3.593971e-05, 2.756687e-06, 3.838532e-06,
  1.066963e-05, 8.007087e-06, 9.977049e-06, 1.209756e-05, 1.543824e-05, 
    1.127807e-05, 1.35192e-05, 1.284742e-05, 3.056371e-05, 1.475671e-05, 
    1.977666e-06, 1.517865e-06, 1.519815e-06, 2.443419e-06, 1.119398e-05,
  7.135384e-06, 1.283155e-05, 1.552539e-05, 8.430788e-06, 7.969756e-06, 
    9.836798e-06, 1.12761e-05, 1.185896e-05, 1.028396e-06, 1.038977e-06, 
    9.419292e-07, 1.087533e-06, 1.37671e-06, 6.946279e-07, 1.300969e-06,
  8.018897e-06, 7.956868e-06, 1.175334e-05, 1.127195e-05, 9.268362e-06, 
    1.274786e-05, 1.061578e-05, 2.362377e-05, 5.700158e-06, 3.325703e-06, 
    2.843947e-06, 1.273033e-05, 9.269547e-06, 8.398388e-07, 1.161125e-06,
  7.260294e-06, 1.287346e-05, 5.244062e-06, 7.12744e-06, 2.558869e-05, 
    2.906482e-05, 2.185196e-05, 2.167275e-05, 1.666684e-05, 1.336236e-05, 
    1.000056e-05, 8.263431e-06, 1.599165e-05, 5.599408e-06, 7.445165e-06,
  9.205727e-06, 8.418494e-06, 9.447005e-06, 9.222465e-06, 2.150868e-05, 
    3.390352e-05, 2.633526e-05, 2.593696e-05, 1.64355e-05, 9.858627e-06, 
    1.67213e-05, 1.644745e-05, 9.913014e-06, 2.228979e-06, 8.454413e-06,
  7.034303e-06, 1.324241e-05, 1.600278e-05, 1.227531e-05, 1.689997e-05, 
    2.053572e-05, 3.457469e-05, 2.366005e-05, 2.544184e-05, 2.39389e-05, 
    2.236074e-05, 2.771132e-05, 1.63688e-05, 2.414649e-05, 6.06189e-06,
  5.541866e-06, 1.265486e-05, 2.418732e-05, 2.259597e-05, 3.616893e-05, 
    3.009817e-05, 3.016064e-05, 3.473171e-05, 2.493363e-05, 3.183183e-05, 
    3.198479e-05, 3.498017e-05, 3.399578e-05, 5.16016e-05, 2.927798e-05,
  2.956217e-06, 2.832548e-06, 3.197896e-06, 3.202902e-06, 2.677439e-06, 
    2.380737e-06, 2.684573e-06, 3.455475e-06, 2.72906e-06, 1.443471e-05, 
    5.076131e-05, 7.541844e-05, 6.577707e-05, 8.337011e-05, 0.0001113745,
  2.807171e-06, 2.637015e-06, 3.634581e-06, 2.552287e-06, 2.320287e-06, 
    2.631488e-06, 2.759919e-06, 3.032095e-06, 1.434911e-05, 4.303771e-05, 
    5.765626e-05, 3.762784e-05, 3.914407e-05, 0.0001119801, 0.0001115027,
  2.424443e-06, 1.996048e-06, 2.673962e-06, 2.632497e-06, 2.13532e-06, 
    1.980947e-06, 3.893097e-06, 1.413299e-05, 1.624984e-05, 4.042223e-05, 
    5.018929e-05, 1.98747e-05, 7.207519e-05, 3.417208e-05, 8.294442e-05,
  2.461652e-06, 2.415293e-06, 1.222857e-06, 1.512798e-06, 2.792232e-06, 
    3.694022e-06, 1.245548e-05, 3.641858e-06, 2.404065e-05, 3.997843e-05, 
    3.236935e-05, 2.055492e-05, 6.479578e-05, 3.065402e-05, 7.314431e-05,
  2.270692e-06, 2.036822e-06, 3.015546e-06, 7.591375e-06, 1.031767e-05, 
    7.846668e-06, 5.70952e-06, 2.483848e-05, 2.289002e-05, 2.987104e-05, 
    1.024587e-05, 1.468283e-05, 1.417334e-05, 1.463992e-05, 5.4933e-05,
  3.104131e-06, 4.469939e-06, 1.207771e-05, 1.210433e-05, 1.445492e-05, 
    1.503229e-05, 2.017277e-05, 2.146851e-05, 2.18432e-05, 1.814848e-05, 
    1.717387e-05, 1.402091e-05, 2.637033e-05, 1.170288e-05, 1.929639e-05,
  3.528751e-06, 5.786589e-06, 8.902693e-06, 9.870863e-06, 1.144372e-05, 
    1.175937e-05, 1.429071e-05, 2.192918e-05, 2.765937e-05, 1.850345e-05, 
    2.137653e-05, 1.564775e-05, 2.048653e-05, 1.175623e-05, 5.22569e-06,
  3.282127e-06, 5.531699e-06, 9.662244e-06, 1.051379e-05, 1.377497e-05, 
    1.211127e-05, 1.06973e-05, 1.596712e-05, 9.684006e-06, 1.44994e-05, 
    2.096997e-05, 1.112616e-05, 1.401905e-05, 2.078352e-05, 4.69011e-06,
  2.140459e-06, 3.272639e-06, 6.009765e-06, 8.978017e-06, 1.312942e-05, 
    1.122255e-05, 1.210285e-05, 1.130738e-05, 1.381967e-05, 1.003886e-05, 
    2.275193e-05, 1.682451e-05, 2.24608e-05, 2.941249e-05, 2.041741e-05,
  3.888519e-06, 4.49645e-06, 7.35117e-06, 1.174117e-05, 1.847147e-05, 
    1.938452e-05, 2.180035e-05, 2.222262e-05, 2.246792e-05, 1.612441e-05, 
    2.556221e-05, 1.244424e-05, 1.943759e-05, 2.525778e-05, 3.021155e-05,
  7.475697e-06, 1.428338e-05, 1.654768e-05, 1.044808e-05, 4.943657e-06, 
    2.388915e-06, 3.425301e-06, 7.955913e-06, 7.49473e-06, 1.474558e-05, 
    2.021528e-05, 1.942483e-05, 1.752667e-05, 1.742511e-05, 1.698477e-05,
  8.174724e-06, 1.031556e-05, 1.587231e-05, 1.108216e-05, 2.486177e-06, 
    1.999958e-06, 3.199325e-06, 5.727809e-06, 6.445163e-06, 6.618495e-06, 
    1.004222e-05, 1.407541e-05, 1.323118e-05, 1.247163e-05, 1.366445e-05,
  1.66731e-06, 7.88189e-06, 1.481367e-05, 1.30246e-05, 3.333117e-06, 
    2.309118e-07, 3.609406e-06, 5.738028e-06, 2.235896e-06, 3.522817e-06, 
    7.786953e-06, 7.386778e-06, 9.175181e-06, 1.00677e-05, 1.149689e-05,
  2.930517e-07, 6.816308e-06, 1.242813e-05, 1.160405e-05, 4.070442e-06, 
    4.610477e-07, 4.737808e-06, 5.097674e-06, 4.721951e-06, 4.26098e-06, 
    4.245205e-06, 4.587092e-06, 4.076752e-06, 5.983098e-06, 7.699136e-06,
  1.290644e-07, 1.517466e-06, 9.314465e-06, 1.488709e-05, 6.752914e-06, 
    4.099002e-06, 4.010833e-06, 5.042628e-06, 5.180897e-06, 2.929917e-06, 
    2.553104e-06, 1.611541e-06, 5.325887e-07, 4.357312e-06, 3.755684e-06,
  1.455445e-08, 4.936239e-07, 4.965336e-06, 1.26318e-05, 1.368173e-05, 
    6.523438e-06, 4.811779e-06, 7.005008e-06, 4.648974e-06, 4.414629e-06, 
    2.952728e-06, 1.973714e-06, 2.675723e-06, 1.637797e-06, 3.786088e-07,
  3.870531e-08, 3.97292e-07, 2.158728e-06, 5.460701e-06, 1.277718e-05, 
    1.280395e-05, 7.787699e-06, 5.309871e-06, 7.314251e-06, 5.636316e-06, 
    5.159164e-06, 5.848035e-06, 2.528142e-06, 2.889408e-06, 2.73035e-06,
  2.32753e-10, 7.587336e-07, 1.624266e-06, 4.086525e-06, 8.35711e-06, 
    1.306145e-05, 8.51496e-06, 7.309629e-06, 1.011247e-05, 8.289532e-06, 
    9.130631e-06, 5.545428e-06, 4.036168e-06, 2.066581e-06, 2.4823e-06,
  7.851741e-10, 8.569498e-07, 2.833565e-06, 4.285607e-06, 1.355198e-05, 
    1.327806e-05, 8.189384e-06, 4.273501e-06, 5.242451e-06, 6.477902e-06, 
    7.298376e-06, 6.791178e-06, 5.275534e-06, 3.455419e-06, 2.618917e-06,
  7.330725e-08, 1.120461e-06, 5.54343e-06, 1.118922e-05, 2.450315e-05, 
    2.239856e-05, 2.051996e-05, 1.656928e-05, 6.835985e-06, 5.227696e-06, 
    4.817572e-06, 5.795554e-06, 8.101633e-06, 4.630745e-06, 2.953248e-06,
  7.05071e-05, 8.231054e-05, 7.848538e-05, 6.231508e-05, 2.489064e-05, 
    2.071834e-05, 9.479182e-06, 9.537096e-06, 7.481636e-06, 1.301243e-05, 
    2.008105e-05, 1.911263e-05, 1.189175e-05, 1.047844e-05, 1.345204e-05,
  6.898233e-05, 6.381347e-05, 8.533394e-05, 7.434322e-05, 3.646713e-05, 
    2.148727e-05, 1.562137e-05, 7.613281e-06, 6.339558e-06, 8.48181e-06, 
    1.071533e-05, 1.793519e-05, 2.101718e-05, 1.471731e-05, 6.1633e-06,
  5.979548e-05, 7.828829e-05, 3.536595e-05, 3.732532e-05, 3.446002e-05, 
    1.058025e-05, 8.378159e-06, 7.283918e-06, 9.191366e-06, 9.725732e-06, 
    6.735903e-06, 9.076969e-06, 1.474555e-05, 1.725713e-05, 1.076044e-05,
  5.604926e-05, 4.735838e-05, 1.275168e-05, 2.845205e-05, 3.532132e-05, 
    9.261299e-06, 6.461857e-06, 8.537787e-06, 6.730837e-06, 5.885002e-06, 
    4.206122e-06, 6.964053e-06, 6.660857e-06, 1.229188e-05, 1.50769e-05,
  2.376387e-05, 1.490296e-05, 1.447754e-06, 1.851218e-05, 2.483056e-05, 
    1.69737e-05, 1.288983e-05, 2.332276e-05, 1.851726e-05, 9.802551e-06, 
    5.332794e-06, 2.689997e-06, 3.967234e-06, 4.4007e-06, 8.552949e-06,
  5.392671e-05, 4.521933e-05, 7.527965e-07, 1.630217e-05, 2.727236e-05, 
    2.312133e-05, 6.340538e-05, 6.197774e-05, 4.377492e-05, 8.927873e-06, 
    5.648e-06, 2.393055e-06, 3.962721e-06, 3.104554e-06, 2.492155e-06,
  0.0001034831, 5.558715e-05, 9.966438e-06, 1.333505e-05, 3.986251e-05, 
    5.808296e-05, 0.0001554178, 0.0001988176, 8.445225e-05, 4.675779e-06, 
    5.657334e-06, 5.062196e-06, 4.714222e-06, 4.360102e-06, 4.382449e-06,
  0.0001665026, 4.051594e-05, 2.638016e-05, 3.897167e-06, 3.821474e-05, 
    0.000132491, 0.0003346043, 0.0002994705, 7.456679e-05, 3.238757e-06, 
    5.719761e-06, 6.831326e-06, 7.551569e-06, 8.138566e-06, 5.801019e-06,
  0.0002192805, 4.716195e-05, 5.02535e-07, 2.236947e-06, 5.011037e-05, 
    0.0001733949, 0.0002003048, 0.0002508091, 4.174048e-05, 6.05653e-06, 
    3.156295e-06, 6.681965e-06, 8.674919e-06, 1.181116e-05, 1.188642e-05,
  7.042636e-05, 4.692257e-06, 4.162278e-07, 8.715107e-06, 6.20954e-05, 
    0.000116913, 0.0001226704, 0.0001089838, 5.167871e-05, 8.107873e-06, 
    4.807139e-07, 2.601733e-06, 6.35359e-06, 8.835446e-06, 7.822268e-06,
  1.062366e-05, 1.962816e-05, 3.206205e-05, 0.0001875991, 0.0001951853, 
    0.0001288452, 0.0001052202, 9.634814e-05, 0.0001219805, 0.0001586655, 
    0.0001258718, 8.171752e-05, 4.778558e-05, 3.57178e-05, 1.75574e-05,
  6.710903e-06, 1.279041e-05, 2.953814e-05, 0.0001897028, 0.0001875647, 
    0.0001266878, 9.307206e-05, 0.0001687983, 0.0001400429, 0.0001697335, 
    9.505416e-05, 0.0001100803, 3.180175e-05, 3.649078e-05, 1.50842e-05,
  1.299393e-05, 3.58945e-05, 0.0001151551, 0.0002152812, 0.0002524677, 
    0.0002098928, 0.000197359, 7.790486e-05, 0.0001293052, 7.806987e-05, 
    0.000111636, 4.944835e-05, 8.972455e-05, 5.927764e-05, 1.655547e-05,
  6.146031e-05, 0.0001586413, 0.0001716388, 0.0001572653, 4.799513e-05, 
    3.59903e-05, 2.371775e-05, 4.576848e-05, 3.408653e-05, 6.030597e-05, 
    0.0001407568, 9.720228e-05, 0.0001108642, 5.309374e-05, 7.754174e-06,
  0.0001921915, 0.0002451233, 0.0001376062, 0.0001141366, 0.0001024587, 
    8.808835e-05, 6.763274e-05, 6.790124e-05, 7.701424e-05, 6.656287e-05, 
    5.683576e-05, 8.269264e-05, 6.629803e-05, 1.794859e-05, 5.075728e-06,
  0.0002227609, 0.0003188555, 0.0003825098, 0.0003723797, 0.0003214547, 
    0.0002616246, 0.0002039467, 0.000157154, 0.0001547038, 4.911309e-05, 
    4.444614e-05, 4.752777e-05, 2.527433e-05, 7.529622e-06, 4.137662e-06,
  0.0002246319, 0.0003128261, 0.000348211, 0.0003318349, 0.0003323211, 
    0.0003922363, 0.0004082982, 0.0003381557, 0.0002939095, 0.000109997, 
    6.778968e-05, 3.864305e-05, 1.575496e-05, 6.340561e-06, 6.543656e-06,
  7.466022e-05, 0.0001586657, 0.0001747467, 0.0002293761, 0.0002532108, 
    0.0002836988, 0.0003294303, 0.000418875, 0.0003090138, 0.0001849475, 
    0.0001128815, 8.729102e-05, 1.76397e-05, 4.432586e-06, 5.320127e-06,
  3.533223e-05, 0.0001526653, 0.0001371524, 9.371398e-05, 0.000135784, 
    0.0001070626, 0.0001507718, 0.0002046779, 0.0001382888, 9.25302e-05, 
    0.0001893568, 7.881987e-05, 5.735347e-05, 1.965698e-05, 7.589499e-06,
  7.654622e-05, 0.0001413491, 0.000136023, 7.396831e-05, 8.740721e-05, 
    6.88342e-05, 7.777121e-05, 8.97718e-05, 0.0001374897, 0.0001623315, 
    0.0001713024, 0.0002156618, 0.0001109335, 3.858068e-05, 9.524851e-06,
  4.705325e-06, 1.506786e-05, 2.286924e-05, 2.119417e-05, 2.959137e-05, 
    2.348137e-05, 2.659843e-05, 3.865463e-05, 6.849728e-05, 3.963753e-05, 
    2.926566e-05, 3.158757e-05, 1.787791e-05, 0.0001192755, 0.0001544378,
  4.830577e-06, 1.173198e-05, 2.145036e-05, 2.428379e-05, 1.877922e-05, 
    1.532949e-05, 1.482628e-05, 2.234405e-05, 2.60205e-05, 1.770318e-05, 
    1.837445e-05, 8.866228e-06, 7.120256e-05, 0.0001437989, 0.0002575255,
  9.419814e-06, 1.459344e-05, 2.690106e-05, 1.730804e-05, 1.022584e-05, 
    1.680391e-05, 1.245958e-05, 1.865006e-05, 1.378004e-05, 7.927662e-06, 
    9.215058e-06, 3.923467e-05, 9.28683e-05, 0.00021613, 0.0003153937,
  1.165576e-05, 2.092859e-05, 2.069347e-05, 1.205003e-05, 1.31293e-05, 
    5.513058e-06, 1.062094e-05, 7.137872e-06, 5.307542e-06, 8.957802e-06, 
    1.904451e-05, 4.161843e-05, 0.0001325114, 0.0002126675, 0.0002145135,
  1.243812e-05, 1.96786e-05, 2.007507e-05, 1.595473e-05, 1.301027e-05, 
    8.755555e-06, 7.214715e-06, 4.218915e-06, 6.886067e-06, 2.187236e-05, 
    2.896565e-05, 5.868716e-05, 0.0001043053, 0.0001136948, 0.0001091401,
  1.264535e-05, 1.690237e-05, 1.450797e-05, 1.755825e-05, 1.72064e-05, 
    1.338883e-05, 1.102278e-05, 1.661034e-05, 7.893323e-05, 0.0001331374, 
    0.0001353181, 0.0001247786, 0.0001126688, 0.0001078305, 9.545283e-05,
  1.008473e-05, 1.163629e-05, 1.75657e-05, 1.880573e-05, 2.061551e-05, 
    1.896277e-05, 1.892487e-05, 9.566016e-05, 0.0001858782, 0.0003997721, 
    0.0001976744, 0.0001080939, 6.004232e-05, 4.068959e-05, 1.715696e-05,
  1.130602e-05, 1.584145e-05, 1.659754e-05, 1.808613e-05, 2.312682e-05, 
    1.997657e-05, 1.933878e-05, 0.0001013987, 0.0002195618, 0.0002491582, 
    0.0001640871, 3.947835e-05, 4.99779e-05, 1.500382e-05, 8.610508e-06,
  1.181837e-05, 1.447514e-05, 1.939078e-05, 2.59408e-05, 2.610607e-05, 
    2.780164e-05, 2.149842e-05, 1.946888e-05, 7.168495e-05, 5.454042e-05, 
    3.090016e-05, 1.657482e-05, 2.48274e-05, 6.815445e-05, 2.515816e-05,
  9.572419e-06, 1.514369e-05, 2.125401e-05, 2.644659e-05, 2.916941e-05, 
    2.965324e-05, 2.347855e-05, 3.132552e-05, 2.10301e-05, 5.519362e-05, 
    4.45335e-05, 2.93478e-05, 6.55729e-05, 8.014822e-05, 4.902951e-05,
  4.481913e-06, 6.981139e-06, 7.853919e-06, 9.3744e-06, 7.478746e-06, 
    9.059583e-06, 9.40905e-06, 8.3601e-06, 8.20201e-06, 9.977492e-06, 
    1.15476e-05, 1.349922e-05, 1.706483e-05, 2.7853e-05, 3.333324e-05,
  2.122825e-06, 3.209999e-06, 5.084078e-06, 6.825822e-06, 7.819342e-06, 
    6.970444e-06, 4.752015e-06, 5.959291e-06, 6.658888e-06, 6.327292e-06, 
    6.334587e-06, 5.349872e-06, 6.240433e-06, 1.017019e-05, 1.424795e-05,
  1.851258e-06, 2.592044e-06, 4.521236e-06, 4.736284e-06, 6.239045e-06, 
    5.434173e-06, 5.787176e-06, 4.609527e-06, 4.446833e-06, 5.15227e-06, 
    5.701106e-06, 3.015457e-06, 3.752104e-06, 4.591596e-06, 6.974622e-06,
  2.106276e-06, 1.789789e-06, 3.284549e-06, 3.6896e-06, 4.498255e-06, 
    4.75809e-06, 5.057532e-06, 5.579982e-06, 7.43423e-06, 6.193487e-06, 
    4.512654e-06, 2.775746e-06, 3.405299e-06, 3.440982e-06, 3.054169e-06,
  2.395258e-06, 2.594007e-06, 2.453995e-06, 2.496249e-06, 4.325373e-06, 
    4.848445e-06, 5.760298e-06, 6.777263e-06, 6.659403e-06, 4.980352e-06, 
    4.225305e-06, 3.666785e-06, 3.411519e-06, 2.616935e-06, 3.30848e-06,
  2.665418e-06, 2.709447e-06, 2.258847e-06, 3.183711e-06, 3.356374e-06, 
    4.688287e-06, 6.068512e-06, 7.624962e-06, 5.3925e-06, 4.323942e-06, 
    3.421872e-06, 3.160259e-06, 3.300373e-06, 2.376979e-06, 2.322322e-06,
  3.328129e-06, 3.465635e-06, 3.883651e-06, 4.749432e-06, 5.604653e-06, 
    6.762544e-06, 8.09951e-06, 6.730691e-06, 5.550998e-06, 4.557706e-06, 
    3.333512e-06, 3.484048e-06, 3.388543e-06, 1.645236e-06, 1.921142e-06,
  4.969034e-06, 4.941896e-06, 6.083526e-06, 7.574944e-06, 1.021416e-05, 
    1.024028e-05, 8.981641e-06, 6.0852e-06, 6.182278e-06, 5.895271e-06, 
    3.41691e-06, 5.575954e-06, 3.782491e-06, 3.697794e-06, 5.605706e-06,
  7.743047e-06, 7.676741e-06, 8.848888e-06, 9.908698e-06, 1.42313e-05, 
    1.297129e-05, 8.914699e-06, 7.615789e-06, 4.863305e-06, 6.414582e-06, 
    9.361185e-06, 7.47393e-06, 6.084303e-06, 7.659193e-06, 1.930738e-05,
  8.696647e-06, 1.086207e-05, 1.082536e-05, 1.206317e-05, 1.45055e-05, 
    1.217444e-05, 9.35289e-06, 8.724439e-06, 1.093217e-05, 1.076393e-05, 
    8.631742e-06, 8.305183e-06, 1.034409e-05, 1.836114e-05, 2.507923e-05,
  5.504486e-06, 6.089473e-06, 7.867449e-06, 5.733615e-06, 6.482814e-06, 
    5.915495e-06, 7.184247e-06, 5.929863e-06, 6.906152e-06, 7.728201e-06, 
    1.169269e-05, 1.719584e-05, 2.217627e-05, 3.159042e-05, 5.630132e-05,
  8.697728e-06, 7.26636e-06, 7.096859e-06, 5.660011e-06, 5.873192e-06, 
    6.838286e-06, 5.904085e-06, 5.939331e-06, 5.627559e-06, 5.935967e-06, 
    7.50489e-06, 9.93239e-06, 1.17184e-05, 1.876342e-05, 2.672207e-05,
  4.758299e-06, 8.22888e-06, 6.023812e-06, 5.811076e-06, 6.352991e-06, 
    7.55208e-06, 7.079347e-06, 7.614694e-06, 6.356695e-06, 6.998084e-06, 
    5.492628e-06, 6.116788e-06, 7.674236e-06, 1.031432e-05, 1.768088e-05,
  3.13766e-06, 3.862873e-06, 6.684385e-06, 5.223937e-06, 5.694831e-06, 
    7.481505e-06, 6.624978e-06, 6.652853e-06, 5.723071e-06, 5.943962e-06, 
    5.030525e-06, 4.653409e-06, 5.856943e-06, 8.105857e-06, 1.034781e-05,
  2.586188e-06, 3.073709e-06, 4.734607e-06, 5.365885e-06, 6.920033e-06, 
    6.218428e-06, 7.204727e-06, 5.828987e-06, 6.865651e-06, 7.041911e-06, 
    5.967275e-06, 5.592768e-06, 7.320128e-06, 7.307075e-06, 7.883556e-06,
  2.256945e-06, 2.420294e-06, 2.274011e-06, 3.789692e-06, 4.526382e-06, 
    6.314993e-06, 7.483318e-06, 8.278311e-06, 6.559924e-06, 5.89379e-06, 
    7.112944e-06, 7.068492e-06, 7.23219e-06, 5.792608e-06, 8.556583e-06,
  1.752878e-06, 1.40208e-06, 2.590611e-06, 1.857749e-06, 2.741227e-06, 
    4.900671e-06, 5.826997e-06, 5.884584e-06, 5.823861e-06, 5.347792e-06, 
    5.280308e-06, 5.971883e-06, 7.394092e-06, 6.462321e-06, 7.482437e-06,
  2.20808e-06, 2.310994e-06, 1.698756e-06, 2.599317e-06, 3.483938e-06, 
    4.080033e-06, 3.385971e-06, 2.784392e-06, 3.61874e-06, 4.159403e-06, 
    5.998657e-06, 5.60012e-06, 5.086672e-06, 5.517829e-06, 5.126663e-06,
  4.870564e-06, 1.88122e-06, 2.234106e-06, 2.538781e-06, 3.300748e-06, 
    3.601399e-06, 2.572919e-06, 3.335623e-06, 4.15455e-06, 4.295725e-06, 
    3.9998e-06, 4.519817e-06, 4.021918e-06, 5.402677e-06, 4.331725e-06,
  4.54748e-06, 1.224583e-06, 2.600231e-06, 3.160927e-06, 3.055134e-06, 
    3.215699e-06, 2.80763e-06, 3.36814e-06, 3.38859e-06, 3.593854e-06, 
    4.142527e-06, 4.129156e-06, 5.396278e-06, 5.205163e-06, 5.548205e-06,
  1.321305e-05, 1.744174e-05, 1.652648e-05, 8.625419e-06, 4.04614e-06, 
    1.471177e-06, 2.747031e-06, 2.449809e-06, 1.389976e-06, 4.938771e-07, 
    4.050877e-06, 3.007102e-06, 4.896609e-06, 9.772174e-06, 1.338943e-05,
  2.177951e-05, 1.311931e-05, 1.747333e-05, 1.030775e-05, 6.634786e-06, 
    3.090791e-08, 6.118576e-08, 9.662539e-08, 5.384172e-07, 7.608573e-08, 
    8.671693e-07, 1.967212e-06, 5.90125e-06, 5.147288e-06, 9.622972e-06,
  1.915935e-05, 1.960824e-05, 1.565275e-05, 1.282635e-05, 5.802517e-06, 
    4.930611e-09, 5.011446e-09, 2.902397e-08, 1.17765e-07, 7.416057e-08, 
    2.229193e-07, 1.234525e-06, 3.40879e-06, 5.583808e-06, 5.833807e-06,
  1.017282e-05, 1.514131e-05, 1.30067e-05, 1.130599e-05, 4.568788e-06, 
    1.534219e-08, 4.409158e-09, 1.829319e-08, 6.040772e-08, 2.436954e-08, 
    3.726299e-08, 2.505365e-07, 9.502494e-07, 1.963907e-06, 3.677158e-06,
  6.879237e-06, 7.505561e-06, 1.046234e-05, 1.266355e-05, 6.230227e-06, 
    2.622926e-06, 4.862606e-09, 3.866929e-09, 7.359866e-09, 5.201339e-09, 
    6.579774e-08, 3.945899e-08, 2.396264e-07, 8.187828e-07, 1.360712e-06,
  5.035715e-06, 4.629509e-06, 4.593496e-06, 7.194723e-06, 8.705663e-06, 
    5.539376e-06, 1.70514e-07, 1.000119e-08, 3.449424e-09, 6.981713e-09, 
    2.712014e-08, 6.3556e-09, 2.337653e-08, 3.037108e-07, 2.918839e-07,
  5.053999e-06, 6.281398e-06, 3.755333e-06, 5.036005e-06, 8.140336e-06, 
    6.927819e-06, 4.024198e-06, 2.535521e-07, 1.110847e-07, 9.072388e-08, 
    1.357263e-08, 6.999723e-09, 2.98807e-09, 1.555402e-08, 2.049976e-07,
  7.154195e-06, 3.809815e-06, 4.631408e-06, 5.233869e-06, 9.78765e-06, 
    1.271619e-05, 7.759254e-06, 1.803187e-06, 1.077795e-06, 1.8126e-07, 
    4.527874e-08, 3.769605e-08, 1.01493e-08, 2.459691e-08, 2.910577e-08,
  6.923123e-06, 3.967211e-06, 4.435297e-06, 5.229585e-06, 6.713726e-06, 
    7.817292e-06, 5.682786e-06, 3.524107e-06, 1.526068e-06, 1.292113e-06, 
    1.073168e-06, 8.312696e-07, 3.910055e-07, 1.938052e-07, 1.697694e-07,
  6.223936e-06, 7.218314e-06, 5.543832e-06, 6.339808e-06, 6.257416e-06, 
    6.413773e-06, 3.302909e-06, 4.153731e-06, 4.061817e-06, 2.695071e-06, 
    1.472843e-06, 9.62188e-07, 1.008231e-06, 4.197601e-07, 5.54844e-07,
  8.612026e-06, 1.290852e-05, 1.747163e-05, 2.773697e-05, 3.578165e-05, 
    5.045422e-05, 7.731669e-05, 7.446212e-05, 7.341951e-05, 2.632306e-05, 
    1.245159e-05, 8.1552e-06, 1.459513e-05, 2.451e-05, 2.850922e-05,
  1.00109e-05, 1.569144e-05, 2.205832e-05, 2.283555e-05, 2.719295e-05, 
    2.863878e-05, 3.847039e-05, 4.321748e-05, 5.519769e-05, 6.269358e-05, 
    5.681935e-05, 1.575409e-05, 1.038937e-05, 1.644933e-05, 2.040002e-05,
  1.420128e-05, 1.528744e-05, 2.734194e-05, 2.719566e-05, 2.454704e-05, 
    1.767107e-05, 2.024016e-05, 1.996737e-05, 2.778188e-05, 4.318262e-05, 
    5.682313e-05, 5.420448e-05, 2.452604e-05, 1.016256e-05, 1.501734e-05,
  1.11602e-05, 1.515742e-05, 2.095581e-05, 1.909534e-05, 1.438137e-05, 
    1.256143e-05, 1.44046e-05, 1.545308e-05, 1.505777e-05, 1.46187e-05, 
    2.1837e-05, 2.315903e-05, 2.443089e-05, 1.749862e-05, 1.246959e-05,
  1.38777e-05, 1.886112e-05, 2.391406e-05, 9.007713e-06, 7.26819e-06, 
    5.204204e-06, 9.033241e-06, 1.700831e-05, 9.975529e-06, 7.076985e-06, 
    1.783436e-07, 1.176074e-06, 4.955098e-06, 1.022822e-05, 1.449674e-05,
  1.083695e-05, 2.101629e-05, 1.297327e-05, 5.776032e-06, 5.336406e-06, 
    6.17472e-06, 1.496639e-05, 2.31023e-05, 1.422441e-05, 1.216356e-06, 
    5.625365e-08, 6.587043e-08, 5.437986e-07, 4.843224e-06, 7.940489e-06,
  1.592583e-05, 1.992783e-05, 1.348411e-05, 8.607741e-06, 3.701983e-06, 
    8.08276e-06, 2.268062e-05, 4.483525e-05, 2.783522e-05, 3.049917e-06, 
    5.078243e-08, 3.466014e-08, 3.672789e-07, 2.332771e-06, 6.067726e-06,
  1.606522e-05, 1.125467e-05, 7.754854e-06, 6.089005e-06, 1.242782e-05, 
    2.297714e-05, 4.004714e-05, 6.067047e-05, 3.598459e-05, 5.256545e-07, 
    1.159495e-09, 1.031359e-08, 7.047419e-08, 1.383087e-06, 3.666714e-06,
  1.040929e-05, 6.307967e-06, 5.725155e-06, 4.508756e-06, 1.162069e-05, 
    2.516957e-05, 3.859007e-05, 4.436561e-05, 1.407431e-05, 8.725679e-10, 
    5.318453e-10, 1.538378e-09, 5.711854e-08, 5.720486e-07, 3.245656e-06,
  7.474433e-06, 6.308729e-06, 5.116894e-06, 4.61521e-06, 7.592511e-06, 
    1.642412e-05, 2.493771e-05, 2.303735e-05, 4.007171e-06, 1.940337e-09, 
    1.962263e-10, 6.546355e-10, 1.808578e-08, 6.855895e-07, 6.930877e-07,
  9.782069e-06, 1.380734e-05, 3.629467e-05, 3.705281e-05, 6.499095e-05, 
    6.404156e-05, 5.570323e-05, 4.268477e-05, 7.025719e-05, 7.501548e-05, 
    8.902473e-05, 7.296717e-05, 5.771866e-05, 6.66311e-05, 4.278877e-05,
  4.951651e-06, 4.578082e-06, 2.957208e-05, 7.03422e-05, 5.997208e-05, 
    6.189446e-05, 7.810658e-05, 8.615366e-05, 6.846791e-05, 7.756102e-05, 
    7.38428e-05, 6.958376e-05, 5.521491e-05, 4.784134e-05, 3.445581e-05,
  2.175673e-06, 4.37642e-06, 1.271379e-05, 8.805275e-05, 6.123198e-05, 
    6.362193e-05, 9.911259e-05, 3.786215e-05, 4.050746e-05, 8.601683e-05, 
    3.392586e-05, 4.999105e-05, 4.98466e-05, 3.150586e-05, 2.706813e-05,
  3.16719e-07, 9.008692e-07, 8.203102e-06, 1.134304e-05, 1.11128e-05, 
    1.450457e-05, 1.949983e-06, 1.72199e-06, 1.19225e-05, 1.453698e-05, 
    2.108828e-05, 3.70525e-05, 4.680817e-05, 3.457862e-05, 2.747329e-05,
  1.70814e-08, 3.997181e-07, 2.492338e-06, 1.592989e-07, 3.883134e-06, 
    2.181964e-06, 5.767622e-07, 1.219525e-06, 1.171693e-05, 1.608271e-05, 
    1.146775e-05, 9.302462e-06, 1.448751e-05, 1.195867e-05, 1.734489e-05,
  1.747273e-06, 4.190215e-06, 6.092414e-06, 1.697967e-06, 5.38028e-08, 
    1.842626e-06, 7.401996e-08, 7.998786e-06, 3.211912e-05, 2.35338e-05, 
    5.952486e-06, 7.755158e-06, 2.47777e-06, 6.647045e-06, 3.261712e-06,
  5.613173e-06, 7.760675e-06, 1.18781e-05, 7.317633e-06, 1.071238e-06, 
    1.786825e-05, 2.258302e-05, 3.592403e-05, 4.719973e-05, 4.36091e-05, 
    1.685125e-05, 9.305352e-06, 3.075642e-07, 6.707845e-08, 3.912173e-07,
  2.468374e-06, 4.723053e-06, 9.163791e-06, 1.280982e-05, 2.146313e-05, 
    3.147029e-05, 5.376465e-05, 7.320639e-05, 7.669611e-05, 2.56127e-05, 
    2.045713e-06, 5.721157e-07, 1.984725e-07, 8.549343e-08, 5.24848e-08,
  2.37129e-06, 4.211536e-06, 8.473629e-06, 1.141262e-05, 1.871869e-05, 
    2.851672e-05, 3.93142e-05, 4.711618e-05, 4.074351e-05, 2.190625e-06, 
    8.886214e-08, 5.573461e-08, 2.792928e-08, 3.479728e-07, 1.29834e-07,
  3.594115e-06, 5.120292e-06, 7.889498e-06, 8.534473e-06, 1.361255e-05, 
    2.073897e-05, 2.261879e-05, 1.847132e-05, 4.03929e-06, 5.765326e-09, 
    9.071741e-09, 4.186744e-08, 6.685879e-09, 3.141031e-08, 2.918696e-07,
  0.0001445243, 0.0001587234, 0.0002007791, 0.0002229728, 0.0001847964, 
    0.0001984701, 0.0002204312, 0.0002191195, 0.0002299382, 0.0002271368, 
    0.0004768007, 0.0003594099, 0.000164144, 0.0002940071, 0.0002491202,
  9.8374e-05, 0.0001063468, 0.0001196725, 0.0001643436, 0.0002169587, 
    0.0002638029, 0.0002925946, 0.0002431245, 0.0002214286, 0.0003855592, 
    0.0003372652, 0.0001592113, 0.0001233192, 0.0001379971, 0.0001676421,
  4.993586e-05, 5.503876e-05, 7.937735e-05, 0.0001112048, 9.69968e-05, 
    0.0001620866, 0.0001600389, 0.0001873701, 0.0001674661, 0.0001274372, 
    0.0001180659, 0.0001400583, 9.439597e-05, 0.0001159654, 0.0001388264,
  7.118061e-06, 3.609542e-05, 2.565611e-05, 1.565937e-05, 8.207017e-05, 
    4.259889e-05, 7.407321e-05, 0.0001227641, 0.0001094938, 0.0001002325, 
    9.745714e-05, 5.953914e-05, 0.0001309943, 9.48104e-05, 0.0001252064,
  1.03112e-05, 1.482368e-05, 1.58077e-05, 2.877922e-05, 2.372825e-05, 
    4.846989e-05, 5.489671e-05, 5.354672e-05, 9.260733e-05, 9.600628e-05, 
    8.967082e-05, 0.0001020022, 9.570585e-05, 7.637237e-05, 8.229313e-05,
  3.029698e-06, 3.08327e-06, 1.430017e-05, 1.686976e-05, 1.406149e-05, 
    4.22751e-05, 5.198003e-05, 0.0001218468, 5.724858e-05, 7.989829e-05, 
    7.930586e-05, 7.459961e-05, 7.8574e-05, 7.330936e-05, 9.598758e-05,
  1.904878e-06, 5.948142e-06, 8.725868e-06, 7.080223e-06, 1.96157e-05, 
    2.527343e-05, 5.57713e-05, 7.522265e-05, 8.245323e-05, 7.709592e-05, 
    0.0001060665, 0.0001541586, 0.0001686554, 7.850328e-05, 0.000157124,
  1.296253e-06, 5.018485e-06, 2.570972e-05, 3.176165e-05, 4.476995e-05, 
    7.216068e-05, 9.09844e-05, 3.736013e-05, 7.727473e-05, 6.000079e-05, 
    0.0001968482, 0.0002609102, 0.0002056647, 0.0002575804, 0.0001157939,
  5.796356e-07, 3.575314e-06, 1.205756e-05, 1.85611e-05, 4.393427e-05, 
    6.192794e-05, 9.663369e-05, 0.0001002428, 0.0001074466, 0.0001609586, 
    0.0002757118, 0.0002671981, 0.0002013177, 0.0001387502, 8.224395e-05,
  3.904934e-07, 2.424795e-06, 8.756162e-06, 1.43061e-05, 2.12483e-05, 
    4.105967e-05, 6.226479e-05, 0.0001421296, 0.0002201037, 0.0002548798, 
    0.0002101776, 0.0002260468, 0.0001760654, 0.0001688807, 3.067186e-05,
  4.612949e-08, 3.164157e-07, 1.950275e-07, 1.861016e-08, 5.076549e-08, 
    1.703222e-07, 1.918927e-06, 1.768529e-06, 2.013887e-06, 2.841792e-06, 
    3.380496e-06, 4.220495e-06, 6.076288e-06, 7.363028e-06, 1.305395e-05,
  2.648665e-08, 1.041308e-08, 6.736578e-08, 2.70683e-09, 6.989728e-09, 
    7.76031e-08, 6.956376e-07, 1.414198e-06, 2.029807e-06, 2.795304e-06, 
    3.006043e-06, 4.235763e-06, 3.961816e-06, 5.185553e-06, 1.147149e-05,
  3.310105e-08, 4.174983e-08, 1.558086e-08, 3.757531e-08, 1.207636e-09, 
    1.946023e-09, 1.435967e-08, 2.305795e-07, 2.866862e-07, 3.012775e-06, 
    2.40105e-06, 2.391023e-06, 3.910048e-06, 6.409609e-06, 1.098374e-05,
  1.523462e-07, 2.112601e-08, 2.815363e-08, 1.849079e-07, 4.784808e-09, 
    3.426552e-10, 1.591979e-09, 1.453783e-07, 1.210503e-07, 1.258447e-06, 
    2.327787e-06, 3.320695e-06, 3.425909e-06, 6.121287e-06, 9.484926e-06,
  9.916794e-08, 3.613825e-08, 4.617229e-08, 1.930634e-07, 1.504983e-07, 
    6.716272e-09, 1.06606e-08, 5.166763e-07, 4.4777e-07, 1.046605e-06, 
    3.999698e-06, 5.258778e-06, 5.016856e-06, 6.228551e-06, 5.709267e-06,
  2.248881e-06, 5.480346e-07, 1.628623e-07, 1.16863e-07, 2.464645e-07, 
    1.815498e-07, 3.474325e-07, 3.736924e-07, 5.505167e-07, 1.0569e-06, 
    1.08663e-06, 2.106061e-06, 4.124268e-06, 5.272228e-06, 5.549428e-06,
  4.340825e-06, 2.897969e-06, 7.168441e-07, 1.857632e-07, 2.176792e-07, 
    3.328691e-07, 4.448385e-07, 6.597177e-07, 7.122448e-07, 1.15997e-06, 
    1.278907e-06, 2.436504e-06, 4.087147e-06, 1.047074e-05, 7.618311e-06,
  6.458733e-06, 4.809267e-06, 4.005714e-06, 9.622888e-07, 2.225671e-07, 
    3.478335e-07, 6.47239e-07, 6.723018e-07, 1.303628e-06, 1.107168e-06, 
    1.378991e-06, 2.999313e-06, 5.026292e-06, 6.797634e-06, 1.203628e-05,
  6.949409e-06, 8.749753e-06, 1.088276e-05, 4.350533e-06, 9.123843e-07, 
    4.344745e-07, 9.96445e-07, 9.100167e-07, 1.346914e-06, 1.635238e-06, 
    2.21228e-06, 3.680142e-06, 4.296452e-06, 8.558191e-06, 9.417437e-05,
  6.977848e-06, 1.010305e-05, 9.598785e-06, 1.16345e-05, 1.58311e-06, 
    3.945772e-07, 3.541601e-07, 8.706447e-07, 1.656162e-06, 1.203943e-06, 
    2.035173e-06, 1.533416e-06, 3.178359e-06, 2.741288e-05, 0.0001338508,
  7.199427e-05, 3.395106e-05, 2.272939e-05, 1.512316e-05, 1.281466e-05, 
    9.567833e-06, 1.059231e-05, 8.503915e-06, 6.433994e-06, 7.627798e-06, 
    1.342985e-05, 9.240278e-06, 8.045474e-06, 7.635332e-06, 8.076276e-06,
  4.715119e-05, 2.828085e-05, 2.273506e-05, 1.479437e-05, 1.084291e-05, 
    6.908885e-06, 7.804239e-06, 5.938537e-06, 4.219213e-06, 4.346457e-06, 
    6.26486e-06, 1.044126e-05, 8.110141e-06, 6.253947e-06, 6.141936e-06,
  3.36592e-05, 1.933307e-05, 2.261569e-05, 1.539101e-05, 9.750092e-06, 
    4.34533e-06, 7.135047e-06, 5.059163e-06, 3.238813e-06, 2.70398e-06, 
    3.779055e-06, 2.81311e-06, 4.033154e-06, 3.836888e-06, 3.990352e-06,
  3.121122e-05, 1.431792e-05, 1.521668e-05, 1.431685e-05, 9.189262e-06, 
    5.27011e-06, 4.422451e-06, 4.356615e-06, 4.646373e-06, 4.329278e-06, 
    3.370877e-06, 4.770176e-06, 4.740929e-06, 5.042682e-06, 2.998543e-06,
  1.913387e-05, 2.074214e-05, 1.191753e-05, 1.541611e-05, 1.180359e-05, 
    5.724748e-06, 5.922309e-06, 5.11635e-06, 4.744571e-06, 4.541068e-06, 
    3.708371e-06, 3.664313e-06, 4.009267e-06, 1.9466e-06, 4.530129e-06,
  2.603557e-05, 1.423309e-05, 1.237942e-05, 1.347311e-05, 1.501725e-05, 
    9.006811e-06, 3.952269e-06, 3.101084e-06, 6.396767e-06, 4.211853e-06, 
    3.155501e-06, 2.110276e-06, 1.349596e-06, 9.611566e-07, 2.000148e-06,
  2.327766e-05, 1.124389e-05, 1.384801e-05, 1.43374e-05, 1.695328e-05, 
    1.563694e-05, 9.499545e-06, 7.619973e-06, 4.099145e-06, 2.76589e-06, 
    3.363022e-06, 2.088347e-06, 1.265833e-06, 6.51438e-07, 1.038397e-06,
  1.532062e-05, 2.28893e-05, 1.512877e-05, 1.885406e-05, 2.825948e-05, 
    3.04948e-05, 2.304763e-05, 1.043198e-05, 7.882487e-06, 4.862335e-06, 
    2.773857e-06, 3.369014e-06, 2.263856e-06, 9.303296e-07, 1.414085e-07,
  1.497756e-05, 1.71665e-05, 1.636382e-05, 2.078333e-05, 3.056131e-05, 
    4.022838e-05, 3.947601e-05, 2.630731e-05, 1.024624e-05, 5.530168e-06, 
    3.734908e-06, 4.753945e-06, 3.082154e-06, 1.737313e-06, 1.197946e-06,
  9.989791e-06, 1.451996e-05, 1.672274e-05, 2.034099e-05, 3.188615e-05, 
    4.263788e-05, 4.770289e-05, 4.019889e-05, 1.825162e-05, 6.824909e-06, 
    4.051459e-06, 3.297297e-06, 3.393407e-06, 2.929899e-06, 2.475236e-06,
  0.0002044186, 0.0002688133, 0.0001832907, 0.0002287974, 0.0002644899, 
    0.0002460546, 0.0002479591, 0.0002813008, 0.0002619504, 0.0004484377, 
    0.0003665588, 0.0001361005, 1.698658e-05, 1.615497e-05, 1.446804e-05,
  0.0002189724, 0.0002115354, 0.0002540314, 0.0002230336, 0.0002001838, 
    0.0001804142, 0.0001864131, 0.0002060387, 0.0002760332, 0.0004542976, 
    0.0002949855, 2.435135e-05, 1.501687e-05, 2.190103e-05, 2.496955e-05,
  0.0002027986, 0.0002219416, 0.0002177032, 0.0002172881, 0.0001707481, 
    9.33482e-05, 0.000102947, 0.000153669, 0.0003444059, 0.0003945399, 
    0.0001273705, 1.43539e-05, 1.749959e-05, 2.987961e-05, 4.197114e-05,
  0.0002603913, 0.00023845, 0.000209431, 0.0001681376, 0.0001574026, 
    0.0001172981, 0.0001338847, 0.0001900928, 0.0003173891, 0.0002685784, 
    4.195514e-05, 3.117963e-05, 8.074542e-05, 0.0001306317, 0.0001236258,
  0.0002099162, 0.0002280671, 0.0002143266, 0.0001348323, 0.0001038399, 
    0.0001508595, 0.000128014, 0.0001696494, 0.0002604678, 0.0001323171, 
    5.533244e-05, 0.0001391911, 0.0002088225, 0.0002419863, 0.0002068707,
  0.0002768669, 0.0003065223, 0.0002649058, 0.0002053155, 0.0001733524, 
    0.0001830426, 0.0001326175, 0.0001469215, 0.0001298466, 0.0001339907, 
    0.0001712656, 0.0002870238, 0.0002914661, 0.0002776052, 0.0002436128,
  0.0002529373, 0.0003466964, 0.0003676173, 0.0003128817, 0.0002151056, 
    0.0001746315, 0.0001409497, 0.0001401526, 0.0001197839, 0.0001770992, 
    0.0002980033, 0.000355243, 0.0003401868, 0.0003109525, 0.0002412347,
  0.0003218532, 0.000359471, 0.000490038, 0.0003311698, 0.0002684153, 
    0.0001682821, 0.0001588094, 0.0001407562, 0.000143676, 0.0002383438, 
    0.0003762198, 0.0004018146, 0.0003645761, 0.0002825749, 0.0001799756,
  0.0003410201, 0.0003905113, 0.0004206176, 0.0003126038, 0.0002607793, 
    0.000177784, 0.0001168594, 0.0001168023, 0.0001535572, 0.0002719169, 
    0.0003945667, 0.0003663701, 0.0002932886, 0.0001992759, 0.0001008054,
  0.0002010836, 0.0002362268, 0.0002725196, 0.0002504244, 0.0001654595, 
    0.0001112852, 8.483479e-05, 7.317238e-05, 0.0002264167, 0.0003295706, 
    0.000369525, 0.0003537418, 0.0001601528, 0.0001065108, 6.890357e-05,
  2.260704e-05, 3.553947e-05, 4.324104e-05, 4.981328e-05, 4.757436e-05, 
    6.034668e-05, 8.43711e-05, 0.0001082105, 0.0001334929, 0.0001549888, 
    0.0001305701, 0.0001106663, 0.000143437, 0.000233777, 0.0002480858,
  3.876815e-05, 3.541448e-05, 4.073699e-05, 4.472182e-05, 4.584124e-05, 
    5.512829e-05, 8.962079e-05, 0.0001257147, 0.0001320342, 0.0001066603, 
    8.350601e-05, 7.205507e-05, 9.985318e-05, 0.0002030234, 0.0003124044,
  3.607335e-05, 3.022473e-05, 3.884813e-05, 4.036328e-05, 5.164244e-05, 
    4.568673e-05, 8.017055e-05, 0.0001030448, 0.0001010227, 6.595923e-05, 
    4.420599e-05, 4.985452e-05, 4.793049e-05, 0.0001239727, 0.0003158545,
  3.28625e-05, 2.909419e-05, 3.701237e-05, 3.981979e-05, 4.348728e-05, 
    4.195396e-05, 5.619639e-05, 9.190739e-05, 6.67227e-05, 3.737918e-05, 
    1.271688e-05, 1.289188e-05, 1.919971e-05, 7.115531e-05, 0.0002964227,
  3.114342e-05, 2.937427e-05, 3.926664e-05, 3.548073e-05, 3.894191e-05, 
    5.435734e-05, 5.768356e-05, 7.726892e-05, 5.79747e-05, 2.155528e-05, 
    4.129981e-06, 1.463953e-05, 5.377732e-06, 3.713512e-05, 0.0002444805,
  2.636893e-05, 2.458919e-05, 3.686595e-05, 3.600617e-05, 3.890043e-05, 
    4.133761e-05, 5.967669e-05, 7.615642e-05, 4.72734e-05, 1.146097e-05, 
    1.390888e-06, 7.424287e-06, 3.392829e-06, 2.042394e-05, 0.0002004911,
  3.026241e-05, 2.924269e-05, 3.407527e-05, 3.907637e-05, 4.647589e-05, 
    4.378752e-05, 4.458509e-05, 5.900518e-05, 3.861483e-05, 9.591929e-06, 
    2.422665e-06, 2.479788e-05, 1.105817e-05, 1.271548e-05, 0.0001562308,
  2.97434e-05, 3.00333e-05, 3.948294e-05, 4.383646e-05, 5.476434e-05, 
    5.409988e-05, 5.072707e-05, 5.724667e-05, 4.526947e-05, 2.218833e-05, 
    4.466309e-06, 6.155603e-05, 2.52991e-05, 4.169102e-05, 0.0001114406,
  3.063683e-05, 3.824157e-05, 4.5926e-05, 4.966953e-05, 7.220826e-05, 
    7.591632e-05, 6.464556e-05, 7.045522e-05, 7.456111e-05, 0.00014761, 
    7.283485e-05, 8.364811e-05, 5.95495e-05, 7.638832e-05, 7.911122e-05,
  4.113189e-05, 5.327422e-05, 7.937397e-05, 0.0001043469, 9.615916e-05, 
    0.0001050123, 0.0001515447, 0.0001019844, 0.0002627923, 0.0003799851, 
    0.0001483467, 6.168705e-05, 6.743301e-05, 4.842681e-05, 5.747826e-05,
  6.968751e-05, 9.094225e-05, 9.673722e-05, 6.275293e-05, 4.690505e-05, 
    2.351075e-05, 4.170873e-05, 4.984066e-05, 2.713376e-05, 5.240462e-05, 
    2.424034e-05, 3.454441e-05, 2.340155e-05, 7.327939e-05, 0.0001996503,
  3.653124e-05, 9.261777e-05, 0.0001249922, 5.620483e-05, 5.969763e-05, 
    2.551618e-05, 3.463622e-05, 4.521841e-05, 2.478544e-05, 1.808364e-05, 
    2.237828e-05, 3.859835e-05, 5.999035e-05, 0.000143508, 0.0002028879,
  2.553774e-05, 3.710627e-05, 3.981426e-05, 7.464008e-05, 4.585972e-05, 
    2.156928e-05, 3.100364e-05, 3.809399e-05, 2.20291e-05, 1.493545e-05, 
    2.046577e-05, 5.102015e-05, 0.0001069482, 0.0002515063, 0.000181273,
  1.100195e-05, 1.462562e-05, 2.546674e-05, 2.78168e-05, 2.60674e-05, 
    1.311701e-05, 2.539159e-05, 2.585568e-05, 2.074376e-05, 1.642916e-05, 
    1.795951e-05, 3.342764e-05, 0.0001496579, 0.0001903401, 0.0001196259,
  5.719758e-07, 2.090493e-06, 8.712153e-06, 1.182506e-05, 1.070504e-05, 
    1.0272e-05, 3.301537e-05, 2.719637e-05, 2.299953e-05, 1.193565e-05, 
    1.305808e-05, 4.75079e-05, 9.300803e-05, 0.0001309955, 0.0001147435,
  2.578316e-07, 1.285668e-06, 1.657602e-06, 3.628079e-06, 5.282155e-06, 
    1.219351e-05, 2.886353e-05, 2.948044e-05, 2.180529e-05, 1.303156e-05, 
    2.614938e-05, 8.276459e-05, 7.112476e-05, 8.289504e-05, 8.065198e-05,
  1.013555e-07, 7.022642e-07, 1.602171e-06, 2.486284e-06, 4.416204e-06, 
    9.911124e-06, 1.941654e-05, 2.511476e-05, 2.339504e-05, 2.061709e-05, 
    3.535393e-05, 7.873643e-05, 6.285172e-05, 5.107913e-05, 0.0001015838,
  1.219094e-07, 3.616711e-07, 1.959407e-06, 1.99787e-06, 3.459681e-06, 
    7.160485e-06, 1.03999e-05, 1.581515e-05, 2.057803e-05, 2.709565e-05, 
    6.537829e-05, 7.142865e-05, 8.187566e-05, 5.119773e-05, 8.371697e-05,
  2.168005e-07, 1.89641e-07, 1.049552e-06, 2.578797e-06, 5.284361e-06, 
    1.042131e-05, 7.654256e-06, 1.204401e-05, 1.715553e-05, 6.490049e-05, 
    0.0001377001, 8.931219e-05, 2.993403e-05, 4.64877e-05, 6.473711e-05,
  4.78651e-07, 2.224954e-07, 1.00709e-06, 3.270486e-06, 7.472651e-06, 
    9.610843e-06, 1.035413e-05, 1.278664e-05, 2.236938e-05, 9.562522e-05, 
    0.0001678604, 4.399818e-05, 4.104942e-05, 2.855835e-05, 3.719843e-05,
  2.766209e-05, 3.741308e-05, 3.514977e-05, 4.438354e-05, 7.604726e-05, 
    0.000108393, 0.0001162587, 0.0001398666, 7.51165e-05, 9.684121e-05, 
    6.636948e-05, 7.269023e-05, 7.756823e-05, 6.777324e-05, 8.621439e-05,
  7.007626e-06, 1.280191e-05, 1.229713e-05, 2.213449e-05, 1.919099e-05, 
    5.034055e-05, 9.181337e-05, 0.0001089926, 8.946531e-05, 0.0001024242, 
    9.122933e-05, 4.384016e-05, 4.628278e-05, 3.202324e-05, 5.685148e-05,
  1.490903e-06, 1.430462e-06, 5.020009e-06, 1.275791e-05, 1.856271e-05, 
    4.734466e-05, 5.280371e-05, 4.980918e-05, 8.231743e-05, 9.931617e-05, 
    6.76405e-05, 4.69216e-05, 4.059715e-05, 2.711846e-05, 4.043e-05,
  7.703935e-08, 4.903108e-07, 1.671332e-06, 4.939893e-06, 1.098742e-05, 
    2.426341e-05, 2.710837e-05, 2.232372e-05, 2.542223e-05, 3.170672e-05, 
    2.456851e-05, 2.192366e-05, 3.377339e-05, 1.773667e-05, 1.672192e-05,
  3.459986e-10, 1.580318e-08, 6.715058e-07, 2.331704e-06, 3.797177e-06, 
    7.743957e-06, 4.943173e-06, 5.434019e-06, 6.963749e-06, 7.362284e-06, 
    4.480567e-06, 3.378399e-06, 1.830081e-05, 6.478393e-06, 1.507652e-05,
  3.516272e-10, 4.472988e-10, 5.27213e-10, 6.89059e-08, 1.305385e-08, 
    2.169817e-06, 6.689106e-06, 4.224941e-06, 1.415572e-06, 2.803347e-06, 
    1.10025e-06, 3.62476e-06, 4.444894e-06, 5.297153e-06, 1.211547e-05,
  8.086965e-11, 9.915432e-11, 1.398105e-10, 1.428722e-10, 1.214155e-10, 
    1.592651e-06, 3.619916e-06, 4.770262e-06, 7.175526e-07, 6.349434e-06, 
    4.0777e-06, 1.179099e-05, 7.383151e-06, 1.10372e-05, 1.296136e-05,
  3.275885e-11, 4.107596e-11, 5.047231e-11, 5.029901e-11, 1.232289e-08, 
    6.884428e-07, 6.930667e-06, 4.459474e-06, 6.249406e-06, 4.987368e-06, 
    9.52683e-06, 8.74701e-06, 1.15035e-05, 1.532682e-05, 1.618866e-05,
  3.772903e-11, 1.053448e-10, 8.984511e-11, 3.734454e-11, 3.473994e-07, 
    3.044607e-06, 4.742579e-06, 7.810059e-06, 4.776432e-06, 1.033346e-05, 
    6.101067e-06, 7.058229e-06, 4.99052e-06, 1.391155e-05, 1.178643e-05,
  1.801291e-11, 1.32801e-10, 5.146708e-11, 4.000433e-07, 3.288544e-06, 
    1.328624e-05, 1.287038e-05, 1.046579e-05, 2.09521e-05, 9.862292e-06, 
    9.596786e-06, 1.434475e-05, 7.495685e-06, 1.479732e-05, 1.117885e-05,
  6.461608e-06, 8.53482e-06, 9.477396e-06, 1.290739e-05, 2.021485e-05, 
    1.728264e-05, 0.0001090054, 6.128335e-05, 3.808838e-05, 3.524283e-05, 
    8.075005e-05, 5.853042e-05, 6.663772e-05, 5.292773e-05, 6.84386e-05,
  7.546909e-07, 9.122467e-07, 9.511388e-07, 6.895668e-06, 7.031984e-06, 
    1.101136e-05, 1.872618e-05, 1.949682e-05, 3.512349e-05, 6.355879e-05, 
    4.187293e-05, 5.237198e-05, 3.637427e-05, 5.065214e-05, 4.16319e-05,
  6.103882e-10, 1.486136e-10, 1.425861e-06, 1.022733e-06, 7.873819e-06, 
    7.266628e-06, 1.162792e-05, 1.31983e-05, 1.649585e-05, 2.27777e-05, 
    2.379945e-05, 2.583941e-05, 9.065642e-06, 1.122853e-05, 1.801451e-05,
  1.816046e-09, 2.589064e-09, 1.760966e-08, 1.072419e-06, 1.035996e-06, 
    6.720476e-06, 8.337517e-06, 9.096812e-06, 1.060555e-05, 1.105181e-05, 
    1.746494e-05, 1.259658e-05, 8.874518e-06, 1.775364e-09, 4.22338e-09,
  5.100951e-10, 6.509517e-10, 1.945167e-10, 1.720627e-08, 1.112874e-10, 
    8.443954e-07, 2.107745e-06, 3.328977e-06, 3.789147e-06, 6.910077e-06, 
    1.015496e-05, 5.030367e-06, 7.373766e-06, 3.448508e-06, 1.904442e-06,
  8.318191e-10, 6.497796e-10, 2.207615e-10, 1.623923e-10, 1.092059e-10, 
    3.503515e-10, 3.93326e-10, 4.736644e-08, 6.606005e-07, 2.294505e-06, 
    2.632642e-06, 3.456019e-06, 5.304246e-06, 4.649903e-06, 3.869131e-06,
  6.091116e-10, 4.968913e-10, 8.92543e-10, 5.862962e-10, 4.904715e-10, 
    1.231806e-09, 6.773376e-10, 2.39589e-10, 3.21164e-08, 4.773942e-07, 
    5.84659e-07, 1.118814e-06, 1.698733e-06, 2.844086e-06, 6.528311e-06,
  1.265697e-10, 5.553715e-10, 1.527025e-08, 2.529645e-07, 8.461522e-07, 
    1.333546e-06, 1.188392e-09, 1.155237e-09, 4.078148e-10, 2.159195e-07, 
    3.211597e-07, 4.789906e-07, 1.16869e-06, 3.68909e-06, 3.91888e-06,
  9.503631e-12, 1.078591e-10, 1.851653e-07, 6.854249e-07, 7.780582e-07, 
    1.489582e-06, 1.782594e-06, 6.404338e-09, 1.218532e-07, 2.123513e-07, 
    6.074484e-07, 4.776172e-06, 1.07065e-06, 8.560019e-07, 2.123629e-06,
  6.231538e-24, 3.243769e-23, 1.76404e-08, 3.614105e-07, 8.531132e-07, 
    2.986444e-06, 3.513429e-06, 3.902041e-06, 4.316325e-06, 8.281839e-07, 
    1.999441e-08, 2.353845e-08, 2.616294e-08, 3.502437e-08, 1.53109e-05,
  4.123742e-08, 3.07107e-09, 3.82413e-09, 1.463287e-08, 8.422351e-08, 
    1.541541e-06, 6.250873e-06, 1.284203e-05, 1.412161e-05, 2.286738e-05, 
    1.090085e-05, 1.205704e-05, 4.460867e-06, 2.425286e-06, 5.252738e-06,
  3.962095e-09, 4.732907e-09, 5.00335e-09, 5.889659e-09, 1.484804e-08, 
    2.444311e-07, 4.464555e-06, 2.508237e-05, 3.015372e-05, 1.11558e-05, 
    2.318338e-05, 1.294765e-05, 4.529194e-06, 7.128534e-06, 7.618258e-06,
  7.701741e-09, 6.237123e-09, 9.938595e-09, 1.2794e-08, 5.37028e-08, 
    6.088513e-07, 4.043394e-06, 6.759076e-06, 7.655137e-06, 1.195738e-05, 
    1.279003e-05, 1.239336e-05, 1.249683e-05, 1.171252e-05, 1.073727e-05,
  4.856459e-09, 4.876139e-09, 3.991156e-09, 1.675478e-08, 1.084087e-07, 
    3.061465e-07, 3.365413e-06, 6.24762e-06, 1.059772e-05, 1.006346e-05, 
    1.092441e-05, 1.033558e-05, 9.174374e-06, 7.955484e-06, 6.931126e-06,
  3.308376e-09, 1.462197e-09, 3.075326e-09, 4.154814e-08, 1.96872e-07, 
    1.597558e-07, 8.739902e-07, 2.229815e-06, 4.67054e-06, 4.95924e-06, 
    4.026554e-06, 2.769632e-06, 1.603044e-06, 1.90567e-06, 5.72975e-06,
  1.01093e-09, 2.254158e-09, 8.996076e-09, 3.094241e-08, 3.131557e-08, 
    1.137962e-07, 5.481546e-07, 1.330631e-07, 3.904783e-07, 1.510053e-07, 
    1.019968e-07, 8.991167e-08, 1.057296e-07, 2.223588e-07, 9.758114e-07,
  4.123739e-11, 2.902209e-09, 1.225573e-08, 1.467279e-08, 1.599022e-08, 
    9.952134e-07, 2.386429e-08, 3.551257e-06, 3.270846e-08, 7.381696e-08, 
    4.183812e-08, 1.449567e-07, 3.712798e-08, 7.518686e-08, 1.249308e-06,
  2.383199e-07, 1.687461e-06, 1.011751e-06, 1.301823e-06, 1.474164e-06, 
    1.826991e-06, 1.625498e-06, 9.044593e-08, 3.472755e-08, 3.898574e-08, 
    5.738545e-07, 2.24823e-07, 8.877549e-08, 5.065953e-08, 6.786327e-09,
  2.593569e-08, 5.806991e-07, 1.407128e-06, 8.520524e-07, 1.838646e-06, 
    2.375608e-06, 5.083177e-06, 2.125499e-07, 7.145511e-07, 9.073489e-07, 
    1.437391e-06, 9.675932e-07, 6.400287e-08, 3.634938e-07, 4.780154e-08,
  8.018383e-09, 4.789435e-07, 1.198623e-06, 1.438402e-07, 1.042049e-06, 
    1.531948e-06, 1.232041e-06, 1.801182e-06, 3.389751e-06, 2.799998e-06, 
    2.951231e-06, 1.63197e-06, 2.030259e-06, 2.705189e-07, 3.23909e-07,
  3.349978e-08, 7.315011e-09, 3.92931e-08, 1.599534e-07, 4.800685e-07, 
    1.883125e-07, 2.341484e-06, 1.184325e-06, 9.671038e-06, 1.25751e-05, 
    3.569972e-05, 5.858354e-05, 1.277407e-05, 2.596545e-05, 2.80408e-05,
  4.78623e-10, 6.340394e-10, 7.368481e-10, 3.100757e-09, 1.533277e-07, 
    5.388559e-07, 4.092676e-06, 1.030976e-05, 2.462775e-05, 3.450659e-05, 
    2.158114e-05, 1.656653e-05, 1.514652e-05, 1.119849e-05, 1.017666e-05,
  7.817751e-10, 1.592307e-09, 4.391655e-09, 5.083583e-07, 1.539412e-07, 
    9.011513e-07, 4.865203e-06, 1.38356e-05, 1.925297e-05, 2.112076e-05, 
    1.524189e-05, 1.088384e-05, 6.105219e-06, 4.383117e-06, 3.606347e-06,
  1.046552e-09, 2.531343e-09, 2.019735e-08, 1.209551e-07, 5.244031e-07, 
    6.61789e-06, 1.013419e-05, 1.0835e-05, 1.184202e-05, 7.988191e-06, 
    3.28289e-06, 2.165465e-06, 2.026962e-06, 2.028527e-06, 2.227713e-06,
  1.149389e-09, 3.34856e-09, 1.318363e-08, 1.393702e-07, 3.529286e-06, 
    8.05311e-06, 1.00679e-05, 7.544736e-06, 2.35684e-06, 1.442801e-07, 
    6.133186e-08, 2.397497e-07, 3.761916e-07, 7.705027e-07, 1.895062e-06,
  1.211226e-09, 6.567351e-10, 4.216705e-08, 1.287376e-07, 1.285559e-06, 
    2.057107e-06, 2.635822e-06, 5.445978e-08, 7.209583e-09, 4.07714e-09, 
    4.947933e-08, 5.309445e-08, 2.310519e-08, 2.318852e-08, 1.382801e-08,
  1.924112e-07, 7.441501e-09, 2.528219e-08, 2.063192e-07, 1.237195e-07, 
    5.604829e-06, 3.339775e-09, 7.156113e-09, 1.126553e-08, 2.37593e-08, 
    3.302084e-07, 8.14128e-07, 3.571314e-07, 1.380583e-07, 2.320957e-07,
  1.046182e-06, 2.093312e-06, 8.874892e-06, 3.484608e-06, 5.239419e-06, 
    6.731432e-06, 8.07778e-09, 9.278763e-09, 1.162178e-08, 3.319263e-07, 
    1.935211e-06, 2.737787e-06, 1.462927e-06, 3.045065e-06, 1.602073e-05,
  1.140793e-07, 3.237306e-06, 1.232771e-05, 1.503482e-05, 6.939412e-06, 
    4.180621e-06, 6.864462e-08, 2.570165e-08, 1.770266e-07, 2.115008e-05, 
    9.823993e-06, 7.689488e-06, 1.997135e-06, 1.452887e-05, 5.820574e-05,
  1.10289e-10, 1.280591e-07, 3.977923e-07, 2.331404e-06, 6.085756e-06, 
    1.578952e-06, 1.170077e-07, 2.289303e-07, 1.037373e-05, 6.275649e-05, 
    3.168913e-05, 8.702325e-06, 6.613288e-06, 2.813808e-05, 8.043232e-05,
  3.668079e-06, 1.110386e-05, 4.291359e-06, 1.063113e-05, 1.600855e-05, 
    1.995693e-05, 2.30992e-05, 6.406284e-06, 1.836385e-05, 2.481245e-05, 
    3.166357e-05, 1.326614e-05, 1.237206e-05, 1.509007e-05, 9.598474e-06,
  4.114837e-06, 3.17422e-06, 5.957034e-06, 1.314255e-05, 1.345758e-05, 
    1.429714e-05, 1.344575e-05, 2.244266e-05, 2.925586e-05, 2.412163e-05, 
    9.134072e-06, 1.299201e-05, 1.188981e-05, 7.29505e-06, 5.051004e-06,
  6.864109e-07, 1.07602e-06, 2.693393e-06, 6.70224e-06, 1.691038e-05, 
    2.267418e-05, 2.118468e-05, 1.945156e-05, 1.171686e-05, 8.901116e-06, 
    8.892091e-06, 7.429004e-06, 2.799351e-06, 3.074177e-06, 3.020495e-06,
  2.355513e-08, 2.404563e-07, 3.132042e-06, 7.12847e-06, 1.315908e-05, 
    1.609078e-05, 1.261546e-05, 7.547921e-06, 5.679726e-06, 5.518181e-06, 
    3.116588e-06, 1.640573e-06, 1.63306e-06, 1.993843e-06, 1.782424e-06,
  1.972205e-08, 2.255589e-07, 1.371503e-06, 4.455299e-06, 6.896581e-06, 
    8.037319e-06, 6.526981e-06, 5.536706e-06, 5.703055e-06, 1.868937e-06, 
    7.460667e-07, 8.144313e-07, 2.166256e-06, 1.646226e-06, 2.400176e-06,
  8.235112e-12, 5.068681e-08, 3.795826e-07, 9.115474e-07, 1.236084e-06, 
    3.611988e-06, 4.141466e-06, 3.31375e-06, 2.054315e-06, 1.053194e-06, 
    4.402325e-07, 3.049432e-06, 1.0866e-06, 2.985322e-06, 6.029951e-06,
  1.971716e-13, 3.603792e-09, 1.087273e-08, 4.328349e-08, 5.40467e-06, 
    4.302779e-06, 7.468754e-08, 4.263404e-07, 1.890361e-07, 3.416412e-07, 
    3.614404e-07, 2.822878e-06, 3.93712e-06, 7.200482e-06, 1.12241e-05,
  3.907556e-07, 8.878831e-07, 2.056246e-09, 2.619178e-08, 2.143062e-05, 
    1.911128e-06, 2.167644e-07, 5.722187e-07, 2.479077e-07, 3.894898e-09, 
    2.953642e-06, 8.951373e-07, 4.019712e-06, 9.218511e-06, 1.016202e-05,
  4.374674e-13, 9.804545e-06, 1.079113e-05, 2.145275e-05, 2.665723e-05, 
    2.727156e-05, 9.670729e-06, 2.268801e-07, 5.675734e-09, 3.859602e-10, 
    5.8735e-06, 8.564388e-06, 3.225066e-06, 5.428793e-06, 5.083873e-06,
  2.328138e-11, 3.510936e-09, 3.519476e-06, 5.426526e-06, 1.079112e-05, 
    1.267931e-05, 5.141582e-06, 4.993012e-09, 7.477041e-10, 3.617449e-06, 
    5.543448e-06, 2.804491e-06, 1.299765e-05, 5.71912e-06, 5.229078e-06,
  2.568067e-05, 3.244695e-05, 3.971667e-05, 6.352551e-05, 6.791102e-05, 
    7.223697e-05, 0.0001034767, 0.0001291768, 0.000133684, 0.0001070496, 
    7.578664e-05, 8.676971e-05, 0.0001006687, 7.940246e-05, 6.690876e-05,
  4.629446e-05, 4.559605e-05, 5.134456e-05, 5.781853e-05, 8.355834e-05, 
    8.358048e-05, 0.0001060774, 0.0001107085, 8.314167e-05, 5.453472e-05, 
    4.978653e-05, 4.066608e-05, 0.0001306344, 0.0001645318, 0.0001091689,
  6.152307e-05, 5.26597e-05, 6.482226e-05, 6.034439e-05, 6.061237e-05, 
    7.922239e-05, 6.065077e-05, 5.229222e-05, 3.842298e-05, 2.153e-05, 
    2.297443e-05, 0.0001787916, 0.0003032418, 0.0002184439, 5.385354e-05,
  5.273195e-05, 5.155441e-05, 5.02169e-05, 4.992313e-05, 4.932197e-05, 
    3.125469e-05, 3.009964e-05, 1.729162e-05, 1.485667e-05, 4.900625e-05, 
    0.0001693426, 0.0002776366, 0.0002119767, 1.174684e-05, 1.506688e-06,
  3.616909e-05, 5.27151e-05, 3.524146e-05, 2.917684e-05, 1.596993e-05, 
    1.584079e-05, 2.286724e-05, 3.093862e-05, 6.847189e-05, 0.0001466899, 
    0.0001686397, 8.795095e-05, 4.038459e-06, 1.217389e-06, 7.780633e-07,
  2.330507e-05, 4.260332e-05, 2.348012e-05, 4.151028e-05, 1.758259e-05, 
    1.898204e-05, 6.989131e-05, 7.975433e-05, 9.597645e-05, 6.976119e-05, 
    1.551555e-05, 1.872382e-06, 5.764417e-07, 1.704942e-07, 2.197834e-07,
  1.796203e-05, 4.416068e-05, 5.211481e-05, 4.502968e-05, 2.745111e-05, 
    5.76645e-05, 5.548801e-05, 5.322732e-05, 3.013406e-05, 6.839885e-06, 
    1.616375e-06, 7.136761e-07, 2.320561e-07, 1.915689e-07, 8.567e-08,
  2.5913e-05, 3.16751e-05, 3.84288e-05, 3.851877e-05, 3.10274e-05, 
    5.52314e-05, 4.423518e-05, 2.615896e-05, 2.690653e-05, 5.214733e-07, 
    2.853334e-07, 1.226361e-07, 5.27182e-08, 4.709748e-08, 9.566582e-08,
  1.878221e-05, 2.041322e-05, 2.298464e-05, 2.02357e-05, 2.027419e-05, 
    2.20067e-05, 6.409099e-06, 1.16875e-05, 9.747504e-08, 7.489514e-08, 
    1.555873e-07, 7.952475e-08, 1.575284e-08, 8.655397e-07, 3.055284e-06,
  1.509881e-05, 1.702319e-05, 2.013606e-05, 1.033976e-05, 2.610255e-05, 
    2.004682e-05, 1.949435e-05, 2.272778e-05, 3.582797e-05, 4.068904e-08, 
    7.046387e-08, 1.961204e-08, 1.477136e-08, 4.849488e-07, 5.898214e-07,
  5.163754e-05, 5.220966e-05, 4.776478e-05, 5.429058e-05, 4.368814e-05, 
    4.837239e-05, 5.355379e-05, 5.466137e-05, 5.395507e-05, 6.974964e-05, 
    7.104505e-05, 7.437626e-05, 0.0001072274, 0.0002775459, 0.0005022784,
  4.61314e-05, 4.574814e-05, 4.625182e-05, 5.065527e-05, 5.305844e-05, 
    5.310098e-05, 5.486339e-05, 6.203431e-05, 6.797541e-05, 7.868002e-05, 
    7.144333e-05, 8.19644e-05, 0.0001820318, 0.0003877467, 0.0004799826,
  3.598186e-05, 3.014207e-05, 4.195402e-05, 4.555515e-05, 5.477922e-05, 
    5.960823e-05, 6.899185e-05, 6.33657e-05, 6.124807e-05, 5.958683e-05, 
    8.51779e-05, 0.0001190033, 0.0002307521, 0.0002959093, 0.0002020193,
  1.725121e-05, 2.414115e-05, 2.675601e-05, 3.15928e-05, 4.570584e-05, 
    3.695678e-05, 3.767383e-05, 5.167543e-05, 5.300556e-05, 6.406201e-05, 
    7.785478e-05, 0.0001137333, 0.0001414836, 0.0001085957, 8.880925e-05,
  2.610167e-06, 6.223133e-06, 1.252486e-05, 1.865403e-05, 2.542784e-05, 
    2.274727e-05, 3.162866e-05, 2.751744e-05, 3.590317e-05, 5.641811e-05, 
    6.628022e-05, 7.127746e-05, 8.199436e-05, 6.507872e-05, 5.960781e-05,
  2.994307e-07, 1.599414e-06, 3.162758e-06, 4.60423e-06, 6.011998e-06, 
    9.853375e-06, 9.849001e-06, 2.352236e-05, 3.974063e-05, 5.274383e-05, 
    3.740653e-05, 3.527777e-05, 3.227833e-05, 2.596971e-05, 2.993102e-05,
  9.490445e-08, 2.456733e-08, 3.613989e-07, 8.177991e-07, 1.487878e-06, 
    3.712144e-06, 6.294709e-06, 1.454857e-05, 2.936381e-05, 4.258343e-05, 
    2.241425e-05, 2.059005e-05, 2.053665e-05, 1.594969e-05, 2.314342e-05,
  5.499689e-09, 4.65397e-09, 4.405656e-08, 1.427638e-07, 9.365333e-07, 
    3.590439e-06, 1.303306e-05, 1.000374e-05, 2.567356e-05, 2.315452e-05, 
    1.864704e-05, 1.969967e-05, 1.230615e-05, 1.652693e-05, 1.264442e-05,
  1.48299e-08, 1.214423e-09, 2.563875e-07, 8.244759e-07, 3.296743e-06, 
    5.005934e-06, 9.70289e-06, 1.256716e-05, 1.04461e-05, 1.116593e-05, 
    4.031647e-06, 1.485832e-05, 3.414071e-06, 5.376376e-06, 3.897893e-06,
  9.053549e-08, 1.131768e-08, 3.5037e-07, 3.377942e-06, 4.706167e-06, 
    6.827085e-06, 1.260572e-05, 1.013897e-05, 8.281475e-06, 1.553956e-05, 
    1.583108e-05, 2.11175e-05, 1.188307e-05, 9.795412e-06, 4.059583e-06,
  7.844037e-06, 9.612505e-06, 1.612049e-05, 2.957114e-05, 4.089591e-05, 
    8.018324e-05, 0.0001974158, 0.0002444626, 0.0001622799, 0.0001167997, 
    0.0001154394, 9.419167e-05, 6.816745e-05, 0.0001308714, 7.659344e-05,
  4.316194e-06, 4.202023e-06, 1.000956e-05, 1.406719e-05, 2.279619e-05, 
    2.223921e-05, 4.559687e-05, 0.0001138648, 0.000194907, 0.000204737, 
    0.0002366781, 0.0001491987, 0.0001232304, 0.000100872, 0.0001103084,
  1.378731e-06, 2.286456e-06, 5.485682e-06, 7.4086e-06, 4.594268e-06, 
    1.101373e-05, 2.152126e-05, 3.006461e-05, 4.965315e-05, 0.0001205272, 
    0.0001246969, 0.0001115828, 9.887251e-05, 0.0001161206, 0.0001547299,
  1.908027e-07, 5.052478e-07, 9.439339e-07, 1.843225e-06, 1.721732e-06, 
    7.751546e-06, 1.371158e-05, 1.731765e-05, 2.395339e-05, 2.796805e-05, 
    1.95246e-05, 6.681204e-05, 4.473063e-05, 3.467158e-05, 5.800661e-05,
  6.884274e-08, 2.799103e-09, 3.750906e-07, 7.887855e-07, 9.16045e-07, 
    2.167459e-06, 6.660605e-06, 1.095474e-05, 1.135655e-05, 1.03715e-05, 
    6.798223e-06, 1.048766e-05, 3.093999e-05, 3.744283e-05, 3.481708e-05,
  4.341947e-10, 2.328982e-08, 1.311812e-07, 6.982406e-07, 7.516379e-07, 
    1.810514e-06, 4.006093e-06, 4.760187e-06, 4.800949e-06, 6.670092e-06, 
    6.394754e-06, 8.420844e-06, 7.63659e-06, 8.750023e-06, 1.845531e-05,
  8.509597e-13, 8.156958e-12, 2.978859e-07, 4.79384e-07, 2.122288e-07, 
    9.703851e-07, 2.196695e-06, 2.473301e-06, 2.464788e-06, 4.733588e-06, 
    4.421416e-06, 3.327005e-06, 6.042928e-06, 4.504764e-06, 1.103562e-05,
  4.195343e-11, 4.392931e-09, 8.482156e-08, 1.665015e-07, 7.834885e-07, 
    6.757808e-07, 6.948463e-07, 9.213099e-07, 1.80468e-06, 2.458094e-06, 
    1.780544e-06, 1.915445e-06, 3.077705e-06, 4.52367e-06, 8.161228e-06,
  7.358255e-10, 1.410812e-09, 3.042247e-08, 5.547865e-07, 7.975836e-07, 
    8.962774e-07, 1.115349e-06, 9.251801e-07, 7.288984e-07, 1.168583e-06, 
    1.570111e-06, 1.520878e-06, 2.208847e-06, 2.758866e-06, 3.104617e-06,
  3.127166e-10, 3.141933e-10, 5.768321e-08, 2.330474e-07, 8.270378e-07, 
    1.092188e-06, 8.851677e-07, 1.790224e-06, 1.64366e-06, 1.647598e-06, 
    6.418299e-07, 1.64416e-06, 1.571199e-06, 1.032758e-06, 2.895941e-06,
  2.357052e-07, 2.703086e-07, 7.457343e-07, 2.594956e-07, 7.602292e-07, 
    7.973055e-06, 4.165926e-05, 5.113052e-05, 3.580314e-05, 2.309012e-05, 
    1.544486e-05, 7.135652e-06, 3.729604e-06, 5.295403e-06, 1.081221e-05,
  1.586225e-07, 1.48718e-07, 1.943752e-07, 5.39009e-07, 1.731093e-07, 
    9.694579e-08, 9.045422e-07, 1.266191e-05, 4.631019e-05, 6.039302e-05, 
    5.971835e-05, 1.510749e-05, 5.646191e-06, 4.074991e-06, 5.65087e-06,
  7.892437e-08, 6.470254e-08, 5.11272e-08, 1.737306e-07, 2.476108e-07, 
    5.384281e-07, 2.561413e-08, 4.67692e-08, 3.266152e-06, 3.174475e-05, 
    3.524578e-05, 2.497925e-05, 7.250619e-05, 1.827639e-05, 2.184503e-05,
  4.902514e-08, 2.49505e-08, 2.993324e-08, 6.379103e-08, 2.582046e-07, 
    3.389218e-07, 7.489464e-08, 8.955008e-08, 3.170092e-07, 7.490494e-07, 
    2.602487e-06, 3.366405e-05, 3.634531e-05, 5.884076e-06, 3.821353e-05,
  1.553179e-08, 2.576288e-08, 3.529836e-08, 1.739305e-07, 1.745248e-07, 
    1.940676e-07, 3.863537e-07, 1.514836e-07, 5.864852e-07, 4.100215e-07, 
    5.192738e-07, 1.881874e-06, 1.242553e-05, 1.765101e-05, 5.000814e-05,
  1.408609e-08, 6.319929e-09, 1.47834e-08, 1.221638e-08, 1.755498e-07, 
    6.618606e-07, 7.315342e-07, 8.508778e-07, 2.088421e-07, 7.06862e-07, 
    3.322074e-08, 1.186932e-06, 2.966554e-06, 6.906964e-06, 1.42211e-05,
  8.245562e-09, 4.017384e-09, 1.508183e-09, 1.23329e-08, 1.213764e-07, 
    3.039593e-07, 6.394767e-07, 4.3009e-07, 2.613235e-07, 5.037928e-07, 
    1.680644e-07, 4.133046e-07, 1.647595e-06, 3.258722e-06, 8.482778e-06,
  3.471368e-09, 9.813092e-09, 4.944831e-09, 4.550854e-09, 2.800202e-07, 
    7.220087e-07, 3.132142e-07, 9.228758e-07, 1.20835e-06, 1.562686e-06, 
    8.172483e-07, 6.431587e-07, 4.180965e-07, 6.544272e-07, 3.492058e-06,
  2.602656e-09, 4.033721e-09, 8.440077e-08, 9.001204e-07, 1.612299e-06, 
    3.537832e-06, 1.827281e-06, 1.273823e-06, 3.948207e-06, 2.969476e-06, 
    3.043174e-06, 2.475044e-06, 3.031369e-06, 2.681873e-06, 2.946447e-06,
  2.152489e-09, 2.159188e-10, 2.155983e-07, 8.602544e-07, 1.568745e-06, 
    3.911495e-06, 4.011791e-06, 4.467357e-06, 4.124401e-06, 1.602462e-06, 
    4.111431e-06, 3.632403e-06, 4.2099e-06, 2.770698e-06, 2.958067e-06,
  7.291227e-06, 1.649069e-06, 1.37113e-06, 3.039515e-06, 5.465977e-06, 
    8.401908e-06, 1.002834e-05, 1.357182e-05, 1.050042e-05, 2.522635e-05, 
    2.908386e-05, 1.911647e-05, 2.032474e-05, 2.132303e-05, 4.275963e-05,
  6.239534e-06, 4.917398e-06, 2.810487e-06, 4.958638e-06, 5.263253e-06, 
    5.21971e-06, 7.111906e-06, 1.189778e-05, 1.459728e-05, 1.347906e-05, 
    2.34281e-05, 2.498097e-05, 1.693184e-05, 3.305166e-05, 3.288344e-05,
  4.618796e-06, 4.281968e-06, 4.800385e-06, 4.915221e-06, 4.426804e-06, 
    5.555708e-06, 5.117941e-06, 7.084046e-06, 7.402748e-06, 6.692881e-06, 
    1.156187e-05, 1.034109e-05, 1.146287e-05, 1.853499e-05, 2.033019e-05,
  1.277773e-06, 1.485797e-06, 2.493029e-06, 3.773473e-06, 4.4979e-06, 
    4.11468e-06, 5.817019e-06, 5.827912e-06, 4.194645e-06, 3.978327e-06, 
    3.974165e-06, 3.718328e-06, 2.946284e-06, 4.38549e-06, 7.675879e-06,
  7.499731e-07, 8.104073e-07, 8.239689e-07, 1.228739e-06, 2.663845e-06, 
    2.200653e-06, 2.851863e-06, 2.420417e-06, 3.874962e-06, 4.2036e-06, 
    3.239179e-06, 3.010392e-06, 3.256393e-06, 2.63382e-06, 1.411635e-06,
  2.239888e-07, 1.560485e-07, 1.569984e-07, 2.66506e-07, 2.304019e-07, 
    5.093967e-07, 1.549194e-06, 3.026359e-06, 7.00841e-06, 1.0155e-05, 
    1.016485e-05, 1.099809e-05, 1.145707e-05, 1.427493e-05, 1.240249e-05,
  1.188372e-07, 7.734611e-08, 8.494975e-08, 3.190795e-08, 5.654249e-08, 
    9.379052e-07, 2.124083e-06, 9.82268e-06, 1.444267e-05, 1.971383e-05, 
    1.761603e-05, 1.31635e-05, 1.35343e-05, 1.91998e-05, 2.183843e-05,
  4.305167e-08, 1.665696e-08, 6.768928e-09, 7.49601e-09, 3.363816e-08, 
    1.951299e-07, 1.25521e-06, 2.808784e-06, 6.32623e-06, 8.341095e-06, 
    6.182853e-06, 8.128954e-06, 7.348294e-06, 6.292498e-06, 7.250143e-06,
  2.605221e-08, 8.309494e-09, 4.422274e-09, 2.943863e-08, 5.324742e-07, 
    2.811612e-07, 4.806218e-07, 1.712353e-06, 1.021721e-06, 4.630499e-07, 
    4.745064e-07, 1.365829e-07, 5.468718e-07, 6.97202e-07, 1.34928e-06,
  1.017093e-08, 1.592009e-08, 8.749996e-09, 9.24816e-08, 8.363752e-07, 
    4.996058e-07, 2.00008e-06, 3.063812e-06, 2.361289e-06, 7.218437e-07, 
    5.616627e-07, 1.809145e-06, 6.156234e-07, 3.321528e-06, 5.83092e-06,
  2.814405e-07, 2.423904e-07, 2.873991e-07, 3.326744e-07, 6.564405e-07, 
    6.414003e-07, 1.240548e-06, 2.91154e-06, 4.96676e-06, 6.436413e-06, 
    9.825545e-06, 1.064066e-05, 1.542241e-05, 2.211081e-05, 1.841949e-05,
  7.838411e-07, 4.072512e-07, 1.985083e-08, 1.931051e-07, 3.257224e-07, 
    7.066184e-07, 1.564219e-06, 1.774436e-06, 2.341809e-06, 3.28172e-06, 
    3.903144e-06, 3.6598e-06, 6.896062e-06, 8.762913e-06, 1.185304e-05,
  9.870396e-07, 1.443783e-06, 1.540456e-06, 1.307074e-06, 1.351314e-06, 
    9.936579e-07, 1.555464e-06, 2.089218e-06, 2.58272e-06, 2.681808e-06, 
    3.0754e-06, 1.989061e-06, 4.03831e-06, 4.901227e-06, 6.877427e-06,
  1.474042e-06, 2.056895e-06, 1.777404e-06, 1.390004e-06, 1.185557e-06, 
    2.162851e-06, 2.028741e-06, 2.231896e-06, 3.29011e-06, 2.103386e-06, 
    2.895959e-06, 2.910579e-06, 3.39284e-06, 3.866565e-06, 3.811203e-06,
  1.552536e-06, 1.16241e-06, 1.362525e-06, 1.514961e-06, 2.060742e-06, 
    3.033078e-06, 4.658381e-06, 4.67032e-06, 4.882166e-06, 4.611429e-06, 
    4.17018e-06, 3.071126e-06, 2.594542e-06, 3.652023e-06, 2.886973e-06,
  1.150193e-06, 2.170266e-06, 2.078768e-06, 1.817833e-06, 3.175757e-06, 
    5.089667e-06, 7.179272e-06, 6.71716e-06, 6.609329e-06, 6.067802e-06, 
    5.468123e-06, 4.750925e-06, 4.033542e-06, 4.389641e-06, 3.512736e-06,
  1.126851e-06, 1.324415e-06, 1.308846e-06, 3.255155e-06, 3.375678e-06, 
    4.818316e-06, 5.399722e-06, 6.659578e-06, 6.517089e-06, 6.311691e-06, 
    9.124672e-06, 1.017963e-05, 1.062184e-05, 1.313904e-05, 1.108681e-05,
  2.829219e-06, 4.15068e-06, 4.400317e-06, 4.944157e-06, 2.929222e-06, 
    5.927254e-06, 3.282142e-06, 3.714301e-06, 7.419117e-06, 9.071928e-06, 
    1.193122e-05, 1.525108e-05, 2.013587e-05, 2.798729e-05, 2.938203e-05,
  3.276855e-06, 4.628043e-06, 3.617913e-06, 5.310936e-06, 9.541994e-06, 
    8.698929e-06, 4.904795e-06, 6.885012e-06, 1.327112e-05, 1.589881e-05, 
    2.237328e-05, 1.916953e-05, 1.928972e-05, 2.750664e-05, 3.458189e-05,
  3.25604e-06, 5.081836e-06, 6.136578e-06, 6.910904e-06, 7.165225e-06, 
    7.022802e-06, 8.301266e-06, 1.017607e-05, 1.318764e-05, 1.224263e-05, 
    8.17693e-06, 9.329724e-06, 2.52513e-05, 2.346219e-05, 2.51639e-05,
  1.384889e-06, 3.416478e-07, 2.099453e-06, 5.073982e-06, 5.978481e-06, 
    5.370668e-06, 5.088131e-06, 2.650982e-06, 3.764502e-06, 3.537277e-06, 
    6.859159e-06, 9.571817e-06, 1.204376e-05, 1.049991e-05, 8.962408e-06,
  2.39746e-06, 9.573532e-07, 7.512988e-07, 5.355615e-06, 5.327955e-06, 
    6.433693e-06, 5.13182e-06, 2.93138e-06, 2.082658e-06, 1.851042e-06, 
    4.055438e-06, 6.583465e-06, 1.017604e-05, 8.127478e-06, 8.818794e-06,
  3.694341e-06, 3.24466e-06, 6.50482e-07, 4.929636e-06, 5.542786e-06, 
    5.619983e-06, 5.643511e-06, 4.782701e-06, 1.677833e-06, 1.551698e-06, 
    1.607931e-06, 4.002512e-06, 3.456139e-06, 5.220417e-06, 1.109085e-05,
  2.82585e-06, 4.835667e-06, 2.574098e-06, 3.474367e-06, 6.416735e-06, 
    6.11903e-06, 5.203577e-06, 5.129768e-06, 2.859966e-06, 1.72402e-06, 
    1.573436e-06, 2.150099e-06, 3.673407e-06, 4.761645e-06, 5.696052e-06,
  5.649486e-06, 5.073679e-06, 6.188491e-06, 2.655487e-06, 2.683676e-06, 
    5.422622e-06, 6.040386e-06, 5.971067e-06, 3.202366e-06, 2.854239e-06, 
    1.879449e-06, 1.583402e-06, 2.687395e-06, 3.990564e-06, 3.870395e-06,
  8.117313e-06, 1.029248e-05, 5.756411e-06, 5.201197e-06, 1.434434e-06, 
    6.745777e-06, 8.29925e-06, 1.010373e-05, 7.276084e-06, 4.97777e-06, 
    2.429482e-06, 2.673053e-06, 2.891808e-06, 3.543063e-06, 5.04912e-06,
  3.274519e-05, 1.440858e-05, 4.970041e-06, 4.188093e-06, 4.804257e-06, 
    6.367652e-07, 8.24025e-06, 8.413665e-06, 8.540045e-06, 6.827651e-06, 
    4.664317e-06, 4.064684e-06, 4.628789e-06, 3.51785e-06, 4.795294e-06,
  6.24155e-05, 2.793057e-05, 8.946718e-06, 1.050057e-05, 5.562736e-06, 
    4.027935e-06, 1.827575e-06, 4.912226e-06, 1.126599e-05, 8.687986e-06, 
    5.932359e-06, 4.393632e-06, 5.014417e-06, 4.530566e-06, 4.957215e-06,
  6.510669e-05, 6.4814e-05, 3.963462e-05, 1.329084e-05, 8.561316e-06, 
    1.254176e-05, 5.757972e-06, 3.085776e-06, 2.363704e-06, 6.398842e-06, 
    6.298271e-06, 6.337384e-06, 6.670532e-06, 6.290919e-06, 5.384605e-06,
  2.63548e-05, 6.331791e-05, 7.629478e-05, 3.939563e-05, 1.112025e-05, 
    6.674799e-06, 1.557396e-05, 4.026107e-06, 1.284401e-06, 3.455131e-06, 
    5.996567e-06, 7.513597e-06, 4.278338e-06, 4.514377e-06, 4.824727e-06,
  7.715227e-05, 6.185432e-05, 4.31136e-05, 2.364694e-05, 1.537312e-05, 
    1.174957e-05, 8.957566e-06, 1.124947e-05, 1.252827e-05, 1.178454e-05, 
    1.027078e-05, 9.987402e-06, 1.307581e-05, 1.365141e-05, 1.434159e-05,
  4.13201e-05, 4.058888e-05, 2.758712e-05, 1.917062e-05, 1.622515e-05, 
    1.552034e-05, 1.063444e-05, 1.005418e-05, 1.178978e-05, 1.315662e-05, 
    1.263652e-05, 1.094542e-05, 1.032387e-05, 1.40299e-05, 1.350568e-05,
  5.61008e-05, 2.828736e-05, 1.418096e-05, 1.247456e-05, 1.354806e-05, 
    1.590294e-05, 1.119298e-05, 8.634195e-06, 1.084168e-05, 1.15605e-05, 
    1.244828e-05, 1.062368e-05, 1.103971e-05, 9.874706e-06, 8.616951e-06,
  3.445094e-05, 1.865377e-05, 7.564589e-06, 6.714574e-06, 8.317059e-06, 
    1.227292e-05, 1.325117e-05, 7.409737e-06, 7.17189e-06, 1.052219e-05, 
    9.570492e-06, 1.040166e-05, 1.071305e-05, 9.230496e-06, 8.432482e-06,
  1.654444e-05, 1.583117e-05, 6.150631e-06, 3.741558e-06, 5.746303e-06, 
    1.141521e-05, 1.312122e-05, 6.236294e-06, 8.001904e-06, 7.977299e-06, 
    8.016498e-06, 8.118724e-06, 1.278368e-05, 1.199846e-05, 1.017106e-05,
  3.393254e-05, 1.758698e-05, 8.484354e-06, 3.417485e-06, 1.471605e-06, 
    9.88177e-06, 1.576651e-05, 7.300576e-06, 7.47788e-06, 1.043659e-05, 
    9.708442e-06, 8.979543e-06, 1.105577e-05, 1.162563e-05, 1.014139e-05,
  5.959867e-05, 1.538405e-05, 2.091834e-05, 6.746766e-06, 1.358828e-05, 
    1.511098e-05, 2.245188e-05, 1.002738e-05, 7.576718e-06, 1.14505e-05, 
    9.42501e-06, 9.978735e-06, 1.102899e-05, 9.779267e-06, 8.949185e-06,
  6.547292e-05, 6.390736e-05, 5.1732e-05, 3.981144e-05, 5.95893e-05, 
    9.490178e-05, 5.017811e-05, 1.949934e-05, 5.11868e-06, 8.966514e-06, 
    1.002757e-05, 1.110541e-05, 8.650268e-06, 1.199434e-05, 9.826598e-06,
  1.750067e-05, 3.693833e-05, 4.375479e-05, 4.354335e-05, 5.934182e-05, 
    0.0001182608, 0.0001046429, 2.364557e-05, 5.009222e-06, 7.144337e-06, 
    1.024271e-05, 1.066718e-05, 1.129305e-05, 1.130847e-05, 1.182132e-05,
  6.169296e-06, 1.436287e-05, 2.150275e-05, 3.42464e-05, 5.447831e-05, 
    0.0001081717, 0.0001896899, 6.388059e-05, 5.313048e-06, 5.167168e-06, 
    6.787965e-06, 1.023328e-05, 1.033264e-05, 1.076493e-05, 1.315297e-05,
  3.160189e-05, 3.599218e-05, 3.622488e-05, 3.044859e-05, 2.906896e-05, 
    4.384352e-05, 8.943214e-05, 0.0001329591, 0.0001674242, 0.0001765619, 
    0.000172393, 0.000153767, 0.0001296452, 0.0001221976, 0.0001067118,
  1.573773e-05, 9.919987e-06, 1.035979e-05, 1.073764e-05, 1.332879e-05, 
    1.538123e-05, 6.676636e-05, 0.0001007385, 0.0001374915, 0.0001554752, 
    0.0001478161, 0.0001370433, 0.0001168987, 0.0001158784, 0.0001144808,
  4.4324e-06, 4.361006e-06, 2.109575e-06, 5.042216e-06, 3.086848e-06, 
    5.159165e-06, 3.200486e-05, 7.723127e-05, 0.0001035336, 0.000110295, 
    0.0001013562, 8.68224e-05, 8.452905e-05, 7.715218e-05, 7.775052e-05,
  7.29654e-08, 5.150483e-07, 7.800752e-07, 3.922244e-06, 1.473961e-06, 
    3.970023e-06, 2.262353e-05, 5.083425e-05, 6.858174e-05, 7.515007e-05, 
    6.58978e-05, 5.977216e-05, 5.234406e-05, 5.921191e-05, 5.858134e-05,
  8.801447e-08, 5.831743e-07, 1.110993e-06, 2.374824e-06, 4.825359e-06, 
    1.026281e-05, 2.023022e-05, 3.769187e-05, 4.395334e-05, 5.20422e-05, 
    5.724725e-05, 5.813734e-05, 6.880522e-05, 9.182346e-05, 0.0001264347,
  2.967036e-05, 1.661184e-05, 1.660852e-06, 3.595517e-06, 4.468467e-06, 
    2.945066e-06, 7.014851e-06, 2.210245e-05, 3.253666e-05, 4.504832e-05, 
    5.078537e-05, 5.73669e-05, 6.649959e-05, 8.792663e-05, 0.0001212513,
  2.016237e-05, 2.178104e-05, 1.047469e-05, 8.513135e-07, 4.306176e-07, 
    3.757908e-07, 1.033634e-05, 1.465737e-05, 2.828109e-05, 3.230509e-05, 
    2.753157e-05, 2.957836e-05, 2.6334e-05, 2.460156e-05, 2.209369e-05,
  0.0001004745, 0.0001038296, 9.472567e-06, 6.904097e-05, 8.093132e-05, 
    4.408589e-05, 9.39342e-06, 2.718577e-05, 2.646144e-05, 1.186656e-05, 
    5.348813e-06, 5.184496e-06, 4.92195e-06, 2.289346e-06, 3.20718e-06,
  0.0001910923, 0.0002170951, 0.0001701015, 0.0001103363, 6.969263e-05, 
    3.5583e-05, 2.056253e-05, 7.508799e-05, 1.115554e-05, 4.242812e-07, 
    3.344653e-07, 2.621203e-07, 4.473709e-07, 1.30998e-06, 2.827226e-06,
  0.0001509041, 0.0002771344, 0.0001675782, 8.05158e-05, 3.943613e-05, 
    3.152575e-05, 5.340769e-05, 0.0001794951, 8.409195e-05, 3.024874e-06, 
    3.351611e-08, 3.522077e-08, 7.801038e-08, 8.886215e-07, 3.111022e-06,
  9.059854e-06, 1.51505e-05, 1.635802e-05, 4.697828e-05, 5.310598e-05, 
    4.255223e-05, 3.639759e-05, 6.012702e-05, 3.92443e-05, 7.394062e-05, 
    6.895795e-05, 1.951345e-05, 2.21421e-05, 3.193992e-05, 4.215202e-05,
  1.913154e-05, 1.325125e-05, 2.432153e-05, 4.27914e-05, 2.877116e-05, 
    3.681135e-05, 4.681623e-05, 2.370332e-05, 2.059328e-05, 1.22572e-05, 
    1.266951e-05, 1.64971e-06, 6.052256e-06, 7.477173e-06, 9.12557e-06,
  1.79281e-05, 2.016768e-05, 3.244247e-05, 3.085758e-05, 1.498914e-05, 
    2.061264e-05, 2.102265e-05, 2.46174e-05, 2.512793e-05, 1.618824e-05, 
    7.24549e-06, 6.912034e-06, 5.453876e-06, 6.161337e-06, 6.551453e-06,
  1.029294e-05, 5.387291e-05, 5.822358e-05, 3.206469e-05, 2.975704e-05, 
    2.683004e-05, 3.059373e-05, 2.041772e-05, 2.43622e-05, 2.440206e-05, 
    1.579943e-05, 1.25681e-05, 5.761057e-06, 6.15555e-06, 7.097105e-06,
  7.954746e-06, 1.188895e-05, 4.263168e-05, 0.0001032962, 3.887582e-05, 
    2.561404e-05, 2.129778e-05, 4.444917e-05, 3.870825e-05, 3.645156e-05, 
    2.400105e-05, 1.396772e-05, 4.421043e-06, 4.099737e-06, 1.109212e-05,
  3.929073e-05, 4.712424e-05, 7.565792e-05, 0.0001524707, 5.177225e-05, 
    1.939082e-05, 1.282745e-05, 1.587775e-05, 2.543591e-05, 2.929162e-05, 
    1.923753e-05, 1.565382e-05, 8.824503e-06, 1.442937e-05, 3.34417e-05,
  7.164243e-05, 8.129657e-05, 0.0001572849, 0.0002384761, 0.0001533466, 
    2.780395e-05, 1.163829e-05, 8.78827e-06, 1.110589e-05, 1.935686e-05, 
    1.561661e-05, 8.919512e-06, 9.084897e-06, 2.545401e-05, 4.614257e-05,
  5.709722e-05, 9.133197e-05, 0.0002621713, 0.0003591096, 0.0001945515, 
    7.766862e-05, 1.131732e-05, 3.648042e-06, 4.654406e-06, 7.575183e-06, 
    9.711988e-06, 6.796836e-06, 1.248645e-05, 1.864527e-05, 2.578975e-05,
  4.265649e-05, 0.0001195521, 0.0002599644, 0.0002679195, 0.0001131211, 
    6.181213e-05, 1.463339e-05, 1.898327e-06, 3.270051e-06, 2.205527e-06, 
    4.707432e-06, 7.566926e-06, 9.081574e-06, 5.700656e-06, 3.453625e-06,
  6.076603e-05, 0.0002599942, 0.0002127248, 0.0002118176, 0.000224316, 
    0.0001180985, 0.0001271919, 7.619636e-05, 9.312366e-05, 4.512926e-06, 
    1.977291e-06, 5.825064e-06, 4.875115e-07, 3.363314e-07, 1.890676e-06,
  8.268365e-05, 7.41434e-05, 4.171468e-05, 2.897459e-05, 2.824002e-05, 
    2.15592e-05, 3.11355e-05, 0.0004319482, 0.0006035798, 0.0002709368, 
    0.0002950319, 0.0002262337, 0.0001116667, 6.174127e-05, 6.177814e-05,
  2.104986e-05, 2.771894e-05, 2.182135e-05, 1.722855e-05, 2.581486e-05, 
    1.6006e-05, 0.0001425484, 0.0006099799, 0.000518002, 0.000297768, 
    0.0003415025, 0.0002564731, 0.000149727, 5.735885e-05, 3.757241e-05,
  3.611318e-06, 7.371529e-06, 7.451675e-06, 1.108446e-05, 1.597049e-05, 
    3.314779e-05, 0.0004993524, 0.0007367745, 0.0003606922, 0.0003217453, 
    0.0002872992, 0.0002218515, 0.00014459, 4.534263e-05, 1.398106e-05,
  2.644362e-07, 1.122475e-06, 3.108882e-06, 1.076279e-05, 1.772146e-05, 
    0.0003122384, 0.0007192654, 0.0006275233, 0.0002818374, 0.0002906989, 
    0.0002640109, 0.0001927841, 0.0001189873, 2.319982e-05, 5.835263e-06,
  1.945138e-07, 6.787182e-06, 3.95977e-06, 2.635404e-05, 0.0002328921, 
    0.0006154625, 0.0007003191, 0.0003844146, 0.0002872507, 0.0002649737, 
    0.0002105114, 0.000187764, 9.617864e-05, 7.541512e-06, 4.853186e-06,
  5.678814e-06, 7.811426e-06, 6.28046e-05, 0.0002298914, 0.000483971, 
    0.0006394529, 0.0004631607, 0.0003112151, 0.0002778316, 0.0002388529, 
    0.0002290911, 0.0001826696, 4.970529e-05, 3.191585e-06, 6.286053e-06,
  3.514001e-05, 0.0001046623, 0.0002722912, 0.0004683933, 0.0006083112, 
    0.0005067665, 0.0003111512, 0.0002606743, 0.0002503032, 0.0002742085, 
    0.0002545168, 0.0001233342, 2.155973e-06, 1.786701e-06, 1.005464e-05,
  0.0003361521, 0.0003070914, 0.00064807, 0.0005742497, 0.0005952363, 
    0.0002605124, 0.0002501713, 0.0002429794, 0.000289678, 0.0003222238, 
    0.0001942651, 1.999532e-05, 2.928596e-07, 2.099223e-07, 6.932886e-06,
  0.0004332392, 0.0004916231, 0.0003886796, 0.0004663936, 0.0002343269, 
    0.0002275772, 0.0002492204, 0.0003068745, 0.0003192532, 0.0002354046, 
    4.70999e-05, 1.090078e-07, 1.808378e-07, 7.868636e-08, 3.121225e-07,
  7.857422e-05, 0.000122225, 0.0001306593, 0.0003318865, 0.0003090689, 
    0.0002254853, 0.0003442023, 0.0004664165, 0.0002355398, 6.44355e-05, 
    2.018165e-07, 5.72206e-08, 1.262634e-07, 3.141374e-08, 7.780476e-08,
  4.374917e-05, 6.880429e-05, 5.914761e-05, 5.560604e-05, 5.776184e-05, 
    5.019133e-05, 4.908666e-05, 6.054365e-05, 5.449961e-05, 5.621844e-05, 
    5.830305e-05, 9.110543e-05, 0.0001207419, 0.0001245904, 6.766429e-05,
  2.927697e-05, 4.1927e-05, 4.347128e-05, 3.876286e-05, 4.841014e-05, 
    4.306703e-05, 4.548527e-05, 4.436059e-05, 4.566537e-05, 4.834081e-05, 
    4.905782e-05, 5.324219e-05, 7.925234e-05, 8.359828e-05, 4.823369e-05,
  2.747209e-05, 2.788986e-05, 2.518671e-05, 2.937758e-05, 3.267101e-05, 
    3.578369e-05, 3.48513e-05, 3.902173e-05, 4.100981e-05, 5.094724e-05, 
    5.244892e-05, 4.009734e-05, 5.387362e-05, 6.672009e-05, 4.494984e-05,
  1.526884e-05, 1.296373e-05, 1.482679e-05, 1.682634e-05, 2.16705e-05, 
    2.585782e-05, 2.609082e-05, 2.826929e-05, 3.273777e-05, 4.786886e-05, 
    3.38225e-05, 2.33929e-05, 3.601353e-05, 7.023648e-05, 7.252979e-05,
  8.063891e-06, 8.260901e-06, 9.071866e-06, 1.033811e-05, 1.346861e-05, 
    1.40609e-05, 1.4483e-05, 1.527406e-05, 3.356473e-05, 2.675202e-05, 
    1.340927e-05, 1.380601e-05, 6.348664e-05, 0.0001136399, 0.000108121,
  2.421484e-06, 3.449853e-06, 4.941805e-06, 5.235045e-06, 6.116952e-06, 
    6.431088e-06, 6.097306e-06, 6.210653e-06, 1.561066e-05, 6.072168e-06, 
    9.55877e-06, 5.801411e-05, 0.0001459237, 0.0001675227, 0.0001533066,
  4.667389e-07, 4.755686e-07, 8.918099e-07, 1.446221e-06, 1.230861e-06, 
    1.764563e-06, 1.507303e-06, 2.10354e-06, 1.782157e-06, 4.88975e-06, 
    5.594853e-05, 0.000163167, 0.0002210345, 0.0001882757, 0.0001725149,
  2.64518e-07, 1.119543e-07, 5.642166e-07, 5.648927e-07, 6.944485e-07, 
    5.114661e-07, 3.041004e-07, 6.044174e-07, 5.602284e-07, 3.319719e-05, 
    0.0001538701, 0.0002450565, 0.0002014858, 0.0001799714, 0.000155831,
  3.954809e-06, 3.085109e-06, 1.016133e-06, 1.262579e-06, 7.452625e-07, 
    8.155489e-07, 3.566122e-07, 4.8249e-07, 1.140218e-05, 9.795668e-05, 
    0.0002144937, 0.0002120022, 0.0001881363, 0.0001669517, 0.0001322308,
  5.816636e-06, 3.771048e-06, 2.740694e-06, 1.073545e-06, 4.033016e-07, 
    5.668408e-07, 3.620446e-07, 2.342645e-06, 4.393888e-05, 0.0001230302, 
    0.0001766504, 0.0001824193, 0.0001514037, 0.0001372223, 0.0001635475,
  1.032456e-05, 2.04482e-05, 2.825934e-05, 4.875478e-05, 6.335574e-05, 
    8.057709e-05, 9.69363e-05, 9.96099e-05, 8.536615e-05, 7.259596e-05, 
    6.13815e-05, 6.158074e-05, 5.521208e-05, 6.687313e-05, 9.596159e-05,
  4.604426e-06, 9.186258e-06, 1.667603e-05, 2.536996e-05, 4.155877e-05, 
    5.459489e-05, 6.587798e-05, 7.522947e-05, 7.353364e-05, 7.13464e-05, 
    7.066652e-05, 6.583605e-05, 6.017652e-05, 7.064984e-05, 7.881548e-05,
  1.89316e-06, 2.893355e-06, 6.343808e-06, 1.490126e-05, 1.992439e-05, 
    3.141423e-05, 4.962654e-05, 5.183195e-05, 6.362708e-05, 7.208247e-05, 
    7.541403e-05, 7.759942e-05, 7.572211e-05, 8.066377e-05, 8.70794e-05,
  3.117446e-06, 2.40675e-06, 3.745968e-06, 5.118362e-06, 1.004986e-05, 
    1.46079e-05, 2.16915e-05, 2.838913e-05, 4.655436e-05, 5.551288e-05, 
    7.685507e-05, 6.950867e-05, 7.141797e-05, 7.460701e-05, 8.009513e-05,
  6.385243e-06, 4.711719e-06, 5.000393e-06, 5.413756e-06, 6.843715e-06, 
    8.027656e-06, 1.256178e-05, 1.75731e-05, 2.494139e-05, 3.436803e-05, 
    4.932861e-05, 4.917486e-05, 5.365186e-05, 6.450892e-05, 6.110875e-05,
  6.71611e-06, 5.780438e-06, 6.204821e-06, 6.631049e-06, 6.884511e-06, 
    8.797185e-06, 8.876258e-06, 1.158939e-05, 1.699397e-05, 1.890174e-05, 
    2.493694e-05, 3.113297e-05, 3.411385e-05, 3.849138e-05, 4.328768e-05,
  4.930846e-06, 5.112332e-06, 5.592796e-06, 5.999576e-06, 6.967745e-06, 
    7.589616e-06, 7.769262e-06, 7.936957e-06, 9.417208e-06, 1.270244e-05, 
    1.364487e-05, 1.760856e-05, 2.389981e-05, 3.232162e-05, 2.824446e-05,
  1.750023e-06, 2.183358e-06, 2.889651e-06, 4.053361e-06, 5.964378e-06, 
    5.865852e-06, 5.80034e-06, 5.647369e-06, 5.842393e-06, 7.520127e-06, 
    9.462021e-06, 1.095025e-05, 1.300448e-05, 2.092173e-05, 1.337856e-05,
  9.621281e-07, 5.882723e-07, 1.855684e-06, 3.081794e-06, 3.639328e-06, 
    3.689465e-06, 4.145201e-06, 4.487028e-06, 3.737214e-06, 3.99545e-06, 
    5.372266e-06, 6.920061e-06, 7.436119e-06, 9.933103e-06, 1.037083e-05,
  1.257279e-06, 7.68721e-07, 7.522727e-07, 1.369388e-06, 1.853869e-06, 
    2.288149e-06, 2.713039e-06, 3.142228e-06, 3.506528e-06, 2.383387e-06, 
    2.404684e-06, 3.007131e-06, 3.703394e-06, 5.053276e-06, 4.83355e-06 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
