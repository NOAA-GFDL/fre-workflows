netcdf atmos_diurnal.orog {
dimensions:
	lon = 288 ;
	bnds = 2 ;
	lat = 180 ;
variables:
	double lon(lon) ;
		lon:standard_name = "longitude" ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_E" ;
		lon:axis = "X" ;
		lon:bounds = "lon_bnds" ;
	double lon_bnds(lon, bnds) ;
	double lat(lat) ;
		lat:standard_name = "latitude" ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_N" ;
		lat:axis = "Y" ;
		lat:bounds = "lat_bnds" ;
	double lat_bnds(lat, bnds) ;
	float orog(lat, lon) ;
		orog:standard_name = "surface_altitude" ;
		orog:long_name = "Surface Altitude" ;
		orog:units = "m" ;
		orog:_FillValue = 1.e+20f ;
		orog:missing_value = 1.e+20f ;
		orog:cell_methods = "time: point" ;
		orog:cell_measures = "area: area" ;
		orog:interp_method = "conserve_order1" ;

// global attributes:
		:CDI = "Climate Data Interface version 2.1.1 (https://mpimet.mpg.de/cdi)" ;
		:Conventions = "CF-1.6" ;
		:title = "c96L65_am5f5b8r0_amip" ;
		:associated_files = "area: 19800101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:code_release_version = "2023.01.02" ;
		:git_hash = "8176c2b45079431f2053ec773253938f8aee4828" ;
		:creationtime = "Sat Mar 23 01:57:39 2024" ;
		:hostname = "pp315" ;
		:history = "Sat Mar 23 01:58:18 2024: cdo --history splitname 19800101.atmos_diurnal.nc /home/Chris.Blanton/cylc-run/c96L65_am5f5b8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/share/cycle/19800101T0000Z/split/regrid-xy/288_180.conserve_order2/19800101.atmos_diurnal.\n",
			"fregrid --debug --standard_dimension --input_mosaic C96_mosaic.nc --input_dir /home/Chris.Blanton/cylc-run/c96L65_am5f5b8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/share/cycle/19800101T0000Z/history/native --input_file 19800101.atmos_diurnal --associated_file_dir /home/Chris.Blanton/cylc-run/c96L65_am5f5b8r0_amip__gfdl.ncrc5-intel23-classic__prod-openmp/share/cycle/19800101T0000Z/history/native --interp_method conserve_order2 --remap_file fregrid_remap_file_288_by_180.nc --nlon 288 --nlat 180 --scalar_field sftlf,orog,tas,evspsbl,hfss,pr,prc,z_Ri_025 --output_file 19800101.atmos_diurnal.nc" ;
		:CDO = "Climate Data Operators version 2.1.1 (https://mpimet.mpg.de/cdo)" ;
data:

 lon = 0.625, 1.875, 3.125, 4.375, 5.625, 6.875, 8.125, 9.375, 10.625, 
    11.875, 13.125, 14.375, 15.625, 16.875, 18.125, 19.375, 20.625, 21.875, 
    23.125, 24.375, 25.625, 26.875, 28.125, 29.375, 30.625, 31.875, 33.125, 
    34.375, 35.625, 36.875, 38.125, 39.375, 40.625, 41.875, 43.125, 44.375, 
    45.625, 46.875, 48.125, 49.375, 50.625, 51.875, 53.125, 54.375, 55.625, 
    56.875, 58.125, 59.375, 60.625, 61.875, 63.125, 64.375, 65.625, 66.875, 
    68.125, 69.375, 70.625, 71.875, 73.125, 74.375, 75.625, 76.875, 78.125, 
    79.375, 80.625, 81.875, 83.125, 84.375, 85.625, 86.875, 88.125, 89.375, 
    90.625, 91.875, 93.125, 94.375, 95.625, 96.875, 98.125, 99.375, 100.625, 
    101.875, 103.125, 104.375, 105.625, 106.875, 108.125, 109.375, 110.625, 
    111.875, 113.125, 114.375, 115.625, 116.875, 118.125, 119.375, 120.625, 
    121.875, 123.125, 124.375, 125.625, 126.875, 128.125, 129.375, 130.625, 
    131.875, 133.125, 134.375, 135.625, 136.875, 138.125, 139.375, 140.625, 
    141.875, 143.125, 144.375, 145.625, 146.875, 148.125, 149.375, 150.625, 
    151.875, 153.125, 154.375, 155.625, 156.875, 158.125, 159.375, 160.625, 
    161.875, 163.125, 164.375, 165.625, 166.875, 168.125, 169.375, 170.625, 
    171.875, 173.125, 174.375, 175.625, 176.875, 178.125, 179.375, 180.625, 
    181.875, 183.125, 184.375, 185.625, 186.875, 188.125, 189.375, 190.625, 
    191.875, 193.125, 194.375, 195.625, 196.875, 198.125, 199.375, 200.625, 
    201.875, 203.125, 204.375, 205.625, 206.875, 208.125, 209.375, 210.625, 
    211.875, 213.125, 214.375, 215.625, 216.875, 218.125, 219.375, 220.625, 
    221.875, 223.125, 224.375, 225.625, 226.875, 228.125, 229.375, 230.625, 
    231.875, 233.125, 234.375, 235.625, 236.875, 238.125, 239.375, 240.625, 
    241.875, 243.125, 244.375, 245.625, 246.875, 248.125, 249.375, 250.625, 
    251.875, 253.125, 254.375, 255.625, 256.875, 258.125, 259.375, 260.625, 
    261.875, 263.125, 264.375, 265.625, 266.875, 268.125, 269.375, 270.625, 
    271.875, 273.125, 274.375, 275.625, 276.875, 278.125, 279.375, 280.625, 
    281.875, 283.125, 284.375, 285.625, 286.875, 288.125, 289.375, 290.625, 
    291.875, 293.125, 294.375, 295.625, 296.875, 298.125, 299.375, 300.625, 
    301.875, 303.125, 304.375, 305.625, 306.875, 308.125, 309.375, 310.625, 
    311.875, 313.125, 314.375, 315.625, 316.875, 318.125, 319.375, 320.625, 
    321.875, 323.125, 324.375, 325.625, 326.875, 328.125, 329.375, 330.625, 
    331.875, 333.125, 334.375, 335.625, 336.875, 338.125, 339.375, 340.625, 
    341.875, 343.125, 344.375, 345.625, 346.875, 348.125, 349.375, 350.625, 
    351.875, 353.125, 354.375, 355.625, 356.875, 358.125, 359.375 ;

 lat = -89.5, -88.5, -87.5, -86.5, -85.5, -84.5, -83.5, -82.5, -81.5, -80.5, 
    -79.5, -78.5, -77.5, -76.5, -75.5, -74.5, -73.5, -72.5, -71.5, -70.5, 
    -69.5, -68.5, -67.5, -66.5, -65.5, -64.5, -63.5, -62.5, -61.5, -60.5, 
    -59.5, -58.5, -57.5, -56.5, -55.5, -54.5, -53.5, -52.5, -51.5, -50.5, 
    -49.5, -48.5, -47.5, -46.5, -45.5, -44.5, -43.5, -42.5, -41.5, -40.5, 
    -39.5, -38.5, -37.5, -36.5, -35.5, -34.5, -33.5, -32.5, -31.5, -30.5, 
    -29.5, -28.5, -27.5, -26.5, -25.5, -24.5, -23.5, -22.5, -21.5, -20.5, 
    -19.5, -18.5, -17.5, -16.5, -15.5, -14.5, -13.5, -12.5, -11.5, -10.5, 
    -9.5, -8.5, -7.5, -6.5, -5.5, -4.5, -3.5, -2.5, -1.5, -0.5, 0.5, 1.5, 
    2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 13.5, 14.5, 
    15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 25.5, 26.5, 
    27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 37.5, 38.5, 
    39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 49.5, 50.5, 
    51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 61.5, 62.5, 
    63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 73.5, 74.5, 
    75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 85.5, 86.5, 
    87.5, 88.5, 89.5 ;

 orog =
  2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 2931.476, 
    2931.476, 2931.476, 2931.476, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 
    2928.302, 2928.302, 2928.302, 2928.302, 2928.302, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 2792.307, 
    2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 2870.053, 
    2870.053,
  2706.976, 2708.441, 2709.924, 2711.426, 2712.948, 2714.488, 2716.048, 
    2717.627, 2719.226, 2720.844, 2722.483, 2724.141, 2725.819, 2727.518, 
    2729.237, 2730.976, 2732.737, 2734.518, 2736.548, 2747.876, 2763.74, 
    2779.185, 2794.216, 2808.835, 2823.048, 2836.857, 2850.265, 2863.276, 
    2874.312, 2883.83, 2893.64, 2903.743, 2914.142, 2924.839, 2935.838, 
    2947.14, 2958.749, 2967.035, 2968.512, 2969.806, 2971.084, 2972.348, 
    2973.597, 2974.831, 2976.05, 2977.255, 2978.445, 2979.62, 2980.782, 
    2981.929, 2983.062, 2984.181, 2985.287, 2986.378, 2987.456, 2988.52, 
    2989.57, 2990.607, 2991.63, 2992.641, 2993.638, 2994.622, 2995.592, 
    2996.55, 3035.946, 3035.155, 3034.353, 3033.541, 3032.717, 3031.883, 
    3031.037, 3030.181, 3029.313, 3028.435, 3027.545, 3026.644, 3025.731, 
    3024.807, 3023.871, 3022.923, 3021.964, 3020.993, 3020.01, 3019.015, 
    3018.009, 3016.99, 3015.958, 3014.915, 3013.858, 3012.79, 3011.766, 
    3013.051, 3015.458, 3017.748, 3019.922, 3021.981, 3023.924, 3025.753, 
    3027.469, 3029.07, 3029.954, 3030.157, 3030.302, 3030.388, 3030.416, 
    3030.386, 3030.297, 3030.149, 3029.943, 3030.229, 3031.534, 3032.849, 
    3034.149, 3035.433, 3036.702, 3037.956, 3039.195, 3040.419, 3041.629, 
    3042.823, 3044.004, 3045.17, 3046.321, 3047.458, 3048.582, 3049.691, 
    3050.786, 3051.867, 3052.935, 3053.988, 3055.029, 3056.055, 3057.068, 
    3058.068, 3059.055, 3060.028, 3037.836, 3037.007, 3036.167, 3035.314, 
    3034.451, 3033.576, 3032.69, 3031.792, 3030.883, 3029.961, 3029.028, 
    3028.083, 3027.126, 3026.157, 3025.176, 3024.183, 3023.177, 3022.159, 
    3021.128, 3020.085, 3019.03, 3017.961, 3016.88, 3015.785, 3014.678, 
    3013.558, 3012.115, 2998.095, 2977.942, 2958.366, 2939.362, 2920.926, 
    2903.052, 2885.737, 2868.976, 2852.766, 2844.424, 2843.606, 2842.818, 
    2842.059, 2841.33, 2840.631, 2839.96, 2839.319, 2838.707, 2837.901, 
    2836.694, 2835.49, 2834.3, 2833.125, 2831.963, 2830.814, 2829.68, 
    2828.559, 2827.452, 2826.358, 2825.278, 2824.21, 2823.156, 2822.115, 
    2821.086, 2820.071, 2819.068, 2818.078, 2817.101, 2816.136, 2815.184, 
    2814.244, 2813.316, 2812.401, 2811.498, 2810.606, 2693.463, 2694.211, 
    2694.97, 2695.739, 2696.518, 2697.307, 2698.107, 2698.917, 2699.738, 
    2700.57, 2701.412, 2702.264, 2703.128, 2704.002, 2704.888, 2705.784, 
    2706.692, 2707.611, 2708.541, 2709.482, 2710.435, 2711.399, 2712.375, 
    2713.362, 2714.361, 2715.372, 2716.104, 2705.031, 2688.208, 2671.944, 
    2656.235, 2641.077, 2626.466, 2612.399, 2598.871, 2585.881, 2583.04, 
    2590.23, 2597.781, 2605.692, 2613.967, 2622.608, 2631.616, 2640.994, 
    2650.745, 2656.768, 2655.133, 2653.331, 2651.549, 2649.789, 2648.049, 
    2646.33, 2644.631, 2642.953, 2641.295, 2639.657, 2638.039, 2636.44, 
    2634.862, 2633.302, 2631.763, 2630.242, 2628.741, 2627.259, 2625.795, 
    2624.35, 2622.924, 2621.517, 2620.128, 2618.757, 2617.404, 2616.07, 
    2695.921, 2697.24, 2698.576, 2699.93, 2701.303, 2702.694, 2704.103, 
    2705.53,
  2616.392, 2617.273, 2618.158, 2619.048, 2619.943, 2620.843, 2621.747, 
    2622.655, 2625.242, 2648.457, 2676.58, 2703.156, 2728.204, 2749.163, 
    2762.994, 2776.313, 2789.418, 2802.31, 2814.865, 2822.017, 2826.455, 
    2830.959, 2835.529, 2840.165, 2844.865, 2849.632, 2854.463, 2864.562, 
    2884.607, 2895.227, 2903.551, 2911.763, 2919.863, 2927.849, 2935.723, 
    2943.483, 2951.13, 2960.719, 2974.247, 2987.969, 3001.793, 3015.721, 
    3029.594, 3040.171, 3049.799, 3059.966, 3070.679, 3079.656, 3081.333, 
    3082.412, 3083.485, 3084.553, 3085.615, 3086.672, 3087.724, 3088.77, 
    3089.81, 3090.844, 3091.874, 3092.898, 3093.916, 3094.929, 3095.936, 
    3096.938, 3097.107, 3096.505, 3095.899, 3095.29, 3094.677, 3094.062, 
    3093.442, 3092.82, 3092.194, 3091.565, 3090.933, 3090.297, 3089.658, 
    3089.016, 3088.37, 3087.721, 3086.918, 3084.25, 3081.138, 3078.166, 
    3075.331, 3073.985, 3075.965, 3078.028, 3080.023, 3081.95, 3083.78, 
    3084.284, 3084.111, 3083.935, 3083.756, 3083.575, 3083.392, 3083.206, 
    3083.017, 3080.883, 3074.548, 3070.135, 3066.166, 3062.25, 3058.388, 
    3054.58, 3050.826, 3047.126, 3043.48, 3039.58, 3035.122, 3030.666, 
    3026.226, 3021.802, 3017.648, 3019.203, 3023.325, 3027.731, 3032.426, 
    3036.207, 3036.153, 3035.789, 3035.427, 3035.067, 3034.708, 3034.352, 
    3033.998, 3033.645, 3033.294, 3032.945, 3032.598, 3032.253, 3031.909, 
    3031.568, 3031.228, 3030.89, 2956.348, 2957.222, 2958.1, 2958.983, 
    2959.871, 2960.764, 2961.662, 2962.564, 2963.471, 2964.384, 2965.301, 
    2966.222, 2967.149, 2968.08, 2969.016, 2969.957, 2967.897, 2928.796, 
    2880.881, 2835.746, 2793.357, 2762.498, 2754.646, 2748.225, 2742.241, 
    2736.693, 2731.746, 2734.142, 2740.325, 2746.601, 2752.969, 2759.428, 
    2765.979, 2772.62, 2779.352, 2762.73, 2756.997, 2767.693, 2757.199, 
    2746.846, 2736.635, 2726.565, 2716.639, 2706.855, 2697.216, 2687.785, 
    2678.614, 2669.573, 2660.66, 2651.876, 2643.676, 2645.808, 2652.588, 
    2659.914, 2667.792, 2673.925, 2672.725, 2670.938, 2669.16, 2667.391, 
    2665.632, 2663.882, 2662.14, 2660.408, 2658.685, 2656.971, 2655.267, 
    2653.571, 2651.885, 2650.208, 2648.54, 2646.881, 2394.907, 2397.965, 
    2401.04, 2404.132, 2407.241, 2410.366, 2413.509, 2416.668, 2419.844, 
    2423.037, 2426.247, 2429.473, 2432.717, 2435.977, 2439.254, 2442.548, 
    2443.66, 2417.692, 2385.279, 2354.901, 2326.535, 2307.414, 2307.181, 
    2308.263, 2309.845, 2311.925, 2314.657, 2324.284, 2337.528, 2350.97, 
    2364.608, 2378.443, 2392.473, 2406.697, 2421.115, 2430.936, 2437.316, 
    2434.09, 2423.859, 2413.765, 2403.81, 2393.993, 2384.315, 2374.777, 
    2365.379, 2358.329, 2355.739, 2353.58, 2351.754, 2350.261, 2349.841, 
    2366.468, 2391.372, 2417.976, 2446.301, 2469.174, 2469.138, 2467.253, 
    2465.377, 2463.51, 2461.654, 2459.807, 2457.969, 2456.142, 2454.323, 
    2452.515, 2450.716, 2448.927, 2447.147, 2445.377, 2443.617, 2441.867, 
    2609.513, 2610.356, 2611.205, 2612.058, 2612.915, 2613.777, 2614.644, 
    2615.516,
  2582.988, 2583.253, 2583.519, 2583.786, 2595.521, 2630.093, 2662.57, 
    2689.178, 2711.952, 2719.18, 2721.893, 2724.634, 2727.404, 2730.203, 
    2733.031, 2735.888, 2738.773, 2746.715, 2769.25, 2796.405, 2826.763, 
    2856.885, 2885.09, 2903.454, 2919.885, 2935.87, 2951.408, 2962.747, 
    2963.64, 2968.408, 2974.942, 2981.664, 2988.574, 2997.808, 3020.722, 
    3045.929, 3071.01, 3092.298, 3108.777, 3118.563, 3125.991, 3133.345, 
    3140.625, 3147.831, 3154.962, 3162.019, 3169.002, 3177.568, 3191.75, 
    3200.878, 3195.187, 3188.354, 3186.815, 3187.933, 3189.047, 3190.156, 
    3191.262, 3192.364, 3193.462, 3194.555, 3195.645, 3196.731, 3197.813, 
    3198.891, 3162.369, 3161.676, 3160.981, 3160.283, 3159.582, 3158.879, 
    3158.173, 3157.464, 3156.753, 3156.04, 3155.324, 3154.605, 3150.023, 
    3137.752, 3126.367, 3120.639, 3117.16, 3115.124, 3113.496, 3111.85, 
    3110.187, 3108.507, 3106.809, 3105.094, 3103.362, 3098.444, 3084.343, 
    3072.186, 3061.927, 3051.776, 3042.211, 3035.488, 3029.354, 3023.388, 
    3017.588, 3013.355, 3013.073, 3012.215, 3011.04, 3009.83, 3008.587, 
    3006.034, 2995.389, 2983.454, 2971.674, 2961.506, 2953.282, 2947.267, 
    2942.05, 2936.884, 2931.77, 2926.708, 2921.699, 2916.742, 2911.837, 
    2907.786, 2906.527, 2898.155, 2869.797, 2838.979, 2826.859, 2824.137, 
    2821.425, 2818.722, 2816.03, 2813.346, 2810.673, 2808.01, 2805.356, 
    2802.712, 2800.077, 2797.453, 2864.33, 2865.305, 2866.284, 2867.267, 
    2868.253, 2869.242, 2870.236, 2871.232, 2872.233, 2873.237, 2874.245, 
    2875.256, 2798.24, 2565.837, 2352.688, 2281.836, 2267.601, 2280.797, 
    2302.173, 2323.778, 2345.609, 2367.668, 2389.954, 2412.467, 2435.206, 
    2406.838, 2230.319, 2141.954, 2131.318, 2124.047, 2110.2, 2042.983, 
    1969.007, 1897.042, 1827.089, 1776.036, 1775.781, 1822.227, 1885.868, 
    1951.338, 2018.639, 2083.223, 2120.932, 2156.036, 2193.689, 2274.409, 
    2402.604, 2423.77, 2408.025, 2392.437, 2377.006, 2361.732, 2346.615, 
    2331.656, 2316.854, 2303.697, 2295.761, 2310.194, 2382.203, 2461.298, 
    2486.398, 2484.39, 2482.389, 2480.396, 2478.409, 2476.43, 2474.457, 
    2472.492, 2470.534, 2468.584, 2466.64, 2464.704, 2101.898, 2104.981, 
    2108.075, 2111.181, 2114.299, 2117.427, 2120.568, 2123.719, 2126.882, 
    2130.057, 2133.243, 2136.44, 2097.523, 1974.723, 1862.217, 1824.545, 
    1817.359, 1830.111, 1848.834, 1867.757, 1886.88, 1906.201, 1925.721, 
    1945.439, 1965.356, 1979.219, 1975.203, 1984.363, 2005.388, 2027.524, 
    2045.519, 2034.652, 2019.56, 2004.878, 1990.606, 1980.191, 1980.475, 
    1996.017, 2017.314, 2039.223, 2061.745, 2083.276, 2095.299, 2106.37, 
    2118.307, 2145.842, 2190.669, 2198.325, 2193.16, 2188.045, 2182.982, 
    2177.971, 2173.011, 2168.104, 2163.247, 2163.411, 2180.639, 2214.85, 
    2289.264, 2369.915, 2396.58, 2396.135, 2395.693, 2395.251, 2394.812, 
    2394.374, 2393.937, 2393.502, 2393.069, 2392.637, 2392.207, 2391.779, 
    2580.903, 2581.161, 2581.419, 2581.678, 2581.938, 2582.199, 2582.461, 
    2582.724,
  2572.232, 2573.315, 2586.612, 2607.861, 2630.823, 2634.508, 2637.59, 
    2640.697, 2643.828, 2646.985, 2650.167, 2653.772, 2668.616, 2690.826, 
    2719.141, 2747.194, 2774.702, 2797.762, 2808.478, 2810.998, 2810.998, 
    2810.998, 2812.313, 2834.287, 2871.53, 2908.28, 2944.53, 2980.279, 
    3015.455, 3050.581, 3085.987, 3121.673, 3157.633, 3180.69, 3182.582, 
    3182.582, 3182.582, 3185.97, 3199.684, 3219.367, 3240.975, 3262.72, 
    3284.31, 3299.129, 3309.324, 3315.379, 3321.243, 3327.061, 3332.833, 
    3338.558, 3344.238, 3349.731, 3350.603, 3344.664, 3338.302, 3339.477, 
    3341.265, 3343.048, 3344.826, 3346.599, 3348.367, 3350.131, 3351.889, 
    3353.643, 3294.686, 3293.157, 3291.624, 3290.087, 3288.546, 3287, 
    3285.451, 3283.897, 3282.339, 3278.427, 3245.819, 3214.572, 3203.504, 
    3199.691, 3196.061, 3192.402, 3188.714, 3184.996, 3181.249, 3176.896, 
    3156.275, 3131.616, 3113.532, 3096.049, 3078.911, 3064.579, 3058.019, 
    3056.479, 3056.479, 3056.479, 3056.105, 3045.913, 3027.202, 3008.831, 
    2990.805, 2973.125, 2956.62, 2941.047, 2925.453, 2909.837, 2894.202, 
    2883.267, 2882.136, 2882.136, 2882.136, 2879.463, 2868.812, 2855.97, 
    2842.571, 2829.205, 2814.933, 2777.971, 2741.862, 2730.966, 2721.041, 
    2711.193, 2701.424, 2691.732, 2682.118, 2672.063, 2645.87, 2614.773, 
    2589.717, 2585.455, 2582.903, 2580.358, 2577.819, 2575.288, 2572.763, 
    2570.246, 2567.735, 2565.231, 2302.347, 2309.09, 2315.851, 2322.63, 
    2329.428, 2336.245, 2343.08, 2349.934, 2356.807, 2339.495, 2026.666, 
    1709.26, 1591.317, 1611.288, 1635.694, 1660.297, 1685.099, 1710.097, 
    1735.294, 1753.235, 1561.479, 1320.545, 1172.337, 1035.045, 905.1483, 
    822.4051, 859.9432, 871.4916, 871.4916, 871.4916, 879.2747, 896.0859, 
    883.2956, 873.3459, 866.2548, 862.0209, 903.0869, 990.0635, 1080.809, 
    1175.324, 1273.574, 1309.332, 1305.293, 1305.293, 1305.293, 1299.384, 
    1281.856, 1351.541, 1455.159, 1563.995, 1680.324, 1857.068, 1996.811, 
    1988.177, 1974.378, 1960.688, 1947.106, 1933.633, 1920.267, 1908.479, 
    1946.522, 2111.525, 2287.59, 2299.054, 2297.043, 2295.038, 2293.039, 
    2291.044, 2289.055, 2287.072, 2285.094, 2283.122, 1987.154, 1988.164, 
    1989.177, 1990.193, 1991.212, 1992.233, 1993.257, 1994.284, 1995.314, 
    1981.148, 1781.403, 1582.754, 1512.199, 1516.823, 1523.793, 1530.82, 
    1537.903, 1545.043, 1552.239, 1556.746, 1483.982, 1412.3, 1419.391, 
    1430.95, 1443.755, 1462.614, 1494.996, 1503.457, 1503.457, 1503.457, 
    1507.567, 1521.691, 1525.743, 1531.028, 1537.553, 1545.317, 1574.778, 
    1626.374, 1679.864, 1735.247, 1792.505, 1816.095, 1814.671, 1814.671, 
    1814.671, 1813.204, 1809.424, 1836.021, 1874.373, 1914.509, 1957.668, 
    2032.656, 2095.127, 2095.787, 2094.263, 2092.752, 2091.252, 2089.764, 
    2088.289, 2088.302, 2136.152, 2248.722, 2357.925, 2365.917, 2365.621, 
    2365.326, 2365.032, 2364.739, 2364.446, 2364.154, 2363.863, 2363.573, 
    2571.575, 2571.656, 2571.738, 2571.82, 2571.902, 2571.984, 2572.066, 
    2572.149,
  2507.865, 2550.77, 2556.477, 2558.917, 2561.373, 2563.845, 2566.333, 
    2568.836, 2574.769, 2590.403, 2611.468, 2632.239, 2643.192, 2649.851, 
    2656.58, 2663.379, 2667.274, 2681.932, 2710.385, 2744.155, 2779.217, 
    2814.806, 2857.302, 2890.027, 2911.18, 2932.724, 2954.665, 2993.996, 
    3053.429, 3091.615, 3116.519, 3140.971, 3164.977, 3197.965, 3238.456, 
    3273.046, 3307.143, 3339.061, 3363.391, 3375.833, 3381.774, 3392.15, 
    3402.418, 3412.578, 3424.243, 3439.459, 3455.768, 3478.595, 3490.129, 
    3496.469, 3502.768, 3509.026, 3515.245, 3521.423, 3525.599, 3520.381, 
    3517.102, 3519.121, 3521.136, 3523.146, 3525.153, 3527.154, 3529.152, 
    3531.145, 3453.831, 3452.036, 3450.237, 3448.435, 3446.628, 3444.818, 
    3443.004, 3441.186, 3400.166, 3342.26, 3329.826, 3325.026, 3320.195, 
    3315.333, 3310.439, 3305.515, 3287.213, 3239.67, 3208.957, 3181.718, 
    3168.715, 3161.957, 3155.126, 3148.225, 3144.272, 3131.434, 3106.626, 
    3078.806, 3050.432, 3023.489, 3001.163, 2985.969, 2977.611, 2969.099, 
    2960.43, 2941.688, 2909.57, 2886.421, 2869.775, 2853.43, 2837.385, 
    2818.593, 2797.607, 2779.112, 2760.877, 2744.654, 2734.706, 2729.707, 
    2722.396, 2709.628, 2696.992, 2684.489, 2662.327, 2618.121, 2571.572, 
    2523.625, 2505.56, 2499.713, 2493.903, 2488.13, 2482.395, 2476.696, 
    2465.276, 2264.471, 2078.934, 2072.39, 2065.861, 2059.345, 2052.844, 
    2046.357, 2039.884, 2033.425, 1324.879, 1336.371, 1347.888, 1359.43, 
    1370.997, 1382.59, 1394.208, 1405.85, 1109.479, 668.9953, 628.1596, 
    665.8774, 703.8411, 742.0505, 780.5058, 819.2067, 829.6528, 733.8724, 
    482.0731, 230.1169, 162.5387, 176.472, 190.5528, 204.7811, 212.9248, 
    193.7189, 158.7268, 153.3229, 159.0761, 160.8323, 132.0868, 129.2712, 
    159.2557, 189.82, 220.9477, 271.3913, 321.7152, 336.9072, 345.4443, 
    353.8268, 362.0825, 427.4072, 541.6088, 626.5125, 709.4601, 801.019, 
    910.6169, 968.3083, 963.6867, 955.6019, 947.6009, 939.6837, 989.4218, 
    1169.603, 1365.752, 1582.781, 1638.927, 1628.308, 1617.757, 1607.274, 
    1596.858, 1586.51, 1619.92, 1885.616, 2067.39, 2064.658, 2061.931, 
    2059.21, 2056.496, 2053.787, 2051.084, 2048.387, 1999.795, 1999.451, 
    1999.108, 1998.763, 1998.417, 1998.071, 1997.724, 1997.377, 1819.175, 
    1542.373, 1491.024, 1488.953, 1486.869, 1484.771, 1482.66, 1480.536, 
    1428.735, 1265.53, 1153.587, 1054.873, 1024.05, 1023.203, 1022.348, 
    1021.484, 1020.986, 1002.777, 969.2682, 957.6859, 954.5271, 955.6179, 
    974.0505, 1007.466, 1054.005, 1101.425, 1149.719, 1191.817, 1259.093, 
    1304.739, 1309.47, 1314.116, 1318.691, 1353.353, 1416.325, 1480.073, 
    1546.065, 1615.728, 1691.401, 1731.007, 1726.137, 1717.624, 1709.199, 
    1700.862, 1716.591, 1786.698, 1866.41, 1978.599, 2009.779, 2005.315, 
    2000.879, 1996.471, 1992.092, 1987.741, 2010.291, 2169.756, 2277.037, 
    2275.842, 2274.649, 2273.459, 2272.272, 2271.087, 2269.905, 2268.725, 
    2462.676, 2464.075, 2465.477, 2466.882, 2468.291, 2469.702, 2471.116, 
    2472.534,
  2417.969, 2423.733, 2429.528, 2435.354, 2441.212, 2448.275, 2498.81, 
    2530.062, 2542.343, 2546.875, 2551.056, 2555.274, 2559.53, 2577.852, 
    2607.827, 2634.506, 2662.848, 2685.807, 2698.749, 2711.889, 2725.225, 
    2757.73, 2821.978, 2883.795, 2943.733, 3001.836, 3042.558, 3063.11, 
    3063.346, 3078.865, 3113.746, 3175.7, 3239.848, 3297.559, 3346.552, 
    3376.785, 3395.66, 3414.256, 3432.573, 3457.488, 3480.301, 3499.673, 
    3525.75, 3550.401, 3563.182, 3575.851, 3588.409, 3601.442, 3626.152, 
    3659.073, 3689.275, 3697.376, 3704.859, 3712.302, 3719.706, 3727.069, 
    3726.403, 3713.486, 3715.319, 3717.549, 3719.775, 3721.997, 3724.215, 
    3726.429, 3612.654, 3610.893, 3609.129, 3607.362, 3605.592, 3603.818, 
    3599.986, 3515.486, 3466.552, 3461.98, 3457.383, 3452.762, 3448.115, 
    3442.305, 3392.832, 3334.671, 3294.689, 3285.035, 3276.819, 3268.53, 
    3260.168, 3233.028, 3193.182, 3158.741, 3123.35, 3101.934, 3093.246, 
    3084.426, 3075.473, 3054.093, 3012.15, 2974.411, 2939.791, 2906.228, 
    2882.542, 2870.549, 2870.421, 2862.922, 2845.144, 2811.172, 2775.96, 
    2739.161, 2700.039, 2675.492, 2659.808, 2644.355, 2629.135, 2608.717, 
    2586.673, 2568.504, 2543.337, 2515.941, 2500.869, 2485.928, 2471.118, 
    2455.059, 2411.356, 2326.164, 2211.967, 2194.804, 2180.319, 2165.91, 
    2151.58, 2137.325, 1901.427, 1449.001, 1430.431, 1423.113, 1415.809, 
    1408.517, 1401.239, 1393.973, 283.5397, 295.1469, 306.7751, 318.4243, 
    330.0944, 341.7856, 352.7019, 279.5561, 88.36246, 97.63815, 106.9651, 
    116.3424, 125.77, 135.2467, 140.6181, 72.1124, 4.407782, 1.312659, 
    1.429233, 1.546839, 1.665475, 4.460826, 11.57062, 17.82682, 27.56687, 
    25.7016, 25.19915, 24.68904, 24.17128, 34.48947, 62.95461, 110.1863, 
    170.8522, 229.7268, 273.4659, 296.1462, 296.3458, 304.208, 322.8071, 
    358.2492, 394.9845, 433.2184, 473.6566, 499.0136, 515.201, 531.1491, 
    546.8578, 595.2074, 663.3764, 735.8531, 816.6348, 863.4515, 872.7776, 
    882.0227, 891.1866, 907.8212, 1076.341, 1311.173, 1469.03, 1471.886, 
    1470.771, 1469.662, 1468.56, 1467.463, 1654.959, 1959.475, 1966.346, 
    1965.803, 1965.261, 1964.72, 1964.18, 1963.641, 1952.149, 1952.88, 
    1953.612, 1954.346, 1955.081, 1955.818, 1950.273, 1688.524, 1515.207, 
    1514.969, 1514.73, 1514.49, 1514.248, 1509.255, 1323.691, 1129.191, 
    1014.88, 1013.563, 1017.898, 1022.271, 1026.683, 953.5953, 790.9396, 
    634.5114, 488.637, 467.1274, 504.8156, 543.0782, 581.9149, 607.1954, 
    609.7045, 640.8179, 693.5481, 743.7175, 743.764, 735.2078, 735.4746, 
    784.8616, 865.8653, 931.783, 998.816, 1088.438, 1207.701, 1243.877, 
    1230.092, 1216.509, 1203.131, 1233.729, 1331.984, 1438.829, 1544.266, 
    1597.374, 1592.83, 1588.325, 1583.859, 1583.464, 1664.207, 1778.368, 
    1849.562, 1845, 1838.537, 1832.108, 1825.713, 1819.353, 1919.26, 
    2076.531, 2077.831, 2075.299, 2072.771, 2070.249, 2067.73, 2065.217, 
    2285.444, 2287.547, 2289.655, 2291.766, 2293.881, 2296, 2299.907, 2373.95,
  2286.4, 2290.566, 2294.752, 2298.958, 2365.091, 2450.854, 2476.203, 
    2480.038, 2483.903, 2487.797, 2509.636, 2549.327, 2583.674, 2603.08, 
    2607.016, 2612.797, 2618.668, 2662.247, 2738.71, 2802.105, 2855.816, 
    2891.822, 2899.201, 2904.123, 2921.436, 2979.917, 3053.518, 3130.385, 
    3194.388, 3246.078, 3290.815, 3311.875, 3318.475, 3341.535, 3374.126, 
    3422.995, 3481.765, 3530.93, 3567.555, 3594.439, 3610.26, 3625.88, 
    3636.355, 3654.066, 3690.511, 3734.728, 3753.662, 3761.404, 3769.087, 
    3776.712, 3794.903, 3839.186, 3869.627, 3874.377, 3879.106, 3883.813, 
    3888.499, 3884.381, 3872.996, 3874.564, 3876.158, 3877.75, 3879.338, 
    3880.925, 3756.281, 3754.721, 3753.159, 3751.594, 3750.027, 3748.246, 
    3651.187, 3596.416, 3591.986, 3587.535, 3583.064, 3578.573, 3533.508, 
    3458.252, 3429.052, 3420.678, 3412.241, 3403.74, 3377.998, 3314.378, 
    3259.929, 3232.676, 3225.683, 3215.359, 3204.897, 3175.019, 3128.163, 
    3080.278, 3031.471, 2993.915, 2974.687, 2961.187, 2953.571, 2929.141, 
    2896.192, 2861.182, 2823.539, 2782.939, 2746.286, 2723.934, 2716.996, 
    2701.252, 2678.974, 2643.965, 2601.194, 2555.446, 2505.41, 2471.348, 
    2455.574, 2440.002, 2429.533, 2405.889, 2356.14, 2281.98, 2225.844, 
    2200.357, 2175.06, 2149.955, 2077.313, 1856.227, 1670.002, 1648.254, 
    1626.605, 1605.055, 1583.604, 1227.222, 484.0244, 470.3725, 458.4476, 
    446.541, 434.6526, 422.7826, 13.05668, 13.63029, 14.20478, 14.78015, 
    15.3564, 15.93352, 10.76648, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04014483, 1.538256, 3.789015, 6.072715, 19.04842, 41.40682, 72.81525, 
    111.0232, 139.232, 151.2006, 159.5457, 169.4505, 202.5452, 248.4973, 
    297.6593, 343.4088, 386.1395, 424.7769, 448.5375, 455.7775, 468.7647, 
    487.1888, 518.8571, 558.6288, 604.6682, 659.3762, 695.4293, 710.1022, 
    724.5844, 734.442, 783.2798, 881.3284, 993.6006, 1034.229, 1047.167, 
    1060.008, 1072.752, 1158.295, 1405.98, 1552.758, 1559.038, 1565.289, 
    1571.512, 1577.707, 1743.583, 2008.169, 2009.589, 2010.456, 2011.322, 
    2012.186, 2013.049, 2010.282, 2009.239, 2008.195, 2007.149, 2006.101, 
    2004.433, 1723.251, 1568.941, 1566.299, 1563.645, 1560.979, 1558.301, 
    1359.241, 1058.275, 970.3054, 969.4023, 968.4924, 967.5755, 896.8425, 
    701.8871, 516.5125, 413.3745, 413.4785, 414.3311, 415.1687, 358.8437, 
    252.8424, 202.9199, 194.9326, 200.6423, 228.1807, 248.0919, 238.6214, 
    208.1117, 222.3655, 251.5968, 301.2507, 371.7545, 449.3096, 541.5269, 
    568.5027, 542.9609, 508.4511, 550.4748, 640.1557, 757.4654, 911.2913, 
    982.7734, 959.7604, 936.99, 922.348, 1036.365, 1234.683, 1431.237, 
    1491.49, 1477.827, 1464.266, 1450.808, 1472.913, 1589.164, 1672.705, 
    1667.06, 1661.44, 1655.846, 1650.278, 1739.077, 1912.045, 1910.833, 
    1909.234, 1907.638, 1906.045, 1904.454, 2098.642, 2100.724, 2102.809, 
    2104.897, 2106.989, 2109.349, 2225.564, 2282.252,
  2231.854, 2232.311, 2248.591, 2395.362, 2457.512, 2454.439, 2451.331, 
    2448.203, 2490.268, 2569.555, 2620.918, 2622.948, 2621.961, 2621.024, 
    2681.026, 2776.42, 2846.989, 2872.887, 2867.472, 2861.983, 2898.416, 
    2976.783, 3053.299, 3129.272, 3180.24, 3188.132, 3194.952, 3237.168, 
    3300.053, 3355.282, 3401.907, 3448.073, 3498.618, 3522.933, 3539.071, 
    3571.407, 3598.016, 3615.508, 3632.765, 3658.817, 3693.5, 3725.508, 
    3749.54, 3760.49, 3766.961, 3768.314, 3796.655, 3839.092, 3862.486, 
    3864.161, 3865.824, 3867.482, 3895.554, 3950.737, 3957.544, 3958.849, 
    3960.148, 3961.442, 3969.173, 3982.054, 3983.094, 3984.134, 3985.172, 
    3986.208, 3886.682, 3885.26, 3883.836, 3882.41, 3880.982, 3818.683, 
    3727.428, 3722.966, 3718.486, 3713.989, 3701.584, 3616.827, 3568.286, 
    3560.719, 3553.11, 3545.451, 3507.352, 3432.329, 3379.485, 3376.698, 
    3369.555, 3357.314, 3317.654, 3261.697, 3209.234, 3175.63, 3157.799, 
    3139.727, 3105.662, 3064.042, 3038.384, 3008.525, 2969.331, 2941.995, 
    2914.637, 2872.983, 2816.354, 2770.259, 2749.49, 2728.799, 2689.823, 
    2647.703, 2610.039, 2559.092, 2515.382, 2497.778, 2480.409, 2448.251, 
    2391.039, 2312.725, 2256.849, 2239.887, 2229.994, 2223.634, 2098.976, 
    1915.242, 1804.945, 1783.02, 1761.239, 1739.565, 1542.357, 1085.254, 
    1015.029, 993.297, 971.6512, 950.0919, 376.4841, 48.82112, 47.15998, 
    45.50104, 43.84432, 42.18981, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.01814248, 1.593398, 4.785732, 24.11693, 40.4681, 
    48.06828, 55.77158, 75.39605, 132.4407, 170.9472, 211.1353, 248.6506, 
    265.9076, 282.61, 299.4491, 334.7076, 372.504, 385.7674, 399.1413, 
    434.5659, 480.9564, 524.3339, 591.0495, 654.6258, 686.2673, 717.4854, 
    765.887, 835.537, 910.5857, 966.0714, 988.5964, 1001.864, 1006.814, 
    1094.294, 1214.589, 1273.185, 1290.946, 1308.591, 1326.151, 1483.391, 
    1704.289, 1727.673, 1733.061, 1738.428, 1743.773, 1959.091, 2099.614, 
    2100.686, 2101.755, 2102.824, 2103.891, 2108.253, 2107.14, 2106.026, 
    2104.911, 2103.794, 1974.508, 1757.134, 1748.729, 1740.291, 1731.819, 
    1684.019, 1281.393, 1067.246, 1054.494, 1041.702, 1028.825, 861.1204, 
    563.6516, 365.8732, 356.9218, 359.6991, 363.4859, 294.4648, 182.3021, 
    79.47626, 32.69877, 33.38852, 34.08763, 30.49054, 22.56217, 14.71135, 
    13.94608, 14.04704, 23.00423, 33.13614, 47.60875, 47.94914, 34.00398, 
    24.16135, 17.10599, 55.43153, 113.6577, 182.9376, 258.152, 252.6471, 
    229.9988, 207.6536, 264.2766, 416.6413, 590.784, 692.7862, 672.5236, 
    659.5286, 666.8179, 849.7219, 1118.225, 1221.978, 1198.721, 1175.617, 
    1152.686, 1225.884, 1482.372, 1508.029, 1502.722, 1497.435, 1492.169, 
    1665.97, 1795.302, 1794.135, 1792.969, 1791.804, 1790.641, 2020.92, 
    2021.375, 2021.83, 2022.286, 2022.742, 2110.518, 2230.944, 2231.398,
  2271.499, 2298.749, 2480.609, 2517.394, 2513.175, 2508.931, 2533.648, 
    2657.216, 2728.562, 2725.188, 2723.473, 2731.69, 2826.094, 2923.154, 
    2950.07, 2940.414, 2931.698, 2978.17, 3058.842, 3138.799, 3180.843, 
    3180.532, 3184.142, 3234.391, 3295.818, 3356.674, 3416.17, 3439.871, 
    3439.871, 3459.615, 3504.06, 3548, 3590.074, 3628.505, 3654.004, 3662.99, 
    3670.084, 3686.816, 3703.394, 3710.503, 3711.141, 3711.664, 3719.972, 
    3744.249, 3768.285, 3772.347, 3772.336, 3763.736, 3786.017, 3836.969, 
    3844.266, 3835.906, 3827.594, 3833.566, 3904.766, 3915.75, 3912.003, 
    3908.27, 3906.904, 3964.8, 3970.384, 3969.691, 3969, 3968.31, 3925.66, 
    3925.618, 3925.576, 3925.533, 3918.118, 3816.224, 3805.838, 3804.154, 
    3802.463, 3790.804, 3709.763, 3683.615, 3677.876, 3672.103, 3650.2, 
    3566.651, 3511.147, 3504.95, 3502.794, 3484.539, 3418.531, 3352.879, 
    3323.903, 3311.276, 3298.064, 3261.986, 3211.943, 3166.115, 3149.236, 
    3141.011, 3116.432, 3067.057, 3012.58, 2963.541, 2915.373, 2894.569, 
    2894.569, 2871.32, 2815.241, 2757.158, 2689.803, 2630.577, 2611.87, 
    2606.375, 2575.163, 2503.093, 2425.539, 2369.596, 2358.584, 2348.563, 
    2313.762, 2178.821, 2025.607, 1986.357, 1982.431, 1991.629, 1856.782, 
    1592.422, 1515.382, 1514.153, 1512.931, 1386.314, 658.9482, 502.4041, 
    488.8896, 475.4227, 420.0609, 22.91726, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.750073, 13.04912, 21.49358, 
    20.28802, 17.88101, 15.44909, 12.81549, 7.463051, 2.387415, 1.250797, 
    13.76716, 51.18564, 126.25, 199.8179, 216.8334, 225.8941, 230.111, 
    230.111, 267.4045, 353.6554, 437.7119, 505.5228, 563.4755, 594.2936, 
    604.7546, 645.7354, 763.8188, 893.3362, 986.5775, 1025.809, 1063.577, 
    1120.356, 1210.241, 1296.074, 1330.288, 1335.872, 1348.319, 1422.991, 
    1527.21, 1555.219, 1566.16, 1577.038, 1634.42, 1820.474, 1847.059, 
    1849.925, 1852.781, 1875.035, 2086.654, 2100.651, 2100.153, 2099.655, 
    2099.157, 2154.697, 2154.415, 2154.133, 2153.851, 2139.569, 1942.92, 
    1921.773, 1917.658, 1913.528, 1848.098, 1418.221, 1301.004, 1285.492, 
    1269.889, 1130.824, 655.5745, 390.891, 389.257, 388.7375, 364.7886, 
    223.2671, 82.52729, 37.23098, 35.86035, 34.2843, 23.64924, 13.47776, 
    4.813199, 0.4541103, 0.5494496, 0.8123864, 1.08686, 3.193648, 14.8494, 
    27.82338, 33.37933, 33.37933, 51.68832, 90.29761, 123.2752, 123.158, 
    121.6044, 140.8415, 148.706, 143.5132, 140.2252, 123.9206, 66.85396, 
    53.33577, 40.97689, 100.2805, 243.8672, 361.2292, 360.3512, 355.2744, 
    347.0272, 517.4183, 812.3451, 870.7962, 860.2645, 849.7943, 919.6375, 
    1246.371, 1287.198, 1277.891, 1268.617, 1279.34, 1662.406, 1698.768, 
    1697.749, 1696.731, 1695.714, 2052.424, 2051.752, 2051.081, 2050.408, 
    2067.328, 2266.995, 2277.197, 2274.353,
  2366.138, 2520.391, 2555.055, 2555.978, 2556.906, 2657.013, 2794.567, 
    2804.754, 2802.877, 2813.933, 2922.885, 3024.623, 3029.926, 3022.394, 
    3034.943, 3109.455, 3185.776, 3209.76, 3207.749, 3220.967, 3274.629, 
    3330.957, 3389.333, 3405.079, 3411.149, 3443.011, 3480.327, 3519.586, 
    3559.834, 3585.301, 3594.92, 3607.459, 3614.139, 3624.028, 3645.081, 
    3665.803, 3685.468, 3690.173, 3683.374, 3670.561, 3662.812, 3638.017, 
    3615.763, 3597.52, 3582.42, 3592.01, 3605.037, 3602.823, 3590.904, 
    3578.25, 3637.44, 3672.881, 3658.95, 3645.092, 3647.829, 3723.11, 
    3723.551, 3714.82, 3706.117, 3737.445, 3771.708, 3768.701, 3765.698, 
    3762.698, 3790.26, 3792.46, 3794.662, 3796.867, 3791.314, 3774.23, 
    3777.106, 3779.992, 3783.815, 3757.279, 3745.794, 3745.465, 3745.135, 
    3710.177, 3632.349, 3618.31, 3614.275, 3603.866, 3535.297, 3467.897, 
    3448.191, 3435.215, 3410.463, 3354.489, 3306.083, 3279.305, 3272.842, 
    3260.622, 3208.74, 3154.413, 3102.054, 3071.901, 3046.416, 3013.574, 
    2993.564, 2960.785, 2913.311, 2869.743, 2834.16, 2794.548, 2775.724, 
    2748.948, 2683.247, 2601.836, 2521.23, 2501.919, 2501.282, 2476.124, 
    2407.83, 2344.289, 2331.412, 2334.416, 2321.449, 2243.98, 2185.951, 
    2183.521, 2185.938, 2152.175, 1772.569, 1571.897, 1586.598, 1601.222, 
    1455.466, 517.4026, 408.7929, 414.7833, 420.7549, 222.803, 1.138203, 
    1.15751, 1.176797, 1.196063, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.471831, 23.60061, 40.66413, 40.26577, 38.37702, 33.56215, 
    25.19385, 26.73575, 28.38287, 29.0506, 46.88717, 119.4331, 187.6333, 
    219.6661, 212.493, 199.6839, 272.3419, 381.0488, 492.0388, 553.6685, 
    541.79, 505.315, 525.5818, 593.9067, 668.2168, 765.5681, 861.2631, 
    950.9992, 971.5608, 999.3796, 1091.441, 1231.762, 1316.017, 1352.862, 
    1383.517, 1420.918, 1489.661, 1550.053, 1562.03, 1566.254, 1580.576, 
    1657.991, 1690.982, 1691.064, 1691.146, 1717.782, 1831.042, 1837.016, 
    1833.877, 1830.748, 1902.864, 1966.609, 1964.597, 1962.588, 1960.58, 
    2032.004, 2034.107, 2036.213, 2038.321, 2017.574, 1974.503, 1974.333, 
    1974.161, 1940.741, 1598.229, 1521.177, 1512.744, 1504.267, 1079.193, 
    444.7661, 377.4638, 373.4092, 354.761, 192.6595, 42.33033, 27.2869, 
    29.56788, 31.71604, 27.00497, 10.22225, 2.464777, 1.332851, 1.205324, 
    0.6701186, 0.2070511, 0.2301773, 0.319214, 0.4209029, 2.492963, 5.062005, 
    10.87739, 64.91257, 145.9952, 206.2483, 255.5906, 261.1143, 259.425, 
    239.2852, 228.173, 219.0093, 216.5157, 202.9371, 143.9775, 38.40372, 
    53.64306, 85.42174, 101.3828, 133.6189, 176.6659, 170.9041, 166.3376, 
    195.3281, 276.5435, 636.1906, 778.5042, 786.293, 794.0412, 857.9529, 
    1201.496, 1248.445, 1254.177, 1259.892, 1484.871, 1692.794, 1693.228, 
    1693.662, 1694.095, 2081.164, 2081.004, 2080.844, 2080.685, 2225.306, 
    2360.557, 2357.84, 2355.115,
  2546.797, 2580.593, 2575.669, 2572.322, 2717.728, 2844.222, 2842.325, 
    2840.932, 2918.557, 3047.806, 3066.964, 3064.836, 3092.071, 3184.888, 
    3244.741, 3244.907, 3244.258, 3293.182, 3354.253, 3397.152, 3397.786, 
    3404.192, 3454.456, 3503.917, 3552.015, 3565.503, 3567.877, 3599.412, 
    3627.309, 3645.214, 3668.81, 3674.098, 3663.96, 3654.023, 3631.226, 
    3622.546, 3618.596, 3611.119, 3591.426, 3576.427, 3555.24, 3533.41, 
    3500.002, 3440.368, 3403.846, 3381.678, 3363.646, 3360.6, 3360.898, 
    3342.601, 3316.917, 3350.625, 3390.941, 3370.715, 3350.022, 3353.577, 
    3410.396, 3399.111, 3386.761, 3382.793, 3456.015, 3453.181, 3449.435, 
    3445.692, 3549.55, 3552.431, 3555.315, 3559.629, 3658.424, 3667.595, 
    3671.739, 3677.038, 3725.807, 3732.916, 3735.197, 3737.462, 3720.787, 
    3697.233, 3696.478, 3695.941, 3647.326, 3564.58, 3544.938, 3536.83, 
    3512.602, 3450.44, 3402.919, 3389.615, 3377.023, 3344.437, 3298.981, 
    3253.353, 3230.847, 3204.957, 3154.413, 3107.031, 3079.201, 3063.486, 
    3036.415, 3001.413, 2952.991, 2902.177, 2884.169, 2866.332, 2819.241, 
    2760.742, 2695.526, 2674.567, 2659.51, 2603.837, 2542.525, 2496.349, 
    2498.196, 2499.968, 2455.242, 2409.906, 2406.204, 2416.076, 2409.376, 
    2300.718, 2232.839, 2242.742, 2256.547, 2063.76, 1850.987, 1866.763, 
    1884.708, 1604.962, 751.5079, 754.6127, 770.6727, 724.9202, 62.7219, 
    55.49179, 56.4132, 57.33372, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 3.384167, 9.939319, 14.75, 19.60527, 19.59743, 13.20769, 15.16736, 
    22.51605, 96.82114, 190.9584, 257.633, 263.8174, 269.9198, 334.3635, 
    490.733, 598.4749, 625.8487, 628.1277, 654.2975, 721.4735, 814.3557, 
    874.6158, 890.0057, 896.0983, 999.3834, 1088.404, 1186.378, 1289.058, 
    1386.368, 1417.83, 1432.344, 1491.051, 1552.476, 1628.461, 1627.451, 
    1632.779, 1658.151, 1683.611, 1666.343, 1647.541, 1648.052, 1648.792, 
    1666.979, 1635.381, 1623.028, 1611.848, 1621.938, 1641.224, 1631.225, 
    1621.296, 1622.626, 1708.576, 1706.182, 1702.864, 1699.549, 1753.088, 
    1756.651, 1760.217, 1764.747, 1833.418, 1844.27, 1851.945, 1857.062, 
    1655.227, 1576.43, 1581.173, 1580.601, 1023.165, 498.2543, 473.5003, 
    456.1139, 344.0132, 153.9532, 112.2552, 99.92363, 67.58768, 14.30644, 
    14.59048, 16.69151, 18.41009, 13.2531, 4.606415, 0.5053398, 0.3747498, 
    0.2324216, 0.01148218, -1.56782e-16, -3.423825e-17, 0.7861331, 3.105798, 
    5.582565, 30.0408, 70.90997, 91.36034, 111.3166, 156.7123, 188.764, 
    198.2682, 173.8806, 143.8394, 91.98463, 34.40762, 5.468679, 15.06332, 
    30.27674, 93.45506, 253.6712, 333.1825, 362.3015, 407.3329, 620.8641, 
    753.7205, 772.492, 798.8773, 881.0955, 1039.544, 1074.414, 1106.56, 
    1238.481, 1461.939, 1472.555, 1481.346, 1527.435, 1806.925, 1811.215, 
    1812.998, 1814.78, 2153.594, 2152.474, 2151.354, 2152.11, 2365.266, 
    2395.218, 2395.135, 2397.866,
  2662.239, 2658.33, 2655.473, 2805.033, 2885.527, 2875.435, 2877.643, 
    3026.779, 3111.224, 3106.622, 3113.283, 3202.281, 3275.048, 3275.655, 
    3280.67, 3340.436, 3406.248, 3420.146, 3418.33, 3461.844, 3523.102, 
    3572.203, 3577.38, 3586.766, 3622.096, 3659.385, 3697.607, 3708.364, 
    3712.104, 3718.875, 3718.814, 3706.963, 3691.234, 3686.558, 3673.686, 
    3637.305, 3590.368, 3547.657, 3532.028, 3511.882, 3468.17, 3400.35, 
    3362.564, 3331.265, 3261.367, 3160.465, 3123.042, 3095.266, 3066.354, 
    3045.612, 3015.966, 2983.613, 2982.402, 2990.806, 2965.59, 2940.376, 
    2974.699, 3015.088, 3001.722, 2988.39, 3091.261, 3128.179, 3124.738, 
    3121.301, 3338.033, 3340.032, 3342.032, 3396.889, 3552.488, 3555.909, 
    3559.338, 3628.592, 3695.964, 3697.66, 3699.495, 3708.008, 3706.336, 
    3705.626, 3700.426, 3638.617, 3598.231, 3594.013, 3581.324, 3510.575, 
    3464.094, 3459.647, 3449.579, 3396.531, 3342.951, 3323.964, 3314.897, 
    3279.691, 3233.677, 3193.955, 3182.426, 3176.94, 3146.214, 3111.095, 
    3075.612, 3046.792, 3035.571, 3019.373, 2971.836, 2908.972, 2844.881, 
    2829.327, 2816.549, 2754.696, 2687.03, 2643.696, 2641.401, 2628.808, 
    2580.316, 2537.577, 2535.655, 2537.175, 2505.764, 2470.516, 2470.271, 
    2474.682, 2448.594, 2404.153, 2394.474, 2387.55, 2252.618, 2012.477, 
    1999.346, 1987.928, 1334.051, 737.2125, 721.4674, 705.7629, 246.7386, 
    131.4117, 132.1874, 132.9624, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.536153, 50.88648, 106.1154, 135.1531, 157.7303, 
    162.4228, 208.2697, 289.1352, 333.3496, 322.2963, 301.9858, 341.721, 
    523.9764, 691.3443, 779.5907, 898.9597, 1050.888, 1260.571, 1466.653, 
    1506.879, 1565.076, 1628.024, 1713.523, 1825.734, 1918.999, 1970.869, 
    1917.67, 1903.234, 1943.994, 1983.559, 1961.555, 1860.895, 1864.8, 
    1884.928, 1817.473, 1665.538, 1641.738, 1627.67, 1550.323, 1427.576, 
    1414.753, 1402.745, 1377.226, 1346.244, 1337.021, 1327.822, 1389.943, 
    1407.859, 1404.628, 1401.4, 1439.486, 1442.84, 1446.196, 1457.743, 
    1507.887, 1521.206, 1534.559, 1523.25, 1460.423, 1469.121, 1475.986, 
    1075.413, 770.6211, 761.2312, 735.3962, 493.1752, 336.6808, 313.7148, 
    280.2278, 174.6711, 94.48317, 65.49535, 45.31432, 32.74599, 41.22555, 
    40.27128, 32.66009, 18.65729, 8.442912, 3.503948, 0.120401, 
    -1.560545e-18, -7.193992e-19, 0.04831598, 0.2237047, 0.3360482, 
    0.3360482, 5.471201, 27.53351, 20.16712, 4.694813, 3.045152, 6.422132, 
    35.70369, 47.81778, 30.76674, 13.63443, 10.22249, 46.37926, 73.56437, 
    68.12915, 66.64082, 210.8164, 513.9006, 571.1777, 590.5852, 768.0147, 
    1051.742, 1070.512, 1068.454, 1210.697, 1435.901, 1435.647, 1434.023, 
    1553.654, 1691.086, 1697.085, 1703.069, 1920.359, 1990.928, 1993.004, 
    1995.079, 2239.434, 2238.596, 2237.757, 2293.984, 2463.75, 2459.928, 
    2456.096, 2546.387,
  2753.314, 2746.197, 2861.879, 2994.902, 2992.817, 3009.696, 3147.906, 
    3179.549, 3172.52, 3216.395, 3313.229, 3321.046, 3314.415, 3361.428, 
    3430.863, 3442.235, 3445.398, 3496.214, 3560.025, 3583.208, 3587.095, 
    3614.95, 3644.241, 3673.042, 3682.039, 3675.093, 3693.946, 3695.918, 
    3704.604, 3716.475, 3707.763, 3701.355, 3680.396, 3651.234, 3632.246, 
    3606.123, 3582.813, 3548.797, 3478.783, 3402.599, 3378.182, 3355.846, 
    3244.15, 3121.462, 3079.84, 3029.427, 2886.241, 2792.249, 2758.186, 
    2715.052, 2639.648, 2591.478, 2551.993, 2531.666, 2535.397, 2511.959, 
    2495.374, 2640.291, 2652.771, 2642.809, 2750.637, 2887.861, 2885.799, 
    2883.739, 3202.071, 3203.231, 3204.393, 3345.075, 3468.01, 3470.322, 
    3489.459, 3644.943, 3656.497, 3659.578, 3687.105, 3708.411, 3710.542, 
    3702.781, 3630.011, 3609.656, 3608.899, 3565.121, 3481.129, 3469.731, 
    3467.204, 3400.318, 3334.201, 3323.474, 3319.893, 3279.141, 3239.67, 
    3230.793, 3232.716, 3223.03, 3206.16, 3184.919, 3171.347, 3159.95, 
    3146.192, 3144.51, 3118.453, 3077.5, 3029.104, 2989.745, 2978.164, 
    2923.694, 2853.62, 2791.712, 2780.985, 2757.138, 2697.078, 2649.388, 
    2644.79, 2636.49, 2588.342, 2550.316, 2547.627, 2539.61, 2491.258, 
    2465.465, 2463.711, 2434.403, 2321.052, 2283.861, 2261.95, 2010.352, 
    1723.236, 1699.246, 1607.263, 431.8068, 299.8416, 287.4518, 171.1071, 
    64.40877, 62.71233, 61.01723, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1.511268, 16.77075, 35.311, 33.29043, 
    34.74964, 44.18677, 36.23867, 36.74366, 39.37407, 59.55199, 103.6159, 
    290.467, 413.8759, 618.7913, 823.7323, 1032.218, 1248.352, 1286.407, 
    1459.059, 1708.111, 1868.642, 1841.524, 1799.369, 1890.107, 2115.529, 
    2159.149, 2140.465, 2049.51, 2064.494, 2034.963, 1975.949, 1865.854, 
    1836.931, 1828.185, 1756.461, 1498.967, 1433.705, 1400.558, 1268.799, 
    1146.864, 1125.336, 1100.394, 1025.334, 1007.175, 994.7917, 1002.008, 
    1011.397, 1006.415, 1001.437, 1063.637, 1068.126, 1072.619, 1114.209, 
    1150.544, 1161.202, 1182.629, 1259.382, 1274.595, 1288.053, 1157.635, 
    920.5621, 899.107, 858.4648, 710.7036, 647.7098, 615.9561, 492.645, 
    316.9719, 280.0913, 268.2321, 375.5646, 366.1596, 355.1998, 320.9935, 
    330.6047, 277.2531, 179.2619, 78.0381, 14.92651, 4.948391, -2.435307e-20, 
    0, 0, 0, 0.001930746, 0.001930746, -2.176492e-16, -3.122068e-16, 
    -2.275466e-16, 0.04297423, 0.1702917, 2.854574e-16, 3.814184e-16, 
    3.01149e-16, 0.09063171, 0.2097051, 0.100082, 0.009018716, 2.370771, 
    16.15766, 19.54172, 15.73925, 66.39478, 234.8315, 225.9868, 177.7843, 
    311.7837, 932.0079, 946.9777, 878.7223, 1001.555, 1169.989, 1129.335, 
    1106.958, 1502.868, 1546.252, 1531.707, 1754.358, 2048.062, 2047.738, 
    2047.415, 2370.361, 2368.602, 2366.843, 2472.43, 2568.448, 2565.264, 
    2581.865, 2750.996,
  2837.594, 2876.796, 3001.012, 3006.747, 3030.758, 3188.445, 3217.064, 
    3215.174, 3296.758, 3369.436, 3367.315, 3379.906, 3440.349, 3462.59, 
    3465.559, 3495.268, 3540.664, 3557.725, 3559.385, 3574.364, 3594.081, 
    3602.45, 3595.33, 3552.338, 3554.084, 3565.32, 3560.413, 3541.179, 
    3544.115, 3568.881, 3575.15, 3568.457, 3567.949, 3573.641, 3559.603, 
    3545.921, 3513.803, 3463.664, 3429.42, 3390.144, 3280.445, 3178.01, 
    3157.048, 3075.183, 2873.38, 2763.525, 2721.041, 2568.434, 2373.436, 
    2329.012, 2278.155, 2123.977, 2063.448, 2020.171, 2088.717, 2136.02, 
    2118.77, 2239.388, 2412.069, 2406.19, 2479.002, 2771.492, 2770.8, 
    2770.108, 3140.152, 3140.506, 3140.86, 3352.605, 3413.554, 3414.891, 
    3507.809, 3591.382, 3595.385, 3617.733, 3669.384, 3675.431, 3672.51, 
    3606.572, 3593.872, 3594.43, 3523.311, 3460.45, 3461.249, 3421.038, 
    3311.031, 3282.596, 3280.567, 3222.2, 3168.129, 3175.654, 3187.144, 
    3186.926, 3180.046, 3179.141, 3186.45, 3198.135, 3208.395, 3213.751, 
    3210.691, 3196.017, 3169.59, 3134.49, 3126.125, 3094.517, 3026.086, 
    2951.991, 2918.808, 2902.287, 2837.136, 2766.636, 2747.644, 2732.067, 
    2673.891, 2624.562, 2618.556, 2596.608, 2542.91, 2522.792, 2517.443, 
    2452.375, 2345.969, 2330.545, 2279.555, 2056.43, 2014.553, 1998.12, 
    1567.78, 1409.899, 1406.404, 813.4013, 117.6464, 117.7202, 92.04891, 
    0.1419247, 0.1382803, 0.1346385, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9100384, 2.98663, 
    4.317764, 2.691871, 2.001092, 28.61652, 151.818, 249.0694, 309.0305, 
    323.4313, 416.4194, 676.0397, 920.04, 933.5768, 948.3104, 1166.477, 
    1327.41, 1250.95, 1139.995, 1320.3, 1536.286, 1479.468, 1354.76, 
    1429.718, 1424.575, 1305.479, 1226.092, 1256.305, 1191.819, 1133.913, 
    1010.09, 940.2251, 877.41, 699.8884, 616.4221, 576.3007, 508.8169, 
    447.5602, 423.8362, 407.5251, 429.3942, 422.3122, 415.2354, 686.8015, 
    690.5506, 694.3024, 902.8237, 953.8391, 956.7819, 1058.525, 1130.373, 
    1129.742, 1136.754, 1147.017, 1144.021, 1117.182, 921.6127, 870.6376, 
    849.3878, 767.6731, 627.1446, 574.0612, 581.8477, 854.0009, 944.5726, 
    947.9935, 1087.469, 1148.428, 987.7026, 810.0967, 514.8839, 292.1046, 
    247.9374, 157.8803, 34.10544, 9.435918, 0.1348292, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, -5.237299e-19, -9.098777e-19, -6.684368e-20, 0, 0, 0, 
    0, 0.5035203, 30.00143, 21.39013, 8.260679, 28.11338, 158.7416, 158.0209, 
    146.4624, 415.0629, 449.9345, 415.9597, 697.8641, 1066.841, 1050.189, 
    1210.723, 1861.519, 1858.385, 1855.253, 2415.562, 2415.87, 2416.178, 
    2638.522, 2690.523, 2685.889, 2760.055, 2838.399,
  2771.246, 2852.542, 2889.931, 2930.052, 3110.294, 3150.304, 3160.999, 
    3278.099, 3338.685, 3346.018, 3359.271, 3405.973, 3428.104, 3431.031, 
    3415.947, 3439.237, 3453.413, 3438.134, 3461.69, 3486.851, 3449.107, 
    3392.323, 3371.352, 3385.813, 3315.745, 3226.369, 3236.144, 3309.581, 
    3348.095, 3322.397, 3336.293, 3398.311, 3435.293, 3399.131, 3380.738, 
    3391.653, 3403.584, 3379.198, 3322.232, 3266.426, 3231.48, 3168.011, 
    2995.177, 2906.601, 2874.648, 2674.45, 2441.211, 2403.175, 2233.888, 
    1863.065, 1803, 1735.715, 1535.865, 1487.517, 1488.326, 1820.868, 
    1837.63, 1848.062, 2262.084, 2283.753, 2292.542, 2695.698, 2705.52, 
    2704.831, 3086.861, 3087.558, 3094.468, 3342.086, 3351.612, 3360.828, 
    3502.846, 3516.427, 3523.831, 3583.112, 3596.997, 3600.461, 3549.857, 
    3538.877, 3541.402, 3475.439, 3439.539, 3441.691, 3354.351, 3258.732, 
    3257.6, 3211.626, 3112.203, 3097.411, 3098.139, 3074.765, 3078.798, 
    3090.521, 3103.447, 3128.877, 3156.34, 3180.174, 3196.723, 3201.128, 
    3209.415, 3215.982, 3212.474, 3200.039, 3160.796, 3112.543, 3064.148, 
    3039.21, 2977.884, 2896.956, 2849.867, 2834.008, 2768.688, 2697.156, 
    2672.214, 2645.423, 2591.708, 2559.613, 2542.914, 2494.979, 2457.104, 
    2446.412, 2380.117, 2262.306, 2251.511, 2178.81, 1932.785, 1950.666, 
    1920.596, 1541.829, 1543.046, 1490.827, 594.5919, 588.3399, 612.8005, 
    25.36505, 0.8091006, 0.8233781, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1702477, 
    0.03521304, 0, 0, 5.689764, 34.75395, 24.19427, 30.84762, 28.84321, 
    210.3864, 184.7929, 142.7398, 145.6204, 384.0143, 405.4324, 257.2557, 
    172.8251, 274.7045, 330.7485, 293.5327, 499.8311, 509.4197, 409.6299, 
    367.9375, 376.9431, 299.5526, 267.9969, 241.7466, 222.8664, 189.7327, 
    99.19085, 90.07831, 78.45374, 41.75248, 38.94295, 38.18476, 126.8187, 
    129.1422, 128.7105, 576.8413, 576.3446, 584.0032, 911.4412, 920.3956, 
    921.5487, 1045.982, 1068.664, 1068.158, 1056.048, 1092.165, 1108.074, 
    977.8293, 960.4396, 946.9863, 786.2373, 734.962, 742.5505, 700.4499, 
    856.8281, 945.7138, 1092.408, 1291.525, 1362.956, 1393.334, 1444.634, 
    1443.993, 1441.241, 1188.418, 748.0234, 441.076, 183.1587, 35.33849, 
    10.5561, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5.97522, 34.5936, 31.87986, 74.67491, 528.4946, 
    522.8108, 529.8214, 1314.979, 1326.723, 1319.439, 2115.295, 2120.305, 
    2138.141, 2574.502, 2593.562, 2611.08, 2742.067, 2759.156,
  2415.972, 2483.922, 2526.433, 2878.701, 3105.384, 3115.629, 3130.344, 
    3170.909, 3191.119, 3162.439, 3201.18, 3234.099, 3163.477, 3110.101, 
    3154.842, 3030.224, 3043.607, 3167.357, 3189.942, 3085.677, 3105.43, 
    3100.532, 2968.514, 2872.607, 2873.791, 2855.831, 2875.115, 2948.975, 
    2962.286, 3020.308, 3096.433, 3142.882, 3138.69, 3158.712, 3177.948, 
    3150.855, 3125.85, 3181.723, 3204.532, 3175.801, 3128.265, 3082.664, 
    3058.29, 2929.802, 2752.448, 2727.149, 2564.764, 2193.406, 2146.279, 
    1917.999, 1389.614, 1347.329, 1233.461, 1006.309, 970.0369, 1231.863, 
    1551.363, 1532.136, 1913.697, 2152.571, 2146.768, 2516.796, 2605.055, 
    2603.765, 2987.046, 2988.309, 3037.129, 3242.978, 3246.954, 3306.535, 
    3408.693, 3415.823, 3455.828, 3494.808, 3504.885, 3476.357, 3464.939, 
    3469.124, 3404.02, 3379.883, 3381.659, 3266.83, 3217.943, 3221.45, 
    3111.068, 3027.604, 3035.078, 2990.705, 2959.509, 2974.492, 2990.015, 
    3000.526, 3027.26, 3050.135, 3076.093, 3098.622, 3111.157, 3133.031, 
    3159.849, 3186.012, 3186.577, 3178.302, 3159.843, 3136.999, 3119.639, 
    3048.174, 2951.736, 2898.843, 2844.09, 2783.857, 2724.894, 2681.269, 
    2601.948, 2552.199, 2529.265, 2495.266, 2442.378, 2417.953, 2382.024, 
    2381.54, 2376.226, 2335.592, 2275.761, 2275.974, 2259.853, 2234.205, 
    2235.945, 2057.624, 1899.165, 1912.445, 1550.265, 1385.948, 1408.692, 
    666.3326, 499.6955, 508.4097, 0.1083049, 0.1064435, 0.0808678, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.66507, 0.632016, 0.7361499, 
    1.947761, 34.09342, 110.5448, 131.6132, 100.5916, 46.10235, 36.95004, 
    52.48995, 55.05325, 38.26681, 37.13551, 22.74773, 6.109411, 12.34699, 
    21.14057, 19.17539, 9.217195, 2.550325, 2.328024, 2.142627, 2.968732, 
    3.143221, 74.13859, 89.21502, 88.80952, 352.2433, 356.4258, 377.3625, 
    505.4632, 529.1852, 545.2026, 583.4738, 629.0906, 607.4274, 579.5976, 
    633.189, 406.9331, 249.412, 293.6666, 261.7129, 277.793, 348.3815, 
    339.9253, 323.0953, 379.9896, 323.6219, 307.0536, 492.6911, 679.5224, 
    962.3381, 1230.187, 1396.819, 1304.049, 1185.052, 1085.873, 680.4366, 
    206.4469, 125.405, 47.82164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04465972, 0.07341602, 
    0.06701668, 138.7616, 208.912, 205.3913, 678.1078, 776.1987, 771.5107, 
    1587.93, 1593.741, 1709.095, 2177.959, 2193.169, 2204.594, 2271.102, 
    2313.644,
  1665.958, 1766.78, 2005.679, 2394.572, 2488.598, 2548.831, 2620.788, 
    2676.98, 2554.492, 2637.584, 2693.163, 2509.039, 2519.025, 2476.923, 
    2172.47, 2256.876, 2312.294, 2181.371, 2129.835, 2247.967, 2128.252, 
    2151.648, 2304.337, 2142.054, 2086.202, 2243.116, 2375.114, 2352.1, 
    2466.932, 2655.219, 2699.21, 2663.854, 2727.155, 2822.879, 2792.528, 
    2810.536, 2905.027, 2901.144, 2939.198, 3037.505, 3059.259, 3033.919, 
    3018.576, 3013.368, 2942.215, 2701.854, 2657.285, 2509.609, 2051.262, 
    2008.253, 1658.086, 1110.942, 1105.329, 750.8151, 513.935, 513.7252, 
    1114.546, 1156.158, 1372.195, 1978.934, 1973.892, 2303.612, 2492.551, 
    2491.487, 2838.077, 2839.777, 2922.018, 3071.783, 3078.158, 3178.127, 
    3229.337, 3247.552, 3318.998, 3338.877, 3340.614, 3325.469, 3341.284, 
    3279.913, 3248.718, 3256.671, 3142.13, 3113.604, 3105.602, 2974.406, 
    2944.068, 2928.405, 2848.21, 2846.127, 2859.88, 2862.795, 2865.661, 
    2886.475, 2889.401, 2918.324, 2946.593, 2936.618, 2959.596, 3015.348, 
    3058.323, 3062.226, 3090.862, 3128.218, 3125, 3088.739, 3039.307, 
    3005.62, 2959.971, 2851.531, 2742.632, 2688.891, 2645.766, 2548.444, 
    2491.884, 2443.985, 2362.357, 2319.173, 2296.961, 2263.582, 2237.225, 
    2223.463, 2248.588, 2233.032, 2235.553, 2277.059, 2263.651, 2223.609, 
    2187.068, 2158.807, 1880.01, 1815.001, 1755.33, 1748.198, 1749.312, 
    1339.698, 1125.587, 1130.47, 59.49807, 58.49676, 34.96015, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20.62126, 22.37635, 
    2.40676, 0, 0, 0, 0, 0, 0, 0.3763808, 0.06727493, 0, 0, 0, 0, 0, 0, 
    1.019751, 2.639158, 2.465536, 52.71156, 81.86205, 82.00864, 181.3399, 
    181.5287, 148.4794, 98.42897, 102.4558, 69.96147, 59.10136, 63.99092, 
    40.4422, 42.56801, 32.82777, 0.0008582778, 2.874529, 19.54268, 23.23581, 
    36.82943, 39.30602, 35.5212, 45.80632, 48.78159, 51.29636, 100.3955, 
    182.744, 191.4607, 268.2026, 553.4864, 712.006, 911.4213, 1193.65, 
    1108.558, 1025.99, 516.4547, 46.01832, 8.978831, 0.2277288, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28.35638, 73.38754, 68.55959, 240.8364, 327.3661, 322.8138, 
    1005.626, 1011.71, 1159.311, 1449.092, 1477.573, 1406.121, 1412.553, 
    1462.306,
  590.6178, 662.6359, 1053.757, 1203.002, 1215.359, 1236.61, 1396.586, 
    1365.813, 1469.478, 1570.504, 1376.477, 1504.337, 1366.796, 1149.165, 
    1284.8, 1115.338, 937.6082, 997.0908, 879.6879, 840.0182, 1058.796, 
    1051.395, 907.0745, 1140.317, 1369.757, 1524.742, 1562.547, 1760.47, 
    1929.115, 1970.816, 2041.452, 2140.007, 2225.932, 2155.486, 2337.718, 
    2527.563, 2531.309, 2634.174, 2760.275, 2763.042, 2843.203, 2943.062, 
    2926.468, 2926.679, 2932.325, 2888.897, 2666.042, 2600.893, 2434.997, 
    2012.942, 1997.785, 1441.056, 1069.745, 990.5055, 237.4895, 174.5968, 
    492.6822, 786.6786, 796.4959, 1712.963, 1752.907, 2029.332, 2327.906, 
    2325.851, 2644.382, 2646.498, 2744.449, 2842.719, 2853.751, 2953.158, 
    2970.993, 3018.172, 3070.997, 3093.23, 3102.927, 3124.529, 3099.013, 
    3050.449, 3068.134, 2968.454, 2949.839, 2944.74, 2834.841, 2836.438, 
    2789.117, 2718.156, 2730.309, 2713.494, 2712.535, 2723.647, 2708.428, 
    2711.292, 2736.988, 2725.589, 2701.114, 2749.15, 2781.971, 2825.808, 
    2840.249, 2897.837, 2944.562, 2953.365, 2960.406, 2950.888, 2924, 
    2865.895, 2821.601, 2760.678, 2715.527, 2616.338, 2508.81, 2483.213, 
    2406.838, 2296.83, 2255.161, 2170.501, 2111.699, 2074.691, 2034.798, 
    1992.096, 1972.95, 2003.922, 1976.837, 2036.613, 2069.728, 2028.094, 
    1870.985, 1816.345, 1509.985, 1170.803, 1137.754, 1280.351, 1259.309, 
    1050.735, 851.3014, 843.5267, 48.9119, 49.71339, 25.8634, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18.57255, 34.3597, 33.47045, 
    66.53275, 68.30042, 44.87642, 17.8591, 19.10402, 1.153011, 0, 0, 0, 0, 0, 
    0, 2.055017e-05, 0, 0, 1.000033, 2.611686, 5.174166, 30.01795, 39.71861, 
    82.20617, 147.1211, 159.7841, 297.3846, 477.1503, 539.5934, 924.3657, 
    1200.882, 1219.114, 978.1096, 675.7386, 429.0988, 65.9558, 6.602714, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38.92105, 74.65038, 73.40634, 355.7201, 
    362.5836, 437.7601, 532.7929, 555.1108, 466.8683, 506.949, 544.5602,
  18.03429, 52.04677, 97.32604, 103.5047, 121.3791, 229.6428, 289.5833, 
    342.2204, 430.679, 294.0422, 329.4568, 258.2624, 261.7762, 387.8197, 
    266.1458, 186.9893, 177.8753, 116.2193, 164.0127, 190.8543, 51.08019, 
    53.65794, 238.8831, 401.6841, 578.6693, 627.7045, 834.0241, 1099.147, 
    1160.757, 1082.903, 1221.892, 1433.147, 1467.003, 1740.799, 2047.28, 
    2106.447, 2302.967, 2393.189, 2396.604, 2546.431, 2599.206, 2611.419, 
    2764.931, 2776.2, 2787.814, 2803.205, 2750.694, 2546.349, 2490.88, 
    2299.481, 2001.043, 1964.201, 1191.131, 1040.329, 585.9238, 81.64281, 
    121.023, 415.9229, 398.7615, 1034.832, 1279.398, 1481.982, 1885.691, 
    1879.85, 2344.911, 2348.394, 2481.111, 2557.897, 2590.554, 2659.466, 
    2675.679, 2736.939, 2765.516, 2808.543, 2848.058, 2865.266, 2830.327, 
    2850.584, 2767.783, 2736.893, 2738.699, 2667.121, 2688.131, 2636.5, 
    2593.343, 2597.347, 2548.82, 2566.686, 2557.27, 2501.946, 2529.648, 
    2480.124, 2446.396, 2457.965, 2458.898, 2486.558, 2557.4, 2560.002, 
    2602.271, 2683.407, 2703.591, 2677.501, 2701.365, 2740.708, 2688.588, 
    2665.173, 2652.263, 2636.06, 2602.061, 2563, 2515.804, 2421.467, 
    2332.681, 2240.587, 2081.742, 2017.474, 1935.613, 1823.498, 1753.269, 
    1667.035, 1600.693, 1582.375, 1615.339, 1579.295, 1683.731, 1637.395, 
    1413.076, 1159.486, 1028.147, 422.2416, 375.9933, 384.0838, 367.8711, 
    294.1305, 207.7352, 202.2109, 6.880322, 7.068289, 2.804695, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1409208, 12.76095, 41.41293, 95.15853, 
    269.8792, 339.5587, 509.6674, 851.3785, 1002.392, 1248.589, 1339.322, 
    1283.846, 609.3582, 112.4164, 13.00174, 3.752836, 0.1854097, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3.97741, 10.02372, 9.757164, 35.74642, 36.72299, 
    48.85838, 59.62074, 52.10133, 13.45668, 14.8341, 16.17722,
  0, 0, 0, 0.0006215409, 4.551234, 12.06382, 9.280968, 13.39801, 2.441525, 
    1.875412e-07, 0.02385139, 7.594793, 32.81744, 12.05854, 3.815145, 
    2.33419, 1.565117, 11.56645, 8.603318, 0, 0.1163873, 1.473388, 
    0.01854268, 0.0226858, 10.1976, 153.724, 318.8033, 283.3621, 321.8593, 
    438.466, 355.332, 323.099, 846.4395, 1358.309, 1529.359, 1875.661, 
    2002.336, 1929.218, 2064.169, 2088.292, 2186.29, 2380.477, 2387.384, 
    2522.057, 2542.292, 2515.692, 2469.048, 2363.97, 2224.501, 2174.826, 
    1896.399, 1687.671, 1461.676, 900.8322, 844.7673, 93.21449, 32.89951, 
    93.50941, 96.13092, 290.0595, 463.8329, 600.5393, 1159.744, 1151.958, 
    1823.603, 1829.568, 2067.961, 2146.225, 2213.968, 2277.84, 2307.905, 
    2358.55, 2399.041, 2498.373, 2540.624, 2562.839, 2588.514, 2551.211, 
    2493.715, 2498.203, 2419.907, 2454.006, 2448.446, 2442.482, 2432.917, 
    2371.105, 2382.124, 2305.938, 2272.796, 2244.818, 2108.124, 2146.387, 
    2113.27, 2035.82, 2122.081, 2164.428, 2159.731, 2237.652, 2327.44, 
    2372.029, 2385.987, 2392.022, 2378.246, 2337.616, 2402.123, 2459.168, 
    2432.999, 2477.983, 2493.586, 2443.446, 2377.018, 2327.428, 2188.934, 
    1953.658, 1816.67, 1587.998, 1436.788, 1362.995, 1281.63, 1166.738, 
    1068.912, 991.3848, 982.0762, 964.8165, 900.6691, 834.6942, 725.2911, 
    376.5895, 328.2077, 74.26664, 8.847977, 4.319468, 0.7749048, 0.5343943, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.207087, 2.702672, 1.804711, 0, 0, 0, 0, 0, 0, 
    0, 0, 5.863971e-05, 7.457768, 13.60514, 31.50537, 136.3042, 192.1596, 
    321.8073, 442.2468, 576.8663, 909.7634, 1210.569, 1054.537, 540.0894, 
    276.8775, 58.62088, 10.00244, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.622982e-05, 0.00443128, 0.0009650817, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6.320719e-06, 0.5922344, 42.28226, 72.99135, 
    58.22504, 23.60832, 0, 15.13064, 159.6497, 352.3127, 425.8737, 882.8994, 
    1143.479, 1185.229, 1303.212, 1210.182, 1387.859, 1710.169, 1774.273, 
    2005.944, 1937.508, 1959.549, 1922.148, 1782.9, 1701.266, 1567.828, 
    1515.942, 1410.279, 1271.513, 1184.542, 789.9104, 616.7271, 282.4797, 
    32.57191, 17.93108, 0, 10.67043, 34.54045, 84.44239, 436.1034, 429.6452, 
    1112.585, 1119.797, 1421.595, 1480.597, 1611.715, 1676.297, 1753.644, 
    1814.261, 1913.22, 2019.553, 2076.499, 2145.025, 2178.324, 2110.019, 
    2141.344, 2011.126, 2059.697, 2119.229, 2182.542, 2184.784, 2148.607, 
    2133.908, 1962.034, 1996.269, 1758.714, 1601.711, 1651.337, 1523.359, 
    1496.405, 1463.38, 1503.414, 1647.811, 1598.424, 1735.264, 1952.526, 
    1893.357, 1910.31, 2004.662, 1874.603, 1864.82, 2009.37, 2000.058, 
    2118.945, 2234.348, 2220.527, 2187.206, 2105.146, 1950.985, 1805.485, 
    1599.598, 1226.019, 1004.874, 743.4344, 581.7036, 530.5262, 473.8739, 
    365.8261, 279.0865, 180.4223, 124.5852, 73.62144, 24.38551, 5.817718, 
    2.254883, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.00148, 3.923336, 
    2.472864, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.008201447, 1.385557, 21.52813, 
    39.11131, 86.46773, 125.4521, 123.5826, 254.6765, 474.9824, 441.8616, 
    374.9601, 279.2499, 57.36595, 0.008567562, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9.531374, 57.01103, 56.65789, 183.2217, 292.1819, 
    289.4909, 483.7878, 573.3635, 762.7877, 1369.411, 1372.442, 1339.54, 
    1188.664, 1010.666, 813.2481, 702.388, 568.6976, 432.3323, 346.8519, 
    213.1217, 181.1843, 162.9754, 155.3973, 116.8555, 5.480179, 4.249075, 0, 
    0, 0, 2.821523, 64.81277, 62.71669, 254.9253, 264.6146, 478.9108, 
    516.3237, 715.197, 772.6674, 942.086, 1017.009, 1192.809, 1288.119, 
    1347.699, 1468.427, 1417.734, 1462.336, 1351.19, 1369.762, 1478.518, 
    1605.944, 1708.53, 1741.777, 1697.67, 1407.042, 1438.41, 1156.374, 
    1081.688, 1061.455, 917.9648, 844.9738, 574.6211, 656.8115, 691.1896, 
    557.1426, 783.5517, 964.7368, 1027.335, 1159.174, 1169.207, 1056.952, 
    1083.887, 1187.73, 1172.633, 1439.059, 1558.977, 1527.176, 1687.071, 
    1581.525, 1454.94, 1375.057, 1188.272, 952.3291, 719.2452, 352.9966, 
    176.3894, 41.06569, 14.55585, 13.81337, 11.61005, 10.02094, 7.039319, 
    2.973443, 0.009719314, 0, 0, 4.544891e-07, 0.0001139448, 0.0001361256, 
    5.083121e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.104511, 44.77611, 57.88408, 159.5562, 465.6332, 
    497.9623, 271.3645, 109.0002, 5.990397, 0.03503641, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4441628, 8.95208, 10.15624, 142.3696, 
    422.4524, 502.968, 847.0935, 779.0596, 455.1889, 229.5041, 56.95454, 
    13.12048, 14.70561, 10.83676, 21.24232, 7.490313, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.9525716, 3.126865, 43.4058, 54.01857, 115.984, 141.7184, 
    216.9358, 263.3754, 357.2512, 375.0049, 337.47, 313.6855, 277.1616, 
    361.28, 381.1482, 520.3611, 665.7684, 826.0345, 966.3919, 945.157, 
    605.7979, 692.4514, 228.8178, 169.3667, 418.4273, 522.0573, 508.7098, 
    338.3628, 237.395, 52.47231, 9.418461, 105.2781, 54.10379, 48.29434, 
    191.0345, 296.2173, 298.335, 203.916, 80.55537, 127.0886, 475.8766, 
    741.3522, 684.0757, 678.3928, 484.1764, 625.67, 551.395, 359.8978, 
    178.812, 119.3686, 157.2741, 92.74212, 14.00688, 1.705264, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.280546, 2.399927, 0.7897938, 0.01014344, 0.002112578, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4.133505, 42.84299, 141.7157, 338.8036, 553.8666, 472.5853, 242.1392, 
    41.90912, 17.81757, 6.743396, 0.3872084, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24.41029, 54.98615, 
    91.36515, 235.9627, 109.852, 8.360318, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.879204, 2.902804, 
    0.4108636, 9.802505, 16.66334, 22.53514, 29.24665, 38.96732, 50.45575, 
    83.07205, 85.1552, 108.0663, 23.45089, 0.0003052703, 25.01204, 92.55255, 
    94.70995, 74.12923, 77.00787, 3.042856, 0, 0.04883529, 0, 0, 0, 0, 0, 
    0.9142088, 2.677619, 0.7438642, 24.3284, 33.94885, 20.43999, 47.7958, 
    43.60358, 67.25209, 1.141844, 2.340516, 3.5237, 4.846861, 0.0003324859, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8787168, 1.860621, 0.7109822, 
    0.004783506, 0.001227291, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02883749, 2.894586, 137.5194, 
    356.6974, 523.2764, 390.2472, 214.6421, 50.61837, 0.09942365, 1.06244, 
    0.3060259, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06062585, 0, 0, 0, 0, 0, 0, 0, 0.2586277, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.158044, 11.94201, 94.69837, 227.4336, 280.281, 281.9613, 292.3566, 
    221.7773, 74.78673, 1.519979, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.579831, 
    23.88888, 106.4477, 140.1274, 136.5105, 139.0071, 99.59026, 55.47078, 
    5.571563, 0.04507341, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.941696, 
    8.889275, 16.29175, 22.22206, 13.32617, 3.939316, 7.839354, 7.839354, 
    0.4093648, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5170894, 7.169375, 15.67392, 10.90475, 4.613606, 4.510818, 3.992095, 
    0.3088567, 0, 0, 0, 0, 1.159464, 1.155876, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04463466, 2.521838, 1.437868, 1.386273, 2.431348, 0.04303304, 0, 0, 0, 
    0.268631, 9.553189, 7.673763, 0.00895416, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01503891, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2362988, 0.936215, 0.243221, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05594731, 2.646427, 1.423687, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03938901, 0.3163572, 0.3907959, 0.003227432, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1311353, 0.6234697, 
    0.8366612, 0.6355648, 0.0134637, 1.669041e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.707685e-06, 0, 0, 0, 
    0.09186153, 0.2376563, 0.3677765, 0.02923858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2720909, 0.3440705, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1702828, 2.740691, 
    21.26693, 127.9737, 51.16943, 7.951087, 1.411934, 0.0310415, 0.1596602, 
    0.01668881, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.8661806, 7.894113, 15.89043, 0.2572514, 0.0001458136, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -1.066399e-05, 0.5691465, 1.350524, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7447463, 0.9990342, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.457745, 12.13834, 202.4566, 257.557, 421.1448, 312.7731, 87.61121, 
    2.04354, 0.4918164, 0.2538341, 0.01294378, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 4.734055e-05, 4.426789e-05, 0.0001989858, 4.580274, 
    67.36448, 39.83454, 4.571144, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -2.817969e-05, -1.136271e-05, 0.0004287733, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01537742, 
    12.07182, 10.18145, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.02885614, 0.279215, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6624289, 9.918129, 213.1098, 291.8737, 
    276.2269, 180.1272, 82.33691, 2.251745, 0.526271, 0.03732056, 
    1.762412e-06, 0, 0, 0.000543329, 0.001995932, 0.0001191641, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.000220222, 0.0001886455, 0.1364876, 7.940151, 
    34.49795, 18.22237, 0.005200748, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.001930204, 0.3654139, 0.02615089, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1148066, 1.277598, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.01135122, 2.741379, 110.6423, 288.4021, 269.8642, 183.8733, 
    97.90216, 13.0034, 0.1822562, 0, 0, 2.499078e-05, 0.001790266, 1.14844, 
    0.5038718, 0.3242314, 0.02052839, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6377345, 4.380006, 0.4495623, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1836666, 9.321361, 
    94.07313, 426.8449, 394.5175, 231.4857, 91.63313, 5.877855, 0.0001054795, 
    0, 0, 0, 0.3998594, 2.582462, 3.550398, 0.9040038, 0.2424715, 
    0.004129146, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.7332023, 13.3652, 1.381984, 0.004339822, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4916189, 
    5.990397, 0.5141228, 0.0002272683, 0, 0, 0, 0, 0, 0, 0, 0.0003262791, 
    0.1033869, 0.001834185, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.9621782, 26.12735, 
    460.8656, 752.9393, 602.0097, 373.9108, 175.6023, 31.15347, 0.3345744, 0, 
    0, 0, 0.03500172, 0.06385407, 0.09471958, 0.08736823, 0.008385038, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.01587494, 20.58621, 77.93482, 15.25101, 0.6093944, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.2767738, 0.03358667, 0.0005778636, 0, 0, 0, 0, 0, 0, 0, 0.01824347, 
    0.2164043, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5495449, 158.7542, 555.2477, 
    967.3378, 719.9592, 450.8792, 230.1222, 108.553, 11.72476, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 14.79329, 27.28531, 10.04026, 0.3682708, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.585245e-05, 
    0.003155032, 0.0006623662, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2.153775, 91.42873, 458.1242, 897.1926, 940.429, 641.3556, 
    453.6378, 228.6973, 37.32151, 1.77637, 0.008350741, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.9845688, 4.140163, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4750706, 
    0.01123958, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0001734606, 3.209494, 8.408097, 3.203027, 0, 0, 0, 0, 0, 0, 
    0.0002626959, 0.0001242783, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1700168, 
    12.46845, 181.8088, 865.7809, 955.9866, 783.1808, 640.0667, 323.3945, 
    129.0697, 14.48532, 0.1598094, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.10743, 5.051364, 0.04059443, 0, 0, 0, 0, 0, 0, 0, 
    0.6077597, 2.885018, 4.573367, 0.9662914, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8.904971, 92.96897, 135.3427, 117.7756, 19.8626, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7158951, 9.649881, 
    268.7047, 840.7597, 953.1501, 696.6509, 503.0017, 263.5447, 36.45748, 
    0.6965974, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1835729, 0.3095913, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13.91417, 265.1042, 
    597.7688, 576.1215, 241.6265, 0.1444124, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.01391995, 3.326213, 108.2358, 613.186, 843.5461, 
    707.7412, 552.3075, 419.6042, 187.6315, 35.40749, 1.740049e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2003551, 
    2.067987, 0.05236836, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7842886, 
    26.15788, 524.2261, 918.0246, 644.9684, 73.27732, 2.588682, 0.003022553, 
    0, 0, 0, 0, 0, 0.05845414, 0.7972198, 0.8584681, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.7304063, 31.35818, 439.0558, 910.0109, 843.0219, 689.4072, 446.666, 
    306.8687, 151.1995, 3.599358, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8459378, 
    63.66971, 127.9097, 11.89414, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 14.02517, 440.8638, 619.5756, 477.8512, 110.7044, 2.002045, 0, 0, 0, 
    0, 0, 0.08374179, 1.813394, 2.268621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4190142, 
    8.151013, 347.1316, 881.4787, 925.9868, 775.559, 534.5961, 286.4486, 
    141.7835, 10.61713, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17.83841, 318.2258, 
    474.5805, 113.4041, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.321118, 124.8607, 677.453, 638.9067, 151.9681, 0.08658671, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003748207, 5.357027, 229.7243, 875.959, 
    947.0231, 1025.9, 946.106, 531.5417, 201.5818, 51.95796, 1.170505, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40.62353, 394.2583, 
    411.6251, 248.5301, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16.63172, 302.3406, 608.2631, 193.2175, 110.3051, 0.01421851, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16.2754, 304.9714, 992.2845, 1139.245, 
    1108.48, 1077.206, 793.1174, 340.5469, 34.45227, 1.693283, 0.1668559, 
    0.0008615133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005833376, 
    0.03323527, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02824904, 15.43679, 
    72.92188, 9.112865, 4.911317, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6.593254, 22.48983, 29.3053, 237.9958, 12.88725, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29.44415, 323.9431, 937.9124, 1022.014, 
    990.0472, 822.2456, 450.804, 183.3924, 58.91031, 35.09547, 5.725437, 
    0.01405082, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03905309, 
    2.225024, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01800254, 0.01278392, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.05530041, 0.6063908, 0.2314757, 1.179664, 1.383117, 0.326624, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.260805, 165.5909, 
    554.0589, 321.4837, 22.20998, 0.005874773, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14.88112, 212.311, 867.2741, 1115.777, 666.8633, 561.7639, 
    255.8239, 177.912, 109.9881, 44.05696, 6.909386, 7.52843, 0.05320534, 
    0.0173502, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5460697, 0.3825809, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.988424, 
    38.65697, 98.13758, 54.36794, 97.04861, 72.65929, 27.73439, 5.29118, 
    0.0002478067, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.6329815, 93.92059, 407.5471, 458.3563, 232.0045, 0.749948, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 35.06068, 255.3221, 830.9753, 1274.318, 745.7563, 
    458.187, 289.5876, 232.1219, 152.137, 113.2261, 156.948, 117.146, 
    63.54305, 20.7716, 0.5308164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.349678, 0.2319917, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.767381e-05, 
    6.239011e-06, 0.4817159, 52.69125, 170.5017, 279.2373, 297.8989, 
    386.1169, 552.4821, 474.2657, 235.7939, 5.684123, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.951542, 154.6919, 163.3024, 163.2682, 
    1.700415, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33.58019, 289.0226, 
    802.3174, 1488.865, 1018.361, 595.573, 304.1579, 277.8465, 206.8251, 
    169.4075, 230.656, 201.0125, 170.5851, 78.90333, 6.181812, 0.03314363, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.747797, 1.918709, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2870086, 0.2879882, 4.695856, 
    76.30035, 153.5668, 170.7645, 193.2896, 268.4077, 530.8789, 862.7049, 
    601.2026, 26.08447, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.175502, 2.391562, 36.16692, 0.04562337, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.3355515, 79.2103, 593.8276, 1900.202, 1630.975, 913.8342, 
    346.4595, 308.5696, 206.9561, 123.7278, 122.4443, 117.0263, 90.11703, 
    26.39464, 1.810491, 0.01115009, 4.265336e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.777052, 0.5013778, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04850387, 0.6324823, 0.9992909, 
    0.01875544, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3.789136, 3.629767, 14.17716, 0, 0, 0.0001789696, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.005426887, 0.1459763, 1.738111, 26.18267, 
    84.66904, 84.72141, 84.63051, 79.82909, 87.23138, 113.6659, 263.565, 
    665.0464, 726.6257, 221.1805, 1.070413, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.02665801, 0.3924785, 0.9974071, 0.4957287, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60.10113, 321.6766, 1886.564, 1899.45, 
    979.9465, 389.7755, 329.0944, 200.0761, 114.2748, 89.23959, 68.02219, 
    40.1021, 15.32402, 3.227205, 1.124794, 0.806437, 0.1284226, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19.63962, 216.7453, 151.3867, 
    49.05574, 85.18954, 72.99554, 4.173137, 1.189671, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5391172, 85.40571, 175.1282, 
    176.2003, 51.98185, 16.16949, 16.46254, 3.358395, 0.1506761, 0, 0, 0, 0, 
    0, 0, 0, 0.1716822, 12.57517, 14.97444, 110.2753, 151.8983, 60.78812, 
    58.35716, 67.02755, 80.66826, 119.3769, 210.6807, 426.7547, 662.723, 
    320.195, 6.133488, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002032076, 0.1506091, 0.5290205, 0.1990197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.4204397, 0.6064368, 0.03898298, 0.001524889, 0, 0, 0, 0.7833207, 
    150.2995, 1699.418, 2189.595, 826.324, 451.2817, 417.6789, 222.0445, 
    128.3999, 100.2722, 66.89939, 33.19941, 23.58981, 46.86787, 80.45917, 
    58.24134, 3.721146, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.10063, 89.40348, 596.3478, 
    666.8564, 591.394, 652.2402, 595.1525, 318.677, 170.95, 6.403108, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2061634, 
    87.07784, 287.6782, 304.671, 277.0926, 190.0759, 152.187, 123.9766, 
    40.03922, 0.5552845, 0.002972871, 0, 0, 0, 4.596487e-07, 0.001911092, 
    7.618953, 103.1634, 136.5377, 208.5589, 252.9298, 95.60206, 63.75122, 
    72.34969, 89.18761, 141.7349, 218.1745, 347.6282, 679.1434, 422.4627, 
    43.80862, 0.2143922, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005062858, 
    0.01175183, 0.0144366, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.230724, 
    0.4888345, 0.1494787, 0.01307711, 0, 0, 0, 0, 99.18201, 1628.889, 
    2441.639, 775.515, 602.6862, 706.2284, 361.2233, 150.8217, 101.9297, 
    55.58748, 21.88517, 40.12035, 96.79882, 143.1583, 86.97305, 10.69366, 
    0.03930662, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03612367, 117.1902, 662.0591, 
    1051.479, 1007.953, 1004.66, 980.3722, 981.061, 904.6642, 469.5939, 
    77.86052, 0.07097008, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 62.64774, 289.7885, 322.4895, 372.0777, 333.6976, 287.9106, 
    232.7851, 138.0785, 38.58958, 24.01395, 5.46848, 1.235958, 0.440236, 
    5.436836, 11.19636, 63.98316, 168.1433, 164.1105, 259.0268, 333.079, 
    178.0129, 116.8504, 82.8353, 105.1621, 192.135, 247.4189, 314.4903, 
    541.7823, 424.2846, 200.4327, 17.4241, 0, 0, 0, 0, 0.0025757, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 46.98773, 1925.962, 2519.025, 824.3611, 572.7868, 814.8135, 
    624.4693, 189.6015, 94.57539, 48.08117, 40.39698, 46.90089, 112.1453, 
    132.2464, 118.2398, 64.30252, 5.560091, 0.05948743, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.885378, 157.7066, 675.8417, 
    1117.676, 1272.397, 1313.217, 1368.889, 1377.063, 1480.051, 1201.435, 
    479.6372, 33.34804, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 89.37342, 269.4676, 328.312, 396.2931, 412.5576, 339.3434, 284.8559, 
    184.8258, 142.0229, 126.5364, 99.82055, 90.46408, 51.68258, 73.10482, 
    93.4927, 137.1221, 151.5809, 117.0362, 193.748, 230.3193, 124.6491, 
    172.9935, 124.9841, 117.9316, 206.8239, 207.5924, 226.6611, 424.3082, 
    559.7695, 577.7419, 59.06447, 0, 0, 0, 0.008436895, 0.07163155, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009679735, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 318.5692, 2255.52, 2513.303, 1105.152, 568.3367, 
    624.6456, 715.6223, 192.3756, 93.49286, 44.98126, 59.40482, 60.02718, 
    146.5208, 176.3745, 174.6166, 189.9253, 58.50751, 1.392609, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001397563, 64.73356, 486.5651, 
    831.4321, 988.1431, 1093.073, 1183.692, 1312.665, 1439.21, 1578.132, 
    1870.992, 1283.831, 279.1647, 0.227633, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.165965, 183.222, 307.0978, 371.689, 421.8028, 
    429.675, 375.4235, 346.1321, 251.7014, 200.066, 204.2942, 186.1086, 
    160.2067, 125.7472, 140.6481, 166.7921, 158.4811, 148.7925, 106.7582, 
    172.5229, 180.4118, 75.12927, 142.5373, 133.1286, 116.0215, 140.7905, 
    145.5771, 163.8873, 308.2479, 600.6851, 801.6199, 160.0717, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.07666183, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 218.2384, 2279.855, 2839.516, 1308.155, 
    679.2444, 435.8649, 535.561, 172.0074, 83.86958, 48.27812, 47.01646, 
    65.52027, 123.0483, 178.9258, 187.4919, 188.2097, 107.9868, 41.37278, 
    0.3784643, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.514285, 178.8383, 691.333, 923.7204, 
    910.9808, 994.0078, 1125.025, 1179.335, 1349.513, 1537.688, 2109.614, 
    1828.657, 753.7578, 48.34106, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0003535612, 4.018133, 220.7036, 323.4764, 391.5331, 445.5506, 
    424.8635, 399.0803, 419.7336, 352.2723, 236.0119, 237.668, 234.9762, 
    225.463, 221.0029, 215.0713, 196.4316, 170.674, 140.3396, 59.97283, 
    73.19926, 80.22798, 74.48715, 129.4444, 123.8968, 127.8858, 132.3327, 
    133.4457, 142.8761, 212.4393, 470.5186, 745.779, 214.3459, 0.004355592, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1931676, 0.04965259, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3005273, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28.39257, 2161.471, 
    3381.285, 1917.059, 865.7023, 361.1256, 247.1886, 171.3001, 76.89898, 
    58.85208, 47.25829, 68.28066, 77.07005, 132.0991, 230.509, 273.0426, 
    279.8915, 377.0726, 78.64452, 1.101563, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 78.93523, 361.0667, 748.3067, 802.6099, 
    848.2653, 995.7048, 1271.416, 1228.839, 1278.11, 1427.784, 1741.449, 
    1711.395, 1021.674, 263.7831, 3.604623, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.3091095, 62.91591, 262.8626, 359.8786, 428.4573, 464.3272, 
    444.5198, 456.5864, 458.874, 407.2716, 331.4111, 339.2321, 337.7972, 
    341.2208, 332.7867, 310.8422, 250.8219, 206.4852, 109.0646, 26.69283, 
    15.96027, 33.70029, 66.94215, 115.2257, 131.5484, 160.6219, 170.2549, 
    165.9246, 174.7384, 208.2959, 332.4551, 538.7546, 197.9195, 0.0467078, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03266417, 0.007956498, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.05223094, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.03820974, 3.000286e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    10.74888, 1458.088, 3761.399, 2842.54, 1377.383, 739.4715, 234.4863, 
    132.0681, 87.18903, 63.88172, 54.47548, 65.4408, 73.71259, 123.355, 
    301.8839, 456.0324, 642.2784, 831.5916, 502.9808, 46.96783, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1894609, 418.4838, 871.1957, 944.6196, 
    945.7229, 869.4675, 984.9916, 1245.592, 1329.606, 1314.505, 1383.642, 
    1568.032, 1653.743, 1231.111, 407.7769, 18.08652, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6.653165e-05, 1.288491, 120.8556, 288.922, 392.183, 
    463.0468, 512.4948, 502.8403, 505.3195, 486.4092, 438.4559, 418.7603, 
    435.1577, 410.1254, 448.9712, 457.8134, 443.2514, 354.0945, 247.9053, 
    115.4568, 37.08583, 22.25363, 35.5222, 66.02837, 112.9075, 151.6104, 
    193.8575, 226.7909, 241.7822, 263.8828, 272.1542, 333.3326, 406.1204, 
    127.5017, 0.002632135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.2783271, 1.544159e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3022502, 0.7625732, 
    0.08615553, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.2726899, 909.5847, 3485.945, 3723.64, 2286.165, 
    1088.172, 277.8031, 151.8562, 122.7472, 79.85472, 63.51342, 63.70974, 
    85.95111, 162.5309, 324.9848, 487.1127, 730.7104, 928.7892, 595.827, 
    66.51587, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.069803, 624.4039, 1194.453, 1049.597, 
    1010.534, 921.7643, 963.5883, 1094.983, 1237.806, 1373.928, 1436.614, 
    1526.442, 1628.834, 1320.716, 393.8683, 19.00888, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.2321375, 0.02614409, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002468355, 1.555462, 85.69622, 
    270.489, 386.5388, 475.1803, 554.0732, 544.3365, 507.5302, 474.027, 
    450.6302, 448.1553, 469.2498, 486.3567, 584.0611, 613.5104, 582.1614, 
    460.8552, 290.631, 134.3587, 59.36531, 29.1989, 40.18928, 80.37932, 
    123.9354, 169.0607, 235.5126, 302.9901, 378.7519, 401.5203, 324.3041, 
    343.4445, 338.9859, 43.72432, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1740191, 0.3604606, 
    0.02819098, 0, 0.0001089571, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.02784524, 0.01332446, 0, 0, 0, 0, 0, 0, 622.9456, 3109.44, 
    4187.303, 3544.686, 1933.761, 441.2773, 201.7201, 157.0204, 107.1256, 
    78.66496, 65.35883, 117.1102, 204.9081, 355.1263, 573.7363, 935.9915, 
    916.3714, 554.4952, 68.27861, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16.53199, 768.9169, 1331.36, 1136.01, 
    1044.142, 995.5248, 1005.116, 1045.59, 1132.859, 1244.613, 1249.77, 
    1275.452, 1411.149, 1230.043, 355.7857, 38.42538, 11.36239, 0.1664333, 0, 
    0, 0, 0, 0, 0, 8.918203, 63.82284, 32.24533, 0.06845794, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002621257, 4.873797, 70.57458, 244.3705, 390.5649, 484.1496, 569.4086, 
    573.7692, 519.7415, 463.3563, 454.0973, 452.4254, 485.5903, 558.1556, 
    658.0222, 615.2677, 554.7277, 466.9654, 315.5821, 167.0048, 102.4408, 
    55.8221, 63.31611, 90.15622, 132.1443, 174.2476, 271.2532, 361.4143, 
    476.5542, 499.5148, 344.0411, 301.3713, 206.5754, 16.46008, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.01711944, 0.00622351, 0.003869146, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.311946e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0172474, 0.01136346, 0, 0, 0, 0, 0, 
    0, 382.8545, 2876.062, 4165.984, 3891.626, 2193.506, 607.6644, 242.2492, 
    172.8224, 125.3955, 95.70429, 75.37946, 140.6825, 238.058, 330.3408, 
    590.7173, 860.9318, 892.1171, 743.56, 130.7965, 2.388815, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 149.1542, 863.8923, 1386.298, 1222.701, 
    1141.65, 1102.65, 1092.354, 1075.796, 1116.129, 1109.456, 1022.57, 
    1177.949, 1161.804, 873.0604, 292.4129, 58.97485, 65.39774, 20.34796, 0, 
    0, 0, 0, 0, 1.710002, 179.1329, 361.7984, 462.2877, 4.185929, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002116192, 8.215295, 93.8396, 260.59, 396.9593, 492.264, 583.0269, 
    577.7393, 511.6616, 437.3181, 434.9788, 429.9127, 447.5896, 503.0964, 
    535.1639, 550.9879, 601.609, 533.6042, 408.2331, 247.6928, 156.6912, 
    95.288, 89.71935, 107.4393, 162.3367, 192.1965, 249.0505, 356.6118, 
    472.8666, 420.214, 277.4969, 241.9379, 120.1581, 5.656234, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05569103, 
    0.007873038, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002160446, 0.01524386, 
    0.01595653, 0.07471912, 0, 8.891283e-05, 0.0005039916, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 313.1699, 2450.393, 3771.613, 
    4009.91, 2647.487, 747.3575, 248.2146, 179.1539, 139.321, 109.0235, 
    82.54051, 126.2465, 250.5499, 341.3198, 477.3122, 682.464, 790.146, 
    777.675, 402.0463, 142.8018, 12.9641, 0.1612704, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 206.0882, 905.4355, 1492.06, 1352.789, 
    1274.61, 1207.498, 1153.37, 1094.322, 1066.59, 1079.198, 961.5387, 
    988.6851, 1025.991, 624.6832, 253.0147, 89.52007, 93.68048, 55.51164, 0, 
    0, 0, 0.0003273949, 0, 16.96347, 324.5697, 698.6456, 671.6307, 10.65277, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10.21097, 82.69306, 241.7677, 373.667, 525.0147, 590.1464, 
    539.6522, 457.6314, 373.2543, 391.3733, 389.4047, 410.9097, 447.8246, 
    477.1811, 592.577, 672.8408, 655.7264, 580.9046, 373.312, 230.2575, 
    152.8479, 129.1694, 142.0154, 175.9838, 214.094, 232.5521, 319.338, 
    369.7514, 272.0832, 169.7341, 75.59463, 3.838568, 0.004566191, 
    1.067821e-05, 1.803288e-05, 0, 0, 0, 0, 0, 0, 0, 0.01736655, 0.05717497, 
    0.02134362, 0.0003499125, 0.0001778217, 0.0008473143, 0.0002311722, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.852015e-06, 0.0005623066, 0.0009736617, 0.06533751, 0.02656565, 
    0.007943218, 0, 0, 0, 0, 0, 0, 0.0004043824, 0.001626686, 0.01220574, 
    0.08809307, 0, 0.000279937, 0.0003478193, 0, 0, 0, 8.663214e-06, 
    9.113139e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    248.9795, 1963.14, 3415.902, 4186.658, 3366.991, 897.4039, 249.4845, 
    192.3507, 152.2305, 115.1808, 90.19453, 160.9946, 318.3405, 337.7122, 
    380.7813, 516.6271, 602.3742, 639.9847, 624.5349, 639.9632, 438.9142, 
    272.7673, 44.73225, 5.146412, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.081696, 245.6028, 968.4772, 1535.874, 
    1536.646, 1396.359, 1235.617, 1136.242, 1031.815, 1013.401, 1089.909, 
    1051.364, 839.1882, 732.7265, 540.6644, 288.8536, 128.5742, 129.3381, 
    30.40051, 0, 0, 0.003471407, 0.01092446, 0, 99.00717, 429.6659, 765.282, 
    735.4365, 56.52505, 0, 0, 0, 0, 0.0009473734, 0.00745804, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.557781, 26.37342, 
    154.109, 402.0398, 565.1448, 510.6704, 452.9216, 389.1734, 315.1229, 
    333.6582, 362.3361, 396.6921, 402.651, 423.4743, 540.3842, 621.2191, 
    623.5266, 571.3902, 417.0475, 279.7386, 195.6605, 196.6405, 220.1435, 
    202.9082, 225.1523, 246.4414, 297.0576, 298.4344, 254.6906, 142.7628, 
    35.38766, 0.2406005, 2.410453e-05, 4.678628e-05, 3.603175e-05, 0, 0, 0, 
    0, 0, 0, 0.02738773, 0.7861398, 1.237422, 0.1430842, 0.007873153, 
    0.0005202456, 0.002570945, 0.0007618599, 0, 0, 0, 0, 0, 0, 0, 
    0.004309868, 0.007082606, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01432367, 
    0.01865591, 0.1351462, 0, 0, 0.0009616442, 0.01069677, 0.04506977, 
    0.09431192, 0.03692892, 0, 0, 0, 0, 0, 0, 5.379522e-05, 0.001917429, 
    0.0009913536, 0.0008271347, 0.008883133, 0.03388457, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 223.7495, 
    1953.551, 3660.128, 4345.27, 3703.139, 1291.774, 338.182, 216.5628, 
    163.2808, 117.8495, 105.1776, 225.6686, 420.6713, 350.7291, 333.3784, 
    388.3565, 468.8985, 556.2679, 625.6486, 830.5468, 973.2249, 764.7795, 
    458.0817, 143.6824, 3.06489, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 63.22075, 447.4166, 1123.125, 1474.772, 
    1519.456, 1404.536, 1225.526, 1118.053, 1005.884, 968.1827, 1014.392, 
    1051.521, 920.0976, 754.5247, 560.9785, 369.7255, 195.4297, 111.9998, 
    1.897617, 0, 0, 0, 0, 0, 30.42347, 262.1609, 608.1423, 1003.023, 
    184.9282, 0.4479533, 0, 0, 0, 0.0320581, 0.2066001, 0.0002376924, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01763733, 
    1.009019, 57.72128, 239.9636, 295.133, 293.6826, 317.2214, 300.0989, 
    286.7005, 311.7386, 339.3264, 382.7134, 380.3221, 399.5885, 471.2103, 
    513.2486, 497.9005, 460.0551, 369.7978, 266.9686, 212.3264, 293.0757, 
    277.8092, 196.2818, 231.2053, 315.2725, 320.841, 263.2466, 301.713, 
    128.7204, 0.2290849, 0.002320653, 6.842137e-05, 0.0002180163, 
    1.34197e-05, 0, 0, 0, 0, 0, 0, 0.4746329, 2.654137, 3.062384, 0.2586081, 
    0.01649346, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008811429, 9.63827e-05, 
    0.001782605, 0.4635037, 0.2798483, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0826657, 0.2926077, 0.07386908, 0, 0, 0.0004918269, 0, 0.02177816, 
    0.08921915, 0, 0, 0, 0, 0, 0.001058054, 0, 0.004293167, 0.001877439, 
    0.0007863464, 0.004625599, 0.01026416, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 188.8455, 2042.651, 
    3833.509, 4083.839, 3578.691, 1705.318, 539.9378, 257.6141, 170.6759, 
    118.6289, 106.4746, 281.8179, 391.9007, 387.6766, 370.0793, 352.657, 
    412.1588, 482.489, 605.4061, 851.1165, 966.4521, 948.9276, 718.8047, 
    279.4622, 54.37357, 0.6717988, 0, 0, 0, 0, 0, 0, 0, 0.005348207, 
    0.004198826, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 1.668972, 216.3955, 749.1286, 1181.931, 
    1425.453, 1380.386, 1286.105, 1125.671, 1005.855, 968.5856, 939.8107, 
    935.4818, 1041.838, 1177.268, 1077.743, 872.0697, 633.3443, 405.0339, 
    84.63959, 0.106948, 0, 0, 0, 0, 0, 1.386793, 105.6473, 545.3414, 
    1230.705, 485.1578, 8.365142, 0, 0, 0, 0.06630934, 0.3088309, 0.3657435, 
    0.1342976, 0, 0, 0, 0.4603773, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5.671914, 41.4291, 42.15157, 94.58195, 156.2347, 204.9556, 
    231.9005, 278.6586, 284.6802, 324.2, 364.0796, 388.0253, 390.4885, 
    386.5884, 371.7647, 383.3232, 309.1913, 248.2855, 244.372, 312.1449, 
    205.5524, 149.9717, 267.6299, 489.7645, 398.223, 240.6597, 198.9537, 
    8.701391, 0.006575745, 0, 2.856021e-05, 0.0001477387, 0, 0, 0, 0, 0, 0, 
    0.05834794, 1.331946, 1.199006, 0.256244, 0.1441629, 0.4216602, 
    0.02553727, 0, 0, 0, 0, 0, 0, 0.004988394, 0.01328979, 0.001315807, 0, 
    0.5707712, 0.4010023, 0.003105322, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02868333, 
    0.1114157, 0.002806145, 0.02299087, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001548231, 
    0.004198918, 0.00378691, 0, 0, 0.004006569, 0.004596448, 0.002391663, 
    0.001764931, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 200.5349, 2205.909, 3754.746, 3880.177, 3527.569, 
    1961.977, 721.6547, 336.5783, 192.6983, 123.5193, 93.65848, 194.1664, 
    280.7815, 462.5269, 428.2898, 372.8152, 406.7669, 484.9255, 633.3601, 
    898.6265, 872.9783, 907.5272, 751.6215, 631.5092, 271.749, 15.36807, 0, 
    0, 0, 0, 0, 0, 0, 0.02276951, 0.01253423, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 59.34797, 545.6973, 1021.1, 1196.811, 1304.559, 
    1314.177, 1216.361, 1126.031, 1004.464, 951.8962, 953.8419, 978.6846, 
    1009.668, 1149.911, 1275.21, 1242.173, 1030.044, 672.7522, 125.4332, 
    12.55386, 0.2692544, 0, 0, 0, 0, 0.001992823, 56.98149, 572.5043, 
    1344.431, 813.0041, 78.45969, 0, 0, 0, 0, 0, 0.1177232, 0.04211174, 0, 0, 
    0, 0.4466666, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003872079, 0.0524085, 0.01861755, 4.812591, 32.89614, 82.01479, 
    163.1112, 188.6211, 216.5176, 306.168, 367.2151, 404.4103, 353.7346, 
    294.749, 290.3604, 295.2501, 241.0304, 244.4243, 254.7502, 206.8943, 
    103.8301, 133.0215, 376.4355, 631.4564, 449.5743, 164.1917, 19.29567, 
    0.002406351, 0, 0, 0, 0, 0, 0, 0.0002727428, 0, 0, 0, 0.2035922, 
    0.3194466, 0, 0, 0, 1.336402, 0.04671611, 0, 0, 0, 0, 0.05879996, 
    0.2017837, 0.1024817, 0.0489494, 0.08602279, 0, 0.3418902, 0.2794547, 
    0.008365069, 0, 0.1863148, 0.07948165, 0, 0, 0, 0, 0, 0, 0.005171813, 
    0.01600509, 0.08009271, 0.005973219, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.220226e-05, 0.0007515773, 2.540459e-05, 0.001626681, 0.004254468, 
    0.002696703, 0.001008588, 0.0001575875, 0.0002195451, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 306.8601, 
    2693.796, 3824.856, 3917.359, 3529.92, 2131.154, 768.7119, 364.644, 
    258.3862, 178.2268, 114.5725, 116.2875, 185.0063, 476.3114, 511.8191, 
    486.7108, 453.4619, 558.2297, 752.1304, 959.8199, 797.8405, 805.2585, 
    739.6364, 492.9413, 275.0653, 26.4997, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 160.6064, 882.3549, 1162.796, 1129.222, 
    1130.997, 1170.312, 1162.814, 1105.061, 1025.301, 965.5159, 965.4726, 
    1006.815, 955.4867, 1029.395, 1119.532, 1314.683, 1294.268, 849.2126, 
    257.5528, 56.19818, 4.743866, 0.02761184, 0, 0, 0, 0.03248502, 143.1412, 
    668.9073, 1128.408, 933.5784, 240.1967, 0.88444, 0, 0, 0, 0, 0, 
    0.0002821074, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2582259, 42.83031, 127.9336, 119.5595, 185.465, 
    324.0564, 385.4601, 395.1321, 335.8682, 249.0504, 248.3894, 240.1774, 
    225.6175, 266.7238, 199.9953, 82.14463, 40.2777, 101.211, 298.5282, 
    541.8779, 402.6116, 40.36655, 0.2139159, 0, 0, 0, 0, 0, 0, 0, 
    5.373165e-06, 0, 0, 0, 0.000217319, 6.01968e-06, 0, 0, 0.2650951, 
    1.019112, 0, 0, 0, 0, 0.002198522, 0.3068771, 0.9770192, 0.3985396, 
    0.4019007, 0.1162169, 0, 0.06322376, 0.3621572, 0.05163841, 0, 0.5162622, 
    0.3049748, 0, 0, 0, 0.0001316561, 0.0005437847, 0, 0.002817692, 
    0.01354941, 0.001151136, 0, 0, 0, 0, 0.0007822034, 0.3503827, 2.89994, 
    0.009312551, 0.001338001, 0, 0, 0.00153209, 0.008564333, 0.01470851, 
    0.002413101, 0.001395677, 0.005249981, 0.00108064, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.706651, 
    514.3159, 3265.038, 3949.23, 3804.174, 3124.612, 1830.161, 670.9692, 
    324.3877, 339.7944, 284.3907, 182.9888, 111.2254, 148.5408, 401.9024, 
    640.1982, 641.5475, 561.7526, 610.8893, 786.5002, 855.7067, 748.66, 
    801.2665, 821.2248, 452.3961, 237.3811, 24.96506, 2.785639e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 424.7021, 1039.75, 1141.513, 1117.404, 1139.51, 
    1153.328, 1141.572, 1100.598, 1039.432, 998.369, 985.0875, 1045.073, 
    944.1666, 808.9749, 1002.354, 1235.806, 1154.99, 756.4064, 317.3525, 
    147.2696, 87.65554, 20.40592, 3.579888, 0, 0.000175195, 0.1095807, 
    140.5684, 464.1875, 625.594, 842.4777, 315.3376, 3.185327, 0, 0, 0, 0, 0, 
    3.164616e-05, 0.000545998, 7.190741e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003644392, 9.271911, 58.43213, 
    85.59987, 275.9697, 419.9669, 377.0512, 320.8733, 281.7533, 223.175, 
    235.4737, 237.4207, 241.1763, 229.585, 114.4579, 19.47482, 7.417144, 
    60.78455, 184.0048, 445.5703, 386.9784, 6.37737, 7.911539e-06, 
    0.0001689458, 8.628888e-05, 0, 0, 0, 3.182994e-05, 1.884119e-05, 0, 0, 0, 
    0, 3.950985e-05, 1.088194e-06, 0, 0.05533992, 0.9281242, 0.2273573, 0, 0, 
    0, 0, 0.006392346, 0.3372472, 0.7412739, 0.9412045, 0.5059027, 
    0.03487262, 0, 0, 0.1156928, 0.0231991, 0, 0, 0, 0, 0, 0, 0.0001576808, 
    0.0008927984, 0, 0, 0, 0, 0, 0, 0.0004816438, 0.000904039, 0.08648013, 
    0.5848449, 29.86509, 0.007331183, 0.001859789, 0.02298578, 0.003762891, 
    0.007122362, 0.006248528, 0.008012623, 0, 0.006553994, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01637446, 
    15.59363, 288.1043, 2023.704, 3927.666, 3956.127, 3483.344, 2494.916, 
    1075.257, 457.6613, 303.1644, 331.8053, 274.7975, 162.8466, 115.3191, 
    152.0384, 448.9722, 690.0363, 750.97, 651.7511, 669.7906, 797.7618, 
    746.9589, 664.2542, 752.8363, 826.8702, 584.7307, 340.8673, 88.10323, 
    0.0003057911, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 139.7007, 878.0717, 1161.137, 1157.316, 
    1191.586, 1196.701, 1185.213, 1131.527, 1051.287, 1026.153, 1071.549, 
    1090.193, 1101.081, 841.0447, 825.4402, 863.6016, 743.7269, 441.5237, 
    290.1812, 418.6487, 338.2615, 195.0542, 63.64782, 1.233794, 0.002424632, 
    0.02704389, 39.07079, 142.9925, 210.215, 616.2933, 488.3251, 57.3394, 0, 
    0, 0.0002915235, 0, 0, 0.0001187494, 0.001512473, 0.0001085015, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1957919, 
    21.82922, 103.8146, 394.6642, 455.5143, 285.3593, 191.844, 198.3348, 
    211.5676, 234.2803, 232.0327, 149.2595, 95.75577, 29.65902, 2.123153, 
    2.030516, 36.09526, 125.5197, 347.8274, 303.9944, 0.2987032, 
    2.795298e-05, 0.0004210524, 0.0001467324, 0, 0, 0, 3.629953e-06, 
    1.339359e-06, 0, 0, 0, 0, 0, 0, 0.004245521, 0.3670297, 1.474632, 
    0.3125433, 0, 0, 0, 0, 0.002137339, 0.115092, 0.5954696, 2.117683, 
    0.7633625, 0, 0, 0, 0.04522271, 0.007462858, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.003122849, 0.0009074097, 1.505878, 1.775292, 0.01853255, 
    0.02877364, 0.006427244, 0.0183768, 0.01764533, 0.009966639, 0.005118342, 
    0.004092733, 0.003947109, 1.161786e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 143.6156, 1006.928, 
    2008.783, 3838.906, 4155.401, 3461.32, 2143.492, 932.2435, 306.7647, 
    274.221, 388.409, 342.5102, 239.047, 148.9487, 141.3877, 234.3398, 
    466.6049, 572.747, 561.063, 573.8524, 791.7665, 905.1641, 782.4678, 
    628.8995, 690.347, 777.0225, 675.2941, 482.3146, 161.034, 0.01123264, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.9148086, 0.1960665, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 92.40324, 783.9673, 1253.813, 1257.313, 1306.73, 
    1290.295, 1238.698, 1167.349, 1070.49, 1047.921, 1122.583, 1132.982, 
    1089.235, 1047.785, 778.2995, 623.4105, 614.2996, 535.6914, 652.0543, 
    703.6795, 664.7524, 473.676, 240.2652, 49.35349, 0.1625683, 1.082343e-05, 
    0.5136233, 10.08208, 36.63795, 363.2193, 600.5404, 92.53114, 0, 0, 
    9.762146e-05, 0, 0, 1.697265e-05, 0.0002031709, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4342294, 
    38.95743, 331.2641, 342.6676, 152.6043, 92.58819, 142.8874, 188.0837, 
    185.9535, 135.5564, 53.18517, 15.3731, 0.4312218, 0.005795754, 1.153572, 
    30.31803, 112.1737, 154.7345, 39.21417, 5.682861e-07, 0, 1.167903e-05, 
    1.955601e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1315296, 1.049161, 
    2.866518, 0.5865215, 0, 0, 0, 0, 0, 0, 0, 0.007800326, 0.003875447, 
    0.06003619, 0.05264203, 0.09403974, 0.01410556, 0.002335062, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002055086, 0, 0.001824039, 7.747502e-05, 
    0.01908099, 0.07046012, 0.0281525, 0.02594023, 0.006462191, 0.001722018, 
    0.00428438, 0.001929154, 0.00182072, 0.0006521175, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6945149, 40.65553, 
    1518.492, 3164.02, 3909.127, 4350.673, 3766.611, 2197.368, 717.933, 
    245.9577, 174.4986, 248.3382, 328.324, 276.2947, 309.8626, 268.0678, 
    269.3501, 385.1758, 547.7411, 477.9313, 365.31, 424.3435, 708.3638, 
    872.3875, 806.0463, 696.9042, 618.964, 689.5978, 760.7966, 561.5822, 
    192.7178, 0.02185223, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.702187, 0.3834732, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 97.44191, 816.2964, 1332.494, 1420.212, 
    1465.397, 1414.752, 1305.217, 1210.457, 1097.196, 1058.122, 1132.157, 
    1166.029, 1153.446, 1139.031, 996.1191, 774.9492, 880.2678, 931.6177, 
    997.2878, 745.6705, 665.7014, 530.7267, 349.6855, 90.39388, 0.2572696, 0, 
    0, 0.01589896, 1.590077, 406.1989, 774.4727, 99.39961, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6.797702e-08, 1.072985, 98.37104, 160.9242, 41.99627, 23.93826, 
    124.2789, 160.5256, 190.5656, 105.1975, 27.10711, 0.5355767, 0.001215189, 
    0, 1.318926, 43.09715, 129.1528, 72.18356, 0.6946584, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2322872, 1.578719, 3.188058, 0.5964511, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.6444468, 0.001260127, 0.004589351, 
    0.0003895785, 1.380291, 12.01374, 1.98469, 0.5416846, 0.03535328, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009007449, 0.01690677, 0.01244818, 
    0.02287822, 0.009786648, 0, 0.003852606, 0.001659558, 0.0028247, 
    0.0008283978, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 16.65062, 819.3293, 3142.764, 4069.355, 4310.026, 4138.791, 
    3028.498, 1302.141, 243.1281, 152.0525, 161.9577, 197.8529, 241.7904, 
    305.0269, 491.4062, 495.6271, 352.8353, 417.0757, 533.1383, 443.0636, 
    304.9228, 305.4563, 502.5239, 701.9562, 745.4413, 762.6639, 609.6328, 
    610.1339, 720.3016, 583.702, 244.3076, 0.001969652, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 60.44611, 569.196, 1242.847, 1595.085, 1550.8, 
    1457.302, 1367.953, 1243.161, 1115.287, 1091.343, 1146.535, 1205.741, 
    1217.304, 1218.542, 1265.714, 1041.938, 821.9119, 1037.91, 793.716, 
    825.8652, 670.2501, 512.3199, 349.7946, 92.08901, 0.02760974, 0, 
    0.02102749, 0.1391274, 0.02398786, 156.1709, 405.765, 55.77312, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0001584216, 1.112368, 22.48359, 0.6684555, 
    6.000947, 61.34658, 131.1282, 247.6988, 168.4841, 52.69407, 1.405685, 
    0.001375962, 0, 1.062894, 43.22084, 142.5586, 23.63516, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05182566, 1.023114, 0.6405272, 0, 0, 0, 
    0, 0, 0.0003461041, 0.01172155, 0, 0, 0, 0, 0.07398921, 0.1301732, 0, 
    8.790442, 36.68662, 1.236627, 0.6211582, 0.04952403, 0, 0, 9.038179e-05, 
    0.000422647, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.97051e-05, 
    5.762122e-05, 0, 0.0001804551, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.09430607, 256.0096, 2240.09, 
    3589.398, 3518.739, 3371.597, 2457.386, 1204.915, 389.7961, 164.63, 
    147.0752, 147.3907, 164.4407, 203.5153, 324.1829, 483.8195, 493, 
    398.0503, 423.4395, 433.023, 383.5118, 306.0105, 254.2152, 369.3506, 
    563.5505, 665.8275, 753.7077, 621.5485, 607.6984, 766.229, 574.882, 
    251.6911, 2.80182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 2.631258, 184.7836, 1037.382, 1613.968, 
    1587.197, 1421.362, 1371.082, 1224.363, 1107.84, 1187.991, 1260.877, 
    1291.597, 1298.282, 1241.88, 1231.665, 1257.576, 887.7167, 1026.194, 
    769.0425, 815.6431, 568.5188, 400.7073, 322.7233, 78.84225, 0.0007804855, 
    0.2038229, 0.3951181, 0.1204067, 0.0004067368, 4.699538, 53.47083, 
    12.35164, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009154984, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003377812, 0, 0, 0, 0, 
    0.2611172, 18.30615, 32.94106, 121.8148, 99.45173, 49.98167, 11.19526, 
    0.003446214, 0, 0.2526211, 26.70875, 37.50763, 1.382225, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.08200728, 0.1866251, 0, 0, 0, 0.06016999, 0.1461664, 
    0.04239536, 0.001928552, 8.152956e-05, 0, 0, 0, 0.0007845775, 0.02830604, 
    0, 0, 0, 0, 0, 0.0008604063, 0, 2.057355, 10.74469, 0, 0, 0, 0, 
    0.000197937, 3.257612e-05, 4.104956e-05, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0009298478, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11.73289, 1080.56, 3511.118, 
    2951.567, 1949.043, 1632.744, 695.0728, 272.4091, 194.3447, 167.1012, 
    151.8194, 159.9302, 182.3958, 243.8948, 354.8651, 407.0592, 348.9862, 
    341.921, 378.308, 354.5844, 330.6007, 306.325, 231.2864, 275.1855, 
    361.7611, 543.5178, 725.8599, 629.7708, 601.614, 849.6011, 568.0197, 
    257.2422, 64.72485, 1.231367, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20.85937, 782.5779, 1498.876, 1451.47, 
    1321.201, 1330.172, 1197.824, 1099.718, 1165.045, 1321.316, 1403.87, 
    1320.554, 1190.967, 1185.801, 1237.166, 1128.338, 1019.333, 795.7546, 
    746.1132, 565.8998, 362.0942, 312.638, 72.44051, 0.004879808, 0.2674159, 
    0.20156, 0.006711525, 0.001859001, 0.03593374, 0.280799, 0.05919315, 0, 
    0, 0, 0.0004575096, 0.0005675748, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003035371, 0, 0, 
    0, 0, 0, 0, 0.1131979, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001520942, 
    0.001476608, 0, 0.1377717, 3.665503e-05, 0, 0, 0, 0.1806471, 13.08924, 
    6.431772, 19.68396, 11.99404, 2.622614, 0.2812903, 0.000233318, 0, 
    0.05158404, 21.95412, 21.74654, 0.01552816, 0, 0, 0, 0.006042699, 
    0.01501778, 0.02881803, 0.4153237, 0.3736666, 0, 0, 0, 0.3674484, 
    0.764245, 0.06223431, 0.01477209, 0.02172371, 0.3360474, 0.4728598, 
    0.07631892, 0.003380621, 0.0001421189, 0, 0, 0, 0, 0, 0, 5.137702e-05, 
    2.271225e-05, 0, 0, 0, 0, 0, 0.0007775159, 0.001250692, 0, 0, 
    0.0006139073, 0.001183125, 0.0001388024, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002403033, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 188.6543, 2135.244, 3513.08, 
    1800.895, 772.4872, 565.9453, 367.2146, 278.4082, 220.9072, 174.0726, 
    156.9657, 197.383, 242.1336, 252.5421, 302.4565, 351.8124, 304.3204, 
    330.0841, 353.2343, 338.0011, 318.5869, 279.1342, 202.8548, 238.3413, 
    334.9028, 549.219, 691.8004, 521.5296, 559.9948, 758.9493, 588.9148, 
    313.9533, 173.4209, 37.48432, 0.2012519, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01666973, 26.16632, 593.6545, 1254.888, 
    1187.172, 1152.983, 1243.4, 1156.376, 1078.201, 1084.911, 1146.937, 
    1275.083, 1219.27, 1168.484, 1235.814, 1298.01, 1281.905, 1135.987, 
    1059.275, 882.8276, 688.4268, 454.46, 305.9841, 37.85909, 0.006671593, 
    0.0321888, 0.009452602, 0.001791614, 0.001540999, 0.004539344, 0, 
    0.0007131108, 0.00452225, 0, 0, 0.001518113, 0.001693755, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0002039297, 0, 0, 0, 0, 0, 0, 0.446679, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.003794376, 0.1531117, 0.2974987, 0.2212669, 34.4014, 48.09744, 0, 0, 
    0, 0.001116863, 0.05740427, 0.1271315, 0.1287978, 0.003256722, 0, 
    0.02469566, 0.0001917199, 0, 0.001534145, 0.8834689, 0.5840206, 
    0.006881718, 0, 3.780504, 198.7262, 312.874, 9.970533, 0.637512, 
    0.4400855, 0.02683332, 0, 0, 0.001624759, 0.03438782, 0.296788, 
    0.4003879, 0.05607034, 0.04936704, 0.6750979, 0.7274987, 0.01126266, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0004224136, 0.0001978505, 0, 0, 0, 0, 0, 
    0.0002318844, 0.0004446706, 0, 0, 0.0009304152, 0.000896834, 0, 0, 0, 
    0.009191659, 0, 0, 0, 0, 0, 0, 0, 0.001371316, 0.0003560028, 0, 0, 0, 0, 
    0, 0, 0, 3.842387, 1.503404, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 565.4529, 3203.447, 2551.167, 937.3546, 375.4412, 
    359.7348, 318.6917, 263.4679, 211.9243, 168.8679, 155.905, 203.9936, 
    230.7551, 203.5252, 214.9235, 268.8992, 300.3767, 311.264, 317.7905, 
    349.8843, 321.2719, 279.9691, 212.0554, 241.2103, 343.1111, 488.3593, 
    612.6195, 500.2083, 504.221, 588.9614, 617.0619, 435.5623, 302.8723, 
    102.7165, 9.055063, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1420867, 45.12899, 409.3235, 997.4451, 
    1001.589, 967.4796, 1109.542, 1063.807, 1036.905, 1027, 1018.944, 
    969.9167, 1134.365, 1203.458, 1226.709, 1380.683, 1391.921, 1374.297, 
    1557.639, 956.9144, 559.1038, 417.6834, 183.3681, 1.125171, 0, 0, 0, 
    0.01918598, 0.01514417, 0.002904604, 0, 0.002400817, 8.188255e-06, 0, 0, 
    0.0009390252, 0.0009730477, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1365849, 0.3070608, 1.240934, 18.78064, 3.259233, 
    0.9229355, 1.260465, 0.5219114, 17.75053, 195.1978, 187.4934, 5.189983, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6576656, 3.770286, 2.580236, 0.09102324, 
    2.409301, 279.3913, 602.9868, 185.6282, 4.259978, 0.4710427, 0.5097216, 
    0.002233235, 0.003105277, 0.04912517, 0.1078833, 0.3050857, 1.062314, 
    0.7734881, 0.04263875, 3.594548e-05, 0.01002609, 0.05076782, 0.024118, 0, 
    0, 0, 0, 0, 0, 0, 0.0002378482, 0.001180097, 0.0004484665, 0, 0, 0, 0, 
    0.000327047, 0.00369656, 0.00174795, 0, 0, 0, 0, 0, 0, 0, 0.0007904948, 
    0, 0.007785264, 0, 0, 0, 0, 0, 0.001523588, 0.0005352268, 0, 0, 0, 0, 0, 
    0, 2.399226, 8.868602, 0.7920406, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8727367, 1527.919, 3210.651, 1479.458, 
    447.3285, 289.2018, 309.1454, 263.265, 221.1709, 187.4926, 157.7339, 
    143.3953, 135.0224, 141.3967, 153.2697, 160.61, 183.1641, 242.4199, 
    272.6623, 340.5567, 387.2139, 324.7878, 329.6567, 249.6499, 238.4274, 
    295.1248, 388.3338, 468.3013, 481.9316, 485.308, 479.7583, 481.3517, 
    432.6334, 373.1745, 308.9651, 109.7373, 0.3743297, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2731493, 81.4484, 468.8848, 991.5443, 
    834.1259, 887.2373, 1063.804, 944.6383, 938.6408, 988.9345, 1028.416, 
    869.2354, 970.5076, 1165.823, 1177.526, 1196.688, 1371.09, 1319.563, 
    1391.155, 1151, 530.2675, 281.886, 67.55002, 0.001599195, 0, 0, 0, 
    0.01429991, 0.009382211, 0, 0, 1.114319e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.002695026, 0.0008894327, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04255218, 1.955136, 
    3.995822, 30.26241, 17.03727, 18.01497, 363.2165, 120.1673, 5.426353, 
    145.382, 240.3315, 8.855088, 2.104571, 1.543891, 2.01486, 39.64231, 
    160.2999, 75.84798, 0.2077301, 0.1807699, 0.1412029, 0.05523544, 0, 0, 0, 
    0, 0.3345877, 1.253838, 15.76354, 26.14391, 14.09119, 5.486448, 104.3638, 
    716.6565, 424.1461, 10.36979, 0.276234, 0.1290997, 0.04641811, 
    0.0001044085, 0.09608363, 0.6743831, 0.8213216, 0.7635866, 0.7947268, 
    0.2155333, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.5395e-05, 0.0005254643, 
    0.001709412, 0.002009305, 0, 0, 0, 0, 0, 0.0002994406, 0.002716592, 
    0.0004319724, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002529571, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.044793, 2.26989, -2.459776e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59.72311, 2465.959, 
    2492.194, 757.6249, 233.7132, 243.0279, 261.1306, 230.3328, 201.3103, 
    176.7246, 139.8282, 123.2135, 99.8299, 92.80446, 106.7481, 130.1343, 
    165.9621, 197.5922, 293.9864, 368.5302, 339.7237, 318.7803, 353.7786, 
    285.0697, 229.3984, 257.1193, 365.2487, 431.3322, 449.2942, 423.2672, 
    391.5136, 454.6512, 437.8264, 479.8955, 569.3419, 292.2216, 3.256101, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04947826, 0.2286389, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 1.75305, 137.12, 559.2642, 955.357, 744.716, 
    866.6011, 952.1718, 790.124, 823.2786, 887.2266, 925.4518, 874.6791, 
    734.7263, 896.0626, 1281.138, 1123.317, 1205.685, 1272.165, 1270.966, 
    1132.69, 731.1902, 251.832, 28.88612, 0.01947437, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003082636, 0.0003462703, 0, 0.002280536, 0.002642102, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0005825761, 0.01119671, 0.003326741, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006385451, 
    30.9361, 225.7328, 165.5352, 207.578, 311.6804, 182.19, 220.0666, 
    58.26403, 1.887577, 0.4186608, 1.073593, 0.04459526, 0.7318642, 
    0.4755288, 0.8065952, 0.4155093, 2.478187, 2.066725, 0.6541026, 
    0.4808548, 0.6047196, 0.2915172, 0, 0.05044046, 0, 0, 2.935481, 15.9624, 
    27.24394, 52.94956, 163.0943, 267.2931, 608.1235, 805.6119, 135.2004, 
    0.0002903433, 0.01897152, 0.01114246, 0.0001635766, 0.02778582, 
    0.3318132, 0.9591927, 0.4629342, 0.3071502, 0.007719098, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7.022802e-05, 0.002482594, 0.00338394, 0.004104684, 0, 
    0, 0, 0, 0, 2.6971e-05, 0.0002750601, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1191253, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001174511, 3.124686, 684.8111, 
    2606.018, 1690.914, 453.2092, 216.8986, 229.8212, 217.2619, 201.0126, 
    175.1401, 161.9311, 128.3158, 103.3088, 84.7302, 76.10276, 83.90617, 
    112.3133, 158.662, 173.4812, 274.657, 287.7389, 284.235, 303.9271, 
    333.7502, 316.6927, 219.1855, 239.2968, 320.8535, 369.6996, 347.3692, 
    295.1655, 320.6506, 517.6194, 525.0957, 480.9168, 528.4131, 309.5065, 
    5.411519, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1528082, 0.6848901, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 13.30163, 187.7791, 544.0811, 801.4567, 
    730.2797, 843.6208, 804.3792, 648.2288, 693.4432, 742.1865, 769.3554, 
    801.8218, 668.6127, 798.9274, 985.9318, 1077.402, 1139.354, 1232.697, 
    1255.429, 1004.778, 904.877, 345.6557, 34.84753, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0005141902, 0.003332616, 0.0006415482, 0.001687007, 0.001496426, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003040906, 0.00371619, 0.0003963878, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.606086, 35.19846, 303.0148, 284.0193, 34.01775, 42.77401, 28.20191, 
    6.155642, 0.8346311, 0.05835645, 0.0006624601, 0.01265507, 0.442468, 
    0.5354704, 0.06963733, 0.1052065, 0.02631074, 0, 0.05270771, 0.02592173, 
    0.2459802, 0.04599865, 0.1861853, 0.1325027, 0.0852237, 0.02484975, 0, 
    3.398033, 21.75287, 64.52866, 292.4435, 973.353, 1208.669, 1291.886, 
    1076.844, 162.7944, 0.1484219, 0.1081316, 0.01406904, 0, 0.216453, 
    1.232409, 0.8691837, 0.05235884, 0.0005418619, 0.0002069957, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0006287425, 0.002636893, 0.0002569956, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003835073, 0.0002237879, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3061398, 46.44129, 1161.355, 2248.184, 
    1257.469, 317.4962, 179.8916, 193.8407, 181.5945, 172.1181, 156.7818, 
    139.4105, 117.2525, 95.80608, 74.27556, 68.58242, 66.50262, 78.61134, 
    118.2647, 153.5741, 223.1534, 260.1624, 262.4831, 269.1656, 274.3157, 
    308.8841, 211.9856, 217.8957, 286.7696, 344.6348, 303.933, 232.5552, 
    329.6046, 489.3919, 377.0792, 297.0201, 336.2711, 207.4011, 2.539395, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 30.90609, 238.7426, 473.7993, 660.1224, 
    657.2318, 670.7422, 638.9839, 555.5311, 569.1903, 612.0215, 643.3967, 
    654.0831, 644.0405, 843.1142, 1067.394, 1143.835, 1126.159, 1198.126, 
    1290.289, 1223.169, 1160.878, 567.2612, 76.55764, 0.01523804, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.004061643, 0.006893082, 0.03300945, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7.744831e-05, 0.006418847, 0.001986018, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2069234, 10.13997, 
    150.8278, 58.55067, 8.022274, 4.573344, 0.1354259, 0.03486525, 
    0.0005235374, 0.06353292, 0.01169681, 0.01822534, 0.002955696, 
    0.01728253, 102.7345, 32.73269, 1.311184, 1.125546, 0.09783464, 0, 
    0.000187077, 0.0009269184, 0.005631806, 0.01757337, 0.3199503, 0.8257626, 
    0.5131206, 3.850443, 25.61097, 80.84402, 245.2973, 550.8616, 874.5777, 
    1486.351, 1235.58, 673.1469, 344.4223, 48.70829, 0.8781251, 1.419754, 
    0.6598847, 0.06283266, 0.3307174, 0.4124692, 4.337736e-05, 0.0004525667, 
    0.004570665, 0.001366328, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002444419, 
    0.0004240095, 0.001356724, 0, 0, 0, 0, 0, 4.371697e-07, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.005757192, 0.00808523, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 5.197316, 217.4259, 1388.577, 1405.166, 683.001, 187.7769, 127.2043, 
    150.5833, 149.509, 144.9751, 148.6489, 131.3339, 107.076, 93.30508, 
    70.20202, 59.02925, 58.33901, 53.72469, 77.98226, 128.6013, 152.542, 
    215.8673, 240.3334, 230.7882, 240.4893, 248.0928, 170.4243, 192.7941, 
    247.5671, 234.574, 178.5971, 161.9675, 274.353, 437.9448, 302.0298, 
    161.3467, 146.6843, 64.82175, 0.2946063, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.5898916, 111.9517, 305.1574, 435.4559, 561.3026, 
    530.6106, 465.0716, 480.7618, 485.0654, 505.3505, 545.4196, 565.3085, 
    560.6644, 616.3363, 920.3812, 1318.535, 1195.16, 1139.82, 1174.354, 
    1282.379, 1434.859, 1179.219, 700.5102, 174.3544, 0.01241766, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0009923651, 0.03986278, 0.2278189, 0.01772633, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.002353815, 71.1639, 407.267, 268.619, 43.60738, 
    0.0007397631, 0.0001781541, 2.783722e-05, 0, 0.003673667, 0.0005656133, 
    0.06202865, 1.346996, 0.03449136, 0.2518563, 157.1279, 56.19671, 
    47.49209, 9.25582, 0.01375156, 0.001978266, 0.2363144, 6.947223e-05, 
    0.05050875, 0.1620802, 0.3321952, 2.479105, 90.26145, 308.0739, 735.6808, 
    1047.08, 1075.36, 877.1577, 648.2787, 593.2044, 316.1261, 76.42161, 
    3.107916, 0.3842088, 0.2479623, 0.381507, 1.917333, 1.248883, 0.1718794, 
    0.004355286, 0.0007304089, 0.0004277528, 0.002812181, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002734331, 0.000784012, 
    0.003332643, 0.001278591, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002749223, 
    0.0004297326, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73.03286, 502.4315, 1591.494, 
    858.8749, 260.321, 138.7338, 123.6117, 131.0815, 126.3469, 115.1181, 
    124.3315, 115.7275, 93.57825, 86.22854, 70.48559, 53.11283, 45.30869, 
    41.7937, 47.76453, 75.49673, 112.3317, 164.0374, 218.3762, 202.8534, 
    195.9872, 170.658, 133.9172, 193.5645, 225.0441, 150.9866, 84.64154, 
    102.412, 221.9939, 347.7148, 240.7158, 74.99409, 26.37796, 4.622642, 0, 
    0.02341218, 0.006792379, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.1089746, 114.2516, 228.0603, 397.3794, 519.8107, 
    538.6803, 420.0827, 359.9961, 389.8728, 433.6115, 477.0428, 517.2871, 
    525.0765, 529.0318, 653.3698, 1213.313, 1796.626, 1394.303, 1198.659, 
    1195.198, 1334.629, 1511.156, 1256.08, 835.1061, 260.3607, 8.089208, 
    0.008692329, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01253636, 0.06614882, 
    0.004457357, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02011364, 0.06364921, 96.26062, 
    331.9776, 105.8796, 11.78483, 0.190508, 0.1254462, 0.05413755, 0.6445878, 
    5.973927, 5.755947, 8.192096, 56.36252, 1.360781, 32.94004, 397.3424, 
    379.235, 404.4186, 29.96267, 0, 0.4564222, 1.037213, 1.696829, 0.6696701, 
    0.2049611, 9.618599, 66.39384, 340.4262, 655.2341, 1221.189, 1303.458, 
    922.1398, 445.5585, 275.2661, 121.2892, 10.47407, 1.289266, 0.01052378, 
    0.001414816, 0.01521934, 0.09898588, 0.8423927, 0.4354649, 0.003644818, 
    0.002919366, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003059794, 
    0.0003337019, 0, 0, 0, 0, 0, 0, 0.0002028311, 5.211068e-05, 0.0007171545, 
    0.0009870795, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005861364, 0.001028904, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5.77535, 234.7662, 1687.067, 1031.744, 
    212.0773, 170.3075, 145.8955, 126.8283, 121.4304, 111.768, 105.4656, 
    95.46949, 79.7555, 74.33288, 62.03932, 50.90968, 42.06267, 39.35836, 
    37.9878, 37.07386, 67.31104, 108.4079, 174.433, 177.452, 133.6716, 
    97.14431, 80.56622, 117.3322, 133.1633, 61.42667, 38.56435, 68.37933, 
    129.7418, 178.2628, 88.03211, 19.35434, 0.1398182, 0, 0, 0.008339822, 
    0.002269029, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 6.316133e-05, 0, 0.001211517, 32.47667, 178.7139, 407.7849, 
    562.4835, 593.824, 515.9315, 359.6717, 325.7104, 345.7159, 404.6574, 
    457.0207, 484.5351, 508.9108, 515.2759, 656.1442, 1183.874, 1789.746, 
    1486.1, 1246.057, 1202.75, 1393.237, 1568.188, 1349.542, 826.2133, 
    228.9758, 35.25034, 1.753862, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.004231e-05, 
    4.949426e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.246728, 26.31503, 466.992, 
    153.4598, 17.12831, 13.00353, 0.4199718, 0.1797053, 3.062753, 28.13944, 
    41.5963, 18.88794, 22.81141, 133.1751, 11.95007, 70.24403, 757.8314, 
    773.8058, 275.1173, 2.699914, 0.162427, 0.2814271, 0.1482745, 0.5079284, 
    0.7801619, 0.531203, 27.59982, 167.2763, 147.9225, 89.21487, 273.7002, 
    325.8502, 225.4896, 92.00645, 74.03867, 27.29289, 0.3883709, 0.05636277, 
    0.3049138, 0.1703929, 0.09322795, 0.3752461, 0.3802719, 0.1178384, 
    2.648361e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001156922, 
    0.004045923, 0.004164221, 0, 0, 0, 0, 0, 0, 5.885246e-07, 8.34694e-05, 
    0.0007280486, 8.583434e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.184395e-05, 0.002480507, 0.001158284, 4.593778e-06, 0, 0, 0, 0, 
    0.2126504, 63.24081, 1396.308, 1475.272, 317.6386, 200.5062, 163.7878, 
    141.4462, 130.2097, 121.3568, 113.694, 96.16393, 70.12643, 63.10063, 
    59.45152, 56.36339, 51.90287, 69.57879, 82.6097, 62.08439, 49.56733, 
    66.17909, 95.61987, 100.4557, 63.5487, 44.90021, 34.90635, 58.42322, 
    82.8493, 42.65065, 21.49964, 23.30479, 25.05639, 29.66952, 5.326797, 
    0.02969019, 0, 0, 0, 0.0004924394, 0.0001289402, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.1178887, 0.02041369, 0.5407167, 36.34067, 228.5949, 499.5704, 
    520.2678, 489.1911, 407.426, 320.2751, 322.0427, 337.5211, 380.7809, 
    416.651, 441.7715, 480.7947, 502.4111, 650.1739, 1091.358, 1755.007, 
    1471.888, 1196.37, 1148.328, 1369.803, 1751.842, 1554.303, 826.7043, 
    243.2057, 61.9791, 8.834237, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001839924, 5.372166e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.236105, 0.4120569, 550.8731, 
    385.8582, 61.23731, 8.090598, 2.326185, 0.0751637, 0.19664, 10.65241, 
    112.6281, 169.1481, 88.56571, 63.88735, 141.7897, 47.92282, 2.334639, 
    396.1944, 651.8465, 483.2636, 161.9579, 0.7453288, 0.4689422, 0.3611927, 
    1.110567, 0.4734879, 3.69716, 135.5391, 555.5262, 168.6813, 3.3654, 
    33.47021, 54.45396, 31.52476, 1.987829, 0.09870031, 0.00811203, 
    0.03148229, 0.02919042, 0.03150873, 0.02558385, 0.2038447, 0.1143135, 
    0.009645865, 0.001527358, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003416854, 
    0.0002372177, 0.0007233825, 0, 0, 0, 0.01609258, 0.01704678, 0.01274895, 
    0, 0, 0, 0, 0, 0, 0, 1.537907e-06, 1.725398e-05, 1.28121e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01534935, 0.07117005, 0.02933446, 
    0.0003689946, 0, 0, 0, 0, 0.9127732, 95.89819, 1221.54, 1813.4, 365.2418, 
    210.3442, 180.887, 163.4755, 145.0576, 124.9977, 119.4905, 101.4201, 
    74.68756, 62.5457, 61.32218, 52.40113, 49.80539, 79.93115, 108.9538, 
    115.115, 85.47103, 110.5713, 182.4664, 108.4687, 33.40051, 21.5051, 
    16.78692, 30.93296, 43.63352, 17.49367, 4.349619, 0.2933085, 0.001500918, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 9.335735e-05, 0.00479588, 0.5197528, 34.59122, 221.2229, 
    424.2921, 426.9743, 446.5049, 364.7774, 316.1198, 324.221, 340.987, 
    365.0652, 401.1288, 436.4665, 457.3676, 493.6926, 653.562, 997.9219, 
    1474.947, 1378.647, 1192.802, 1135.426, 1326.291, 2040.261, 1976.624, 
    891.6703, 277.4091, 106.1988, 26.64102, 0.5096122, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005805817, 
    0.0001638428, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01236409, 0.2743727, 17.52411, 380.459, 143.6283, 20.05356, 1.634894, 
    0.13894, 0.0007495523, 0.01723105, 21.82663, 130.0445, 218.9798, 
    302.4652, 221.0393, 119.5289, 44.28259, 4.371171, 61.51543, 90.55502, 
    150.9951, 77.03284, 0.2165833, 0, 1.703179, 2.842183, 1.017624, 4.810229, 
    42.54254, 143.7156, 39.82099, 1.241978, 0.4909528, 0.3809555, 0.01515961, 
    0, 0.000364433, 0.0007033322, 0.002693928, 0.003673581, 3.57866e-05, 
    0.0003873771, 0.0058369, 0.002246894, 2.535222e-06, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.009074074, 0.006229228, 0.01861874, 0, 0, 0, 0.009641227, 
    0.002136417, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002817247, 0.0009464882, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5514262, 0.8107207, 
    0.1884509, 0.013205, 0, 0, 0, 0, 0.07393015, 91.3456, 952.8455, 2343.415, 
    600.5396, 208.8347, 195.3803, 194.6314, 180.151, 155.8788, 136.3115, 
    106.7206, 84.38576, 77.97706, 52.48299, 45.35494, 47.48174, 86.74055, 
    147.7259, 177.4688, 160.5796, 279.6231, 331.3211, 195.2143, 69.41557, 
    16.32039, 9.593863, 5.895026, 6.228228, 1.298795, 0.04732686, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.6144081, 0.1201005, 68.11377, 354.8523, 479.4304, 
    513.9052, 499.9954, 401.3651, 332.1432, 326.9913, 347.9315, 376.2162, 
    417.6304, 461.9634, 450.7137, 489.9835, 621.4665, 800.0215, 1186.147, 
    1275.254, 1189.215, 1136.365, 1434.438, 1822.868, 1602.677, 783.5375, 
    272.0565, 121.5143, 45.10757, 19.01457, 2.194686, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01663288, 0.0004693873, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04156717, 9.526273, 
    274.0584, 294.3758, 31.09721, 11.58998, 1.843844, 0.09464782, 0.0499364, 
    0.1618054, 61.13998, 86.30412, 137.3605, 432.8288, 554.4264, 360.2327, 
    133.7913, 29.33884, 0.7256588, 0.8119102, 0.4245986, 120.2096, 248.3328, 
    0.4880391, 0.3305904, 1.617507, 0.3854961, 0.1228008, 0.01078547, 0, 
    0.001883394, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005414573, 0.03179919, 0.01515976, 0, 0, 0, 
    0, 0, 5.543395e-05, 0.0006995233, 0.0005609203, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.330508e-05, 0.00161523, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.08077211, 0.1219026, 
    0.0121253, 0, 0, 0, 0, 0, 0, 8.772388, 365.1465, 2004.132, 1050.409, 
    294.367, 215.5472, 231.9195, 216.0225, 203.2227, 151.2273, 110.9351, 
    137.5822, 264.0167, 150.0225, 80.09899, 60.13586, 90.18864, 192.0183, 
    259.091, 256.1421, 345.3578, 357.4713, 260.5684, 132.1062, 24.24519, 
    0.5306289, 0.0004064651, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.3822465, 0.07691711, 143.7374, 525.5913, 607.3804, 
    551.1872, 531.7218, 459.0758, 362.167, 335.537, 349.8652, 382.8549, 
    421.6853, 441.6607, 462.9118, 501.9698, 592.3005, 748.838, 1001.76, 
    1213.788, 1063.905, 1077.55, 1394.281, 1326.745, 1068.913, 549.7512, 
    284.5153, 200.979, 123.5475, 96.48351, 39.7753, 15.11369, 0.2131498, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01044296, 
    0.0002949031, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0007954999, 1.670932, 160.7741, 389.6662, 95.69798, 14.89198, 22.86562, 
    13.43475, 0.07823121, 0.1197338, 0.105126, 53.14258, 86.77338, 132.0584, 
    401.2292, 704.707, 768.317, 375.4507, 86.21048, 1.002381, 0.637751, 
    0.8032964, 2.94895, 149.8206, 1.17133, 0.2826535, 1.441549, 0.2252018, 
    0.005584534, 0.001965774, 0, 0.001689953, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0004838968, 0.0007354502, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.01101913, 0.02524117, 0.005818065, 0, 0, 0, 0, 0, 8.067823e-07, 
    7.925751e-06, 4.334839e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002307725, 0.030837, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00821214, 0.02833684, 0.00312682, 
    0.0002740621, 0, 0, 0, 0, 0, 0, 0.028745, 18.45026, 914.7099, 1677.321, 
    914.4962, 310.2044, 251.87, 237.9297, 212.4214, 172.178, 131.0494, 
    147.4902, 343.974, 390.7285, 251.5964, 133.0766, 125.8294, 252.0677, 
    322.9473, 294.009, 361.7983, 332.1922, 261.6464, 150.3966, 33.95244, 
    0.3918128, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.09843657, 91.97388, 453.6148, 638.7762, 619.6926, 
    580.2405, 497.8364, 421.7378, 366.9922, 367.3934, 394.8164, 428.218, 
    454.0583, 485.7609, 560.8041, 655.0854, 788.3849, 980.5639, 1170.239, 
    988.6096, 1076.626, 1198.109, 801.9147, 683.6693, 522.9745, 445.783, 
    381.2975, 296.2165, 247.4656, 168.6503, 85.78122, 17.57448, 0.008626499, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01544856, 
    0.000435621, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003996762, 
    0.4524872, 34.0896, 536.0942, 545.1519, 53.72488, 41.52142, 72.55209, 
    24.63595, 0.1727179, 0.2386063, 0.06103327, 0.482772, 1.329854, 37.25333, 
    207.4293, 567.8538, 829.7704, 344.6922, 23.98134, 0.01000843, 0, 0, 0, 
    0.5020146, 0.6617018, 0.07367955, 0.7041492, 0.1237348, 0.00050432, 
    0.0001705237, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.358736e-06, 7.052271e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003671642, 0.005973968, 0.0003965028, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005954421, 0.05153333, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005108805, 
    0.001554958, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02223296, 247.5312, 1567.859, 
    1643.202, 739.0755, 250.4235, 211.7799, 194.1617, 173.4507, 138.696, 
    110.8374, 235.9538, 563.2759, 439.9135, 201.3896, 120.9113, 207.2445, 
    247.1065, 281.3922, 355.0748, 270.4271, 211.5824, 132.3754, 23.47147, 
    0.1184077, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.004217431, 0.2635228, 7.893483, 59.35656, 377.5584, 646.8165, 
    675.9363, 639.3987, 571.4305, 513.9129, 419.3131, 401.6645, 425.2153, 
    451.0465, 495.2184, 525.1556, 610.6055, 676.3268, 732.7196, 840.8959, 
    992.0549, 834.4886, 1069.691, 1074.612, 588.6633, 590.4393, 827.1808, 
    810.6704, 599.5052, 357.4285, 359.3475, 353.7646, 177.5368, 95.99923, 
    1.708315, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0007933234, 0.006911415, 0.0001889592, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5.48637e-06, 1.572862, 132.3509, 626.3925, 179.5571, 
    20.40353, 236.1403, 82.22805, 1.333986, 0.5002958, 0.5961782, 0.1997266, 
    0.03270302, 0.01405512, 1.421707, 61.59838, 317.1569, 820.7129, 265.0794, 
    12.40273, 0.0001557115, 0.0002069142, 0, 0, 0, 0.3371323, 0.1971543, 
    0.04139023, 0.0191645, 0.0001969625, 7.399264e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007675897, 0.001161112, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.002959132, 0.004310356, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001315948, 0.006940145, 0.001528074, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.831687e-05, 0.0001161013, 0, 
    96.33672, 1073.487, 1597.302, 1339.139, 409.7873, 185.086, 176.6566, 
    153.9536, 119.1987, 154.6582, 429.0158, 770.9375, 541.5338, 275.6819, 
    124.3149, 177.4132, 170.2561, 238.8468, 222.3157, 180.9762, 173.0793, 
    82.7534, 8.063197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.9356636, 11.11353, 98.49442, 306.4701, 510.7628, 652.8757, 
    687.6468, 691.2292, 627.6771, 599.4415, 495.4888, 438.5882, 458.6964, 
    500.5348, 535.2602, 576.1835, 627.6067, 672.3499, 690.8812, 751.8135, 
    757.9091, 665.0533, 809.0765, 712.5627, 568.9345, 801.8674, 1250.082, 
    1156.263, 855.7318, 389.9433, 408.8398, 431.4234, 254.5267, 178.1464, 
    74.96397, 0.06013983, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.810041e-05, 0.00907093, 0.0002546076, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.03228528, 268.1548, 811.538, 282.7054, 0.5783633, 130.3572, 
    417.1314, 158.9361, 1.58552, 0, 0.02557044, 0.1628458, 0.02197797, 0, 
    0.0004203951, 5.260473, 96.06978, 685.5736, 444.6298, 156.5452, 
    0.6586325, 0.06921662, 0, 0, 0, 0.06805296, 0.4576773, 0, 0, 0, 
    0.0008097811, 0.0005997634, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002018141, 4.117844e-05, 1.976423e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.003336009, 0.0008498723, 0, 0.0004391342, 0.0006323908, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009980927, 0.007733, 
    0.001445114, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0008487213, 
    0.001407053, 0, 18.64006, 568.6592, 1542.742, 1748.931, 982.3562, 
    261.7751, 145.1952, 131.0685, 130.1353, 348.3577, 573.196, 768.6476, 
    575.1424, 658.439, 619.8652, 354.6944, 114.9397, 146.0238, 119.4428, 
    125.1135, 117.3902, 27.45313, 0.523582, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.592173, 
    28.81653, 37.75988, 2.365597, 0.1322388, 0.7540843, 1.663811, 0.2238849,
  28.48198, 0.3221889, 0, 0.7876517, 15.59501, 57.29479, 137.7144, 540.459, 
    922.596, 781.4624, 759.4465, 829.9693, 772.8839, 668.2366, 564.2856, 
    487.0963, 506.9308, 564.4177, 589.8097, 609.2275, 638.1862, 651.7763, 
    608.2402, 608.0028, 555.4704, 474.4733, 487.9842, 582.956, 719.3857, 
    1093.142, 1570.934, 1405.136, 974.9818, 554.3302, 459.7365, 396.1888, 
    337.882, 228.3336, 113.2856, 1.834241, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.01985261, 0.0005583716, 0, 0, 0, 0, 5.726098, 
    0.2308279, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.483737, 8.7814, 21.33413, 
    1.912896, 1.018441, 187.1211, 363.3875, 107.3548, 0.3020935, 0, 
    0.001335935, 0.02663925, 0.003909053, 0, 0, 0.07829803, 6.565096, 
    179.8289, 406.9817, 76.20972, 1.033353, 0.3010974, 0.1298247, 0.00195613, 
    23.00312, 28.48724, 0.02563323, 0, 0, 0, 0.002201876, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4.294276e-05, 0.0005016982, 0, 0, 0.0058836, 
    0.004324966, 0, 0.001538357, 0.0002214866, 0, 0, 0, 0.0618443, 
    0.001734049, 0, 0, 0.003026105, 0.007889727, 0.0008332449, 0.004080439, 
    0.001180813, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001018301, 0.001118449, 0.007544341, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01422359, 0.09879134, 0, 0, 0, 0, 0, 0, 24.59497, 504.9599, 1407.995, 
    1517.119, 1747.302, 712.1491, 127.4513, 106.1332, 109.724, 460.315, 
    654.3185, 476.4819, 533.6478, 890.1335, 803.3425, 319.2018, 67.28496, 
    37.45008, 31.44653, 47.56361, 33.41845, 0.9784247, 9.807763e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.385951, 98.3731, 161.0315, 150.272, 106.8229, 65.70918, 
    87.25622, 102.009, 99.4771,
  142.2409, 58.5175, 39.11346, 61.07827, 117.6677, 120.9079, 141.2118, 
    464.5714, 950.2702, 971.881, 933.2386, 993.1581, 888.9403, 626.9457, 
    526.6959, 506.179, 548.0914, 619.2492, 659.0546, 663.9831, 675.3394, 
    615.7237, 531.5067, 485.425, 450.0066, 428.0992, 426.7666, 589.5253, 
    1183.673, 1428.737, 1901.277, 2082.662, 1320.023, 721.663, 564.5012, 
    556.967, 484.8531, 332.1138, 167.2313, 30.73286, 0.02773762, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001738021, 0.0269049, 
    0.0007565845, 0, 0, 0, 2.500434, 294.1236, 97.01492, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.043905, 0.08929022, 0.002691046, 0.0007603669, 0.2270243, 12.67626, 
    107.5273, 113.7621, 1.693966, 0, 0, 0, 0, 0, 0, 0, 6.88282e-06, 
    1.333677e-05, 78.0378, 230.4481, 18.74833, 0.004727178, 0.1272831, 
    0.3513788, 2.367951, 269.7895, 346.9709, 35.66251, 0, 0, 0, 0, 0, 
    0.1150766, 0, 0, 0, 0, 0, 0, 0.0008184621, 0.001400569, 0.0001733794, 
    0.0004490871, 0.0003057205, 0.003002651, 0.005329432, 0.01818698, 
    0.003029905, 1.13548e-06, 0, 0.0001054172, 0.1415813, 0.0005295637, 
    0.002168681, 0.0008962362, 0.01303638, 0.0003813234, 0, 0, 0.0006177669, 
    0.003519957, 0.004156905, 0.01521258, 0.0003090867, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009965184, 0.0009707269, 
    9.238986e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001170971, 0.00676976, 0, 0, 
    0.02225824, 0.5781473, 0.688782, 0.002876182, 35.12899, 545.9062, 
    1202.37, 884.5132, 1741.207, 1096.982, 137.7199, 90.72253, 73.31557, 
    250.2422, 392.959, 300.0186, 421.3236, 461.0554, 362.62, 132.7506, 
    32.3471, 1.977075, 0.1556128, 0.1352257, 0.3216732, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.189352, 80.38451, 216.3247, 261.5845, 233.1123, 189.6998, 140.4133, 
    181.6356, 214.8796, 198.4153,
  252.1725, 171.851, 161.2775, 269.3723, 318.7035, 207.9336, 173.3849, 
    203.2355, 481.1755, 836.9971, 861.7103, 867.8267, 724.3207, 504.5536, 
    443.2747, 452.1268, 541.174, 671.712, 729.8811, 730.2318, 689.915, 
    569.5302, 473.6154, 420.299, 410.6874, 413.4931, 413.1507, 582.8369, 
    1687.1, 1843.39, 1979.237, 2298.16, 1623.208, 956.2333, 873.2465, 
    856.9896, 654.0795, 534.8378, 429.1031, 149.5503, 3.065235, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.851034e-05, 0.005708157, 
    0.0001667178, 0, 0.8102365, 0.5540461, 3.135247, 232.9329, 68.10558, 0, 
    0, 0, 0, 0, 0, 0, 0.005906864, 0.2979069, 0.4578249, 2.618528e-06, 
    0.02129698, 5.316709, 65.49004, 34.45197, 0.6580219, 0, 0.01128094, 
    0.002282921, 0, 0, 0, 0, 5.633888e-06, 6.423807e-05, 8.295042e-05, 
    0.5456263, 2.256658, 0.336203, 1.303343e-05, 0.002366495, 1.661705, 
    113.5126, 429.9062, 457.05, 111.4405, 0, 0, 0, 0, 0, 0.3038842, 0, 
    2.122937e-05, 1.140674e-05, 0, 0, 0, 0.0006652306, 0.001456426, 
    0.0003083536, 0.0009400716, 0.0003889856, 0.003066359, 0.03201295, 
    0.1623753, 0.01771627, 0.001624284, 0.002425614, 0, 0.01565143, 
    8.517144e-05, 0.0003986394, 0.0001845766, 0, 0, 0, 0, 0.00950619, 
    0.003932912, 0.00178012, 0.006202288, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.06594879, 26.86364, 62.05737, 32.63319, 0.9462222, 77.27602, 401.1042, 
    737.3174, 520.0771, 1172.242, 1032.835, 264.6966, 77.33611, 58.71748, 
    69.29409, 116.5409, 156.2841, 236.7241, 242.6088, 144.6283, 53.43567, 
    8.560749, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01609659, 10.2879, 70.72753, 
    238.5741, 402.2285, 425.1013, 331.0837, 256.2188, 207.7381, 244.1325, 
    229.7893, 167.2121,
  271.1909, 280.6147, 305.7315, 332.8787, 252.9022, 205.3805, 271.9508, 
    258.5124, 233.695, 453.5862, 467.2225, 489.5421, 476.4453, 421.786, 
    398.0763, 408.3026, 510.3663, 651.957, 775.6343, 760.5718, 631.5822, 
    502.6142, 427.9246, 397.6864, 400.5818, 405.0021, 411.7556, 798.8644, 
    1678.138, 1875.841, 2127.046, 2029.668, 1525.409, 1300.674, 1240.042, 
    1086.694, 835.6548, 712.444, 631.8665, 440.707, 60.93268, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002498722, 6.972792e-05, 1.529409, 
    90.82018, 64.90834, 2.459643, 93.00716, 14.62878, 0, 0, 0, 0, 0, 0, 0, 
    0.02396147, 0.248873, 0.138524, 0, 0.130176, 35.48887, 106.2803, 
    25.34982, 0.00138829, 0.01617281, 0.04477547, 0.06100203, 0.1747074, 0, 
    0, 0, 4.950247e-05, 0, 0, 0, 0.207136, 0.08613342, 0.003588234, 
    0.0001411147, 1.761624, 102.5032, 348.9734, 340.802, 53.18185, 0, 0, 0, 
    0, 0, 0.02667209, 0, 8.929685e-05, 0.01882303, 2.820102e-06, 
    0.0006965794, 0, 0, 0.000288884, 6.943857e-05, 0.0001046995, 1.60713e-05, 
    0.000683044, 0.001332266, 0.001621558, 0.0002755124, 0.000461814, 
    3.787291e-05, 0, 1.194358e-05, 0, 0, 0, 0, 0.0002516212, 0.001573769, 
    0.00485307, 0.006381406, 0.001770964, 0.004054758, 0.003760318, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.001423343, 26.9012, 412.6746, 413.1584, 139.5305, 
    43.4004, 164.5255, 146.8178, 144.5157, 266.1757, 575.4769, 803.7107, 
    938.4072, 202.8317, 74.48077, 95.55794, 108.1834, 147.2102, 139.5167, 
    121.3799, 31.22051, 3.729389, 0.002843817, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5128328, 28.77927, 185.2033, 410.6761, 582.509, 540.1542, 390.3307, 
    317.1128, 275.0884, 276.0371, 198.5125, 141.3501,
  246.1753, 352.6752, 350.3407, 262.0777, 190.3082, 350.8808, 646.1453, 
    627.691, 344.8603, 342.941, 380.5563, 380.7798, 373.1366, 369.2466, 
    379.5113, 392.1536, 417.7881, 482.3943, 631.5909, 632.6683, 530.5132, 
    445.5339, 410.3927, 401.993, 407.0577, 399.0364, 441.1349, 1022.751, 
    1428.385, 1742.936, 2135.097, 2070.855, 1194.018, 1436.676, 1480.258, 
    1142.292, 931.7062, 853.1913, 854.1656, 669.9532, 295.7026, 0.001168092, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002600568, 0.002716534, 
    7.45994e-05, 29.09718, 265.5758, 218.9747, 19.02556, 18.33483, 0.350748, 
    0, 0, 0, 0, 0, 0, 0, 0.005508803, 0.03894449, 0.004375981, 0, 0.1236557, 
    46.80601, 79.87657, 1.632096, 0.002008923, 0.2392406, 0.7460181, 
    0.6653972, 0.2312042, 0.002383319, 0.005942997, 0, 0, 0, 0, 0, 
    0.02866103, 0.5441989, 0.4410607, 0.00583145, 2.000534, 178.7628, 
    5.172748, 9.298877, 2.336139, 0, 0, 0, 0, 0, 0, 0, 0, 0.05762449, 
    0.0004356665, 0.003173247, 0, 0, 0.0001647425, 2.060104e-05, 0, 0, 
    0.0001603405, 0.0003043673, 0, 0, 0, 0, 0, 0, 0, 0.0009082176, 
    0.0007458362, 0, 9.197873e-05, 0.001946518, 0.005071888, 0.001853016, 
    0.007676827, 0.00722508, 0.00133122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001383478, 
    11.88878, 646.7948, 883.3793, 26.15314, 3.937066, 94.84592, 101.1212, 
    11.97805, 52.49405, 132.369, 372.2394, 520.1495, 859.1444, 538.0435, 
    270.9929, 304.0543, 181.1423, 221.3815, 135.453, 16.63721, 3.064498, 
    6.080413e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06904958, 26.03698, 140.9845, 
    327.9371, 464.5642, 532.6739, 494.3611, 402.8531, 350.8956, 305.3644, 
    296.0944, 217.3465, 161.3094,
  225.7294, 341.2296, 313.972, 262.6939, 302.8044, 499.9109, 708.6488, 
    660.1754, 450.3249, 399.3658, 464.6774, 408.7065, 333.6264, 343.3682, 
    387.6309, 420.563, 426.6206, 456.2177, 535.9461, 524.0982, 464.9332, 
    431.7157, 433.2836, 458.7855, 486.7282, 423.7115, 443.1367, 801.36, 
    1145.982, 1784.052, 2191.227, 2167.639, 888.1638, 717.0386, 666.2883, 
    241.6991, 273.7101, 761.2507, 1007.772, 763.251, 356.4659, 0.7562128, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004910638, 0.007967938, 
    0.043763, 87.9554, 377.9861, 278.619, 45.30785, 0.3442256, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.02145035, 0.1408187, 0, 0, 0.2095862, 43.08374, 70.98579, 
    0.7649364, 0.4206844, 40.92967, 52.13824, 4.659302, 34.06265, 57.93167, 
    7.28483, 0, 0, 0, 0.000343531, 6.250646e-05, 0, 0.3558991, 1.365733, 
    0.2331577, 43.40847, 167.596, 3.089865, 2.148132, 0.07875401, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.001677954, 0.0005306152, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0002353485, 0.0002094212, 0, 0, 0.001254711, 
    0.003052011, 0.0007321349, 0.007233372, 0.002682855, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.0002835374, 0.0002323918, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1.588999, 129.5983, 400.5421, 79.17206, 0, 0, 
    0, 0, 0.0004815274, 22.39184, 336.6852, 894.7394, 278.4767, 393.8267, 
    503.286, 308.6811, 204.6909, 60.25893, 116.4038, 208.232, 9.192997, 
    0.5124927, 1.032356e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002817643, 5.772889, 
    92.11348, 351.7063, 557.7882, 490.7862, 430.6049, 410.9663, 378.1926, 
    375.972, 339.9221, 303.2899, 254.3626, 209.0624,
  244.6317, 259.7936, 242.9138, 248.9483, 371.091, 554.5114, 592.5891, 
    493.2202, 418.8201, 393.7914, 391.6306, 340.0166, 314.1319, 337.1869, 
    418.7542, 458.5742, 462.8698, 517.7924, 626.5951, 624.1047, 507.8369, 
    467.7977, 491.4613, 582.9401, 643.0062, 495.2027, 456.0114, 570.5004, 
    857.7321, 1724.711, 2209.393, 2123.341, 780.9756, 500.6788, 284.5303, 
    5.407286, 5.066408, 181.6497, 409.3565, 484.8989, 356.6444, 1.264237, 
    0.01013122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00221296, 
    0.004024901, 3.93992, 218.506, 596.283, 407.7119, 105.4132, 0.0231447, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.2170925, 1.062111, 2.101756e-05, 0, 0.2954868, 
    47.3016, 119.7318, 26.3369, 30.80848, 233.3162, 144.9064, 27.63708, 
    181.0965, 476.2475, 63.77523, 0, 0, 0, 0.0001767295, 2.565738e-05, 0, 
    0.08221614, 0.9285621, 0.589502, 92.40862, 61.61262, 19.3667, 94.27132, 
    0.005529609, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.001580631, 0.0004886921, 0.0006181647, 
    0.003231038, 0.001967551, 0.0008305749, 0.001923599, 0.0001776486, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.773742e-05, 6.938761e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006362479, 5.45014, 89.04519, 
    140.3022, 14.99106, 0.007751393, 0, 0, 0, 0, 1.975018, 73.17046, 
    131.2607, 45.77481, 49.86932, 148.0228, 25.83098, 3.085815, 0.4943291, 
    0.6179842, 1.371737, 0.822658, 0.5385996, 0.06584774, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1286031, 16.60693, 95.55524, 360.2158, 563.2491, 473.0604, 
    402.618, 377.8559, 354.4522, 359.443, 343.3145, 303.7542, 291.3494, 
    268.0665,
  273.551, 247.4509, 225.945, 245.3163, 320.0762, 453.3221, 486.6381, 
    399.5902, 364.985, 346.8224, 312.672, 294.1594, 295.2102, 306.8427, 
    371.1595, 431.8765, 489.2334, 623.9288, 833.0327, 945.118, 640.8551, 
    532.572, 540.8651, 608.8138, 581.1937, 470.5955, 432.1893, 467.1785, 
    637.0756, 1355.838, 2012.643, 1913.786, 598.4062, 415.1297, 286.339, 
    189.7078, 55.29903, 1.301162, 0, 0, 3.326062, 0.1890756, 0.9552103, 
    0.7668002, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002169714, 
    0.0005184109, 47.47632, 475.759, 784.1389, 610.8682, 209.7725, 1.90487, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.182212, 1.218657, 0.04285526, 0, 0.319639, 
    71.00726, 230.1253, 63.11058, 88.78484, 200.3864, 84.10485, 58.48127, 
    239.2285, 558.2792, 80.89851, 0, 0, 0, 0, 0, 0, 0.00167165, 0.3881946, 
    0.7936602, 2.156414, 11.81752, 63.19553, 52.83117, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.0003998104, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0005424285, 0.0001804351, 0.0002907554, 0.00142767, 0.0006168838, 
    0.0003399592, 0, 0.000101912, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10.65846, 176.2071, 
    321.4464, 135.287, 8.192966, 0.04106788, 0.02578112, 0, 0, 0, 0, 
    0.4189152, 0.6167089, 39.85301, 6.72672, 2.304676, 0.1184766, 
    0.001979818, 6.171127e-05, 0.01694601, 0, 0.2057259, 0.15534, 0.04143865, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6376932, 26.32191, 60.53218, 179.2166, 
    305.0039, 341.3399, 376.6859, 382.518, 337.6631, 324.2889, 322.7919, 
    299.9324, 308.294, 297.9937,
  272.5043, 246.0535, 242.8784, 264.7136, 311.8349, 389.9047, 445.8358, 
    415.0854, 371.5056, 333.6163, 308.8101, 303.4797, 299.2106, 295.8722, 
    323.2004, 384.5279, 515.8166, 763.3062, 933.0347, 1087.135, 793.7239, 
    636.2261, 597.5938, 587.3589, 495.6666, 416.0666, 418.7581, 447.545, 
    575.5629, 957.5547, 1669.331, 1767.901, 437.7619, 233.5887, 304.4022, 
    1028.852, 685.6425, 199.27, 12.50759, 0.9788944, 0, 0, 0, 0.0201377, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 92.43568, 616.1606, 755.6024, 
    635.3912, 258.9823, 3.111485, 0, 0, 0, 0, 0, 0, 0, 0, 0.05177718, 
    0.3728021, 0.07056196, 0, 0.4876086, 117.3619, 259.2785, 44.25626, 
    127.2613, 104.081, 72.21581, 102.2262, 232.2458, 511.0663, 72.79794, 0, 
    0, 0, 0, 0, 0, 0, 0.01618654, 3.927418, 7.774903, 25.26597, 28.21404, 
    0.1011353, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1890707, 
    0.1380272, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0775262, 10.00533, 34.09544, 277.0591, 417.3987, 631.4203, 
    552.2681, 151.3372, 7.581177, 0.0317313, 0.05037785, 0, 0, 0, 0, 0, 0, 0, 
    0.00210742, 0.006124891, 0, 0, 0, 0, 0, 0.1600898, 0.4355638, 0.03862382, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.005684737, 0.008212242, 1.457667e-05, 0, 0, 0, 0, 1.289548, 
    28.62348, 45.58126, 77.36942, 146.2352, 238.0009, 317.8664, 359.4682, 
    322.9961, 295.7401, 304.6233, 302.7278, 314.2467, 301.6702,
  269.4134, 264.0243, 267.0051, 297.0068, 376.5886, 413.2691, 452.8355, 
    460.8797, 413.1158, 356.1818, 329.415, 329.1801, 322.5341, 295.0854, 
    309.4218, 369.8365, 522.3846, 841.9219, 913.445, 998.2731, 919.2898, 
    764.2678, 618.4883, 540.7355, 481.2132, 416.4601, 411.7217, 465.1177, 
    537.5942, 781.7757, 1360.016, 1553.332, 227.1851, 31.32765, 425.9471, 
    1723.69, 1464.588, 1066.761, 805.2874, 318.4906, 14.54321, 1.316028, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 281.1864, 609.5691, 
    585.7905, 442.2675, 212.9697, 2.124233, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.00701096, 0.04654004, 0.01405342, 0.006106328, 6.249868, 191.5606, 
    275.8269, 69.67093, 216.6441, 157.9642, 145.9508, 183.1009, 442.4663, 
    616.7739, 71.27069, 0, 0, 0, 0, 0, 0, 0, 0.3457654, 131.92, 124.4837, 
    1.267306, 0.3921685, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04109782, 0.2183067, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0003228024, 0.001227101, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0577864, 105.1874, 736.0284, 
    1013.626, 904.2305, 943.0919, 899.6609, 534.7457, 157.6137, 10.07536, 
    1.174714e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1291069, 
    0.3769271, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.06047232, 0.2303476, 0.06931562, 0, 0, 0, 0.04560825, 
    15.91871, 37.80263, 47.21033, 60.89336, 103.556, 198.5162, 277.6467, 
    309.5074, 300.5234, 283.0021, 291.8886, 335.5964, 306.7596, 291.1651,
  286.0087, 297.9822, 293.3438, 337.2775, 432.5783, 468.2872, 485.4957, 
    482.743, 431.2424, 387.9859, 356.8474, 343.9968, 316.3823, 281.0254, 
    286.9683, 359.8213, 469.9019, 739.0521, 867.1476, 863.3544, 923.9834, 
    823.1363, 587.2379, 498.8038, 520.5927, 438.3772, 429.3544, 463.2368, 
    465.3976, 647.3158, 1112.234, 756.5065, 26.56112, 6.327219, 592.6151, 
    1801.058, 1218.418, 1016.118, 1097.353, 922.6254, 554.9397, 172.7158, 
    3.420658, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.641541, 
    471.6668, 583.4884, 476.6479, 366.4258, 202.9763, 12.70359, 0.382387, 0, 
    0, 0, 0, 0, 0, 0, 0.0002396297, 0.005740316, 0.8337327, 1.235669, 
    16.7155, 305.6983, 343.1118, 110.8247, 266.2481, 176.0089, 150.9703, 
    258.4717, 635.3505, 444.1225, 26.29065, 2.257066e-05, 0.0004921884, 
    0.0004309834, 0, 0, 0, 0, 1.961774, 242.1081, 215.4397, 0.3758883, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02175775, 0.124502, 
    0.01398297, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000206616, 
    0.0008030056, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.077333, 22.11679, 366.2747, 235.5744, 24.29204, 582.5753, 
    1215.269, 1053.085, 545.3748, 447.7611, 665.1036, 437.8134, 118.7977, 
    4.763635, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2207959, 
    0.2595457, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0431494, 0.6089277, 0.3538128, 0.005043821, 0, 0, 
    0.01602322, 7.562269, 36.78865, 47.1722, 58.38185, 110.9552, 193.3285, 
    231.3686, 259.443, 284.4503, 284.5642, 278.3307, 304.9255, 297.4643, 
    292.0335,
  302.6207, 339.3106, 339.2228, 347.3996, 406.412, 464.0841, 521.7245, 
    532.5322, 445.3678, 414.6734, 400.7646, 363.7216, 291.3575, 241.1544, 
    235.2483, 329.4935, 449.7739, 693.416, 904.8916, 734.8011, 711.8109, 
    674.0491, 504.289, 429.5331, 470.8, 424.4445, 434.5703, 404.9462, 
    411.7881, 514.295, 888.8229, 217.6543, 0.0496018, 19.51473, 712.4717, 
    1524.78, 1094.935, 911.7666, 926.4045, 875.9518, 783.0676, 560.0543, 
    364.6401, 177.8449, 2.722338, 0.006191599, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 17.8776, 562.6617, 561.9768, 469.015, 438.5215, 240.1023, 58.02099, 
    26.80125, 4.020744, 0, 0, 0, 0, 0, 0, 0, 0.1227398, 10.55638, 12.59825, 
    28.60055, 264.416, 317.7123, 246.1967, 376.9386, 188.8591, 177.5715, 
    268.2654, 390.2843, 102.2048, 0.9617385, 0.0001816397, 0.002689644, 
    0.001550132, 0, 0, 0, 0, 3.112105, 543.4355, 463.5655, 43.52797, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02281672, 0.1436173, 
    0.008473383, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1872346, 
    22.35824, 382.712, 737.0875, 1230.265, 692.6126, 358.5822, 899.4208, 
    1074.586, 526.9075, 305.9666, 59.5534, 4.745547, 1.596353, 0.3754177, 
    0.0004647044, 0, 0, 0, 0, 0.0001097662, 4.525879e-06, 0, 0, 0, 0, 0, 0, 
    0, 4.288131e-06, 2.984277e-06, 0.003444677, 0.2710683, 0.08078705, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.09098491, 0.2416508, 0.2446091, 0.0258337, 0, 0, 0, 0.614411, 
    26.6793, 44.56842, 70.33549, 157.2269, 218.1267, 209.0873, 233.3854, 
    280.9228, 286.8992, 275.8937, 276.5295, 285.7892, 292.773,
  336.5605, 388.4893, 371.7686, 349.2026, 366.9693, 417.8056, 607.3262, 
    671.5993, 468.1905, 421.5582, 446.4085, 428.6386, 335.3652, 281.8749, 
    258.8414, 309.0987, 440.8155, 649.1459, 863.405, 707.3972, 594.5748, 
    563.7395, 456.5911, 386.5415, 364.001, 379.5974, 432.2464, 381.2984, 
    472.6903, 529.6396, 524.6491, 110.0916, 0.07860577, 175.8245, 1196.177, 
    1471.891, 944.1703, 792.47, 708.6677, 650.6479, 678.2939, 656.6821, 
    596.7901, 457.6963, 67.61382, 8.986737, 0.0001029148, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 179.6408, 628.394, 556.7366, 522.1905, 504.994, 294.1256, 
    160.7078, 239.0964, 156.294, 4.691788, 0, 0, 0, 0, 0, 0, 0.1278733, 
    45.09846, 73.84791, 163.7064, 410.5311, 383.8885, 387.0884, 374.3583, 
    216.1455, 274.0125, 332.5461, 102.272, 2.552336, 17.22299, 0.7804462, 
    0.00171211, 0.0005605019, 0, 0, 0, 0, 0, 501.6506, 338.8492, 23.27959, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01209556, 0.1526054, 
    0.1189834, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.6207879, 14.50541, 
    287.6835, 613.8293, 1068.171, 1441.231, 1470.93, 547.6572, 212.4256, 
    366.9689, 347.8215, 182.1785, 178.7135, 20.04454, 0.000886209, 0, 
    0.0004331574, 7.106494e-05, 0, 0, 0, 0.02318693, 0.08432053, 0.0392032, 
    0.0477153, 0.7327814, 6.548978, 38.41692, 2.65917, 0.2318266, 0.0392304, 
    0.01456798, 0.02600013, 0.05620825, 0.04757133, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2052089, 
    0.3281586, 3.570601e-05, 0.0002343726, 0, 0, 0, 0.07401764, 23.21715, 
    46.79993, 94.43826, 234.8688, 266.0873, 233.1717, 251.4387, 293.1315, 
    297.0283, 288.4081, 276.55, 286.6156, 309.5938,
  392.8387, 488.4619, 451.8623, 387.8266, 370.9583, 414.1181, 685.2869, 
    766.1441, 485.4588, 422.6774, 455.2672, 467.7984, 430.3447, 416.1889, 
    408.9105, 397.4004, 457.034, 579.6365, 743.8334, 684.6434, 567.9512, 
    583.4536, 459.5831, 326.9791, 273.1903, 336.2808, 414.9611, 385.2764, 
    569.3871, 609.2947, 81.50208, 2.31834, 9.107849, 733.1556, 1717.862, 
    1321.356, 856.6255, 681.8816, 520.926, 415.0989, 382.7523, 382.5836, 
    333.1183, 276.241, 209.8208, 75.84883, 1.448402, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 267.8995, 639.0126, 566.5193, 513.6498, 445.1369, 278.2933, 
    264.7586, 481.6906, 394.5965, 72.73242, 1.590796, 0, 0, 0, 0, 
    0.0001962664, 6.500215, 123.3904, 205.7507, 460.6655, 666.9761, 563.4114, 
    513.0554, 458.7825, 492.8423, 544.6861, 271.7018, 4.7952, 1.690305, 
    217.9864, 40.03231, 0.0009057468, 0, 0, 0, 0, 0, 0, 62.97356, 64.35432, 
    0.6435035, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04623526, 
    0.2439728, 0.0118202, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0009476076, 0.001472293, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.247151e-05, 0.008020438, 
    0.001698805, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04228287, 0.3603409, 0, 0, 0, 
    2.168875, 158.9779, 519.3859, 763.6636, 1088.271, 1725.398, 1879.986, 
    1212.513, 193.7943, 23.89315, 39.49089, 41.06394, 90.03802, 150.1664, 
    28.52693, 0.01583713, 0, 0, 0, 0.009915893, 0.01817705, 0, 0.7669531, 
    0.3689948, 0.145493, 1.339995, 147.7285, 527.2662, 509.4995, 61.3713, 
    17.10321, 0.3450269, 0.06363642, 0.03238298, 0.01596504, 0.0002242184, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02224105, 17.85421, 50.62142, 109.2327, 
    273.463, 352.6526, 320.499, 314.5677, 322.3184, 313.0258, 295.2324, 
    278.9248, 303.0909, 354.4732,
  442.1884, 594.8954, 565.0418, 473.9255, 430.8, 453.0199, 678.4496, 
    725.6027, 478.1048, 420.944, 451.6833, 471.7825, 522.8627, 634.4751, 
    830.35, 613.0457, 511.5908, 583.1832, 724.1978, 702.6869, 596.9265, 
    580.4724, 436.6388, 300.9694, 269.1624, 352.4041, 364.6159, 397.8628, 
    607.5164, 524.5532, 2.677896, 8.552654, 173.4247, 1041.965, 1364.173, 
    1057.956, 755.9166, 598.735, 432.5325, 337.5475, 267.133, 219.405, 
    185.0309, 151.62, 156.9159, 128.6733, 19.4975, 0.0003201329, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2788907, 232.2169, 599.0657, 543.3879, 472.7634, 
    373.7747, 249.6898, 348.4809, 536.6453, 481.3254, 248.5191, 32.9144, 
    0.05858242, 0, 0, 0, 0.5034162, 60.42842, 222.9653, 249.5043, 748.5638, 
    825.8325, 702.5027, 669.645, 806.3397, 984.3977, 804.0445, 168.8752, 
    0.2731855, 2.55718, 179.2389, 63.265, 0.2272948, 0, 0, 0, 0, 0, 0, 
    0.1574813, 0.4466992, 0.02788611, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.633844e-05, 4.296753e-05, 0, 0, 0, 0, 0, 0.0414133, 0.2298532, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004690373, 0.0007632322, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.028617e-08, 0.0008502072, 0.02139687, 0.003350336, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0008639033, 0.01942277, 0, 0, 0, 98.26613, 799.9084, 1338.724, 
    1566.699, 1786.769, 2271.628, 2020.339, 867.1221, 42.82516, 0.5412122, 
    0.617964, 2.27297, 47.38787, 98.56119, 27.48889, 0.2292078, 0, 0, 0, 
    0.008091097, 0.03084766, 0.01090882, 3.738859, 48.30343, 108.953, 
    20.27916, 144.7063, 395.8853, 354.0694, 57.11306, 8.065199, 0.005187009, 
    0, 0.003291111, 6.925846e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3200984, 40.53148, 93.36845, 187.2274, 311.3822, 388.1231, 380.9445, 
    357.2439, 334.3976, 312.7577, 292.5607, 282.8434, 307.418, 367.4654,
  433.6788, 584.0782, 632.6719, 582.8133, 534.3633, 524.5817, 642.4552, 
    644.3318, 486.6131, 465.3286, 513.8397, 491.6873, 645.2102, 1165.927, 
    1490.865, 880.6786, 572.1805, 566.6507, 656.6595, 704.7193, 660.4354, 
    559.1111, 430.4431, 333.536, 297.2576, 401.751, 385.7295, 468.3943, 
    570.5828, 461.8753, 6.677346e-05, 92.4138, 779.812, 1268.696, 1040.591, 
    830.1586, 670.9812, 521.1519, 359.7496, 293.7569, 221.2079, 159.9023, 
    130.2733, 101.2735, 108.7102, 117.6302, 37.40805, 3.637927, 0, 0, 0, 0, 
    0, 0, 0.003272676, 0.1988616, 1.901062, 1.564504, 175.4867, 494.2085, 
    413.5671, 408.0959, 359.1264, 271.3205, 354.3282, 404.985, 352.5789, 
    265.249, 107.6353, 7.511302, 0, 0, 0.001996831, 10.16993, 228.5949, 
    395.2381, 271.0521, 935.3456, 950.8614, 837.0136, 803.4595, 837.9974, 
    924.0099, 798.7273, 176.7633, 17.92126, 17.55314, 10.96611, 25.35751, 
    0.2104844, 0.0001917089, 0, 2.373737e-05, 7.919414e-05, 0, 0, 0.01933366, 
    0.3090232, 0.04494533, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.415525e-05, 
    7.552401e-05, 0, 0, 0, 0, 0, 0.01105835, 0.06624987, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00446184, 0.03680261, 
    0.05273988, 0.000618885, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.996364e-07, 0, 0, 
    0, 169.5894, 1188.897, 1678.436, 1932.674, 2075.635, 1893.702, 1131.728, 
    293.5961, 4.660101, 0, 0, 0.02112457, 15.45765, 33.72306, 21.61042, 
    2.09625, 0, 0, 0, 0.0008054632, 0.005477813, 0.1139135, 27.04513, 
    139.0768, 136.8829, 13.60453, 3.55424, 1.563738, 4.366129, 0.1587394, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.280176, 83.67439, 
    146.4108, 271.435, 388.7099, 398.4128, 387.6514, 366.7695, 329.8819, 
    293.9612, 283.0529, 295.4122, 314.1487, 356.7084,
  385.3872, 467.1063, 566.7316, 635.1995, 696.1035, 642.6764, 667.5192, 
    644.1702, 548.7966, 599.477, 638.0853, 544.095, 784.7689, 1236.086, 
    1365.508, 983.0353, 629.7867, 561.2454, 591.3522, 619.5994, 654.6503, 
    517.0252, 361.8463, 312.3237, 306.5308, 386.0362, 398.7388, 497.4073, 
    559.1677, 194.5806, 0.0110149, 235.6834, 1071.164, 1169.659, 965.8761, 
    894.2181, 718.1039, 540.6868, 321.2563, 245.3778, 181.7317, 123.5689, 
    111.2619, 94.61058, 90.59763, 142.0693, 156.6311, 100.8379, 0.002723826, 
    0, 0, 0, 0, 0, 0.08167609, 21.06773, 98.65578, 69.05093, 94.03746, 
    337.3383, 347.865, 396.7599, 468.4401, 422.9413, 412.3752, 328.6121, 
    277.2164, 286.8415, 309.7477, 118.8827, 3.51354, 0.3581138, 0.3971047, 
    53.71002, 537.6266, 570.0897, 249.7113, 862.8484, 1014.729, 1075.184, 
    1050.708, 956.9249, 898.9056, 693.8036, 219.3473, 228.9355, 128.288, 
    40.48083, 40.30056, 45.25633, 2.451566, 0.4187425, 0.07963315, 
    0.0001135752, 0, 0, 0.9117342, 0.06830423, 0.004861436, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007765052, 0.005222111, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007159747, 0.02713225, 
    0.02171584, 0.03361443, 0.0219075, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.004686189, 0.001498268, 0, 0.02123462, 175.3923, 1249.576, 1826.983, 
    2040.793, 1889.158, 1066.356, 266.5604, 25.96716, 0.001682877, 0, 0, 0, 
    0.7125385, 1.146391, 11.38518, 6.322751, 0.001389394, 0.01513089, 
    0.9665338, 0.1141217, 0.8551149, 11.98856, 41.17868, 36.94483, 15.10526, 
    0.3599645, 0.09444457, 0.05254441, 0.008791648, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22.23146, 139.9023, 198.9718, 285.9604, 
    380.5653, 388.1768, 364.6595, 352.3565, 325.2652, 289.1691, 280.3953, 
    299.6466, 323.289, 343.1569,
  369.5396, 426.7726, 535.4895, 727.5086, 1060.43, 949.231, 843.377, 
    728.7923, 699.6417, 782.7468, 742.4287, 652.9568, 805.9807, 782.2319, 
    832.4222, 887.9604, 619.0436, 546.4369, 536.7662, 581.5966, 685.4443, 
    532.7081, 324.4635, 254.6589, 232.1319, 275.3878, 325.0322, 465.5066, 
    347.7954, 56.35401, 1.796414, 357.0097, 1016.861, 986.6382, 963.8297, 
    932.3816, 764.2728, 607.9679, 329.3198, 212.4263, 145.5647, 96.49953, 
    113.3514, 111.7538, 145.127, 366.5991, 401.9952, 189.0011, 1.376681, 0, 
    0, 0, 0, 0, 1.143042, 26.03098, 85.61213, 64.62746, 73.29227, 302.0042, 
    417.8035, 426.0746, 477.8091, 493.5544, 548.0378, 507.4896, 464.5604, 
    454.8298, 379.5999, 131.5459, 13.19003, 4.547818, 4.318508, 122.1453, 
    699.2319, 575.9889, 238.9398, 768.6223, 1021.295, 1245.33, 1266.03, 
    1162.191, 1098.365, 868.7346, 567.8272, 393.3605, 201.9774, 129.8717, 
    215.9289, 178.3175, 37.46669, 45.02709, 60.36355, 2.315857, 0.1704768, 
    0.07761195, 135.5906, 12.82555, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.001651182, 0.002441915, 1.112597e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.04787361, 8.83361, 10.63809, 0, 0.08243045, 435.7784, 1614.9, 
    2058.435, 2109.95, 1731.388, 805.4063, 86.96317, 1.348529, 0, 0, 0, 0, 
    0.0008430668, 0, 0, 0, 0.002104231, 0.5691509, 45.12806, 40.15918, 
    59.46983, 75.78097, 15.58626, 0.2125522, 0.008140751, 0.0306171, 
    0.0240708, 0.0546331, 0.006026743, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6.253698, 175.4863, 259.7228, 299.4385, 317.7915, 
    308.9187, 295.955, 315.1865, 316.5243, 293.2056, 272.7305, 275.879, 
    320.2354, 341.0206,
  347.7965, 418.966, 562.2552, 820.5015, 1296.992, 1267.295, 1064.166, 
    890.6819, 895.5107, 883.4277, 731.1903, 624.9171, 671.4522, 579.5031, 
    566.8748, 680.0339, 554.6023, 506.3958, 476.0154, 514.2544, 758.626, 
    641.5605, 359.8482, 257.0115, 204.9982, 295.3142, 299.809, 429.156, 
    188.9319, 2.458954, 71.56561, 559.0994, 984.5283, 970.0492, 971.8855, 
    930.9053, 773.0588, 635.3317, 384.079, 223.4312, 123.9919, 60.27688, 
    90.43548, 113.4848, 258.6255, 452.4994, 337.419, 12.32377, 0, 0, 0, 0, 0, 
    0.6491734, 5.815516, 50.48944, 38.23403, 55.62584, 166.4128, 308.7408, 
    451.749, 444.122, 458.1162, 445.0182, 485.1528, 512.0165, 529.7402, 
    534.6834, 409.0287, 152.1849, 32.07852, 9.111447, 7.842384, 157.3577, 
    686.8823, 585.9794, 270.8879, 575.1855, 1139.568, 1437.505, 1514.373, 
    1449.192, 1521.215, 1386.076, 985.5462, 559.175, 310.4663, 178.2047, 
    239.9393, 234.778, 149.6889, 199.7453, 221.5135, 120.0964, 22.21674, 
    2.505514, 582.1814, 494.4689, 0.05743101, 0.1109339, 0, 0, 0, 0, 
    5.749473e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.185825e-05, 6.287817e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.396619e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.545735, 113.2851, 198.1115, 
    0.09477463, 44.32423, 1323.019, 2099.929, 2131.979, 2065.898, 1835.858, 
    973.0184, 158.9147, 1.69403, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3942727, 
    18.1228, 7.187973, 0.6999193, 0.1121183, 0.03581052, 0.02583415, 
    0.03022727, 0.009135123, 0.0003793728, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2830645, 138.2685, 267.4936, 298.505, 
    268.9037, 251.0459, 256.5389, 302.3259, 316.7485, 301.4261, 281.5891, 
    279.3524, 285.0648, 314.7705,
  323.2668, 389.2768, 560.0039, 830.4731, 1148.94, 1210.315, 1162.682, 
    1076.238, 945.5571, 849.8019, 678.9407, 570.0232, 563.3746, 501.6432, 
    449.9756, 478.9751, 435.5788, 406.5974, 415.4569, 458.3391, 642.5176, 
    575.6868, 388.3315, 293.3578, 231.1781, 381.2743, 260.8145, 423.3539, 
    82.39389, 41.37816, 405.6402, 770.9765, 941.6445, 936.3031, 940.8395, 
    892.1792, 765.5028, 634.5041, 424.9675, 248.0303, 101.8705, 12.73724, 
    26.73048, 43.31859, 232.4138, 225.3723, 26.30726, 1.461209, 5.5785, 
    2.708922, 0.02225682, 0.2463678, 0.3156092, 40.62003, 25.33394, 25.03576, 
    49.54607, 130.2422, 396.1015, 442.762, 423.5359, 403.6569, 406.033, 
    351.4386, 340.5537, 319.5878, 302.7865, 278.9697, 255.9653, 162.0942, 
    55.60219, 17.67499, 64.36505, 249.0641, 623.581, 724.6849, 375.6157, 
    413.5169, 1302.89, 1715.619, 1792.989, 1746.485, 1823.301, 1517.055, 
    991.2774, 675.8403, 454.7752, 302.1877, 366.0927, 437.0839, 392.9335, 
    356.6635, 348.0479, 401.7336, 215.2848, 30.34251, 355.4783, 498.5672, 
    0.4986214, 0.5007799, 0.1329389, 0, 0, 0, 0.00101586, 0.0003732887, 0, 0, 
    0, 0, 0, 0, 0.009260939, 0.05226945, 0, 0, 0, 0, 0, 0, 0, 0, 
    8.446827e-05, 0.0004581793, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32.32329, 84.06284, 5.961504, 31.71557, 
    549.7613, 2008.809, 2070.353, 1845.099, 1891.462, 1862.213, 746.8804, 
    134.2319, 2.000803, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00217568, 0.0256771, 
    0.05994255, 0.01601593, 0.1703317, 0.04478687, 0.03659392, 0.01946149, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35.46974, 
    199.5, 269.6945, 270.2229, 270.5895, 285.7962, 338.67, 342.202, 300.8127, 
    280.632, 280.3313, 274.273, 291.2681,
  263.2462, 284.5884, 468.1183, 770.9202, 974.9459, 1133.144, 1217.117, 
    998.2538, 773.7898, 777.1089, 620.0529, 514.5913, 522.9897, 489.9959, 
    408.1004, 347.7855, 306.4745, 277.9374, 351.1268, 400.5291, 432.5822, 
    421.2414, 309.0428, 300.5629, 308.1246, 349.6395, 301.6355, 331.7687, 
    1.202404, 129.5541, 615.0019, 928.7737, 1071.859, 900.7906, 818.7495, 
    748.8444, 705.5492, 603.1695, 385.4343, 196.4225, 55.19749, 1.221395, 
    0.0115012, 1.261582, 87.73291, 125.2576, 137.0045, 142.1483, 178.5234, 
    145.3288, 166.8964, 267.4174, 194.4118, 208.5532, 89.00009, 39.60981, 
    111.2856, 160.0921, 294.9518, 440.5912, 347.4731, 324.3401, 295.2901, 
    206.3315, 156.9781, 126.9081, 102.0809, 77.15842, 58.93751, 50.31418, 
    35.45154, 49.30099, 196.6609, 410.6617, 535.1404, 893.442, 646.5032, 
    500.6869, 1418.796, 2123.046, 2099.64, 1939.927, 2094.616, 1820.554, 
    1186.311, 929.059, 762.2305, 512.7437, 529.1393, 490.1915, 473.8611, 
    443.9379, 399.5623, 547.7155, 507.7973, 160.667, 39.65385, 69.58859, 
    0.02925806, 0.03310997, 0.02806808, 0.09657825, 0.01626927, 0, 
    0.01859221, 0.004631748, 0, 0, 0, 0, 0, 0, 0.005736903, 0.04095821, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.877666e-05, 0.0001420318, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001997955, 3.722127e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.835136, 135.7174, 4.789517, 19.04744, 318.4999, 1460.709, 2136.959, 
    1700.521, 1392.469, 1482.793, 1386.474, 335.7827, 66.42863, 3.190663, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002973209, 0.6352931, 2.491891, 0.8138618, 
    0.09514129, 0.02720593, 0.01066479, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16.59806, 135.7921, 243.3941, 344.9666, 
    371.6502, 359.6897, 378.103, 381.3317, 355.234, 325.2544, 296.1037, 
    279.9285, 269.3434,
  236.5887, 253.1677, 358.7563, 571.0236, 731.3325, 722.4735, 743.4526, 
    666.7219, 599.2096, 618.8971, 518.6953, 456.6857, 486.6131, 543.8828, 
    439.4839, 280.6839, 229.2171, 192.6122, 255.1076, 271.4104, 281.6126, 
    275.7565, 229.7789, 278.2134, 275.7716, 304.1842, 392.3536, 139.4066, 
    33.0128, 458.8552, 920.1097, 1038.114, 1118.127, 960.3683, 776.2888, 
    635.3617, 591.0509, 477.8755, 253.2336, 97.80558, 9.85123, 1.627402, 
    12.09361, 198.4388, 113.6606, 238.1357, 561.9626, 556.5967, 715.9232, 
    785.4809, 757.7484, 819.5304, 745.1021, 536.9188, 124.041, 57.69806, 
    153.2543, 213.1749, 262.9545, 374.214, 340.574, 269.8781, 201.2071, 
    147.1432, 116.1977, 91.175, 73.2971, 76.68616, 149.6286, 400.8653, 
    555.6998, 654.2615, 733.0278, 800.9901, 494.8335, 606.881, 707.8926, 
    810.878, 1538.385, 2588.938, 2419.166, 1956.064, 2172.053, 1974.549, 
    1446.878, 1130.417, 891.0532, 625.531, 543.0157, 328.1959, 328.7752, 
    363.0545, 317.9218, 486.5319, 505.6643, 321.8582, 29.09856, 0.005329356, 
    0.004316996, 0.002581715, 0, 0.2576422, 0.8647975, 0.05479293, 
    0.01254045, 0.006202601, 0, 0, 0, 0, 0, 0, 6.259618e-05, 0.1009142, 
    0.09139892, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.698674e-05, 3.883299e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.007198914, 
    3.749324, 120.5373, 151.8816, 7.438391, 142.0757, 896.3428, 2011.567, 
    1952.657, 1446.296, 1233.643, 1159.563, 777.6533, 169.2422, 50.12192, 
    2.106122, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2809023, 6.430042, 10.00201, 
    2.291929, 0.0206799, 0.0321942, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.002652701, 0.0007121718, 0.376531, 35.60808, 
    157.8771, 269.2775, 378.3774, 445.4393, 410.4814, 386.3655, 401.5077, 
    428.1593, 378.8305, 305.6711, 254.8196,
  311.7992, 395.5877, 432.8708, 488.1894, 491.9596, 455.8698, 498.9413, 
    533.1855, 540.7218, 513.9946, 471.9363, 465.892, 505.0617, 617.8649, 
    434.1176, 244.8432, 187.6783, 138.5197, 168.3429, 175.1707, 185.2439, 
    171.4601, 184.4823, 212.1878, 178.8987, 424.5008, 399.632, 79.02595, 
    258.169, 930.0715, 1029.974, 1008.649, 986.2982, 932.3816, 734.9354, 
    569.3074, 450.8971, 349.6758, 146.0535, 18.6776, 12.29715, 133.0716, 
    429.519, 747.2996, 631.5124, 552.8401, 651.7254, 752.6821, 1130.893, 
    1229.507, 880.8947, 959.7202, 1213.855, 934.8705, 142.4921, 70.70444, 
    125.7273, 185.8272, 252.5484, 341.6752, 388.0057, 279.1929, 180.2787, 
    146.0737, 121.422, 199.4011, 442.9223, 723.985, 1486.055, 2640.339, 
    2907.246, 2975.658, 2887.232, 2814.498, 1827.834, 752.6064, 552.7391, 
    1709.945, 2333.681, 3089.403, 2958.684, 2422.924, 2234.675, 1704.245, 
    1291.295, 1053.173, 876.6812, 560.3719, 461.3859, 291.2385, 192.4786, 
    214.8734, 200.1322, 318.3211, 508.591, 622.4544, 184.5554, 2.089956, 0, 
    0, 0, 0.01264686, 0.327778, 0.2354753, 4.464748e-05, 0, 0, 0, 0, 0, 0, 0, 
    4.832438e-05, 0.09589284, 0.1123158, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001072123, 
    0.0007945669, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0001484985, 0.6429842, 50.72206, 261.5746, 49.39819, 93.00819, 
    483.3765, 1486.976, 2011.244, 1570.817, 1394.617, 1305.851, 961.0363, 
    405.7976, 151.1119, 81.06501, 8.738538, 0.08169014, 0.0008955649, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.953568, 21.78077, 12.24485, 1.07415, 0.001584131, 
    6.819148e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.4064472, 1.186353, 0.4749914, 1.063456, 59.91799, 195.2914, 
    379.2884, 478.5082, 433.806, 398.6985, 404.2307, 419.3512, 389.7552, 
    317.8314, 266.4668,
  356.137, 488.0196, 525.0481, 462.7664, 380.1859, 385.0742, 458.4339, 
    558.608, 610.413, 571.0131, 562.7314, 531.9318, 505.2505, 413.2031, 
    281.4167, 186.6899, 138.8866, 93.84417, 122.1802, 118.3982, 114.7902, 
    90.79964, 151.9827, 175.2933, 149.4086, 412.1827, 473.1306, 653.015, 
    827.5731, 978.5537, 909.1771, 885.0692, 863.3699, 767.186, 642.1213, 
    500.9229, 373.5085, 294.3045, 101.8269, 1.344416, 53.2753, 651.5987, 
    1130.408, 1340.512, 1481.681, 1559.811, 1164.816, 848.5647, 1316.412, 
    1165.666, 840.2272, 898.7839, 1274.809, 1223.543, 277.6357, 207.368, 
    122.2911, 125.0566, 184.17, 247.2821, 273.3881, 231.3729, 193.7136, 
    248.106, 443.2143, 1301.328, 2565.46, 3295.099, 4205.998, 4937.032, 
    4773.964, 4663.778, 4548.939, 4451.055, 3627.58, 2251.264, 2021.805, 
    3307.607, 3677.913, 3751.295, 3659.55, 3060.447, 2020.194, 956.3508, 
    714.6304, 900.0114, 881.4429, 565.386, 406.1902, 192.5201, 132.7902, 
    274.0363, 131.1107, 146.5069, 377.0321, 492.1361, 324.5735, 49.08009, 
    0.09172285, 0, 0, 0, 0.01012682, 2.276415, 0.04390513, 0, 0, 0, 0, 0, 0, 
    0, 7.504402e-07, 5.558774e-05, 6.749376e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.481087e-05, 0.0003173137, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3.536257, 0.4066131, 12.77594, 190.7889, 177.2399, 
    77.3595, 297.2285, 849.544, 1832.184, 2035.107, 1417.24, 1315.898, 
    1276.046, 898.1604, 382.3683, 183.029, 99.14983, 29.08071, 4.887974, 
    0.5308673, 0.001209072, 0.02379014, 0.04125052, 0.01250304, 0.0005235381, 
    0, 0.004013969, 0.008801949, 3.331747, 27.98007, 9.583447, 0.0455796, 
    4.645122e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1.591726, 4.157285, 2.159603, 0.8029898, 0.8287141, 10.66547, 
    223.1661, 491.9315, 493.4645, 483.2839, 479.5422, 454.4722, 418.1563, 
    363.4709, 303.4126,
  389.5554, 450.7025, 444.3544, 342.9534, 291.2544, 292.5314, 359.7049, 
    466.8882, 578.2619, 633.2922, 594.0996, 474.4345, 343.1389, 285.8849, 
    226.5928, 103.2897, 50.01753, 51.91085, 81.64977, 76.43392, 94.65741, 
    31.67269, 68.29819, 146.7406, 148.9659, 328.6473, 498.6185, 702.2924, 
    918.2619, 942.1927, 766.6232, 758.2426, 720.8044, 605.1721, 509.771, 
    395.8156, 280.1597, 200.4158, 49.00248, 6.755203, 270.7791, 1279.518, 
    1807.523, 1838.696, 1993.026, 2182.023, 1265.656, 870.415, 1151.028, 
    867.8135, 849.8157, 997.5562, 1204.195, 1417.743, 764.2448, 645.3609, 
    294.3994, 122.3237, 154.7317, 193.7708, 214.4495, 242.906, 451.1191, 
    1113.341, 2119.173, 3344.29, 4568.095, 5045.683, 5142.618, 5122.815, 
    4951.682, 4914.965, 4824.239, 4790.269, 4620.173, 3893.588, 3743.627, 
    4400.479, 4285.227, 4192.585, 4154.279, 3466.801, 1550.915, 499.6396, 
    378.9887, 591.3363, 843.33, 818.22, 599.7932, 154.1871, 88.30436, 
    223.5071, 136.845, 128.7726, 322.8817, 338.9769, 235.237, 74.55579, 
    0.3836409, 0, 0, 0, 0.001294891, 0.4691729, 0.07526001, 0, 0, 0, 0, 0, 0, 
    0, 0.009360115, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.858257, 2.275796, 156.8928, 
    438.1283, 144.3511, 332.8229, 644.2934, 1112.633, 1770.227, 1851.317, 
    1377.889, 1208.554, 1110.734, 786.8075, 484.2887, 366.3296, 211.0903, 
    85.38182, 33.58828, 9.976434, 3.913893, 3.041174, 2.865082, 0.9683344, 
    0.04279455, 0.101553, 3.341461, 7.3607, 13.22865, 23.80757, 3.048281, 
    0.001522384, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.005946, 0.3337682, 0.005045555, 0.2996472, 0.481748, 0, 
    16.33418, 642.7941, 784.2194, 700.0764, 637.8699, 567.3324, 537.2572, 
    472.8118, 404.4005,
  501.8302, 469.2212, 394.8275, 271.4163, 217.2644, 213.8383, 249.5955, 
    323.6784, 477.7948, 605.2174, 541.8069, 309.9892, 182.302, 168.8128, 
    114.8026, 22.32053, 37.94635, 71.16721, 95.46755, 134.0202, 176.4655, 
    140.4458, 85.07382, 81.91493, 59.90077, 84.98973, 258.9031, 388.967, 
    721.7232, 837.8447, 678.611, 750.3956, 664.6459, 468.2991, 371.142, 
    271.4374, 124.6812, 65.89428, 7.602152, 124.1765, 989.6096, 2003.132, 
    2043.672, 1871.768, 1870.07, 1804.669, 794.097, 822.407, 942.0609, 
    591.2064, 739.2117, 944.7733, 1168.432, 1733.64, 1700.623, 1238.064, 
    508.2286, 143.446, 159.6475, 191.3692, 236.3782, 613.3393, 1667.213, 
    3066.058, 4324.365, 4945.152, 5141.235, 5196.927, 5175.205, 5119.337, 
    5073.023, 5025.966, 4892.131, 4874.926, 4949.278, 4573.41, 4439.014, 
    4543.262, 4350.15, 4316.033, 4160.53, 3570.559, 1925.418, 587.246, 
    362.684, 444.8941, 727.0997, 1051.035, 843.4271, 225.7823, 53.28727, 
    64.3373, 206.3961, 214.1255, 226.1105, 205.7556, 63.55518, 6.526137, 
    0.2235134, 0, 0, 0, 0, 0.6133821, 8.17198, 0.2726674, 0, 0, 0, 0, 0, 0, 
    0.05000988, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43.01835, 393.615, 277.4615, 
    121.3069, 547.8228, 1048.834, 1345.56, 1571.768, 1466.603, 1363.507, 
    1274.228, 1055.451, 780.6288, 656.064, 545.8841, 325.0826, 141.6882, 
    76.06046, 48.22424, 30.88945, 23.45646, 36.71673, 38.30359, 32.82429, 
    40.43208, 43.54045, 45.29679, 42.35429, 21.88343, 0.3880563, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.008802585, 0, 0, 0, 0, 675.0645, 1229.676, 1285.706, 1009.838, 
    735.5142, 673.9868, 596.0688, 561.3186,
  638.5468, 560.7847, 477.7018, 294.9648, 179.9539, 160.1006, 188.9391, 
    282.493, 419.4265, 514.0278, 492.7635, 211.3374, 49.51121, 30.31546, 
    3.770097, 12.51885, 112.3752, 178.5331, 148.6629, 125.5913, 92.01548, 
    107.0294, 33.9228, 4.764598, 2.675157, 5.054149, 23.91264, 133.9689, 
    505.7111, 720.3843, 723.8868, 818.0924, 672.5475, 410.331, 261.2775, 
    130.658, 21.59456, 9.977982, 61.48394, 500.2758, 1732.223, 2163.91, 
    1930.653, 1692.791, 1509.105, 1264.759, 728.9548, 1149.75, 948.2756, 
    575.9856, 724.7413, 982.3719, 1258.69, 1807.795, 2083.264, 1473.739, 
    558.8896, 171.6812, 178.2504, 199.0143, 465.3789, 1747.295, 3547.844, 
    4636.691, 5003.326, 5156.62, 5119.51, 4979.202, 4934.622, 4927.064, 
    4890.21, 4831.018, 4828.838, 4846.267, 4868.908, 4779.819, 4606.044, 
    4387.175, 4302.932, 4284.744, 4149.509, 3824.068, 3021.584, 1381.967, 
    574.1375, 558.4055, 798.3796, 1097.277, 1015.926, 385.0119, 123.4571, 
    132.1938, 243.8716, 112.4656, 56.71554, 37.44977, 8.20632, 1.903286, 
    0.01685685, 0, 0, 0, 0.01115504, 2.323969, 148.8537, 40.25793, 0, 0, 0, 
    0, 0, 7.943687e-05, 9.743791e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.000316862, 
    3.351332e-05, 108.9396, 627.876, 216.552, 264.3029, 775.5563, 1286.718, 
    1423.597, 1414.49, 1309.496, 1338.367, 1212.802, 954.1245, 811.7097, 
    694.0857, 522.5944, 340.141, 171.0701, 113.4646, 92.62653, 60.20259, 
    45.51564, 78.87679, 90.9756, 66.1013, 82.39753, 92.41844, 93.56767, 
    72.66559, 28.25791, 1.857119, 0.04283325, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0007546035, 0.001170857, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 474.17, 1027.907, 1430.493, 1542.452, 1107.297, 885.4199, 
    809.3794, 747.9736,
  883.4425, 737.2343, 611.8303, 384.4641, 172.8423, 119.4213, 138.5042, 
    242.9925, 260.4172, 191.402, 214.7129, 101.8246, 6.125151, 0, 0, 4.44872, 
    111.9656, 339.4658, 124.209, 3.618974, 0.9812769, 0, 0, 0, 0.004050649, 
    0.002791513, 0.02354521, 4.427878, 450.583, 767.4369, 754.4727, 809.8924, 
    655.1429, 394.2546, 174.1188, 50.06233, 72.33865, 244.7708, 607.683, 
    1398.816, 2134.434, 1855.941, 1529.018, 1318.995, 1173.078, 1040.517, 
    1007.168, 1545.558, 1140.663, 797.8842, 1160.718, 1585.277, 1698.333, 
    2127.591, 2229.236, 1780.801, 710.8757, 327.8267, 286.2559, 465.263, 
    1443.105, 3374.885, 4673.201, 4921.816, 4955.859, 4901.027, 4859.34, 
    4906.292, 4981.888, 4972.1, 4963.509, 4892.282, 4898.973, 4940.325, 
    4873.853, 4821.554, 4660.395, 4430.995, 4417.738, 4341.409, 4174.481, 
    3830.322, 3541.61, 2239.179, 1098.264, 1067.492, 1110.55, 1053.703, 
    711.0447, 279.4009, 159.6272, 112.0721, 66.18526, 35.84005, 37.72205, 
    14.1381, 3.197068, 0.5661116, 0, 0, 0.02646444, 0.004196592, 0.4673782, 
    7.541445, 218.5171, 95.47695, 4.138704, 0.4294933, 0, 0, 0, 0.08882221, 
    0.01487839, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01015859, 0.06481439, 1.590909, 386.5612, 
    423.8417, 185.4996, 351.5635, 634.8568, 1135.92, 1439.783, 1530.094, 
    1504.5, 1495.302, 1229.605, 1024.243, 871.163, 673.3406, 479.423, 
    329.9606, 193.3948, 136.8842, 103.0376, 69.0667, 45.88047, 70.47123, 
    111.1198, 83.07092, 112.5653, 162.7183, 161.994, 107.1, 56.84745, 
    18.48079, 2.352574, 0.01919217, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0009955933, 
    0.01022608, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004755442, 2.01799, 
    0.0546252, 0, 0, 0, 0, 58.31841, 361.321, 865.2963, 1518.639, 1445.205, 
    1221.712, 1169.723, 1055.812,
  1138.206, 1031.542, 798.9409, 491.9923, 161.3743, 58.14927, 96.90028, 
    169.3542, 88.08627, 10.73665, 0.3908091, 0.1588924, 0.0005378498, 0, 0, 
    0.02123698, 2.667614, 80.56416, 2.195054, 0, 0, 0, 0, 0, 0, 0, 
    0.002272809, 0.2845615, 460.1474, 877.2943, 712.2029, 679.8596, 530.2719, 
    337.3198, 116.6949, 51.26495, 382.4921, 1056.949, 1498.34, 1982.197, 
    2078.604, 1579.255, 1242.086, 1050.485, 938.3414, 1019.39, 1213.076, 
    1440.212, 1071.705, 1154.472, 1902.855, 2353.223, 2378.783, 2747.496, 
    2702.435, 2155.808, 1168.12, 565.398, 685.2184, 1640.354, 2973.905, 
    4407.279, 5010.863, 5079.21, 4995.299, 5025.908, 5005.139, 5018.24, 
    5057.439, 5076.51, 5134.964, 5131.24, 5150.346, 5019.635, 4794.578, 
    4773.021, 4691.179, 4526.166, 4496.824, 4406.292, 4202.837, 3751.894, 
    3462.172, 2578.806, 1484.944, 1260.712, 1121.709, 1028.017, 819.6217, 
    619.2815, 215.0901, 70.48732, 36.00191, 31.62999, 24.77269, 6.440446, 
    0.807209, 0.001755709, 0, 0, 0.1832342, 0.5934557, 0.04965257, 17.20242, 
    185.5353, 240.396, 293.856, 120.0528, 7.910353, 1.602257, 0.2335676, 
    0.3628228, 0.09872898, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004150902, 0.8579534, 10.77422, 
    122.1946, 651.1418, 418.1667, 310.4165, 507.0439, 741.2247, 1374.22, 
    1889.529, 2045.289, 1758.825, 1675.004, 1311.627, 1164.982, 973.3635, 
    679.0792, 419.1391, 305.7583, 221.5198, 158.1814, 121.2048, 84.55401, 
    52.9109, 57.2296, 100.5746, 119.8476, 184.5681, 246.9068, 256.8273, 
    173.4739, 106.7709, 54.65792, 15.56574, 1.09397, 0.05631513, 0, 0, 0, 0, 
    0, 0, 0, 0, 2.98584e-08, 0.0001462239, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.0008045597, 0.5715503, 0.01843894, 0, 0, 0, 0, 10.77944, 91.3958, 
    343.5856, 930.7227, 1321.466, 1175.285, 1166.477, 1162.554,
  1004.063, 1091.845, 939.7188, 635.8847, 243.0298, 288.0198, 447.8493, 
    297.6858, 55.81105, 0.5823933, 2.103457e-06, 0, 0.0003742431, 0, 0, 0, 0, 
    0, 0.03916743, 1.3382, 2.635849, 0.1669747, 0.05606115, 0, 0, 0.07838815, 
    0.1538332, 0.07272846, 303.3431, 817.912, 667.8759, 461.569, 310.2956, 
    263.948, 139.738, 164.9977, 745.8502, 1545.667, 1840.542, 1914.154, 
    1498.626, 1038.622, 908.1901, 814.3898, 759.5587, 908.0797, 1173.823, 
    1188.469, 1000.288, 1071.988, 1773.319, 2474.708, 2821.639, 3103.517, 
    3020.794, 2470.411, 1754.292, 1221.998, 1699.614, 2815.908, 3872.931, 
    4582.173, 5143.252, 5308.689, 5255.828, 5270.184, 5196.197, 5124.953, 
    5160.559, 5079.649, 5071.878, 5095.899, 5071.76, 4860.334, 4688.228, 
    4665.793, 4639.809, 4568.932, 4475.201, 4340.038, 4032.643, 3667.444, 
    3226.101, 2485.286, 1729.571, 1471.297, 1089.785, 825.2815, 812.0996, 
    649.4391, 248.7007, 78.42821, 46.15985, 51.71777, 51.22176, 17.32959, 
    0.186287, 0, 0, 0.008878704, 2.126103, 43.58032, 32.47812, 7.377217, 
    10.29517, 308.0126, 359.7991, 331.877, 236.2701, 141.4134, 114.9502, 
    4.1093, 0.1245182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.343631, 145.3042, 446.411, 672.5553, 
    929.6007, 635.9108, 636.684, 1070.611, 1433.741, 1769.073, 2049.272, 
    2187.267, 1905.526, 1801.605, 1439.334, 1259.708, 1051.37, 717.6959, 
    442.6573, 347.7022, 274.3106, 230.787, 258.9068, 184.7397, 90.33492, 
    65.87028, 109.6813, 164.0763, 237.5283, 302.2311, 401.8707, 401.7029, 
    220.2157, 114.113, 55.01257, 19.48724, 3.224457, 0.09818311, 
    9.276117e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.02179831, 2.024759, 55.57354, 345.5167, 725.6252, 
    676.2259, 819.7528, 962.77,
  533.136, 808.4719, 821.8669, 701.4637, 834.045, 947.1924, 826.0302, 
    468.552, 108.6253, 2.46531, 0.03890883, 0.1578468, 0.03584212, 0, 0, 0, 
    0, 0.0004631333, 0.8614438, 4.918919, 2.227592, 0.9925623, 1.058668, 
    3.265363, 20.65328, 3.438323, 5.87819, 0.6499826, 120.1984, 432.2348, 
    446.9734, 396.187, 278.4805, 245.8839, 221.1151, 433.9104, 1155.477, 
    1754.306, 1885.722, 1798.436, 1544.127, 1542.336, 1482.027, 1196.203, 
    945.9153, 989.442, 1270.374, 1455.62, 1095.746, 773.6746, 937.6028, 
    1641.641, 2335.161, 2614.873, 2491.024, 2671.889, 3219.281, 3111.022, 
    3284.736, 3563.545, 4307.58, 4980.42, 5343.886, 5250.076, 5233.35, 
    5191.366, 5082.385, 5030.96, 5118.875, 5041.934, 5022.34, 5011.443, 
    5018.072, 4864.628, 4655.928, 4501.825, 4330.26, 4182.997, 4146.882, 
    4085.304, 3616.214, 3329.208, 2700.405, 2153.664, 1860.559, 1541.81, 
    1264.337, 1010.502, 839.8696, 803.7663, 604.913, 220.8288, 46.89907, 
    100.4269, 177.4602, 91.5861, 9.258026, 0.007925773, 0, 0.02519359, 
    0.713772, 133.5067, 260.2882, 89.02231, 0, 60.87315, 228.1951, 146.3748, 
    223.1976, 480.6541, 852.3915, 267.9036, 8.180346, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25.11929, 
    345.4952, 620.2737, 1041.796, 966.2831, 884.076, 1010.437, 1472.149, 
    1751.677, 1779.012, 1963.424, 2108.116, 2078.134, 2042.505, 1619.692, 
    1292.49, 1071.784, 828.94, 561.9624, 404.3633, 295.3569, 238.5847, 
    287.1863, 276.2054, 159.8089, 87.40935, 110.5844, 173.6794, 257.0661, 
    349.3106, 506.4634, 666.3746, 481.9912, 247.4246, 136.2632, 56.22471, 
    12.78049, 1.750744, 0.006582987, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.536611, 278.9793, 
    85.00391, 15.20952, 124.8453, 330.4664,
  92.62735, 224.9857, 514.1376, 563.8992, 551.3384, 559.6557, 476.2484, 
    290.8705, 50.06903, 0.291686, 6.071148, 78.53983, 16.34308, 9.357828e-08, 
    0, 0, 0.007064464, 8.637155, 42.71983, 1.024719, 1.168388, 1.83171, 
    166.0009, 748.8835, 463.161, 440.6506, 900.9833, 557.688, 153.3299, 
    448.5606, 458.4509, 424.1318, 409.631, 441.6748, 550.0775, 1032.487, 
    1562.998, 1880.185, 1728.373, 1514.935, 1594.192, 1080.639, 901.5258, 
    1086.826, 1149.5, 1178.278, 1429.155, 1263.548, 673.6068, 442.3354, 
    524.1259, 613.4094, 690.2988, 1001.505, 1082.829, 1640.867, 3229.411, 
    3996.772, 4211.185, 4251.675, 4642.146, 4565.518, 4254.31, 3445.069, 
    2703.806, 2868.204, 3644.158, 4202.787, 4680.157, 4908.223, 4893.001, 
    4768.883, 4718.43, 4346.809, 3755.799, 3301.89, 3332.336, 3326.023, 
    3516.489, 3597.291, 3327.479, 2942.935, 2370.944, 1920.848, 1802.706, 
    1589.39, 1445.557, 1212.221, 1034.074, 1099.461, 958.3051, 360.7209, 
    43.27131, 123.7093, 205.6238, 73.54734, 36.61703, 14.14034, 0.1713255, 
    1.377384e-06, 8.600493, 122.1276, 301.5171, 259.4481, 0, 0.02519498, 
    0.7334027, 1.424428, 7.766448, 398.3439, 960.6716, 547.6946, 163.6535, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.1042083, 131.1837, 342.8325, 866.9229, 1492.76, 1177.958, 
    1114.048, 1149.951, 1522.847, 1785.231, 1748.308, 1874.776, 2057.966, 
    2382.843, 2433.188, 1962.085, 1487.279, 1100.362, 852.3791, 600.9429, 
    412.2162, 308.4789, 257.3823, 328.1452, 372.9504, 257.9034, 145.9283, 
    110.8266, 153.2345, 206.6768, 298.0198, 388.5441, 554.5134, 674.4021, 
    514.6151, 254.1146, 91.08628, 23.67842, 3.256741, 0.002150735, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04581926, 0.05429609, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4.728824, 27.6183, 27.00719, 229.8114, 202.5654, 
    337.5815, 168.5277, 6.976211,
  0.5517738, 4.567273, 2.20096, 3.175112, 10.09219, 84.83028, 42.51904, 
    4.969155, 1.45377, 1.626421, 120.8795, 404.1806, 71.52944, 1.297614, 0, 
    0.08654193, 5.740495, 393.6379, 362.3304, 7.257306, 1.757145, 34.62215, 
    506.4038, 1066.577, 1156.896, 1268.78, 1281.743, 1273.224, 916.1531, 
    970.4074, 847.1556, 749.6002, 745.4739, 943.8871, 1651.098, 1835.928, 
    1670.005, 1843.557, 1613.487, 708.126, 219.4308, -17.70356, -1.228317, 
    237.5716, 740.6729, 1210.737, 1261.4, 694.7611, 273.9698, 229.1583, 
    313.5432, 305.3273, 388.0406, 600.0505, 596.6004, 1015.485, 2594.182, 
    3940.926, 4462.644, 4441.323, 4032.217, 2831.896, 2035.072, 1546.722, 
    1310.755, 1335.621, 1559.156, 2119.01, 2941.616, 3871.328, 4326.727, 
    4253.578, 4093.514, 3429.374, 2819.071, 2883.427, 3393.673, 3687.75, 
    3875.096, 3793.733, 3556.442, 3079.378, 2229.497, 1687.628, 1493.1, 
    1463.086, 1443.055, 1221.478, 1131.022, 1237.433, 1085.7, 410.4431, 
    27.14528, 23.44693, 23.59412, 20.75784, 66.93874, 41.28713, 1.04267, 
    0.7734949, 9.972763, 109.714, 424.3781, 311.5717, 0, 9.578144e-05, 0, 0, 
    0, 9.431116, 212.359, 548.6569, 368.7649, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02470839, 13.6237, 
    173.7171, 524.9833, 1656.775, 1990.083, 1609.395, 1545.539, 1548.465, 
    1828.763, 1992.08, 1682.587, 1855.338, 2371.117, 2819.758, 2515.049, 
    1926.636, 1446.021, 1101.767, 854.6114, 626.3507, 463.8761, 372.9386, 
    306.1991, 301.629, 337.2941, 313.9757, 230.396, 150.8373, 137.3752, 
    164.8011, 235.8853, 306.9848, 398.2675, 554.8317, 642.8994, 439.2258, 
    131.188, 24.26292, 0.9274922, 0.02712296, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.07046242, 0.07160228, 0.1259949, 0.82448, 0.2724308, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 26.99575, 163.8403, 194.4064, 308.4962, 536.4026, 
    909.1552, 581.7653, 87.90736,
  5.524603, 0.2106795, 0.06117468, 0, 0, 0.001106707, 0.9858552, 2.084524, 
    0.007250982, 0.09791268, 8.467163, 148.3891, 40.20041, 133.1353, 
    1.050158, 0.698374, 95.08443, 603.4061, 346.568, 89.21722, 5.784426, 
    163.0823, 528.9404, 964.2617, 1224.283, 1145.506, 1083.035, 1260.024, 
    1514.948, 1620.2, 1329.965, 1212.592, 1243.346, 1558.333, 2080.932, 
    2112.273, 1593.904, 1573.761, 1264.198, 414.7022, -26.95219, -27.01832, 
    -25.83902, 43.31358, 289.6681, 545.9663, 370.5658, 162.3376, 137.683, 
    173.8771, 201.8835, 236.6482, 425.6211, 1204.362, 1562.504, 1771.867, 
    2764.249, 3997.256, 4503.231, 4179.479, 3119.117, 1704.98, 1232.164, 
    1188.176, 1179.922, 1170.334, 1163.777, 1190.092, 1321.959, 1878.314, 
    2652.745, 3296.654, 3190.252, 2823.26, 2837.28, 3232.735, 3871.69, 
    4173.316, 4095.113, 3523.542, 2740.75, 2067.219, 1480.583, 1389.877, 
    1357.177, 1341.039, 1356.684, 1236.902, 1205.911, 1409.923, 1086.137, 
    544.6427, 64.09715, 2.986501, 1.098339, 0.03515919, 0.5443146, 0.2935042, 
    0.1116209, 2.064476, 93.45126, 327.3704, 439.9635, 27.09679, 0, 0, 0, 0, 
    0, 0.0001652613, 1.751321, 135.4655, 314.1498, 14.58603, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.10488, 
    151.3687, 170.5209, 931.7928, 1869.477, 1960.295, 1962.794, 1915.189, 
    1871.135, 1854.007, 2212.921, 1781.809, 1864.471, 2385.011, 2960.157, 
    2591.642, 1815.004, 1382.749, 1117.803, 875.6705, 643.7021, 493.1649, 
    404.8751, 332.596, 276.7064, 264.625, 251.4656, 204.077, 158.8481, 
    146.3607, 171.6961, 223.1383, 256.2638, 267.8089, 332.9873, 573.2709, 
    628.1931, 245.8801, 51.25586, 9.667789, 1.074436, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.2100399, 1.297667, 0.4601581, 0.4224695, 0.1398023, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22.19897, 165.5422, 321.2482, 423.059, 574.9679, 
    813.0876, 775.3345, 253.5308,
  58.11911, 0.7057103, 2.670072, 0.1470038, 0, 0.005912722, 52.86464, 
    106.4483, 2.176097, 0.004030939, 0.01187678, 1.031699, 228.7305, 
    333.9132, 3.76192, 48.43727, 541.084, 665.0948, 76.33877, 1.491659, 
    27.94194, 270.8664, 549.6534, 931.3119, 1043.812, 1003.341, 1018.624, 
    1086.353, 1296.111, 1549.642, 1639.799, 1739.572, 1920.742, 1988.016, 
    1998.598, 1916.395, 1697.463, 1064.629, 351.8004, 33.46852, -26.99023, 
    -26.8875, 5.593151, 101.6692, 143.3968, 108.7655, 75.84795, 113.7356, 
    154.064, 173.8141, 184.0363, 239.2291, 425.3186, 1018.35, 1852.241, 
    2371.946, 2745.551, 3319.402, 3895.318, 3595.382, 2506.817, 1448.958, 
    1242.326, 1139.346, 1095.955, 1083.396, 1064.625, 1042.256, 1002.766, 
    940.4321, 977.5721, 1223.459, 1702.5, 1982.643, 2176.302, 2535.301, 
    3080.215, 3210.591, 2801.211, 2042.444, 1593.551, 1422.776, 1395.5, 
    1358.87, 1308.801, 1280.701, 1360.659, 1328.895, 1242.51, 1364.062, 
    1277.841, 1032.782, 431.9879, 40.43332, 36.72766, 32.49629, 11.74588, 
    54.25412, 36.6941, 26.17514, 171.8639, 416.9406, 188.8346, 0.003624032, 
    0, 0, 0, 0, 0, 0, 0, 7.249073, 330.5634, 245.694, 0.05019144, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1649839, 
    145.1682, 510.1442, 529.9858, 1373.305, 1634.407, 1616.854, 1965.759, 
    2036.208, 1918.154, 1634.574, 1946.693, 2036.997, 1901.531, 2226.949, 
    2786.348, 2683.617, 1752.335, 1401.295, 1125.746, 868.0985, 630.2976, 
    491.4984, 408.6, 335.9684, 282.6106, 240.715, 222.628, 189.7259, 
    184.9627, 189.7317, 209.8403, 258.7171, 280.8723, 273.613, 278.6961, 
    408.6448, 557.483, 305.4668, 138.5156, 58.12975, 14.19541, 0, 
    0.005009213, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03660801, 0.4714771, 0, 0.05864692, 
    0.008815271, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33.93098, 237.0571, 
    357.8159, 475.6015, 654.2646, 746.6953, 831.3919, 457.4333,
  267.8268, 13.05982, 1.384734, 0.0336902, 0, 0.1878956, 113.6884, 194.9467, 
    2.784834, 0.01134931, 5.906986, 107.6644, 543.8798, 267.7023, 43.91636, 
    142.7146, 880.8245, 668.0551, 191.1742, 96.54187, 79.51864, 164.2434, 
    178.9664, 387.0932, 672.4397, 1043.803, 1144.392, 1029.023, 976.5187, 
    1069.547, 1244.301, 1478.154, 1674.255, 2012.59, 1957.021, 1764.997, 
    1413.883, 738.8796, 437.0512, 115.4106, -25.63052, -26.77975, 6.702291, 
    120.8965, 158.2908, 87.91772, 85.55163, 124.0735, 144.6419, 163.9215, 
    194.0623, 271.6707, 454.1007, 569.8901, 570.1832, 886.5468, 1240.862, 
    1247.89, 1950.485, 3061.844, 2976.08, 2755.273, 2214.088, 1471.647, 
    1051.596, 993.2522, 966.7453, 938.7783, 916.3094, 925.144, 950.0883, 
    928.0298, 914.9496, 1071.79, 1252.155, 1377.319, 1549.455, 1775.616, 
    1551.019, 1333.115, 1171.915, 1219.383, 1375.59, 1337.319, 1262.59, 
    1230.977, 1223.931, 1321.175, 1302.679, 1394.339, 1378.148, 1211.746, 
    927.4117, 530.68, 421.3707, 365.48, 144.321, 52.77738, 193.9884, 
    288.5882, 477.8009, 953.6931, 890.5428, 311.8702, 4.768425, 0, 0, 0, 0, 
    0, 0, 2.971209, 255.346, 150.6877, 0.005446199, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5605842, 254.6885, 
    828.3015, 973.5774, 1576.689, 1508.777, 1474.373, 1709.781, 1908.645, 
    1738.698, 1497.87, 1873.77, 2274.448, 2016.283, 2112.831, 2522.752, 
    2471.199, 1593.402, 1312.828, 1083.33, 871.1516, 676.7658, 538.2769, 
    423.4112, 341.4968, 321.0897, 276.0688, 225.1823, 195.4746, 202.3975, 
    209.4864, 225.1591, 265.0031, 282.5084, 286.6417, 313.5991, 345.6582, 
    457.1176, 405.8619, 260.2231, 208.7539, 96.03938, 9.261443, 6.126817, 
    0.04181948, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 45.63474, 375.6396, 649.5263, 872.9135, 899.4869, 903.0366, 
    1095.192, 855.6779,
  445.0233, 351.4266, 38.30792, 0, 0, 0.1069812, 15.80168, 10.06809, 
    0.07949385, 30.06709, 334.9966, 506.3568, 290.8213, 12.22177, 0.2526761, 
    349.1699, 877.3591, 780.1846, 753.3016, 764.3349, 363.9612, 191.9262, 
    146.9533, 38.18995, 75.95718, 426.9885, 706.8687, 798.8369, 532.4489, 
    247.3566, 38.58874, 26.42688, 75.90255, 1111.113, 1620.344, 1350.999, 
    817.8193, 1236.167, 1223.355, 84.08205, -26.7035, -26.53172, -3.520207, 
    115.547, 165.4659, 90.80605, 69.04671, 93.5676, 108.3082, 126.1647, 
    198.4504, 275.4567, 263.6366, 277.3696, 272.9379, 846.3119, 1830.184, 
    1743.231, 1997.451, 2628.03, 2951.896, 3352.311, 3441.553, 2545.961, 
    1961.267, 1495.057, 1292.205, 1244.402, 1187.478, 1165.582, 1246.284, 
    1091.097, 955.6137, 1015.147, 1080.842, 1304.608, 1733.759, 1808.71, 
    1456.903, 1191.69, 1013.015, 1027.011, 1106.232, 1123.168, 1152.848, 
    1318.058, 1308.928, 1368.847, 1472.844, 1558.173, 1505.434, 1425.074, 
    1378.366, 1131.84, 898.5392, 647.2119, 309.5749, 91.7403, 130.3822, 
    366.4246, 588.8074, 860.438, 1172.794, 775.4387, 24.20318, 0.03165207, 
    1.964692e-05, 0, 0, 0, 0.1016023, 1.368763, 22.33897, 3.686608, 2.202234, 
    0.1302575, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.4327105, 278.1408, 1021.393, 1332.78, 1614.042, 1669.783, 
    1553.26, 1668.652, 1838.495, 1722.452, 1498.633, 1840.985, 2303.281, 
    2190.186, 2135.167, 2317.307, 2197.683, 1563.423, 1293.316, 1107.979, 
    928.3901, 725.1545, 563.6961, 431.3708, 373.5779, 349.8875, 283.476, 
    241.8707, 221.9501, 220.9182, 212.5661, 217.9307, 253.4073, 258.6729, 
    224.7961, 233.2203, 329.9741, 459.4734, 521.5692, 435.6661, 396.3931, 
    272.622, 156.6265, 70.35706, 15.06063, 0.1001706, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57.15924, 447.7066, 
    728.2842, 807.1526, 886.8223, 1057.768, 922.2719, 611.8473,
  1185.601, 1075.845, 253.8555, 0.3205906, 0.1802309, 1.888118, 0.1392453, 
    0.4834277, 8.630255, 321.5133, 594.8525, 250.4044, 19.79789, 14.29809, 
    405.394, 850.6742, 895.6686, 771.8899, 889.6099, 654.85, 445.857, 
    247.8456, 50.42672, 0.06561425, 0, 0.04161381, 11.48845, 8.107579, 
    6.262373, 0, 0, 0, 141.3629, 722.8207, 1543.16, 1645.606, 1591.569, 
    1533.112, 511.8043, -20.16574, -27.00284, 2.159925, 84.06423, 138.6476, 
    162.7526, 119.8016, 85.98859, 76.00282, 91.5968, 107.9918, 194.1754, 
    264.5587, 223.5369, 199.5766, 249.1336, 642.5747, 1418.234, 1740.475, 
    1847.636, 2013.859, 2290.76, 2693.301, 2895.988, 2929.51, 3072.078, 
    2562.047, 2377.528, 2421.979, 2456.333, 2114.605, 1433.238, 1013.753, 
    915.5472, 793.4993, 944.1635, 1421.511, 1579.745, 1507.955, 1295.6, 
    1159.868, 1106.175, 1209.779, 1293.367, 1320.985, 1202.004, 1099.803, 
    1159.94, 1207.144, 1184.125, 1199.408, 1223.053, 1255.663, 1328.157, 
    1350.471, 1151.386, 665.4273, 436.4703, 230.356, 126.5837, 253.5839, 
    424.1454, 606.5503, 820.1623, 631.6375, 171.5208, 39.03421, 95.25896, 
    14.42945, 0.01480233, 0, 0.003400196, 3.222284, 64.84809, 152.0146, 
    172.1592, 40.11589, 0.3631265, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.8056216, 286.8983, 820.6075, 1408.043, 
    1595.236, 1589.162, 1507.651, 1523.362, 1459.125, 1535.912, 1564.839, 
    1840.154, 2311.229, 2240.042, 2052.285, 1974.945, 1832.499, 1422.568, 
    1221.401, 1075.178, 893.7475, 680.9863, 529.2756, 431.7417, 401.8191, 
    359.3887, 321.6649, 294.0847, 276.5602, 264.9191, 241.834, 191.1283, 
    247.5713, 261.2683, 226.9597, 196.604, 261.0652, 345.585, 434.86, 
    370.0406, 422.851, 394.8878, 309.2286, 185.3647, 34.64439, 0.1407993, 0, 
    9.415688e-05, 0.0006615912, 8.456256e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 69.2422, 497.5997, 839.9404, 945.6211, 
    913.7177, 848.2019, 697.5277, 883.2184,
  325.7719, 389.6647, 366.6138, 170.5247, 286.1557, 350.3175, 27.14322, 
    4.930077, 157.9842, 383.1822, 301.3425, 15.31997, 145.7745, 533.2792, 
    860.9586, 962.8611, 729.6182, 503.8995, 427.0553, 289.4353, 216.7994, 
    225.476, 124.4237, 1.019406, 0, 0, 0.001557372, 0.05312407, 0, 0, 0, 
    279.2541, 1210.337, 1751.807, 1364.346, 682.6356, 379.4771, 135.9984, 
    -11.6577, -26.98977, -9.718063, 72.4333, 158.9611, 156.7875, 184.3431, 
    154.4228, 109.7353, 64.25401, 61.09314, 72.82911, 127.2696, 170.9054, 
    172.7442, 195.3659, 353.7366, 458.7604, 534.1633, 612.3792, 738.5699, 
    923.3236, 1088.91, 1325.916, 1430.023, 1399.115, 1513.199, 1719.383, 
    2224.956, 2811.51, 2849.411, 2167.947, 1620.381, 1313.227, 1219.847, 
    1241.146, 1430.529, 1401.99, 1035.019, 1255.08, 1272.251, 1211.268, 
    1359.349, 1538.417, 1574.35, 1589.597, 1468.608, 1209.066, 979.7721, 
    1010.157, 1041.08, 1037.924, 1042.378, 1094.071, 1200.066, 1282.567, 
    1038.127, 630.5131, 343.8075, 221.8435, 160.7519, 189.7369, 293.0468, 
    441.797, 590.9557, 559.6724, 453.6119, 300.0871, 407.3008, 433.2998, 
    96.88019, 1.46743, 0, 0.8922319, 140.732, 341.529, 416.4601, 176.4161, 
    7.827775, 0.2349445, 0.01798946, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.208533, 128.4021, 628.1529, 1293.599, 1466.538, 
    1467.676, 1360.863, 1146.859, 1498.528, 1869.94, 1736.707, 1803.207, 
    2405.826, 2367.827, 1854.521, 1755.475, 1548.718, 1361, 1130.83, 
    880.1629, 721.251, 558.7914, 463.0948, 449.2039, 434.8761, 366.6079, 
    360.2966, 335.5677, 305.4737, 286.3239, 253.7291, 193.3935, 260.425, 
    245.9069, 214.7218, 224.1293, 304.7106, 192.1682, 154.5506, 138.489, 
    312.5544, 434.146, 375.9181, 324.3535, 135.5652, 18.72083, 0.3908859, 
    4.178871, 21.68737, 1.068586, 0.04165883, 0, 2.302622e-05, 0.000318967, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25.86181, 181.0313, 
    324.3846, 368.098, 288.4367, 168.3377, 149.3321, 269.4598,
  134.7829, 383.3967, 751.2313, 616.4398, 948.6702, 1276.596, 479.7618, 
    325.3689, 323.8741, 201.3069, 72.01556, 167.9449, 407.1801, 650.3666, 
    556.2456, 370.9961, 256.1597, 351.5567, 307.9527, 238.6851, 204.8227, 
    87.6537, 54.47084, 12.21142, 0.04147403, 0.0936074, 5.353564, 25.28491, 
    1.579029, 1.649322, 88.01975, 380.4411, 529.6, 575.6082, 416.7852, 
    163.9062, 29.59988, -18.3385, -26.71364, -26.81509, -6.779469, 55.93732, 
    80.90195, 109.7946, 131.4983, 156.0971, 143.4567, 37.21712, 41.79709, 
    66.11372, 88.39603, 108.0333, 131.4864, 183.6172, 300.5077, 309.0844, 
    312.2074, 337.2733, 406.8892, 506.1661, 480.3888, 566.5581, 985.7548, 
    1719.474, 1873.253, 1391.59, 1125.062, 1051.788, 731.9938, 530.9971, 
    659.5547, 845.972, 1076.787, 1334.669, 1314.29, 1201.588, 1428.955, 
    1555.712, 1675.069, 1713.571, 1542.403, 1488.172, 1371.695, 1288.64, 
    1306.404, 1200.959, 1098.898, 952.856, 952.5204, 1062.195, 1148.485, 
    1181.134, 1108.441, 1078.962, 1075.35, 827.2219, 459.4761, 212.3748, 
    156.4711, 174.78, 195.3211, 298.1235, 511.4929, 546.0997, 458.4923, 
    248.5788, 264.8895, 461.7291, 364.6042, 78.57813, 0.130757, 0, 2.51242, 
    137.8275, 73.93156, 29.94359, 2.122291, 1.151326, 0.4277129, 0.0282865, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01295927, 
    33.24023, 392.3328, 1000.464, 1125.371, 1295.121, 1356.886, 1306.639, 
    1829.415, 2189.526, 2142.537, 2038.699, 2414.614, 2220.198, 1697.196, 
    1618.274, 1323.614, 1244.735, 1006.082, 736.7032, 595.5756, 517.9122, 
    467.2306, 467.5121, 392.7173, 317.6983, 311.0505, 317.7751, 333.4388, 
    328.5473, 249.2917, 193.0846, 285.6727, 300.2908, 209.6806, 178.5817, 
    298.3004, 291.2953, 256.2574, 158.7208, 162.479, 355.959, 337.4423, 
    418.3747, 338.9467, 119.6824, 46.85309, 24.59101, 64.62159, 71.26684, 
    39.46763, 6.434648, 0.2060366, 0.0007213038, 1.44927e-05, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1687387, 1.76992, 3.556161, 3.130101, 
    1.38521, 0.2365721, 16.18559, 64.20919,
  198.5991, 513.2113, 706.6056, 582.6232, 820.0352, 1709.845, 902.1078, 
    573.4025, 628.8603, 291.3704, 231.4335, 471.0799, 364.6606, 195.7161, 
    165.8737, 98.94559, 108.8485, 364.8844, 691.4595, 759.3024, 653.2693, 
    400.0212, 90.88813, 29.91551, 2.056026, 2.457185, 57.52008, 72.7826, 
    2.53535, 6.038398, 24.17636, 58.83421, 112.778, 187.0657, 168.954, 
    98.36449, 11.12561, -20.56032, -26.30639, -26.99186, -25.81065, -22.9365, 
    -20.77874, 5.6212, 63.99236, 105.8428, 118.9219, 41.40837, 37.70866, 
    62.69654, 88.21542, 111.4256, 134.1934, 159.343, 212.6318, 260.1141, 
    323.3558, 394.4828, 446.9649, 381.2402, 356.7253, 383.8136, 508.8347, 
    998.1973, 1568.436, 1380.85, 1055.252, 769.7596, 414.7127, 427.1404, 
    653.4495, 906.3173, 1187.628, 1423.794, 1745.533, 1805.913, 1899.968, 
    2023.965, 2007.942, 1825.254, 1764.472, 1708.418, 1487.05, 1358.287, 
    1345.907, 1268.355, 1168.33, 1059.39, 1016.202, 1017.433, 1119.964, 
    1242.388, 1085.921, 959.4313, 947.9687, 928.6378, 663.5068, 319.8902, 
    159.1487, 135.6131, 155.1372, 196.0303, 276.0444, 376.324, 343.4353, 
    201.4925, 133.8106, 305.9968, 565.4852, 311.8119, 42.69448, 0.04077369, 
    0.6807221, 1.09381, 0.06465454, 0.005266901, 0, 0.5601527, 2.024031, 
    1.411731, 0.6386642, 0.04973439, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.05632153, 86.15315, 288.2992, 646.9312, 769.1035, 746.407, 
    1086.887, 1312.366, 1677.646, 1946.63, 2020.579, 1931.543, 2009.922, 
    1664.603, 1315.809, 1141.892, 1023.728, 997.9595, 879.2858, 726.4648, 
    598.501, 543.4471, 450.1937, 405.8009, 362.7404, 343.9048, 309.5486, 
    346.8863, 413.1714, 444.4728, 336.5836, 212.6304, 197.2327, 241.4291, 
    195.5558, 185.1576, 209.467, 313.4066, 342.7289, 245.5191, 184.3604, 
    153.5431, 117.784, 295.8724, 445.2908, 297.1679, 156.8097, 106.7463, 
    107.714, 111.64, 106.2599, 92.36662, 22.72518, 1.638889, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0004705076, 5.859629, 
    54.95887,
  153.1524, 282.0642, 365.8515, 357.7076, 540.0745, 1189.793, 1465.544, 
    1557.793, 1650.682, 1476.673, 1084.294, 837.059, 483.3738, 202.0709, 
    151.347, 111.004, 96.51801, 252.1635, 535.3167, 678.3774, 698.8224, 
    450.3364, 170.493, 91.76162, 34.39745, 18.04377, 26.07745, 31.38563, 
    31.87274, 8.058367, 10.27361, 38.7353, 64.00056, 74.72749, 86.04457, 
    66.1438, 6.460943, -14.82185, -20.84778, -23.86658, -25.58394, -26.80298, 
    -23.79078, 1.873433, 55.98904, 105.269, 135.2005, 113.2983, 89.9667, 
    79.32413, 100.5755, 126.9466, 162.0791, 231.5735, 261.4696, 318.9235, 
    426.7239, 502.1569, 495.2846, 418.2052, 390.8795, 414.4824, 434.062, 
    442.893, 543.8828, 743.8888, 1086.514, 1229.295, 1004.674, 680.251, 
    665.8293, 1017.3, 1776.176, 2193.851, 2130.682, 1879.952, 1860.84, 
    2093.249, 2183.176, 2157.849, 2272.139, 2177.936, 1765.554, 1538.141, 
    1443.227, 1404.861, 1322.967, 1240.981, 1168.145, 1108.121, 1035.654, 
    984.2963, 895.5591, 828.546, 892.6108, 989.7599, 845.5907, 466.0449, 
    207.6372, 140.435, 156.4812, 180.6231, 262.96, 301.4807, 225.4205, 
    133.5546, 133.4378, 204.3734, 464.5609, 675.4373, 239.2331, 3.794266, 
    0.07450061, 0.2229451, 0.3089383, 0.130912, 0, 0, 0.1550962, 0.7067999, 
    0.932089, 0.8703596, 0.1680117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1565143, 60.53839, 331.5735, 751.3165, 744.5818, 429.5865, 
    572.5468, 901.7349, 1331.926, 1643.574, 1789.187, 1660.139, 1668.764, 
    1337.937, 1026.51, 917.7629, 868.0641, 859.9366, 814.2829, 697.3281, 
    593.4163, 558.0633, 417.3791, 348.2489, 386.9695, 399.5235, 366.4043, 
    355.6556, 369.4089, 402.4993, 357.6656, 244.9649, 219.8819, 280.3364, 
    337.7258, 331.6732, 287.1907, 307.7718, 340.4637, 315.8674, 323.7686, 
    363.6587, 254.7796, 220.4984, 327.1406, 347.2398, 252.6705, 213.0592, 
    111.2491, 34.6552, 7.621826, 26.68723, 144.1777, 8.461684, 0.001237476, 
    0.2612488, 0.8080437, 2.007894, 0.9289774, 0.1346615, 0.0009252121, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04167476, 25.30412, 77.0424,
  109.2693, 137.8501, 205.5703, 313.439, 320.2293, 529.5438, 747.915, 
    979.4609, 1234.923, 1255.769, 1217.286, 1052.158, 647.5029, 252.7099, 
    178.4732, 179.3629, 131.0711, 166.9237, 373.0456, 688.7805, 677.8123, 
    328.6298, 164.0024, 143.9124, 113.7872, 94.8535, 82.46211, 79.49993, 
    95.83374, 133.3086, 99.34294, 93.74997, 74.08489, 67.71928, 85.51957, 
    61.66181, 11.11381, -7.539976, -12.29743, -16.15827, -18.99532, 
    -20.94397, -11.43562, 35.05849, 110.7344, 147.3769, 201.0651, 197.6199, 
    145.2554, 87.56669, 85.93134, 126.8988, 246.3241, 378.7465, 354.4667, 
    368.2503, 476.5359, 630.2359, 667.1591, 604.4746, 566.3921, 593.0729, 
    606.2556, 561.368, 677.4869, 898.1255, 879.7053, 964.821, 974.934, 
    868.2034, 1068.178, 1840.587, 2423.719, 2145.945, 1629.781, 1540.773, 
    1735.503, 2207.301, 2549.122, 2488.623, 2228.458, 1826.002, 1508.05, 
    1334.651, 1338.239, 1490.489, 1497.013, 1373.759, 1225.087, 1105.78, 
    1012.007, 865.905, 730.3913, 653.7793, 722.3007, 922.6825, 972.0062, 
    645.337, 281.5837, 175.0263, 198.771, 250.4568, 361.6537, 392.6619, 
    205.9537, 78.29983, 64.51853, 112.582, 307.3622, 675.9061, 652.8943, 
    149.5045, 3.725435, 0.3590779, 0.4722362, 0.007159858, 3.080651e-06, 0, 
    0, 0, 0.08578687, 1.846867, 0.5791237, 0.00559359, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.698241, 93.83714, 401.8361, 659.1234, 922.0559, 
    611.1923, 661.2104, 887.2751, 1258.764, 1389.879, 1643.886, 1349.247, 
    1242.34, 1047.991, 886.8261, 813.6723, 773.3261, 735.2281, 711.2335, 
    642.8856, 558.7678, 508.3784, 411.021, 314.9867, 378.224, 413.6927, 
    412.9915, 439.1799, 304.6605, 207.3989, 183.205, 179.3029, 189.8379, 
    391.1242, 440.8367, 404.01, 351.9052, 300.9068, 334.468, 377.8862, 
    412.4525, 449.847, 419.4991, 469.8304, 428.1302, 306.8965, 312.2477, 
    290.9785, 147.2815, 10.9004, 0.03723383, 0.03549428, 0.1414406, 6.996796, 
    124.846, 59.08067, 113.4522, 96.42812, 93.694, 7.924925, 9.195313e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01162703, 1.734384, 26.52215, 54.8782, 
    82.08762,
  142.3178, 130.4512, 133.4851, 203.8016, 278.6282, 345.01, 429.7573, 
    523.0563, 517.8198, 534.1415, 583.5115, 567.5313, 468.8252, 326.0786, 
    334.3853, 468.4581, 402.1276, 305.6375, 512.864, 632.5613, 419.8971, 
    246.6624, 228.2628, 211.8145, 184.6159, 157.7082, 137.1225, 105.3211, 
    120.6595, 143.6004, 157.1687, 153.8044, 118.5471, 107.4489, 98.0548, 
    65.00665, 19.89009, 3.944678, 0.105921, -6.533163, -9.39222, -6.86598, 
    9.422341, 73.79856, 153.5831, 218.1455, 272.2792, 252.624, 171.2262, 
    109.0305, 99.97236, 151.3901, 284.1615, 442.0058, 460.5809, 424.026, 
    471.3872, 589.5248, 719.0064, 826.4303, 841.942, 816.5634, 777.521, 
    753.3342, 745.238, 750.7159, 590.8809, 764.2705, 1175.475, 1658.203, 
    2217.382, 2441.069, 2252.371, 1752.251, 1352.165, 1472.647, 1858.281, 
    2133.639, 2239.722, 2144.459, 1869.276, 1608.337, 1424.721, 1203.038, 
    1142.748, 1422.119, 1655.942, 1500.4, 1279.54, 1091.823, 949.7327, 
    798.5269, 718.2721, 644.5741, 638.3768, 757.2607, 905.2473, 781.3608, 
    468.7405, 278.3626, 277.8269, 340.9755, 390.8184, 372.8437, 292.4178, 
    225.0815, 138.0792, 67.86915, 124.9117, 453.0229, 721.0461, 555.2239, 
    155.6841, 21.86419, 8.730263, 0.7218965, 0.0008120779, 0, 0, 0, 0, 
    0.1688487, 0.5500224, 0.5095904, 0.1417561, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1.393449, 22.25437, 354.1327, 515.7268, 827.9959, 1168.326, 
    1064.139, 956.5106, 1098.677, 1281.468, 1450.56, 1442.861, 1148.374, 
    983.0171, 928.001, 847.0422, 791.1342, 750.2274, 683.267, 662.6528, 
    591.2401, 499.2674, 479.2394, 402.3772, 287.5651, 342.9493, 365.4809, 
    388.0802, 437.3572, 459.0589, 358.643, 235.0905, 242.1442, 351.9156, 
    382.6072, 352.2855, 323.7015, 310.036, 307.3141, 317.7708, 358.8003, 
    421.9719, 452.568, 414.5871, 399.4982, 466.2424, 320.7542, 202.3461, 
    334.6939, 289.0134, 79.38692, 1.849855, 0.005193034, 0.02077778, 
    17.88385, 245.8173, 317.0123, 214.2401, 137.7892, 25.72491, 0.4853109, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8479855, 36.25705, 99.17735, 84.4957, 
    119.1772,
  62.87701, 118.0103, 108.4703, 175.6332, 303.9168, 306.817, 252.5901, 
    329.449, 414.6758, 479.0469, 511.3866, 474.5561, 423.2299, 406.1709, 
    401.9231, 561.6601, 557.7254, 389.787, 368.4766, 348.583, 319.0773, 
    287.6952, 272.9836, 231.125, 183.0162, 140.632, 110.0775, 119.4187, 
    137.2057, 140.2922, 142.3265, 137.8181, 141.4195, 133.079, 126.9698, 
    97.08437, 52.76869, 24.86823, 16.72916, 6.681043, 1.103742, 5.227499, 
    36.38683, 109.372, 183.0074, 263.3933, 319.1121, 299.4172, 226.264, 
    159.8448, 127.9879, 143.6917, 225.7771, 412.8821, 469.8937, 410.8768, 
    433.6516, 503.0591, 617.9167, 732.0046, 801.3393, 753.6541, 591.4202, 
    465.1469, 446.1022, 565.3156, 802.3586, 1062.787, 1670.608, 2156.022, 
    2500.713, 2417.878, 2072.402, 1807.993, 1350.391, 1421.16, 1728.899, 
    1978.551, 2038.647, 1897.298, 1665.599, 1449.603, 1309.755, 1145.813, 
    978.3882, 1039.86, 1290.916, 1457.758, 1417.414, 1206.094, 974.1864, 
    800.8099, 703.1967, 691.4738, 660.6443, 675.6011, 778.5321, 814.866, 
    609.2058, 388.8049, 362.1662, 367.7457, 257.1624, 213.0947, 320.0247, 
    444.534, 418.0684, 311.0552, 184.6308, 228.825, 537.2193, 585.6755, 
    233.2688, 192.6097, 224.1531, 39.27412, 0.1964533, 0, 0, 0, 0, 0, 
    0.2488128, 1.523081, 0.5462044, 0.01051013, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02214108, 7.466173, 313.21, 434.3052, 607.8076, 753.3428, 1079.435, 
    1312.072, 1285.051, 1323.413, 1505.258, 1537.162, 1557.59, 1129.629, 
    935.6879, 922.4156, 913.1953, 860.5278, 810.3507, 739.6919, 658.9257, 
    619.9458, 564.9073, 487.7058, 425.2112, 320.0811, 262.0454, 324.9103, 
    361.2815, 389.5933, 418.6406, 450.1284, 409.5188, 346.2076, 344.7409, 
    304.8754, 275.0458, 249.2003, 243.0425, 274.7803, 283.5438, 287.1927, 
    316.4399, 370.9124, 409.6602, 400.5841, 402.0221, 465.1623, 410.8765, 
    243.9812, 198.312, 85.20193, 47.56075, 5.244726, 4.087999, 4.323982, 
    1.389558, 118.9203, 213.591, 73.54279, 22.31983, 6.615984, 0.01501575, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001105127, 0.01574967, 0.3731294, 1.408006, 
    0.7327028, 12.36994, 51.13934,
  2.496701, 56.47428, 67.3052, 134.3256, 236.7472, 283.3006, 297.1014, 
    321.1642, 374.1868, 426.1517, 442.9759, 357.7471, 395.6037, 376.1304, 
    296.0233, 281.6389, 256.8011, 239.3192, 230.0778, 232.7337, 227.1398, 
    230.698, 216.167, 181.7157, 137.8015, 125.5255, 137.2948, 150.386, 
    170.2027, 177.3434, 166.3967, 157.8046, 147.7821, 136.5725, 134.4278, 
    149.0592, 111.9832, 56.63974, 43.25705, 30.75291, 22.94107, 40.6287, 
    81.01137, 142.7441, 191.9426, 265.1708, 321.9136, 309.4189, 280.8097, 
    236.9384, 186.9155, 164.3916, 204.4578, 303.1568, 331.4703, 341.3737, 
    373.5767, 437.0652, 517.2995, 521.5381, 505.0607, 409.2562, 291.2585, 
    252.2856, 286.6728, 403.5825, 820.5607, 1288.641, 1583.237, 1858.465, 
    2120.359, 2305.981, 2002.771, 1417.134, 1102.36, 1222.863, 1556.939, 
    1840.42, 1989.827, 2013.498, 1853.452, 1559.529, 1452.16, 1284.551, 
    944.7426, 854.6462, 979.381, 1144.847, 1253.435, 1237.704, 1003.507, 
    808.721, 735.7459, 782.2019, 760.3269, 694.5384, 790.4561, 861.2177, 
    712.9924, 522.0662, 427.1132, 332.0608, 215.898, 246.2131, 372.9935, 
    523.418, 674.3666, 853.593, 527.9724, 333.238, 391.3175, 471.9327, 
    115.2076, 94.95418, 188.1124, 8.46489, 0.03515024, 0, 0, 0, 0, 0, 
    0.01253535, 0.2055177, 0.5415505, 0.7795085, 0.8468797, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01696419, 0.0234534, 0.002375286, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002031238, 0.1419092, 114.2471, 
    479.0662, 786.2939, 1173.355, 1488.77, 1342.881, 1201.569, 1209.84, 
    1434.139, 1680.65, 1746.331, 1527.47, 984.627, 787.7053, 770.4208, 
    763.9011, 735.5531, 688.8949, 625.7838, 603.2035, 609.0561, 552.9663, 
    509.5374, 370.9828, 265.0435, 240.4553, 303.8818, 369.0324, 393.3753, 
    403.44, 413.787, 377.8459, 331.9669, 290.3476, 210.9386, 163.0418, 
    142.3099, 129.1365, 146.474, 173.871, 225.6789, 283.9551, 342.0289, 
    398.8251, 466.3244, 514.8624, 550.3365, 540.9114, 486.1489, 402.7083, 
    343.3196, 258.5035, 183.5906, 161.7388, 129.7702, 47.80243, 59.13809, 
    203.2783, 48.43516, 0.05176627, 0.01542342, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02726323, 0.000588363, 0.0147949, 0.6816624, 85.19174, 64.90533, 
    49.62014, 9.959903,
  32.80307, 7.98277, 5.168087, 19.52959, 48.15039, 114.1893, 241.8551, 
    263.4387, 265.8207, 195.31, 167.5222, 178.9858, 166.7894, 139.4841, 
    157.5792, 178.5267, 180.3525, 174.2237, 172.9613, 170.9986, 162.9474, 
    160.7891, 159.3648, 145.4607, 126.892, 134.1567, 149.6773, 173.2433, 
    194.7241, 206.9443, 184.6305, 153.8452, 144.0511, 140.9794, 155.5726, 
    183.1039, 159.2662, 94.48742, 68.51237, 77.47488, 86.63057, 91.22647, 
    109.4375, 151.3914, 186.838, 280.7965, 324.8289, 318.7262, 312.5193, 
    267.868, 232.0612, 189.1541, 236.293, 287.5121, 315.8879, 333.0435, 
    351.8202, 369.1386, 369.0467, 310.4318, 246.0696, 178.6416, 159.8972, 
    182.2894, 243.0864, 317.7323, 570.7515, 862.8789, 967.5267, 1198.933, 
    1629.652, 1804.37, 1549.987, 1379.818, 1285.188, 1221.166, 1338.393, 
    1609.639, 1911.138, 2070.336, 1997.709, 1690.824, 1356.69, 1095.801, 
    956.0564, 823.9498, 863.5275, 944.6961, 1017.248, 1027.37, 948.0721, 
    839.8313, 767.9204, 811.2511, 819.8428, 785.5138, 812.5242, 876.9158, 
    857.1652, 650.3183, 466.8417, 296.4872, 234.0867, 238.503, 398.3628, 
    608.6905, 781.9844, 831.3923, 540.4121, 273.7153, 315.2288, 271.1372, 
    116.3179, 44.71602, 121.1515, 13.66153, 0, 0, 0, 0, 0, 0, 0, 0.04417975, 
    0.7995526, 73.27557, 36.45834, 2.02336, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.3590926, 0.7031543, 0.4019015, 0.5328932, 0.9531209, 1.510096, 
    1.552819, 0.5022201, 0.05853625, 0.08055027, 0.0227679, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.07241476, 0.4991371, 2.517156, 173.3939, 763.7124, 1414.628, 1499.819, 
    1455.987, 1261.048, 1178.42, 1317.442, 1683.426, 1930.743, 1779.641, 
    1261.818, 920.3959, 795.5938, 737.7306, 691.3679, 641.2322, 589.3427, 
    566.7949, 568.4863, 572.6649, 520.2504, 467.4853, 299.2236, 251.0989, 
    242.6156, 302.4815, 365.5584, 396.1295, 402.2466, 383.4164, 345.4184, 
    298.8433, 240.6213, 176.6061, 125.182, 82.32549, 58.15251, 23.40827, 
    42.75769, 130.3623, 233.3544, 307.3527, 362.999, 462.8122, 571.1421, 
    611.3059, 596.0009, 597.5264, 616.5421, 606.6191, 610.8198, 516.1464, 
    422.0352, 355.8859, 269.934, 205.9718, 197.3346, 98.00138, 1.487198, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.1164714, 2.149752, 81.73408, 10.18455, 
    1.231145, 2.270527, 158.2819, 144.1404, 115.0255, 80.37354,
  30.25532, 15.22529, 0.05774624, 0.5911842, 6.755296, 23.15621, 62.50331, 
    92.66872, 96.67418, 72.09167, 59.09659, 67.65337, 75.2924, 90.40241, 
    97.29047, 108.9601, 120.2069, 129.2026, 150.1645, 155.3292, 155.1979, 
    150.6721, 141.9426, 138.1929, 136.4271, 151.1962, 170.1705, 189.2829, 
    207.9605, 211.88, 197.2425, 164.0269, 151.9234, 158.4813, 180.417, 
    204.455, 209.0111, 182.1513, 121.6905, 95.39534, 105.0443, 124.1743, 
    160.6243, 199.5449, 248.7912, 376.4545, 465.8036, 376.5368, 308.0159, 
    249.9769, 206.0722, 184.5465, 217.6384, 271.2474, 336.8931, 346.9473, 
    323.7444, 263.5324, 191.4721, 142.6588, 124.904, 117.0247, 128.5519, 
    142.0424, 193.5832, 215.9247, 246.0654, 300.1264, 354.4006, 492.1281, 
    755.2769, 1022.38, 1090.596, 1099.709, 1157.982, 1194.312, 1254.268, 
    1455.788, 1766.926, 1941.656, 1782.409, 1254.401, 793.8506, 688.838, 
    701.832, 784.8435, 912.9474, 984.9802, 1033.975, 1033.87, 1014.515, 
    942.2949, 843.1401, 761.8826, 757.4646, 717.6158, 703.0925, 731.7596, 
    700.3924, 546.201, 384.6826, 300.0076, 282.5623, 273.2426, 375.3759, 
    552.0548, 892.2322, 978.8475, 624.9924, 291.8902, 261.8087, 216.2638, 
    153.5658, 98.59215, 38.25227, 1.961729, 0, 0, 0, 0, 0, 0, 0, 
    1.982099e-06, 13.43534, 241.5155, 230.8685, 37.0118, 1.989155, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.6743881, 1.812494, 0.5765836, 0.07700097, 0.2077032, 
    0.174242, 0.1472005, 0.4762342, 1.132957, 1.511994, 0.8909723, 1.494937, 
    0.9272659, 0.4672569, 0.7380159, 1.100274, 0.4356244, 0.2224446, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.5607325, 5.209057, 3.908259, 84.57672, 487.4668, 1081.089, 1322.505, 
    1292.228, 1100.757, 1051.505, 1442.053, 1669.606, 1819.919, 1803.941, 
    1396.308, 969.9709, 817.9538, 741.9974, 691.8995, 652.3807, 609.4356, 
    556.4875, 526.7487, 524.3944, 513.6147, 473.0761, 361.2754, 259.5472, 
    226.2071, 248.5821, 299.0684, 334.5462, 348.5111, 350.0092, 334.2562, 
    296.7508, 256.1983, 207.6281, 158.5576, 112.5472, 57.24558, 24.61476, 
    6.21199, 13.57706, 100.3118, 211.8075, 297.1721, 371.2862, 455.0604, 
    547.5605, 631.9322, 635.8278, 636.6499, 597.9122, 587.1418, 554.1342, 
    509.644, 445.5923, 405.0834, 395.6985, 344.6743, 274.5173, 103.2803, 
    0.9090499, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.08440799, 1.223302, 110.108, 
    86.23002, 88.89346, 27.88332, 166.7321, 192.7967, 124.4891, 72.08824,
  2.412836, 0.2777807, 0.02403365, 0.05077571, 0.8098862, 3.15499, 7.584254, 
    23.98851, 34.31339, 38.25267, 41.14117, 41.33563, 82.49149, 99.42232, 
    112.7692, 111.0558, 118.8645, 131.5201, 138.3541, 150.9029, 171.4604, 
    187.6689, 173.6623, 163.331, 161.5032, 173.1302, 187.479, 196.2933, 
    205.9576, 216.4906, 204.9883, 174.7445, 149.2208, 153.461, 179.1279, 
    206.1786, 225.746, 222.5263, 174.9161, 118.1781, 104.2182, 144.9896, 
    191.7793, 237.5705, 261.6089, 430.6682, 527.5412, 452.6647, 319.951, 
    219.3656, 180.719, 164.1551, 172.7692, 202.7945, 245.6591, 251.8852, 
    209.7664, 151.3411, 111.9648, 100.5483, 102.6594, 104.9545, 115.2192, 
    135.8635, 172.4194, 187.154, 186.6964, 221.1685, 272.1998, 365.7198, 
    563.9398, 806.9812, 616.8997, 591.6264, 758.2245, 1015.611, 1321.008, 
    1507.668, 1454.292, 1383.16, 994.1575, 671.1288, 579.9672, 701.8064, 
    792.7704, 860.5122, 974.8707, 1027.509, 1188.503, 1199.935, 1087.761, 
    1020.579, 955.3137, 930.0458, 878.968, 785.0318, 671.4976, 612.8235, 
    497.7969, 458.9165, 400.6777, 383.7278, 377.0617, 422.1144, 484.0882, 
    555.1851, 690.944, 815.8306, 553.3707, 284.0944, 199.8105, 129.5959, 
    102.3608, 44.64846, 21.42765, 0.2175567, 0, 0, 0, 0, 0, 0, 0, 0, 
    116.4937, 387.2163, 621.8568, 251.8127, 11.16654, 1.124135, 0.09560291, 
    0, 0.01010601, 0.02667685, 0.01857915, 0, 0, 0.1285264, 0.2653117, 
    0.07926562, 0.001047007, 0, 0, 0, 0, 0, 0, 0.0008430172, 0.0001090577, 0, 
    0.06230972, 0.2783441, 1.301513, 2.332806, 3.847753, 0.8005066, 
    0.1766222, 0.0005744135, 0, 6.072785e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1084164, 5.786307, 9.918187, 81.89671, 
    421.8526, 869.0035, 1072.843, 1098.982, 1028.264, 934.2908, 1099.104, 
    1440.995, 1708.009, 1530.735, 1181.759, 936.9722, 790.071, 707.3079, 
    663.4688, 631.2878, 608.8522, 599.3853, 558.9546, 505.3079, 441.8009, 
    374.5419, 353.1812, 280.9854, 255.2099, 222.1815, 246.0928, 268.0079, 
    273.7544, 273.4182, 271.3401, 257.6674, 224.2582, 187.507, 152.6027, 
    124.9871, 95.54329, 56.34914, 8.645053, 0.4116594, 10.82566, 103.4201, 
    195.7967, 265.0341, 354.1939, 427.669, 486.439, 550.0139, 609.0536, 
    613.6898, 592.6232, 536.5614, 503.3919, 490.2436, 418.2097, 358.0248, 
    344.2176, 269.6707, 159.2626, 53.46779, 0.06294316, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.1002379, 0.7881545, 78.7939, 101.2808, 105.4847, 40.10086, 
    8.459635, 64.73666, 142.2411, 65.43371,
  4.919068, 0.008572195, 0, 0, 0.0002187628, 0.00431326, 6.148, 16.33585, 
    15.66748, 5.173548, 10.69731, 4.673275, 18.46478, 45.79006, 75.92396, 
    71.44189, 56.51721, 86.52747, 105.3328, 126.6551, 164.041, 181.166, 
    186.6069, 176.6074, 186.9285, 198.4358, 211.4073, 209.9819, 203.8876, 
    199.4759, 187.7478, 150.5249, 132.5192, 131.1255, 156.5745, 173.4979, 
    185.5967, 180.0389, 156.4083, 121.3786, 134.7526, 168.165, 217.4006, 
    197.5112, 198.3453, 311.4803, 531.9188, 499.1912, 342.132, 222.703, 
    165.2046, 141.3972, 143.4367, 149.5323, 149.404, 142.2128, 128.5719, 
    111.0091, 105.2806, 103.9649, 102.9193, 103.553, 110.3417, 129.583, 
    166.0531, 182.2675, 214.1717, 251.4292, 281.8083, 341.4292, 573.1824, 
    707.696, 532.2667, 497.1506, 615.3599, 831.8939, 1081.983, 1166.839, 
    980.8156, 775.3804, 565.5085, 525.0767, 592.2892, 705.9196, 777.0842, 
    791.7678, 970.9343, 1069.026, 1215.237, 1373.24, 1243.177, 1066.545, 
    975.698, 948.8546, 947.9986, 891.0973, 797.1302, 752.4106, 689.6935, 
    644.1699, 626.1002, 532.0483, 501.56, 518.7145, 664.5046, 715.5826, 
    701.2019, 568.9152, 288.5578, 133.1576, 20.68132, 16.51421, 3.367378, 
    0.7943002, 0.5845824, 0.1529268, 0, 0, 0, 0, 0, 0, 0, 0.1154558, 
    120.0936, 508.8923, 664.7625, 539.5366, 305.3639, 187.4475, 13.09079, 0, 
    0.3642445, 1.18932, 1.970586, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.153782, 2.533659, 1.764091, 1.927123, 3.139146, 1.642686, 
    2.61611, 0.7462649, 0.1985903, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.3051782, 5.45147, 12.82297, 208.9811, 718.5417, 966.3851, 
    1027.382, 995.5499, 942.6932, 921.7947, 1076.374, 1253.036, 1161.514, 
    1020.949, 888.6792, 825.8789, 706.2319, 646.436, 630.6771, 623.3245, 
    600.0434, 527.0399, 518.0312, 488.1535, 426.0578, 356.9651, 307.1834, 
    288.2178, 254.5977, 224.986, 220.6133, 218.2315, 212.5904, 205.7119, 
    195.1549, 175.6493, 150.7557, 130.4452, 115.8835, 101.3156, 91.00654, 
    43.06038, 9.543821, 1.118416, 18.94706, 120.7411, 213.5428, 285.8357, 
    349.4542, 406.6175, 465.2273, 510.2496, 552.565, 579.3892, 553.5745, 
    516.3127, 508.3579, 493.2723, 378.5906, 268.1178, 213.3669, 105.2307, 
    13.67198, 0.04563162, 0.002884715, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01308964, 
    0.08465132, 6.248717, 84.94481, 93.49541, 63.73012, 56.04049, 100.8483, 
    205.1813, 49.52119,
  0.1037096, 0, 0, 0, 0, 0.3173788, 5.081631, 37.65478, 12.67908, 12.49209, 
    31.55777, 10.09756, 12.90577, 1.015718, 0.7561651, 0.2891517, 17.88934, 
    67.70225, 75.22325, 93.72872, 129.6724, 148.4861, 150.205, 160.0022, 
    177.4912, 199.5753, 217.1373, 220.6155, 207.082, 189.2652, 162.5883, 
    142.2003, 127.5409, 124.413, 134.0152, 147.9355, 140.0433, 136.2423, 
    123.7013, 126.6482, 128.4287, 143.5078, 148.3034, 151.5911, 151.0044, 
    281.4285, 369.0809, 407.7724, 333.2746, 197.3605, 153.2443, 132.6341, 
    124.9474, 128.3281, 129.0838, 124.65, 120.2516, 114.6961, 105.0679, 
    103.9084, 106.5016, 109.9837, 115.9913, 127.0985, 140.8714, 145.0928, 
    158.9637, 180.0543, 212.8158, 260.795, 429.4057, 422.0957, 405.9527, 
    430.4442, 473.4073, 483.8292, 486.8795, 509.0421, 505.5709, 462.8823, 
    469.8702, 504.4337, 550.015, 664.2174, 737.6888, 764.5994, 847.0208, 
    1107.857, 1235.461, 1316.507, 1343.689, 1254.597, 1108.379, 1060.965, 
    1116.571, 1003.154, 864.9898, 765.1527, 769.2305, 829.1945, 796.061, 
    780.2474, 773.0483, 937.1343, 1037.196, 1111.925, 1004.564, 835.8282, 
    590.8559, 264.5349, 29.83088, 0.2726912, 0, 0.02562582, 0.04808182, 
    9.400145e-05, 0, 0, 0, 0, 0, 0, 0, 3.01363, 37.46404, 450.6561, 694.5378, 
    673.2141, 568.6823, 398.3767, 6.833825, 0.452408, 0.7848065, 0.8307315, 
    0.0872502, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006008104, 
    0.01198069, 0, 0.01239326, 0.01249807, 0.2853698, 23.23273, 146.7104, 
    87.58156, 152.6909, 3.490258, 0.3605898, 0.1024441, 0.01298359, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3504601, 7.460026, 67.67462, 251.675, 
    597.1992, 863.3519, 979.736, 1121.721, 1147.21, 1143.594, 1104.271, 
    998.4769, 935.9226, 765.0177, 682.182, 696.1772, 712.803, 684.9299, 
    622.6885, 629.6263, 601.7662, 548.705, 475.4591, 455.9382, 457.167, 
    418.3767, 373.6586, 336.3819, 312.1499, 273.731, 233.5184, 212.9149, 
    193.5791, 168.3653, 141.0569, 135.6687, 132.6844, 115.6048, 88.78099, 
    67.37737, 36.77668, 25.84525, 13.39029, 3.856152, 0.06285892, 1.190556, 
    78.06513, 198.1698, 277.3407, 338.2536, 376.6179, 427.2278, 463.383, 
    471.4552, 472.8181, 496.7475, 487.7807, 485.2014, 458.3683, 329.3343, 
    115.338, 21.35109, 2.886387, 0.512166, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.06230798, 2.719209, 7.505898, 82.74612, 213.9138, 218.9389, 
    118.0055, 21.40057,
  0, 0, 0, 0, 0, 0.03378252, 18.81201, 29.97211, 23.0547, 10.57135, 79.77882, 
    121.7605, 95.52518, 21.46502, 0.4486876, 0.0959833, 24.78417, 61.02703, 
    67.8613, 69.37209, 97.49801, 126.3562, 133.4255, 139.0697, 155.4775, 
    194.8082, 225.3066, 218.9407, 186.0535, 167.7975, 161.3444, 152.2095, 
    132.6878, 118.9827, 117.2522, 112.5718, 112.6843, 114.8091, 129.0433, 
    136.543, 140.8296, 145.4046, 141.5063, 144.2454, 187.1087, 243.6195, 
    305.897, 360.7583, 300.14, 202.7668, 135.2522, 112.797, 101.8629, 
    101.8292, 114.083, 107.9538, 104.1766, 101.1058, 97.41016, 101.5928, 
    114.0993, 120.589, 125.3507, 130.5241, 134.1557, 127.9121, 123.2517, 
    130.5993, 164.637, 182.2455, 213.0129, 233.9451, 259.553, 305.8153, 
    288.3746, 296.3653, 302.3282, 303.9196, 335.5743, 377.8776, 430.7833, 
    477.0864, 503.1766, 550.5393, 611.0358, 620.2182, 757.0104, 1041.451, 
    1151.438, 1187.371, 1197.201, 1156.392, 1099.938, 1256.038, 1406.226, 
    1340.49, 1062.711, 925.06, 951.6456, 978.8389, 980.806, 1024.956, 
    1094.22, 1063.015, 1035.187, 1027.827, 996.1818, 810.6388, 728.9537, 
    692.5972, 281.21, 17.06039, 0.4778104, 0.00291224, 0.0001943904, 
    3.102328e-05, 0, 0, 0, 0, 0, 0, 0, 0.2945038, 36.02558, 156.2673, 
    517.385, 586.1339, 457.1775, 293.554, 101.1336, 0.09928098, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.675433e-05, 0.07447594, 
    0.07733262, 0, 0, 0, 0.004361894, 0.02733142, 7.511605, 28.21364, 
    206.001, 122.4869, 4.642686, 1.843176, 36.55193, 27.35227, 0.002855681, 
    0.002366547, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.173499, 9.088313, 83.18864, 
    262.4997, 735.6247, 1027.532, 1145.21, 1248.557, 1329.559, 1373.352, 
    1345.353, 1189.152, 894.141, 751.7992, 727.2402, 688.4752, 608.1703, 
    618.981, 613.402, 590.2661, 538.4998, 498.6893, 482.7774, 473.2635, 
    484.6255, 499.4903, 442.742, 394.8707, 355.0567, 327.7505, 289.6916, 
    263.109, 230.213, 191.7849, 145.2503, 85.44183, 85.81218, 82.24927, 
    65.18149, 8.231372, 0.5482306, 0.008331239, 0, 0, 0, 0.5473455, 
    0.9744639, 2.641841, 141.3694, 221.0411, 285.196, 334.4658, 361.3416, 
    367.6213, 343.7043, 327.5902, 373.1913, 438.3948, 484.3891, 414.238, 
    209.683, 14.4057, 0.5565194, 1.689482e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.1809491, 7.94604, 85.88988, 342.8634, 257.2502, 
    80.55859, 0.9219272,
  6.990595e-05, 0, 0, 0.009281853, 1.1239, 1.35835, 7.845103, 0.9874427, 
    3.416009, 41.66479, 145.9707, 203.5287, 134.4015, 34.97104, 1.751759, 
    0.233736, 3.440017, 31.16527, 29.31215, 52.83877, 95.20691, 112.1423, 
    98.16907, 91.96889, 95.02732, 126.7443, 193.1268, 197.1006, 169.6435, 
    155.1846, 147.5441, 142.1195, 132.9599, 131.0143, 132.655, 130.4676, 
    125.7518, 128.0106, 136.0226, 143.8916, 153.8184, 163.7278, 186.7656, 
    184.4975, 195.8315, 219.3869, 288.883, 327.4375, 248.1454, 164.3483, 
    120.7269, 96.92941, 74.03613, 67.82533, 68.54214, 71.55963, 82.29095, 
    89.25205, 97.24905, 110.2552, 119.5475, 121.8304, 122.2665, 121.2867, 
    116.4663, 106.4772, 100.837, 102.4518, 135.1196, 146.8853, 160.2789, 
    173.9389, 186.945, 210.8533, 222.505, 237.3573, 282.8452, 291.3376, 
    302.9503, 327.3851, 387.0242, 415.1717, 451.4163, 472.7819, 503.7173, 
    500.5816, 478.9549, 672.6696, 811.6451, 866.2441, 921.9512, 950.8438, 
    1007.77, 1102.233, 1172.452, 1080.532, 1002.075, 925.6157, 859.1212, 
    881.7025, 967.954, 1010.343, 999.9883, 967.6564, 879.1035, 827.8918, 
    728.5366, 622.3107, 574.9156, 652.7604, 665.9392, 464.7997, 163.0975, 
    21.60582, 0, 0, 0, 0, 0, 0, 0, 0.002459203, 0, 0, 2.281191, 71.77944, 
    181.9072, 317.2759, 442.9366, 288.3585, 132.0369, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.02147744, 0.06122907, 0.003346619, 0, 
    0, 0, 0, 0, 0.02759107, 0.145356, 11.60702, 90.63374, 78.20203, 60.09513, 
    205.5446, 249.456, 86.93553, 0.03397703, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.8666349, 7.99083, 175.073, 350.6861, 842.5231, 1115.008, 1235.441, 
    1381.784, 1506.417, 1503.537, 1518.813, 1473.253, 1064.393, 814.9124, 
    703.2771, 728.2607, 599.1451, 527.5717, 523.2224, 546.0634, 525.3589, 
    491.8752, 421.4688, 487.4109, 503.3438, 508.286, 500.1369, 449.3311, 
    406.633, 376.3765, 361.4974, 307.8099, 289.7761, 253.7083, 201.0309, 
    111.7332, 42.38031, 17.57482, 10.66569, 3.342806, 0.0005948858, 0, 0, 0, 
    0, 7.807768e-07, 0.001381822, 0.0417408, 3.365059, 30.81227, 191.9259, 
    247.4304, 281.1032, 305.8344, 283.9044, 232.532, 210.0196, 241.5411, 
    423.8283, 515.58, 431.389, 143.1918, 9.261302, 0.01894015, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0560388, 0.7403216, 7.951338, 45.77325, 
    326.0547, 149.943, 40.49091, 0.02273438,
  6.285479e-06, 0, 0, 1.490214, 177.1755, 394.339, 315.3454, 118.8556, 
    17.12551, 74.21546, 134.2317, 141.9279, 114.013, 31.51116, 2.011319, 
    0.4660435, 0.07483213, 0.3289439, 7.344112, 34.49738, 62.77875, 76.89153, 
    85.68703, 76.42637, 67.38309, 83.20906, 130.7097, 159.5729, 158.5045, 
    148.4201, 147.8027, 144.8745, 144.7205, 151.8467, 155.1361, 150.4327, 
    152.1391, 147.9245, 147.6059, 159.4093, 170.8969, 207.0426, 213.514, 
    205.8838, 185.1706, 220.3727, 303.4626, 299.5644, 223.6671, 123.9137, 
    99.25799, 87.20428, 74.3191, 56.3315, 61.44574, 71.28058, 83.8583, 
    90.11916, 95.62988, 102.3417, 106.0017, 103.9473, 100.118, 94.58632, 
    87.34202, 84.32126, 86.3202, 96.16251, 117.5621, 131.9892, 144.5497, 
    151.2478, 162.5047, 196.1069, 261.776, 309.8452, 329.3697, 318.0027, 
    292.9229, 302.0037, 313.4496, 332.784, 405.2306, 456.5325, 505.3469, 
    483.7405, 456.811, 428.1185, 497.2188, 537.6924, 730.7077, 889.8257, 
    897.8648, 849.8069, 684.1327, 640.1942, 584.7154, 603.0042, 663.1209, 
    712.4156, 727.9242, 728.8314, 681.1443, 615.1197, 612.6753, 570.6259, 
    522.2361, 500.8903, 525.886, 593.348, 681.0267, 640.1781, 478.6458, 
    96.10685, 4.705627, 0.7714889, 4.021969, 0.2261302, 0.02494026, 
    0.8467315, 3.417147, 2.058573, 1.713983, 1.022477, 0.2797411, 2.18481, 
    52.22627, 164.6862, 464.1557, 321.2085, 153.0177, 3.664359, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7905962, 
    12.08585, 39.81963, 50.31289, 26.83269, 115.5742, 263.5135, 440.9554, 
    223.5525, 36.29975, 1.476148, 0.06730157, 0.003832217, 0.001505081, 0, 0, 
    0, 0, 0.8266903, 5.843782, 91.68998, 551.5381, 561.364, 914.154, 
    1053.676, 1162.834, 1261.185, 1318.149, 1363.154, 1395.952, 1447.754, 
    1075.267, 841.7789, 542.7595, 551.5369, 526.2366, 442.997, 462.1343, 
    483.5762, 489.9306, 371.7027, 309.8163, 285.908, 365.5909, 422.7384, 
    428.3295, 420.3303, 416.6738, 408.2287, 391.545, 371.3323, 309.914, 
    283.9654, 236.5979, 151.896, 53.84359, 18.70917, 0.6324576, 0.01533817, 
    5.997697e-05, 0, 0, 0, 0, 0, 0.003037961, 0.007704118, 2.666646, 
    40.34323, 108.7473, 162.0983, 213.3329, 236.9303, 239.9766, 210.3202, 
    149.2632, 93.44909, 158.2182, 321.6055, 486.9341, 261.5333, 43.32835, 
    0.3786546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001964956, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.04539995, 0.3973858, 1.861022, 4.39137, 75.7228, 27.85487, 2.136931, 
    0.001607413,
  0.000485088, 0, 0, 15.60826, 109.6726, 828.3698, 696.0719, 489.5445, 
    150.7604, 166.8067, 167.8064, 152.9492, 130.6891, 51.74954, 16.34865, 
    2.361931, 0.2884878, 1.639599, 6.479568, 31.35585, 55.31397, 44.66693, 
    27.78062, 54.56249, 57.35855, 59.07015, 86.24779, 133.3726, 160.1804, 
    154.7875, 147.3788, 150.7191, 156.2221, 165.9632, 168.4068, 180.8379, 
    171.8393, 174.2765, 175.3024, 174.642, 181.7714, 188.4763, 201.4641, 
    185.6017, 176.3486, 227.5092, 328.7459, 366.1854, 171.3452, 111.5206, 
    82.99934, 74.11316, 65.81149, 54.21898, 49.75399, 60.85712, 72.62536, 
    82.83826, 85.45224, 87.27561, 89.44934, 86.80495, 79.92211, 70.88648, 
    75.55956, 87.62287, 101.455, 125.0653, 134.2894, 139.1541, 140.6684, 
    141.3033, 193.3456, 276.3874, 410.5264, 425.0551, 426.7878, 392.8753, 
    355.5762, 326.4843, 313.2398, 330.9117, 362.6911, 432.2075, 445.5331, 
    443.6434, 425.0182, 417.2193, 404.0916, 441.2396, 509.8215, 681.8781, 
    802.3056, 610.0692, 464.1464, 393.0627, 402.3937, 451.2505, 502.0411, 
    515.427, 521.9349, 522.9614, 472.5158, 397.127, 339.8048, 332.6423, 
    366.4758, 381.1311, 467.7882, 603.1166, 699.1341, 694.8555, 551.1594, 
    382.6274, 206.6408, 215.4341, 141.7952, 169.5575, 169.1414, 158.2998, 
    192.459, 202.4881, 242.4227, 35.21797, 9.042901, 0, 0, 13.23063, 
    61.15136, 393.7112, 144.1485, 11.97594, 2.622757, 1.13881, 0.6200418, 
    0.3004147, 1.810146, 0.7663906, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.002402687, 0.02916033, 0, 0, 0.03871302, 0.1174289, 0.2317475, 
    0.8005022, 3.538009, 123.0752, 227.675, 201.7235, 175.1833, 125.1719, 
    250.8978, 295.6898, 207.6078, 28.8371, 52.37325, 9.258338, 6.067081, 
    1.74902, 6.066913, 20.01941, 20.3201, 69.3385, 63.36699, 399.117, 
    906.2566, 1070.019, 1160.485, 1098.04, 1113.135, 1179.21, 1215.758, 
    1108.652, 1042.706, 990.644, 947.2479, 758.5189, 504.7683, 501.6226, 
    514.3629, 502.3148, 472.9703, 451.7628, 482.619, 408.9817, 307.0132, 
    238.6153, 277.3391, 318.1176, 388.6982, 399.9906, 405.2738, 407.2638, 
    408.4838, 390.1241, 363.4594, 305.5353, 270.8763, 222.3424, 108.2813, 
    29.74055, 2.095462, 0.007033782, 0, 0, 0, 0, 0, 0, 0, 0.02696288, 
    0.05046848, 0.01513994, 33.80931, 76.48997, 151.0632, 193.2209, 221.7352, 
    219.6982, 186.103, 65.00166, 6.271983, 3.192534, 182.7761, 342.0524, 
    61.69406, 4.945493, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.94174e-05, 0.2316896, 
    0.2696269, 16.19537, 11.6254, 0.4879676, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.214889e-05, 0.02950715, 
    0.1218954, 1.484969, 0.9002973, 0.3741933, 0.06643537,
  0.002089362, 0, 1.412099, 26.46473, 490.6368, 888.3039, 1135.971, 709.175, 
    534.5035, 355.5736, 330.3836, 309.3834, 197.7856, 113.4243, 8.748651, 
    2.184844, 2.557522, 32.08658, 53.47832, 61.61737, 61.77125, 30.52585, 
    42.68884, 35.54211, 26.26413, 10.52586, 57.40441, 134.2131, 156.6786, 
    156.7883, 158.2699, 158.8308, 164.9652, 157.9505, 155.4321, 153.5848, 
    156.4442, 153.1837, 155.5327, 164.734, 173.5995, 182.6821, 178.5456, 
    169.5983, 165.4698, 210.9651, 348.5778, 322.2212, 227.3903, 99.48459, 
    80.63308, 73.28908, 68.85529, 55.97015, 44.73322, 53.9101, 58.34581, 
    62.13969, 62.22141, 63.91478, 65.12193, 63.32931, 63.88552, 63.9667, 
    85.60952, 97.93639, 110.2092, 130.7943, 137.0216, 141.3263, 137.5219, 
    168.7466, 213.6295, 354.2611, 402.6772, 428.3887, 433.8965, 420.1635, 
    409.1618, 367.8534, 360.9081, 351.4519, 375.3124, 390.8479, 389.126, 
    375.8873, 360.2204, 385.7919, 404.6116, 404.389, 412.3467, 400.9159, 
    385.2873, 391.0082, 350.8959, 340.8138, 352.6799, 404.1559, 426.472, 
    438.9901, 434.1502, 424.6885, 416.6674, 340.0075, 309.9525, 294.1677, 
    282.8733, 285.1135, 384.4936, 671.5599, 823.5674, 925.6255, 852.2806, 
    742.6212, 721.0127, 693.4877, 669.465, 620.8027, 634.554, 664.8117, 
    693.1401, 808.8724, 739.8962, 581.1383, 376.3603, 154.5647, 0.6796251, 
    4.982354, 64.11263, 142.5318, 108.1566, 149.5249, 204.1944, 211.7184, 
    208.7517, 208.467, 288.7601, 140.705, 4.269242, 9.153877e-05, 0, 0, 0, 0, 
    0, 0, 0, 0.005518374, 0.1355343, 0.2826844, 0.3221478, 0.01058123, 0, 
    0.001992178, 0.4520722, 0.9488499, 6.779386, 16.57067, 40.10801, 
    255.6327, 344.4668, 265.1516, 232.6011, 400.0099, 586.2018, 695.2791, 
    563.507, 464.1432, 361.5622, 113.9375, 323.1818, 506.1862, 547.4941, 
    894.0842, 1285.52, 1484.35, 1735.863, 1358.374, 1231.392, 1152.969, 
    1131.283, 1152.331, 1170.065, 1158.371, 1089.12, 1003.844, 1009.017, 
    954.9542, 729.5635, 589.0408, 496.241, 444.6862, 450.0207, 394.0024, 
    345.4459, 307.3172, 243.5889, 229.6464, 215.4986, 325.458, 376.5272, 
    435.0629, 457.4943, 440.2969, 414.7746, 388.1772, 372.1166, 354.8122, 
    301.541, 254.2812, 204.0881, 88.55573, 36.70787, 0.3222319, 0.002726495, 
    0, 0, 0, 0, 0, 0, 0, 0.004336663, 0.04531058, 1.227226, 7.522099, 
    100.8121, 187.4572, 296.865, 329.1426, 274.8387, 133.0592, 47.23021, 
    1.316583, 0.9129715, 1.553727, 7.258464, 1.342638, 0.201636, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3.251589, 23.10911, 98.81904, 503.6058, 517.3815, 
    327.3233, 30.79667, 0.3835053, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006569692, 0.2195214, 
    1.876615, 0.6393616,
  0, 0, 1.828225, 19.26351, 448.8344, 835.2745, 1141.588, 1032.039, 786.5547, 
    654.9902, 588.2164, 412.7137, 308.6151, 68.38618, 12.06376, 0.06471667, 
    18.41938, 61.81321, 104.4949, 125.8387, 118.5854, 108.4666, 84.79565, 
    76.40121, 59.19922, 78.75513, 98.56306, 115.2247, 134.3331, 145.9909, 
    151.77, 151.7498, 152.8904, 142.5491, 136.7288, 135.7318, 128.0627, 
    140.0998, 143.6488, 146.3888, 149.8231, 156.6393, 161.7421, 162.2298, 
    164.8261, 217.8509, 291.1935, 348.3962, 195.8417, 129.083, 114.5032, 
    105.5355, 95.45203, 61.35595, 54.60228, 55.04914, 56.48923, 55.82372, 
    54.56919, 55.73862, 57.38455, 68.16464, 69.42513, 70.68404, 84.55488, 
    95.45844, 107.8621, 133.5746, 139.8783, 145.4366, 147.4661, 171.0951, 
    226.8824, 321.1786, 370.2545, 437.2687, 446.555, 451.0341, 429.5266, 
    412.8637, 391.1489, 395.1011, 408.7996, 399.6818, 382.3647, 346.0877, 
    339.6265, 341.1089, 371.4463, 382.2886, 372.0459, 353.894, 321.5528, 
    286.9143, 272.5866, 281.252, 310.7381, 334.1094, 351.0113, 327.032, 
    311.4084, 304.4399, 280.9602, 265.0073, 236.722, 243.8755, 241.4891, 
    261.6405, 407.1862, 663.1442, 1011.532, 1167.707, 1236.869, 1285.631, 
    1263.503, 1149.885, 1082.739, 1000.507, 916.3446, 896.2212, 843.7785, 
    853.3328, 777.1346, 774.0334, 728.1268, 439.2752, 263.6532, 163.5337, 
    222.7859, 251.3487, 95.91259, 169.9095, 229.9653, 309.1035, 429.4353, 
    532.8344, 671.1013, 520.1642, 353.9319, 37.26283, 15.31902, 1.765467, 
    0.6663253, 0.1177541, 0, 0, 0, 0, 0.01669307, 0.002175942, 0, 0, 0, 
    0.02214206, 0.1799842, 4.561895, 12.91159, 25.73379, 40.63332, 75.03893, 
    217.1985, 213.8127, 237.9688, 365.2299, 780.1066, 906.6393, 712.6368, 
    606.8312, 747.8552, 970.0857, 998.6761, 1011.284, 1095.941, 1398.026, 
    1817.498, 1761.355, 1421.368, 1276.808, 1116.542, 1089.972, 1107.633, 
    1178.089, 1242.351, 1232.495, 1234.801, 1316.746, 1304.597, 1103.827, 
    904.4067, 460.6985, 392.8093, 328.2285, 316.8165, 286.4761, 197.7343, 
    183.4523, 169.3739, 182.7746, 222.6871, 324.1719, 385.2672, 415.2478, 
    424.0601, 403.8041, 389.3885, 355.7688, 340.3573, 326.4505, 285.5766, 
    241.9037, 192.1936, 90.21161, 52.75986, 7.89742, 2.043197, 0.009632749, 
    0, 0, 0, 0, 0, 0.08570033, 0.08687565, 0.2519769, 2.217057, 72.71382, 
    169.2529, 317.6039, 368.3998, 408.8689, 227.5118, 18.7586, 3.276534, 
    2.33082, 47.43875, 4.772794, 2.553824, 0.1766333, 0.004686403, 0, 0, 0, 
    0, 0, 0, 0, 0.1143011, 15.10792, 57.493, 503.3056, 1195.094, 1424.029, 
    1637.78, 1029.436, 99.19889, 11.66397, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7659043, 1.689617, 0.1253343, 
    0, 0, 0.06345863, 0.04394071,
  0, 0, 0, 9.18603, 67.33627, 652.2083, 698.2867, 903.2977, 791.1568, 
    821.2966, 652.2013, 535.5381, 325.3865, 216.1812, 18.25854, 6.78636, 
    2.77748, 53.08744, 124.7553, 139.4932, 148.5916, 135.4449, 125.3183, 
    126.9657, 142.3426, 157.2012, 142.0184, 128.6603, 129.407, 134.6527, 
    141.8521, 132.4218, 110.4533, 104.7861, 106.7858, 107.0216, 136.0108, 
    159.6768, 163.2655, 156.4141, 148.5422, 147.0514, 161.0536, 162.2215, 
    161.4925, 182.1215, 275.0815, 265.3517, 173.3195, 98.77954, 81.69308, 
    73.50078, 83.55206, 85.846, 84.78377, 83.22816, 86.88531, 83.45903, 
    80.20251, 81.64954, 82.38533, 86.15968, 91.05025, 94.42326, 120.4377, 
    123.6299, 127.9127, 133.1319, 131.3258, 120.3571, 145.1299, 176.2902, 
    285.127, 348.2451, 446.7507, 466.7538, 466.9656, 457.1467, 440.4509, 
    410.6824, 399.9454, 398.3544, 402.3503, 388.5353, 354.7975, 332.7445, 
    323.295, 330.8784, 332.9599, 340.5439, 340.3431, 316.3052, 250.7962, 
    216.2447, 207.9207, 236.2964, 270.3356, 271.1327, 281.8501, 263.7443, 
    246.2528, 235.041, 189.72, 183.1059, 165.6444, 180.943, 195.0492, 
    184.0648, 349.6989, 553.5489, 972.6125, 1291.18, 1421.197, 1497.029, 
    1237.482, 1217.527, 1138.105, 1061.736, 923.1717, 818.9904, 704.847, 
    599.6451, 557.6539, 670.0704, 719.3553, 722.7904, 670.9245, 582.5764, 
    406.9142, 346.8488, 278.6282, 256.195, 239.0234, 211.3936, 382.6976, 
    500.9314, 720.5585, 609.0164, 448.009, 298.562, 220.2226, 54.00721, 
    32.91389, 3.113513, 0.4547248, 0, 0, 0, 0, 0.03715197, 0.1058386, 
    0.1689842, 0.1235006, 0.007738656, 0.1990487, 2.824826, 32.01704, 
    59.08257, 126.8133, 146.7751, 141.567, 188.4334, 251.0966, 342.7206, 
    454.9237, 611.2901, 909.9222, 996.2937, 1010.439, 1039.88, 1024.344, 
    1035.421, 1225.468, 1282.719, 1047.796, 937.444, 921.0512, 949.0565, 
    946.207, 901.6165, 1020.892, 1128.21, 1188.953, 1223.496, 1412.944, 
    1507.547, 1400.053, 1244.998, 638.0379, 473.8077, 316.8543, 316.7606, 
    324.2363, 285.3842, 260.8806, 207.7252, 220.4391, 248.7498, 307.9653, 
    340.2007, 381.2327, 386.924, 393.2863, 356.0091, 342.5364, 320.4373, 
    299.2019, 284.6974, 247.4959, 212.9148, 161.3572, 109.587, 86.55267, 
    44.18631, 20.04325, 1.685035, 0.2694115, 0.001934427, 0.009342462, 
    0.01149242, 0.1277481, 1.344178, 0.9477215, 0.06420656, 2.531306, 
    13.23086, 225.1991, 230.0539, 190.0253, 96.81186, 21.50346, 82.57745, 
    238.3149, 352.9399, 368.0467, 194.4866, 11.7522, 2.031744, 0.001181567, 
    0, 0, 0, 0, 0, 0, 0.06388535, 5.58617, 128.1033, 912.9094, 1518.721, 
    2110.982, 2481.025, 2132.609, 1414.114, 484.4178, 30.76768, 1.54477, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005166661, 0.3623523, 2.201925, 
    1.430301, 0.8634878, 0.07886008, 0, 0, 0, 0, 0, 2.467292, 6.077, 
    1.148987, 0, 0, 0, 0,
  0, 0, 0, 0.4990054, 0.4105075, 16.4118, 30.50377, 319.1797, 399.7182, 
    576.643, 592.1636, 459.3603, 398.4318, 284.2472, 209.5148, 57.34949, 
    70.75203, 17.37498, 43.04565, 121.5067, 130.4336, 140.5459, 156.2209, 
    173.6517, 185.9281, 180.9441, 153.4432, 127.9112, 119.9615, 132.0899, 
    116.8609, 88.48421, 79.63129, 75.38411, 85.86076, 111.0442, 135.5131, 
    154.0528, 162.3629, 174.6046, 170.0756, 168.9717, 166.2372, 149.558, 
    155.8482, 194.058, 233.2592, 279.8633, 206.2282, 90.39473, 61.77412, 
    51.8238, 55.83362, 66.18795, 85.0791, 94.89624, 104.686, 99.4508, 
    98.42764, 96.52757, 90.28058, 77.16055, 76.74628, 76.66355, 101.0403, 
    100.3977, 100.0436, 97.41985, 95.20831, 73.1783, 124.6243, 258.6244, 
    337.6291, 382.1798, 424.1999, 415.7608, 422.9675, 432.1186, 449.5258, 
    434.0693, 429.2796, 419.7672, 413.4257, 376.6487, 376.8708, 347.6423, 
    347.3596, 353.7901, 368.4431, 367.3064, 356.8146, 304.6212, 264.2978, 
    198.3714, 183.5134, 178.0944, 171.1256, 193.8708, 169.418, 171.4767, 
    160.59, 153.83, 271.3834, 214.4951, 322.3955, 409.8011, 364.5263, 
    605.6127, 555.0153, 802.5508, 1014.164, 1203.025, 1288.973, 1081.302, 
    1032.944, 1146.767, 1159.82, 1169.949, 1054.652, 761.6836, 619.8669, 
    486.295, 477.4393, 482.5888, 600.5913, 668.1846, 809.5635, 764.5266, 
    663.7883, 625.8642, 597.3387, 499.2648, 433.516, 312.4686, 262.843, 
    240.825, 322.2652, 327.7585, 338.623, 306.9521, 283.5958, 176.864, 
    110.5663, 4.941168, 1.403517, 0, 0, 0, 0.1360559, 1.096909, 0.3120382, 
    0.2519662, 0.1819621, 0.01765274, 0.2073749, 0.5467369, 9.687221, 
    18.14567, 54.46339, 180.5516, 173.0188, 148.8622, 184.7714, 267.147, 
    312.3334, 392.5854, 463.3264, 807.8792, 960.6965, 905.6902, 1072.808, 
    1026.749, 916.2828, 867.8626, 852.2236, 802.7931, 840.2682, 856.4594, 
    848.0734, 980.8599, 1014.717, 1127.941, 1205.185, 1440.98, 1520.958, 
    1438.045, 1351.211, 752.0334, 580.1899, 411.7906, 366.1327, 327.8392, 
    321.8054, 293.748, 268.8281, 248.8851, 332.558, 350.3996, 410.0892, 
    404.3516, 400.5793, 391.6209, 387.9602, 327.0846, 314.2092, 295.0971, 
    273.101, 262.0161, 220.7047, 193.3422, 139.1538, 114.4612, 100.9127, 
    71.0108, 57.66841, 31.5654, 19.15824, 4.611352, 19.68997, 23.90316, 
    12.82197, 30.50539, 22.5677, 17.31053, 0.3391515, 3.474163, 10.88561, 
    9.502873, 2.376641, 11.08148, 81.42273, 282.0594, 355.9471, 449.2821, 
    441.8114, 267.1641, 72.81113, 5.423061, 0.01384602, 0, 0, 0, 0, 0, 0, 
    2.228677, 112.5068, 656.6617, 1131.168, 1937.853, 2362.118, 2597.015, 
    2500.656, 1824.832, 1167.206, 138.9148, 18.45758, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2.598965, 12.72333, 110.1043, 185.5357, 246.7095, 218.1962, 
    159.5719, 78.65945, 0.2450386, 0.06335586, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.006711138, 0.4642611, 15.49415, 210.3725, 274.8661, 
    556.0378, 584.5959, 461.9076, 436.8904, 341.9686, 289.6991, 113.7131, 
    33.07074, 5.939446, 15.70688, 91.06759, 133.7827, 175.9086, 195.419, 
    196.4113, 167.8823, 119.3239, 82.73615, 47.22521, 35.94244, 65.74197, 
    67.93156, 58.86282, 64.24126, 70.37502, 82.21825, 104.7593, 128.4086, 
    158.7193, 172.8007, 197.0037, 198.6317, 132.9266, 124.7694, 128.5104, 
    156.0846, 300.5825, 341.3086, 327.2441, 225.6438, 111.7088, 69.47119, 
    36.01659, 49.88657, 61.31368, 75.10065, 82.15571, 73.43854, 74.03111, 
    72.68026, 63.95351, 53.51602, 43.87702, 40.58201, 52.25, 60.52992, 
    84.52159, 83.98617, 83.63194, 95.8566, 112.0164, 342.0878, 367.5606, 
    395.9712, 392.8885, 384.3166, 427.4104, 471.1263, 494.9181, 495.573, 
    464.0248, 458.752, 470.0241, 478.5758, 459.2749, 466.4923, 450.6083, 
    453.846, 436.6663, 439.5466, 395.4367, 360.7103, 279.4871, 227.9757, 
    198.8707, 179.1181, 172.8613, 154.538, 141.8269, 126.4755, 238.588, 
    407.1594, 553.9539, 851.4879, 899.8338, 872.8414, 1098.375, 947.5765, 
    915.9656, 961.4484, 1078.228, 1140.825, 1126.576, 1077.586, 1102.926, 
    1144.051, 1237.868, 1230.951, 878.9684, 738.7202, 345.855, 349.7968, 
    337.6898, 359.5725, 405.3323, 514.2386, 611.831, 627.7592, 647.9431, 
    731.343, 719.1741, 661.5468, 605.7673, 551.1049, 371.3813, 309.8194, 
    152.4344, 158.0018, 171.2113, 150.7313, 131.6786, 72.96445, 59.19989, 
    7.159949, 3.730352, 0, 1.61262, 4.895032, 13.13506, 39.44074, 25.06428, 
    0.2390079, 0.1075483, 0.286315, 11.65734, 48.24539, 97.97038, 138.7014, 
    68.57406, 113.1445, 193.342, 195.0805, 210.8494, 234.041, 271.1232, 
    272.3607, 301.2755, 262.5467, 362.0172, 561.8752, 574.761, 677.5664, 
    802.9904, 834.3304, 864.3197, 906.5961, 921.4742, 1009.76, 1183.24, 
    1094.674, 1135.249, 1228.71, 1386.295, 1405.771, 1272.237, 1251.558, 
    696.1383, 536.7278, 360.8228, 337.9231, 303.7456, 307.6464, 323.558, 
    324.3554, 311.1708, 345.7896, 397.8962, 419.6172, 440.2093, 442.2453, 
    435.8681, 391.2493, 372.918, 321.2558, 279.2823, 234.0026, 210.5916, 
    202.4526, 162.4054, 151.3109, 120.1705, 116.4772, 117.6743, 133.9828, 
    147.2711, 151.5799, 148.9824, 85.92712, 95.84363, 96.8592, 168.0968, 
    183.4117, 67.15431, 34.58618, 2.304035, 13.49032, 111.5204, 88.934, 
    48.49368, 87.72391, 195.7094, 247.2929, 375.258, 435.4196, 500.3941, 
    336.9578, 29.66164, 2.046304, 0.4911519, 0.0429709, 0, 0, 0, 0, 1.055858, 
    14.98069, 146.1425, 609.2309, 1146.736, 1832.361, 2328.555, 2519.978, 
    2538.643, 2305.819, 1302.339, 570.7617, 38.91841, 0.8063998, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.4486028, 1.00745, 120.6145, 171.389, 424.6237, 511.5233, 
    813.5204, 800.3188, 730.7539, 381.4832, 4.793127, 1.075142, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 1.347272e-07, 0.0001361489, 37.51786, 175.727, 284.4844, 
    694.9128, 708.0693, 520.4041, 465.8637, 316.0654, 233.6545, 62.24868, 
    9.48611, 29.91223, 76.69086, 151.5849, 207.9153, 219.8867, 187.6858, 
    149.7711, 99.36585, 25.97108, 6.33916, 6.367791, 1.163611, 16.67007, 
    47.54528, 63.75716, 56.35788, 56.74799, 67.11382, 86.57465, 116.4754, 
    148.0896, 153.6746, 113.4161, 106.4274, 97.36552, 95.56422, 101.2792, 
    139.6314, 275.5676, 351.634, 262.3784, 225.8972, 82.46924, 54.58767, 
    36.34371, 39.45193, 45.44073, 45.95538, 43.69976, 49.66986, 53.45878, 
    52.55042, 51.74163, 39.70052, 37.15316, 33.45551, 38.14437, 59.3439, 
    61.84409, 67.27757, 99.1234, 133.6192, 295.1877, 372.2892, 414.1317, 
    432.824, 499.0305, 532.5197, 588.6198, 590.1069, 526.7081, 515.1794, 
    518.9926, 532.0958, 540.3781, 526.0691, 520.2847, 525.6962, 516.3216, 
    512.2423, 479.6503, 462.7082, 384.529, 332.7986, 289.3895, 233.8969, 
    217.3762, 194.1487, 174.2845, 136.5615, 167.7772, 276.2465, 633.751, 
    976.7137, 1004.534, 973.0449, 923.1946, 804.5515, 799.7959, 878.4363, 
    933.6313, 1050.739, 1225.329, 1229.779, 1112.806, 1069.981, 1011.641, 
    1088.693, 939.9855, 854.4355, 338.7952, 229.8596, 249.6738, 280.5648, 
    367.5424, 381.9058, 426.1577, 440.5712, 455.7285, 527.3271, 668.6664, 
    710.9661, 751.7974, 710.6614, 684.816, 497.2051, 453.7836, 208.265, 
    198.7328, 137.993, 141.5616, 149.3726, 154.0697, 159.0402, 114.372, 
    99.60052, 127.5794, 154.1215, 183.9193, 202.1122, 199.4518, 175.3651, 
    13.74603, 4.271924, 4.655563, 38.85456, 160.4745, 159.278, 198.0601, 
    208.3912, 226.4971, 209.4362, 181.2745, 179.0735, 237.8724, 286.9208, 
    305.2715, 322.5107, 334.449, 356.3649, 375.376, 401.2977, 465.7788, 
    505.5878, 608.4302, 723.4133, 775.6861, 863.5701, 917.6834, 769.8234, 
    809.4301, 843.2911, 817.2551, 840.1667, 671.4922, 711.0405, 381.4118, 
    361.3168, 307.768, 251.3904, 185.3133, 183.5058, 213.0909, 246.8515, 
    299.9273, 311.6287, 414.7622, 427.8901, 464.3052, 466.2618, 476.9598, 
    443.5532, 386.5794, 341.7771, 296.8773, 255.8785, 233.7073, 208.091, 
    202.9507, 166.4952, 163.3595, 149.9456, 173.0595, 224.1687, 250.5235, 
    276.8417, 280.893, 283.1165, 174.1232, 145.2362, 101.971, 89.04053, 
    12.18463, 3.210024, 0.04258642, 0.5493788, 1.318359, 10.33986, 39.29594, 
    40.1795, 87.56113, 112.4894, 214.6106, 223.2263, 195.1201, 64.40204, 
    162.8817, 323.6455, 362.2034, 58.3152, 0.6101816, 0, 0, 0, 0, 99.52487, 
    405.8163, 579.289, 792.6241, 1344.384, 1746.299, 2120.452, 2370.221, 
    2426.624, 2226.688, 1874.045, 898.3805, 324.2918, 66.64768, 44.92525, 
    32.82828, 14.68513, 0.7619895, 0, 0, 0, 0, 0.08936542, 2.159183, 
    35.51629, 287.9611, 269.1317, 315.2691, 439.2047, 639.2167, 577.2025, 
    495.0344, 187.6143, 13.4638, 2.529191, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.002259135, 0.01595649, 105.2375, 416.09, 442.685, 
    767.1923, 771.5544, 543.311, 478.036, 293.0749, 211.3671, 159.5722, 
    123.008, 154.7472, 204.7672, 236.2515, 242.6722, 216.8267, 181.006, 
    126.3164, 104.4388, 79.56461, 74.01538, 143.5681, 127.7467, 64.73118, 
    9.851611, 17.18855, 28.9307, 41.56158, 63.17545, 90.73561, 107.0801, 
    107.9633, 102.7107, 82.67222, 85.89304, 95.33595, 93.48545, 108.5007, 
    137.0855, 160.7206, 174.0978, 193.6842, 196.0486, 156.7319, 125.8291, 
    58.17311, 34.16951, 27.3774, 25.29839, 40.88158, 46.35728, 47.01036, 
    47.81719, 36.20993, 35.09203, 31.48751, 32.81653, 47.93762, 50.72215, 
    63.30566, 90.21721, 181.3236, 248.4462, 385.9447, 438.3613, 553.597, 
    595.6282, 654.1422, 660.9266, 656.1749, 617.4047, 505.4219, 503.6128, 
    506.8136, 492.4366, 488.7919, 481.8042, 515.6224, 513.8269, 476.1539, 
    447.0326, 400.5003, 379.7177, 349.5628, 311.4319, 295.8653, 252.5856, 
    204.662, 174.4188, 136.6998, 222.3898, 406.6851, 707.4203, 937.2181, 
    984.2191, 807.518, 544.1436, 539.5954, 573.7524, 673.0231, 740.77, 
    914.4822, 1037.061, 996.9357, 957.6771, 747.974, 724.6053, 590.9419, 
    602.5323, 346.9653, 206.6231, 147.7196, 141.8199, 212.5911, 278.7321, 
    289.5333, 300.0507, 314.9635, 327.5019, 381.8064, 431.429, 499.5403, 
    530.7937, 618.2186, 628.9042, 618.3481, 614.7897, 476.62, 461.5242, 
    300.1651, 312.3365, 365.5695, 375.0411, 390.6438, 373.2717, 293.0935, 
    289.5076, 238.1081, 217.5476, 160.9597, 155.2435, 146.0707, 59.21703, 
    2.262186, 1.335201, 1.552167, 26.59651, 73.97087, 62.77603, 86.91489, 
    99.57547, 184.4053, 208.4254, 233.6914, 277.5439, 406.2749, 378.8096, 
    340.575, 450.9275, 441.0685, 430.9128, 380.654, 236.7385, 257.6009, 
    393.0115, 473.8694, 576.2799, 620.2967, 510.6674, 514.9241, 445.6316, 
    365.553, 285.0936, 193.4123, 228.264, 156.0837, 180.1685, 271.13, 
    279.7873, 304.1648, 306.4915, 277.1075, 251.3765, 284.0485, 308.1748, 
    364.0248, 425.8113, 458.0905, 474.9592, 451.0251, 448.5496, 358.8801, 
    328.0173, 268.541, 249.7715, 206.5758, 199.6689, 162.8162, 160.0171, 
    130.4523, 129.2327, 122.2571, 144.7552, 268.3323, 279.6682, 329.1225, 
    325.6839, 321.4922, 267.2283, 166.4881, 157.6386, 150.7869, 108.0233, 
    3.595343, 3.821032, 0.01575174, 0.07150077, 0.01421785, 0.8260033, 
    3.974015, 15.74647, 56.65681, 79.79868, 198.6406, 337.2138, 505.0964, 
    700.6447, 716.2372, 625.3304, 548.1509, 140.4764, 0, 0, 0.05033042, 
    0.4008242, 222.7403, 578.9071, 663.5074, 827.0086, 1187.04, 1605.778, 
    1871.908, 2231.532, 2362.803, 2384.707, 2175.984, 1976.378, 1731.382, 
    1507.728, 1216.511, 796.019, 342.3664, 56.85593, 4.048094, 0, 0, 0, 0, 
    0.003348448, 15.89278, 63.10171, 66.52153, 53.53075, 144.2148, 222.9382, 
    200.7522, 195.5594, 40.97123, 0.3134854, 0.03178433, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.3656524, 1.127182, 23.69072, 52.15788, 199.0073, 
    766.5958, 829.2528, 598.1196, 492.7027, 370.3959, 254.2298, 246.5821, 
    232.486, 243.9458, 269.9175, 273.8295, 255.3689, 228.7763, 225.1672, 
    216.461, 213.9356, 219.078, 213.3036, 205.7209, 181.8624, 65.29639, 
    1.183293, 1.838517, 2.839956, 17.69183, 40.47035, 71.1405, 78.3233, 
    56.54005, 59.72765, 80.44005, 99.22546, 109.3633, 109.3479, 103.3906, 
    108.2728, 128.0868, 172.8262, 207.3248, 306.6412, 253.9211, 70.71107, 
    59.91978, 26.77586, 24.5469, 24.31629, 27.07642, 31.32004, 31.52451, 
    28.17364, 28.07833, 38.65579, 39.05622, 60.66639, 61.49097, 83.99942, 
    89.35865, 238.791, 256.9483, 465.0884, 505.7355, 693.5392, 744.2326, 
    753.9547, 765.2906, 717.2798, 656.6039, 516.7385, 364.3393, 367.0169, 
    401.8732, 388.4323, 379.1184, 352.6762, 349.6031, 343.3075, 341.0069, 
    340.8878, 326.6531, 309.365, 288.933, 268.9826, 271.733, 235.8535, 
    167.6273, 131.0547, 204.8647, 500.2416, 782.6526, 930.733, 879.1979, 
    711.9934, 508.3092, 387.061, 372.2128, 395.7212, 481.8896, 709.8532, 
    776.7864, 676.0043, 453.798, 459.4369, 266.1626, 236.5406, 232.8728, 
    207.8306, 147.7249, 76.80683, 69.03156, 77.53581, 87.02776, 114.8945, 
    140.2177, 182.6259, 192.1268, 189.0047, 205.5229, 293.0704, 307.8033, 
    567.8621, 574.3477, 634.1666, 637.0754, 479.2057, 475.036, 448.7006, 
    455.1898, 613.9545, 634.6318, 634.5217, 638.7372, 350.4454, 297.3259, 
    126.7011, 75.49828, 14.90806, 2.061996, 2.343309, 1.962267, 0.3435362, 0, 
    0.1002045, 31.6623, 79.22138, 169.8461, 246.501, 285.096, 339.5764, 
    421.0346, 639.3541, 737.2427, 699.7647, 803.9453, 812.3242, 767.8734, 
    861.3438, 797.1647, 642.563, 631.2531, 530.3723, 409.9285, 469.0479, 
    513.139, 503.0063, 520.9756, 494.7627, 379.593, 175.7493, 126.0577, 
    164.158, 200.3353, 210.7177, 233.7815, 251.5634, 289.9112, 310.6765, 
    386.4908, 403.5676, 409.3076, 421.9493, 353.82, 323.1745, 329.6454, 
    312.8285, 293.1825, 144.1744, 175.2397, 126.8912, 143.4108, 140.2193, 
    142.4148, 90.33322, 92.78184, 63.48882, 63.97128, 49.74289, 49.01741, 
    42.16023, 43.36867, 188.3387, 189.5222, 264.3434, 260.4239, 250.3447, 
    236.8311, 229.5279, 245.1393, 255.3059, 251.0064, 81.69176, 5.208412, 
    1.30707, 0.4630101, 0.429015, 1.930142, 5.58512, 63.26179, 108.4616, 
    228.3357, 316.8307, 482.1983, 759.7762, 837.28, 626.9067, 354.7968, 
    65.11899, 0.1608328, 0, 0, 0.03733866, 0.5234969, 164.6818, 357.1854, 
    399.8932, 635.7303, 932.9971, 1411.621, 1836.409, 2074.039, 2328.994, 
    2397.195, 2477.567, 2421.971, 2461.883, 2530.302, 2348.885, 2006.908, 
    1744.191, 616.3108, 61.99642, 36.09983, 20.63045, 12.69927, 6.687611, 
    1.666052, 0.2396921, 0.6683463, 0.05483739, 7.549096e-06, 0.00189263, 
    0.002261056, 8.443099e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.007547835, 1.226913, 2.148309, 16.50055, 
    39.61559, 136.2474, 617.611, 707.5878, 582.7769, 480.6999, 446.4436, 
    351.2215, 311.8399, 282.2197, 239.4662, 220.2822, 222.3295, 206.7987, 
    189.6968, 202.2691, 212.9107, 210.6333, 196.719, 108.0036, 11.58493, 
    0.07383566, 0.3977811, 1.037106, 0.9561975, 0.6481953, 0.8595715, 
    1.186568, 3.491535, 13.9642, 24.33522, 34.10968, 51.74074, 65.73071, 
    61.4578, 54.07482, 75.10642, 121.9366, 126.3054, 153.6963, 177.8387, 
    80.79975, 27.65865, 33.24729, 27.32014, 20.027, 5.261846, 9.860478, 
    25.9965, 27.0378, 34.50664, 34.38958, 51.90482, 51.88333, 62.17891, 
    62.975, 97.73689, 109.6041, 232.0181, 303.3775, 485.8334, 696.6212, 
    782.4447, 933.1644, 929.2718, 860.6365, 839.7463, 609.233, 540.0855, 
    372.2006, 284.8974, 301.0556, 328.8521, 341.0661, 315.4924, 295.3959, 
    299.6176, 278.9605, 272.5433, 239.9059, 220.9089, 222.2962, 243.0059, 
    244.9916, 215.6221, 161.5913, 138.4761, 195.9038, 395.994, 619.5784, 
    811.3644, 865.7681, 686.0972, 548.7072, 337.5479, 300.0822, 349.8788, 
    520.9444, 640.5895, 616.5434, 506.7898, 410.6275, 154.8251, 90.1037, 
    78.50664, 94.77409, 113.2795, 87.85806, 81.0833, 45.1387, 40.7375, 
    33.17309, 35.83529, 53.86729, 69.96172, 73.46383, 73.56248, 148.9393, 
    261.0967, 300.1353, 459.2666, 451.8837, 378.3816, 381.5088, 223.3205, 
    222.2062, 411.6593, 428.8239, 606.3873, 646.042, 568.9038, 505.55, 
    286.0656, 77.14314, 33.64837, 3.297961, 0, 0, 0, 0, 0, 2.244151, 
    4.955801, 76.38129, 232.1501, 266.3062, 434.145, 537.2087, 521.9823, 
    501.6171, 498.3094, 694.6164, 745.0554, 659.7027, 736.7501, 746.5898, 
    840.2108, 1043.364, 1072.436, 954.7706, 938.1902, 997.8647, 794.3143, 
    547.4996, 522.418, 468.9143, 248.3354, 150.5022, 135.2536, 103.227, 
    142.1164, 173.2986, 193.5094, 204.3717, 229.5863, 246.3172, 349.0729, 
    435.2317, 470.9053, 519.4272, 440.7462, 167.9265, 176.4665, 118.0878, 
    105.2228, 106.8183, 80.91109, 76.35849, 67.92683, 66.1326, 79.67149, 
    66.00079, 20.31273, 17.01694, 1.251958, 1.248565, 2.463363, 2.461658, 
    7.309391, 8.078649, 92.17517, 115.1139, 144.2589, 151.412, 118.2376, 
    68.0869, 118.6906, 270.4812, 258.5865, 187.1602, 142.96, 6.64469, 
    0.530213, 1.703685, 3.35584, 24.6284, 82.64381, 148.3832, 294.4089, 
    380.8008, 462.8892, 331.4127, 240.3512, 75.6171, 5.088551, 2.245178, 
    0.6060866, 0.03932895, 0, 0, 0.09076539, 2.075815, 5.305223, 30.22727, 
    158.8696, 522.1571, 985.0793, 1278.453, 1799.415, 2071.377, 2213.394, 
    2478.286, 2554.209, 2705.74, 2811.148, 2797.423, 2736.203, 2649.412, 
    2008.828, 1506.005, 1299.481, 1079.392, 813.7376, 568.7231, 332.5755, 
    81.91461, 3.301734, 0.7938613, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03154628, 0.3789333, 0.3444321, 7.950816, 
    24.87913, 49.29084, 390.3186, 594.7308, 447.4154, 368.8598, 398.8063, 
    338.315, 270.3526, 241.387, 205.6563, 176.4805, 123.5913, 61.56374, 
    15.44266, 15.56335, 56.58781, 8.468238, 0, 1.796336e-05, 0.0006869612, 
    0.001124317, 0.01055821, 0.02066588, 0.03830245, 0.1681912, 0.2666223, 
    0.2917418, 0.3418891, 0.5433533, 0.2971823, 0.02433836, 5.124776, 
    7.893463, 12.15825, 49.70943, 74.98185, 46.69952, 9.025408, 15.42976, 
    2.974206, 4.438713, 25.80215, 27.13311, 19.2051, 14.42138, 21.81066, 
    31.39333, 33.05875, 40.77766, 40.82666, 45.46812, 45.327, 51.01239, 
    52.68832, 83.11696, 107.1431, 181.584, 378.6721, 421.731, 828.4736, 
    861.0936, 929.9279, 912.6763, 805.2579, 723.7541, 621.0345, 434.2353, 
    406.8522, 360.4369, 363.0312, 380.0546, 439.9548, 485.7769, 433.1863, 
    364.0832, 314.2047, 222.3677, 178.0845, 167.7645, 183.327, 189.2155, 
    201.8522, 203.6375, 189.0745, 150.6317, 148.3065, 190.365, 424.351, 
    653.6736, 734.6793, 530.0281, 340.081, 293.0231, 289.106, 327.0493, 
    365.7855, 414.6701, 477.0976, 394.9033, 233.6338, 191.9619, 103.6808, 
    87.72089, 94.26156, 99.17967, 96.47917, 76.82737, 63.83407, 39.89161, 
    28.82531, 27.36924, 26.99343, 27.91049, 14.74314, 16.02878, 87.80204, 
    144.849, 177.0999, 216.8299, 201.9129, 106.2522, 107.8484, 97.20303, 
    95.81694, 172.7919, 184.7578, 240.4851, 262.9055, 211.1424, 143.4771, 
    96.4643, 2.598303, 1.590208, 0.0003302291, 0, 0, 0, 0, 0, 0.07487243, 
    0.5991578, 0.3164599, 76.11843, 190.2822, 154.6285, 213.987, 244.9862, 
    227.3406, 234.2985, 162.5105, 166.7688, 224.4832, 178.2304, 236.3184, 
    305.8531, 307.9664, 515.9438, 763.0024, 748.7387, 476.8637, 449.2079, 
    523.4851, 252.5942, 25.70342, 13.1048, 8.255834, 15.2962, 31.99196, 
    38.55797, 45.29905, 70.70924, 111.1557, 137.0989, 134.4492, 152.9733, 
    133.8783, 151.4449, 234.5652, 90.4547, 19.38882, 110.2923, 163.7444, 
    166.4156, 181.8149, 169.5413, 123.5023, 120.8614, 108.8013, 102.8274, 
    81.56038, 55.92279, 42.51873, 2.188808, 2.169256, 2.072838, 2.065073, 
    54.10918, 76.51178, 104.74, 119.9372, 107.2853, 47.28667, 33.63344, 
    6.695425, 5.491694, 157.6829, 204.3569, 123.8495, 36.0322, 41.39146, 
    16.19439, 14.742, 107.2656, 198.7973, 293.0785, 414.6164, 503.9863, 
    582.4972, 571.0978, 342.6558, 24.59849, 5.812427, 0.04916823, 0, 0, 0, 0, 
    0, 2.510435, 13.08559, 102.933, 309.4117, 311.289, 336.6183, 956.1763, 
    1514.321, 1759.311, 2124.267, 2355.015, 2477.191, 2718.728, 2795.241, 
    2884.71, 2958.656, 2928.309, 2706.93, 2519.901, 2403.424, 2261.878, 
    2089.283, 1715.032, 1714.814, 1390.384, 1152.663, 818.5399, 26.06024, 
    21.87491, 0.6267257, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002092206, 0.001939588, 0, 2.819104, 
    9.690909, 5.271636, 24.36625, 39.51894, 37.93415, 157.1319, 282.6814, 
    285.1447, 177.3352, 88.31767, 22.28932, 4.861166, 1.651045, 0.6387532, 
    0.04711117, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.004518855, 0, 0.1763545, 
    0.4217878, 0.3235425, 0.4687419, 0.4716088, 0.3968025, 0.9134799, 
    1.80685, 1.636135, 0.004995908, 0.050259, 1.222592, 1.331428, 15.4485, 
    30.87122, 29.60788, 21.91109, 21.85745, 28.17197, 31.78283, 32.42678, 
    32.93935, 33.06306, 36.26751, 36.27071, 47.28019, 53.69877, 63.214, 
    79.20971, 83.28892, 228.5654, 212.5577, 331.3946, 380.9676, 333.4686, 
    339.6719, 308.5343, 336.3013, 326.097, 274.8481, 324.4986, 325.631, 
    385.9315, 431.9165, 434.4316, 487.9322, 486.5526, 400.3533, 245.0974, 
    200.6815, 154.3405, 151.3657, 151.4391, 155.4274, 175.9959, 180.8223, 
    173.2802, 176.8732, 204.2144, 254.1561, 309.9952, 323.8235, 311.4831, 
    296.2622, 193.0391, 118.1543, 124.0405, 129.5596, 141.5291, 173.0228, 
    112.8414, 104.8128, 135.3307, 68.3383, 51.34541, 43.41431, 34.96099, 
    47.87151, 59.26896, 69.63024, 64.44456, 33.1958, 36.64656, 21.6995, 
    19.35295, 11.57213, 2.025564, 2.066754, 2.140966, 2.390357, 0.9228081, 
    0.04845978, 0.5238637, 1.526923, 1.551503, 3.597259, 3.540267, 4.051646, 
    4.134736, 3.874677, 3.522335, 3.058172, 1.397464, 1.801649, 1.047549, 
    0.01079319, 0.0102589, 0.0005264333, 0, 0, 0, 0, 0, 0.001922293, 
    0.00178207, 0, 8.375636, 29.09653, 16.32615, 16.75998, 29.20182, 
    24.24881, 33.91481, 22.92115, 16.94414, 26.68329, 21.80264, 10.35773, 
    50.98469, 78.03835, 34.58555, 13.90501, 27.04267, 16.99714, 1.40201, 
    1.181303, 1.302434, 0.09386167, 0.1357837, 0.4293264, 0.1738737, 
    0.2109183, 1.627126, 14.17181, 27.59934, 8.696632, 0.8427662, 1.552283, 
    3.795937, 6.648767, 4.023899, 0.1551903, 79.74555, 220.7675, 218.9723, 
    212.1464, 210.2332, 202.2739, 183.759, 170.005, 118.8666, 118.5001, 
    86.83704, 74.59409, 49.59726, 2.182123, 2.216111, 2.378325, 2.400676, 
    128.0434, 198.1301, 170.5441, 77.01752, 68.20455, 6.45439, 5.802142, 
    56.76884, 125.1982, 147.0988, 186.8056, 186.4057, 130.5452, 137.1374, 
    153.4046, 286.1644, 365.6142, 514.752, 598.7678, 613.9243, 626.4379, 
    615.8188, 446.4618, 77.3811, 22.78111, 3.1545, 0, 0, 0, 0, 0, 0.04979563, 
    5.979289, 21.3531, 159.0094, 510.1664, 853.342, 1055.414, 1253.785, 
    1753.205, 2160.003, 2246.039, 2513.329, 2704.582, 2755.863, 2932.31, 
    3016.341, 3037.975, 3047.114, 3019.234, 2912.649, 2759.285, 2647.919, 
    2023.611, 1825.246, 1547.427, 1114.831, 1052.746, 211.6943, 55.54091, 
    28.37744, 2.475487, 1.877739, 0, 0, 0, 0, 0, 0, 0, 0.3526169, 0.3622502, 
    0.1437407, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01129005, 0.1611016, 
    0.06155959, 0.4921079, 5.060236, 5.207859, 17.15756, 13.14007, 4.885071, 
    3.622243, 2.130565, 0.2201799, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1787895, 3.932854, 4.457644, 11.37424, 28.88712, 11.34025, 8.519149, 
    0.6693207, 0.003544852, 0.003998959, 0.0002094754, 0, 0.08596522, 
    0.2173533, 2.606282, 25.19457, 27.44424, 24.71391, 20.91696, 20.43615, 
    13.4305, 14.16753, 18.22003, 21.61632, 21.71048, 41.18727, 41.31262, 
    51.81037, 61.47624, 61.67217, 57.14131, 56.32438, 69.31666, 73.45463, 
    76.45298, 92.85718, 70.31824, 56.37527, 56.41111, 59.07753, 103.3043, 
    98.79597, 121.0133, 217.7656, 215.3082, 266.8255, 322.9419, 288.6444, 
    272.9561, 211.9056, 174.7396, 135.5964, 113.9947, 100.8502, 98.2429, 
    105.6102, 103.1117, 125.4043, 165.4013, 182.4245, 181.3254, 196.6318, 
    219.4795, 184.3903, 110.5088, 18.0648, 12.13951, 10.73613, 12.80105, 
    15.29695, 16.43588, 8.230871, 14.02425, 29.97926, 18.9857, 17.19992, 
    13.57385, 11.9585, 13.96772, 15.67309, 17.41601, 15.55453, 1.138336, 
    0.5249552, 0.2522034, 1.117105, 2.89572, 1.061528, 0.429966, 0.3459461, 
    0.0584243, 0.06521162, 0.006037702, 0, 0, 0, 0, 0, 0, 0, 0, 0.007331935, 
    0.07919028, 0.07094805, 0.7040008, 0.9484876, 0.6517554, 0.08337514, 
    0.08449063, 0.05158331, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05168371, 0.7374926, 
    0.281808, 0.1113399, 1.144884, 1.178283, 1.324282, 0.5852334, 
    0.007794229, 0.09388787, 0.8850846, 0.1114421, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.01200662, 0.03142135, 0.002202018, 0.1051138, 3.979558, 
    6.822487, 22.51176, 114.2097, 96.30473, 86.12609, 215.217, 228.5573, 
    249.6619, 259.3207, 257.4472, 273.1035, 267.1587, 188.6571, 121.506, 
    118.285, 45.40639, 44.63829, 24.91634, 0.8000367, 0.7811642, 25.08729, 
    25.65315, 99.69847, 158.1651, 143.1783, 8.971331, 6.455906, 45.75987, 
    109.7733, 126.6494, 150.2144, 149.8375, 163.6934, 202.3132, 230.638, 
    314.8452, 391.4384, 471.4848, 590.6155, 633.5729, 592.3283, 476.7102, 
    349.9024, 210.2554, 70.44303, 0, 0, 0, 0, 0, 0, 0, 0.1180359, 0.6959985, 
    46.13397, 241.5387, 552.2518, 798.3338, 1021.076, 1505.645, 1911.168, 
    2030.748, 2313.179, 2593.792, 2648.057, 2799.521, 2964.745, 2989.76, 
    3079.987, 3145.748, 3140.752, 3035.65, 2944.971, 2874.79, 2425.133, 
    2223.165, 1961.893, 1372.86, 1315.992, 941.4403, 668.8401, 543.3569, 
    22.38679, 7.188397, 3.226073, 0, 0, 0, 0, 0, 0, 0, 0.5936147, 0.5838628, 
    0.2639203, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.222931, 4.045791, 17.66833, 
    190.1475, 276.2941, 205.8335, 17.72166, 4.453807, 1.871546, 0, 0, 0, 
    0.0005139163, 0.01102649, 2.212696, 6.647302, 8.516181, 8.935127, 
    9.631841, 8.518692, 1.167861, 1.230512, 6.584564, 10.09186, 10.24222, 
    88.80971, 89.85795, 87.86716, 80.09071, 81.24897, 65.47025, 57.66935, 
    58.32288, 59.93869, 60.66782, 61.17618, 60.83096, 61.84586, 63.68441, 
    62.52337, 65.01978, 63.80158, 60.49374, 75.17582, 95.71252, 89.244, 
    98.28877, 129.5862, 106.2904, 80.90521, 67.88238, 67.50985, 63.0274, 
    61.95506, 53.85669, 48.25773, 59.18442, 78.51715, 95.57832, 111.432, 
    126.8992, 99.6559, 47.39682, 13.95193, 7.93328, 2.531019, 0.2855781, 
    0.195429, 0.4145107, 0.1178853, 0.004632963, 0.5218551, 4.111443, 
    9.41853, 12.84089, 11.24326, 11.4791, 9.510685, 3.396277, 4.476577, 
    5.605963, 0.5311937, 0, 0, 8.986265e-07, 1.928077e-05, 2.421524e-05, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01141747, 0.0510072, 
    0.03926415, 0.0204257, 0.006693385, 0.0003119613, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1109728, 2.019629, 2.98962, 23.1324, 109.9083, 142.0233, 
    162.0974, 171.9164, 174.5698, 177.7691, 179.0678, 185.2206, 103.8108, 
    88.6438, 108.4814, 65.1298, 58.60521, 52.19173, 9.137685, 9.466018, 
    5.32811, 2.488425, 2.474161, 71.36252, 71.6726, 78.72453, 94.28048, 
    96.39909, 42.77224, 20.26212, 35.71169, 179.1062, 189.2056, 223.6339, 
    313.6664, 322.9731, 357.8791, 427.1599, 448.0221, 566.5837, 614.1494, 
    610.5718, 200.8218, 29.15558, 19.69228, 1.124561, 0.03185803, 
    0.009629801, 0, 0, 0, 0, 0, 0, 0, 2.388714, 6.551964, 118.5045, 401.7821, 
    872.049, 1244.778, 1525.437, 1769.169, 2165.147, 2457.867, 2519.709, 
    2665.992, 2851.917, 2916.329, 2972.409, 3090.935, 3135.112, 3146.467, 
    3134.068, 3129.205, 3067.647, 2822.815, 2700.761, 2435.037, 1776.444, 
    1679.342, 1380.52, 1001.4, 977.777, 340.6629, 32.21367, 28.20054, 
    1.174744, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01179634, 0.04708815, 0.07419837, 
    0.01054658, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 2.240142, 9.766609, 12.89995, 139.6428, 258.3532, 209.2642, 
    82.53162, 6.526961, 4.355578, 0.9824101, 0, 0, 0.002805444, 0.08720528, 
    0.1227466, 0.2120782, 0.3827887, 0.433799, 0.2434374, 0.05201669, 
    0.05510908, 0.6176274, 0.7952771, 0.8090361, 91.48752, 89.93144, 
    82.08043, 59.35839, 56.40231, 57.9114, 81.94021, 83.83617, 95.32581, 
    111.8587, 116.8681, 116.0498, 117.0316, 123.0536, 102.1179, 87.48694, 
    90.6963, 79.69112, 72.14815, 75.06802, 60.81072, 50.16665, 57.95893, 
    62.57076, 39.14536, 32.39653, 32.91811, 35.34062, 27.59287, 18.54519, 
    9.269301, 3.216528, 3.273, 26.12562, 28.22354, 5.484312, 4.244867, 
    6.14327, 4.36779, 0.1858002, 0.135806, 0.05512104, 4.609846e-05, 0, 
    0.03907336, 0.1077177, 0.2710443, 0.4431338, 0.7359222, 0.6231779, 
    0.5750374, 0.6297355, 0.3331494, 0.02107608, 0.02803148, 0.002250044, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.2120616, 37.14077, 
    90.51804, 97.17203, 116.4439, 148.1465, 150.8921, 140.4983, 153.0829, 
    163.0369, 106.4638, 3.813895, 5.360915, 5.575981, 3.13886, 3.540877, 
    2.858114, 2.056646, 2.154571, 2.093306, 2.090781, 2.122128, 55.34973, 
    54.44934, 61.88563, 95.88373, 93.28148, 64.64935, 26.90603, 26.02836, 
    84.78682, 122.3019, 114.3728, 82.20609, 34.6462, 40.25586, 339.1881, 
    375.7428, 318.3542, 306.8981, 216.5912, 102.2038, 2.628926, 0.01052289, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.520032, 17.23043, 308.8558, 763.782, 
    886.7283, 1344.556, 1832.335, 2145.398, 2229.79, 2437.827, 2663.058, 
    2747.33, 2830.091, 2933.559, 3006.813, 3032.917, 3057.595, 3086.901, 
    3111.37, 3072.974, 2990.737, 2964.883, 2785.823, 2279.39, 2190.454, 
    1895.644, 1283.424, 1227.946, 972.3361, 477.4972, 436.7985, 182.3153, 
    4.480132, 4.089619, 1.075562, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05557533, 0.1646548, 0.1493024, 
    0.09278907, 0.002164904, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.9336478, 7.411664, 41.60417, 95.73727, 317.6706, 
    232.5497, 173.0507, 122.3771, 63.25102, 12.75279, 0, 0, 0, 0, 
    0.001389323, 0.001859275, 0.00210628, 0.0001985218, 0, 5.418133e-05, 
    0.005538261, 0.005813877, 0.005882056, 0.6067846, 0.5978108, 0.7293981, 
    4.943247, 4.897565, 8.702167, 109.9428, 119.8533, 123.598, 193.4414, 
    212.6801, 220.1418, 215.2512, 213.5384, 204.8573, 138.8045, 129.0788, 
    135.8481, 130.4676, 133.9239, 145.39, 137.5194, 121.7656, 145.1316, 
    173.1348, 125.5979, 15.28961, 3.666978, 2.438305, 0.634334, 0.2872208, 
    0.1584578, 0.01006543, 0.01618255, 0.01405334, 0.1417449, 0.1371105, 
    0.003695087, 0.004254925, 0.002196203, 0.002814987, 0.000758863, 
    0.04109916, 0.2294971, 0.3546463, 1.868769, 21.28282, 24.20964, 14.95845, 
    4.327038, 0.4296601, 0.2333619, 0.2143899, 0.6819046, 0.6715913, 
    0.490374, 0.1191704, 0.01071954, 0.002174542, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.04936326, 0.560281, 10.34224, 24.25971, 41.89407, 
    77.56198, 95.58471, 89.28447, 9.651242, 5.870116, 13.89363, 18.90882, 
    14.23514, 21.07078, 59.20262, 54.5088, 44.32864, 1.765566, 1.689814, 
    1.560099, 0.7811324, 0.7663231, 0.7542508, 5.117553, 5.17467, 6.373254, 
    70.62938, 74.79388, 75.21275, 136.981, 158.3989, 174.6631, 238.0255, 
    259.5518, 268.5905, 99.78564, 68.35471, 130.9524, 118.9935, 5.144613, 
    5.366468, 4.648913, 1.298131, 0.4915803, 0.01020095, 0, 0, 0, 0, 0, 
    5.384322e-09, 0.0005678148, 0.003186632, 0.01071409, 0.5558234, 12.55716, 
    118.2128, 481.7009, 872.0417, 1355.529, 1583.724, 1931.469, 2184.438, 
    2412.677, 2489.609, 2629.494, 2778.32, 2860.146, 2877.822, 2916.651, 
    2938.978, 2953.437, 2949.673, 2889.044, 2872.304, 2891.84, 2802.748, 
    2610.654, 2592.362, 2399.76, 1933.123, 1875.986, 1719.967, 1177.459, 
    1098.186, 916.819, 74.72463, 41.18377, 34.30184, 0.3727727, 0.05190104, 
    0.045563, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5357471, 2.205235, 
    92.98683, 239.7468, 301.0392, 374.0191, 454.6314, 507.3063, 458.7791, 
    53.8313, 12.63579, 11.37172, 1.905521, 0.01028968, 0.009408246, 
    0.003799471, 0, 0, 0.0001934955, 0.00114702, 0.001167644, 0.001188253, 
    0.07917888, 0.07890601, 0.07863294, 1.380615, 1.561287, 1.469311, 
    43.48175, 59.74667, 52.72649, 81.74112, 186.0909, 182.3164, 175.199, 
    152.8103, 140.47, 126.8701, 127.5607, 172.0223, 174.8016, 181.5547, 
    288.812, 354.6961, 363.3152, 307.6111, 246.1477, 216.5513, 162.7621, 
    69.10014, 10.8606, 0.000637603, 0.0003880932, 3.247865e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0041799, 0.04994637, 0.08205749, 0.2246587, 0.9661701, 
    13.1025, 27.81066, 36.92868, 28.9245, 14.03368, 12.40912, 8.098943, 
    0.9150675, 0.8121813, 0.9752111, 0.8326262, 0.1372756, 0.1049813, 
    0.07810283, 0.007014627, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0283257, 0.2362645, 0.5450493, 0.4114659, 0.5390032, 15.30516, 
    17.62284, 13.09427, 49.59177, 233.8266, 233.6767, 212.0992, 62.45203, 
    45.45558, 49.37403, 34.40012, 3.546567, 3.520004, 15.36721, 43.74399, 
    42.65796, 41.5727, 51.63267, 52.80175, 53.97166, 77.87831, 76.59154, 
    74.72577, 153.4844, 218.1336, 214.9467, 214.3591, 189.6485, 177.8799, 
    205.5759, 648.4339, 707.6396, 650.8654, 228.6538, 4.791981, 3.121726, 
    1.182703, 9.185826e-06, 0, 0.1296413, 1.76468, 7.309915, 13.709, 18.8829, 
    13.11192, 2.077553, 88.60844, 290.7913, 503.5753, 747.1946, 902.8733, 
    982.1814, 1329.531, 1697.469, 2043.089, 2124.555, 2234.162, 2453.85, 
    2629.587, 2706.326, 2728.552, 2781.351, 2837.633, 2855.92, 2858.01, 
    2796.351, 2738.549, 2742.208, 2724.089, 2620.878, 2601.473, 2619.706, 
    2483.29, 2293.212, 2297.128, 2184.901, 1581.49, 1486.295, 1456.603, 
    691.3157, 359.9765, 334.6231, 144.1276, 0.05618618, 0.05972808, 
    0.05222262, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.001426624, 0.01460581, 0.0302564, 0.04648033, 3.440905, 
    5.827036, 7.234798, 5.981942, 0.8777148, 0.09301718, 1.032225, 2.164865, 
    1.147877, 0.4090886, 0.5181287, 0.3877728, 0.1295732, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01004246, 0.3965914, 0.586934, 
    0.7525305, 5.299744, 9.776836, 10.99831, 9.87161, 5.004268, 2.501522, 
    3.625032, 3.557288, 0.1849987, 0.1710271, 0.1436844, 0.002441007, 0, 0, 
    0, 0, 0, 0, 0.04312435, 0.0425566, 0.0419884, 0.02430446, 0.01282243, 
    0.01300719, 0.4823851, 2.447163, 2.157392, 1.863459, 37.7792, 35.81408, 
    22.30786, 9.078338, 8.555648, 9.463291, 8.81891, 59.89272, 148.5211, 
    152.8116, 148.8401, 191.1424, 206.6446, 205.1475, 175.6409, 118.6692, 
    76.7033, 47.69171, 15.64608, 0.003145314, 0.001050897, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3.888616e-05, 0.2036168, 0.6161619, 0.9910291, 0.8916858, 
    0.2230152, 0.170504, 0.5991708, 2.386358, 0.2942748, 0.08226383, 
    0.1054736, 0.1747609, 0.2409313, 0.271032, 0.2393046, 0.02802818, 
    0.0001524652, 0.0001387611, 5.082736e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.005839299, 0.2306025, 0.3412793, 0.4984955, 23.45761, 45.93927, 
    51.59719, 48.20545, 25.99992, 44.4984, 65.13246, 63.64747, 6.434772, 
    7.478892, 8.521506, 3.32242, 2.138077, 2.261718, 26.98445, 62.59423, 
    63.6945, 64.79391, 74.82629, 73.59109, 72.35491, 46.68488, 28.78313, 
    27.59867, 40.13461, 203.2337, 216.3601, 218.4263, 283.4612, 409.8898, 
    435.1038, 441.5143, 277.9224, 254.1241, 280.9964, 239.5807, 46.33988, 
    0.01307672, 0.01622247, 3.497178, 11.90642, 21.50144, 103.3568, 210.4543, 
    462.8162, 710.8943, 908.8584, 986.4906, 981.0486, 1152.949, 1373.562, 
    1605.391, 1840.322, 1881.446, 1988.466, 2138.724, 2337.409, 2473.307, 
    2518.889, 2592.893, 2654.042, 2712.351, 2739.296, 2747.47, 2710.292, 
    2659.928, 2662.509, 2644.108, 2526.91, 2442.899, 2456.033, 2440.237, 
    2264.281, 2193.865, 2212.104, 2073.221, 1503.094, 1434.337, 1443.261, 
    944.0771, 435.0457, 442.9765, 431.7877, 49.08904, 1.453248, 1.355054, 
    0.580736, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.006956431, 0.2062109, 3.375202, 6.319607, 9.975802, 
    46.45114, 184.3265, 233.0237, 272.1836, 182.1654, 41.50302, 7.461129, 
    7.693655, 6.090354, 3.187601, 0.4279502, 0.003152691, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.009802716, 
    0.07145939, 0.1403449, 0.2005274, 0.08574645, 0.09865205, 0.1136614, 
    0.07822511, 0, 0, 0, 0, 0, 0, 0, 0.00640714, 0.006298584, 0.006189934, 
    0.007141049, 0.009181336, 0.008660956, 0.00813923, 0.03071029, 
    0.05141057, 0.04897726, 0.05547363, 0.5894982, 0.4170122, 0.2176536, 
    0.2024886, 2.409217, 3.429365, 3.21738, 10.99365, 63.85539, 57.12791, 
    40.22962, 26.27605, 6.838318, 0.1246243, 1.300339e-05, 5.030922e-05, 
    0.001430663, 0.001748683, 0.0007391122, 2.556974e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005153902, 0.006861422, 0, 0, 0, 0, 0, 
    0, 0, 1.986132e-06, 1.447841e-05, 2.843534e-05, 3.986978e-05, 
    6.430818e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05151607, 
    0.4027379, 0.5123837, 0.5792509, 0.4532813, 0.2880868, 1.283971, 
    2.424161, 3.441849, 0.3049393, 0.2390548, 0.2258121, 0.1254682, 
    0.09780917, 0.1005514, 0.1032866, 0.4840156, 0.6404728, 0.6476363, 
    0.6547936, 2.075105, 2.04694, 2.018751, 3.821675, 11.00225, 11.19729, 
    11.39284, 87.80696, 146.0516, 137.8936, 130.5992, 336.3596, 498.3266, 
    500.8633, 502.8024, 502.1459, 509.3895, 521.5548, 501.7248, 247.5447, 
    37.51022, 33.83801, 48.75304, 303.4308, 581.4425, 720.5878, 830.6633, 
    1051.559, 1348.561, 1639.971, 1764.883, 1775.662, 1814.732, 1894.278, 
    2066.865, 2183.192, 2229.28, 2275.125, 2332.704, 2421.136, 2510.328, 
    2527.803, 2552.099, 2577.989, 2578.809, 2564.435, 2580.133, 2565.348, 
    2458.017, 2362.439, 2356.441, 2357.422, 2219.42, 2043.028, 2029.376, 
    2038.213, 1825.052, 1447.724, 1419.741, 1419.873, 1090.46, 519.3366, 
    505.0762, 494.7145, 210.3396, 3.672246, 3.630306, 3.588475, 0.8144104, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0.1287415, 0.3172891, 0.3479449, 0.3722797, 10.56052, 65.70064, 
    142.8756, 198.0492, 298.9736, 428.8633, 412.8532, 426.3073, 432.9524, 
    303.4384, 124.8179, 12.56132, 5.847012, 4.042201, 0.9580768, 0.4456456, 
    0.0973577, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005695687, 0.02639321, 
    0.0001360721, 0, 0, 0, 0, 0, 0, 0, 0.002370212, 0.001869377, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003928374, 
    0.08108247, 0.1344825, 0.1440853, 0.1535809, 0.929767, 2.072308, 
    2.271417, 2.412489, 2.2374, 1.807042, 1.626911, 1.643325, 1.599138, 
    1.152941, 0.4125512, 0.2083259, 0.04646346, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.000232557, 0.006165095, 0.01451066, 0.03215735, 0.1054334, 0.1244902, 
    0.1419155, 0.1541189, 0.0453755, 0.04299615, 0.04384283, 0.09926861, 
    0.3893085, 0.3864437, 0.3819688, 0.3774982, 2.552748, 2.618662, 2.684638, 
    2.878389, 172.0949, 229.592, 245.8772, 263.04, 291.8297, 300.7723, 
    321.2553, 344.7227, 530.7786, 639.3574, 652.5028, 661.8023, 642.9116, 
    589.7772, 540.2611, 504.1966, 383.6034, 212.0956, 319.5726, 379.4252, 
    451.0999, 724.3992, 1023.614, 1247.62, 1246.781, 1251.871, 1408.681, 
    1639.161, 1840.118, 1893.542, 1894.781, 1960.823, 2053.795, 2152.521, 
    2237.837, 2266.712, 2276.358, 2327.453, 2363.889, 2401.005, 2438.543, 
    2435.173, 2377.748, 2326.692, 2325.413, 2320.757, 2218.384, 2040.828, 
    1979.04, 1973.371, 1920.312, 1596.571, 1401.126, 1402.163, 1403.469, 
    1081.443, 642.2661, 631.3812, 626.3508, 470.2769, 20.52407, 13.12794, 
    12.50861, 9.902725, 0.03938184, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 2.715043, 11.06731, 12.93291, 13.58595, 42.35035, 290.6929, 
    443.8628, 390.705, 333.6344, 264.6847, 227.8168, 316.1471, 337.666, 
    330.4012, 295.9265, 149.9556, 19.19813, 1.103439, 0.4753256, 0.2431479, 
    0.07273453, 0.0504125, 0.0273634, 0.008040211, 1.422252e-05, 0, 0, 0, 
    0.04101518, 0.2196053, 0.288527, 0.3350638, 0.3482242, 0.3263857, 
    0.3780928, 0.6107955, 0.6081859, 0.4810702, 0.3552586, 0.3442105, 
    0.4162166, 0.1639412, 0.05783106, 0.05497336, 0.04689931, 0.0112797, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.03761934, 0.1100873, 
    0.1190885, 0.1281182, 0.155638, 0.6966067, 0.9120213, 0.9789689, 
    1.046267, 2.328794, 4.91506, 5.412734, 5.568405, 5.190845, 2.982296, 
    1.412528, 1.210466, 1.019898, 0.6404744, 0.01668925, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0006850042, 0.00475585, 0.005730734, 0.006700537, 0.007665573, 
    0.01341315, 0.01549972, 0.01646852, 0.01743427, 0.1815393, 0.4146287, 
    0.4216131, 0.4285902, 0.43556, 11.94207, 12.12021, 12.29853, 12.47705, 
    276.8579, 551.6715, 555.0493, 558.4377, 556.1412, 483.3958, 467.3722, 
    469.2356, 471.1088, 528.1255, 576.0696, 573.0675, 568.4356, 566.2015, 
    464.5845, 398.3296, 452.895, 516.6287, 599.9387, 581.1104, 260.9912, 
    110.6626, 87.96307, 182.7001, 575.9969, 949.1753, 1131.477, 1159.289, 
    1160.141, 1293.476, 1471.611, 1656.019, 1810.608, 1874.807, 1876.74, 
    1930.521, 2004.637, 2075.738, 2136.705, 2178.917, 2214.01, 2221.167, 
    2227.531, 2219.942, 2169.858, 2063.915, 2027.799, 2024.554, 1997.257, 
    1777.84, 1540.355, 1511.441, 1505.985, 1452.708, 990.6351, 702.422, 
    699.2285, 696.0515, 659.313, 305.7498, 232.8826, 218.1033, 203.3706, 
    73.1849, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 1.220672, 1.897079, 0.730031, 0.01352223, 0.005471562, 
    1.750542, 13.01954, 20.54317, 17.84661, 14.72392, 12.97755, 69.10082, 
    47.49574, 10.46627, 8.365177, 7.910889, 6.519576, 3.429114, 0.424764, 
    0.06006074, 0.07370005, 0.07887015, 0.07887015, 0.06521574, 0.03325738, 
    0.04208241, 0.3361335, 0.6429934, 0.7804227, 0.8253127, 0.9020664, 
    1.004314, 1.126716, 1.282406, 1.261147, 1.236411, 1.254922, 2.111853, 
    3.261815, 3.571327, 3.603491, 3.407994, 2.201626, 0.7744544, 0.6315035, 
    0.5804571, 0.5297082, 0.3426896, 0.0001249023, 0, 0, 0, 0.009108757, 
    0.05517057, 0.053444, 0.05171876, 0.04999556, 0.04827438, 0.00679071, 
    0.007032826, 0.007275227, 0.007517915, 0.02772184, 0.3676009, 0.4146693, 
    0.4264466, 0.4382655, 0.582739, 0.9716326, 0.9321774, 0.8897934, 
    0.8471609, 1.159998, 0.9906637, 0.2989971, 0.003263349, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.21797e-06, 
    0.001667419, 0.00190949, 0.001940763, 0.001972, 0.0020032, 17.35738, 
    17.15617, 16.95473, 16.75305, 59.73064, 483.5388, 492.9182, 482.9938, 
    473.0343, 447.1481, 493.087, 540.082, 545.8145, 551.5806, 579.1081, 
    808.6615, 991.8098, 1016.818, 1016.505, 1003.987, 937.4294, 867.9664, 
    839.8329, 834.4373, 825.3773, 653.8682, 566.0832, 509.4825, 461.3206, 
    471.7638, 513.4021, 694.1004, 898.5355, 1050.159, 1191.467, 1248.269, 
    1248.269, 1282.863, 1348.145, 1416.86, 1534.719, 1661.981, 1792.671, 
    1841.193, 1831.78, 1852.078, 1872.838, 1869.398, 1902.115, 1935.263, 
    1893.966, 1721.401, 1558.323, 1556.19, 1562.187, 1557.007, 1283.158, 
    836.3808, 737.9418, 736.3299, 734.7275, 695.1374, 515.7474, 484.6891, 
    483.5938, 482.5024, 452.333, 39.81796, 5.27846, 5.108065, 4.937871, 
    4.767877, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0.0006340447, 0.0004262023, 3.244795e-05, 0, 0, 
    0.001555371, 0.1366034, 0.3431902, 0.3539955, 0.2830954, 0.211238, 
    0.1384057, 0.571364, 0.01348354, 0, 0, 0, 0, 0.0001097373, 0.01071619, 
    0.01071619, 0.0001097373, 0, 0, 0, 0, 0.001330174, 0.1026088, 0.3169448, 
    0.4837286, 0.6482798, 0.8106388, 0.9756802, 1.151473, 1.308381, 1.433665, 
    1.508515, 1.512465, 1.460184, 1.245418, 0.8710833, 0.8713894, 0.8716936, 
    0.8719339, 0.5884401, 0.05271416, 0, 0, 0, 0, 0.05080159, 0.1079803, 
    0.1097089, 0.1114351, 0.1131591, 0.1148808, 0.01616017, 0.01591798, 
    0.01567547, 0.01543264, 0.01518948, 0.2251997, 0.4008483, 0.3799295, 
    0.3589267, 0.33784, 0.3177203, 0.2982312, 0.2610804, 0.2231608, 
    0.1849888, 0.1465647, 0.03132969, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.211508, 3.163378, 
    3.115185, 3.066927, 3.018604, 113.2713, 214.9425, 205.7149, 196.4502, 
    187.1485, 193.7552, 465.4679, 732.3383, 747.5858, 762.8777, 778.2706, 
    859.3322, 937.0265, 979.9967, 981.7647, 974.6553, 962.3436, 911.6583, 
    836.9488, 738.0264, 669.4912, 637.5822, 605.2402, 555.7598, 586.077, 
    612.426, 620.5324, 611.9226, 577.7778, 541.6816, 583.987, 641.3745, 
    687.9949, 772.8642, 854.6941, 900.5398, 888.3361, 851.9426, 903.4217, 
    1011.029, 1128.077, 1243.558, 1355.037, 1385.324, 1228.758, 1138.356, 
    1172.027, 1193.069, 1187.329, 1033.27, 789.8279, 648.0201, 655.5637, 
    663.0577, 670.4598, 488.6609, 279.2194, 280.7811, 296.9535, 313.0615, 
    329.1051, 181.1632, 10.66936, 10.83993, 11.01027, 11.18038, 11.35027, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05519296, 
    0.1500467, 0.1642616, 0.2175887, 0.2705155, 0.323042, 0.3752258, 
    0.2609232, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05381548, 
    20.3433, 24.96029, 23.67924, 22.39228, 21.09941, 19.80063, 259.6, 
    391.3439, 357.1784, 311.0936, 264.6576, 217.8704, 217.2504, 440.4203, 
    694.8979, 836.5892, 790.4825, 720.2473, 649.1129, 532.4799, 376.2482, 
    272.4058, 206.7003, 139.728, 71.36232, 22.56477, 43.25294, 118.5302, 
    192.4339, 263.9384, 271.8977, 216.3804, 157.1932, 91.80734, 74.65115, 
    141.4928, 235.1301, 326.3662, 415.5618, 490.5019, 547.5551, 606.3943, 
    667.4617, 727.7755, 767.8253, 747.7278, 724.7731, 695.1131, 648.8344, 
    646.5984, 644.3792, 642.1767, 540.2988, 214.6301, 22.26856, 22.22654, 
    22.18472, 22.14309, 22.10165, 14.11911, 0.04053276, 0.0101087, 
    0.01026339, 0.01041783, 0.01057204, 0.01072601, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.6338732, 24.33825, 30.77678, 26.22121, 21.63318, 17.00451, 
    12.33489, 7.624318, 20.25182, 7.180273, 11.79697, 16.05005, 16.12449, 
    14.49078, 12.83217, 11.14867, 9.655749, 8.490761, 6.332207, 3.422223, 
    0.6367931, 0, 0, 0, 0, 2.218234, 11.92113, 22.0579, 29.78627, 34.34187, 
    39.8235, 45.837, 51.76162, 57.59729, 60.37043, 54.58566, 47.29338, 
    60.6195, 99.94553, 139.5351, 178.7807, 217.682, 255.8241, 285.2885, 
    220.4157, 17.25861, 12.59692, 13.3699, 14.13877, 14.90351, 15.66412, 
    12.8525, 0.3425127, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.001286788, 0.004872708, 0.004556906, 0.00375653, 
    0.002949522, 0.002134513, 0.001310874, 0.0004786106, 2.112361e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.006153398, 
    1.394213, 3.818633, 6.217928, 8.592085, 10.94293, 13.27446, 14.20905, 
    3.897211, 0.2053401, 0.2195868, 0.2337431, 0.2478088, 0.2617841, 
    0.2756689, 0.2893474, 0.1457981, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
