netcdf \00010101.river_month.tile4.rv_o_h2o {
dimensions:
	time = UNLIMITED ; // (12 currently)
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float rv_o_h2o(time, grid_yt, grid_xt) ;
		rv_o_h2o:_FillValue = -1.e+08f ;
		rv_o_h2o:missing_value = -1.e+08f ;
		rv_o_h2o:units = "kg/m2/s" ;
		rv_o_h2o:long_name = "river outflow, h2o mass" ;
		rv_o_h2o:cell_methods = "time: mean" ;
		rv_o_h2o:time_avg_info = "average_T1,average_T2,average_DT" ;
		rv_o_h2o:coordinates = "geolon_t geolat_t" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "areacellr: 00010101.river_static_cmip.nc land_area: 00010101.river_static.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Fri Aug 29 14:00:38 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 /work/cew/scratch//00010101.river_month.tile4.nc -O /work/cew/scratch/workflow-test/river_month//ncks_out//00010101.river_month.tile4.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 31, 28, 31, 30, 31, 30, 31, 31, 30, 31, 30, 31 ;

 average_T1 = 0, 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334 ;

 average_T2 = 31, 59, 90, 120, 151, 181, 212, 243, 273, 304, 334, 365 ;

 rv_o_h2o =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.74502e-05, 9.674058e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.098879e-05, 2.476873e-05, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  1.485455e-05, 5.204221e-05, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 3.175799e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.056132e-05, 1.309405e-05, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.530168e-05, 1.548065e-05, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  1.532359e-05, 1.031035e-05, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 3.727606e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  6.598997e-06, 1.223693e-05, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.453134e-05, 1.324237e-05, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  1.413814e-05, 9.732708e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 3.038601e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  4.381469e-06, 6.427172e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.162161e-05, 8.946614e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  6.275175e-06, 6.760555e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 3.195718e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  2.200511e-06, 4.019693e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  7.306505e-06, 5.575252e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  3.264305e-06, 3.463285e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 3.455353e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  9.212015e-07, 2.085745e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  4.753859e-06, 3.42161e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  8.686408e-07, 2.607322e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 9.589613e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  7.144151e-06, 2.065638e-05, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  2.922873e-05, 6.780586e-05, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  4.709338e-05, 6.781388e-05, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 4.925493e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  2.570043e-06, 3.81459e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.381133e-05, 5.872985e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  3.276348e-06, 3.924609e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 2.522243e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.779718e-06, 2.402312e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  6.324061e-06, 3.543022e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  1.536248e-06, 2.114138e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 2.114569e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  9.04955e-07, 1.353036e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  3.649247e-06, 2.290774e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  1.013921e-06, 1.223131e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 2.176797e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  7.366036e-07, 1.184777e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  2.608617e-06, 2.309598e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  1.987395e-06, 1.270411e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 2.235563e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  1.370563e-06, 2.060396e-06, 0, 0, _, _, _, _, _, _, _, _, _, _, _,
  2.697007e-06, 4.11645e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  2.142113e-06, 3.98037e-06, 0, _, _, _, _, _, _, _, _, _, _, 0, _,
  0, 0, 0, 0, _, 0, 0, _, _, _, _, 0, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 2.70476e-05, 0, 0, 0, _, _, _, _, _,
  _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _,
  _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _ ;

 time_bnds =
  0, 31,
  31, 59,
  59, 90,
  90, 120,
  120, 151,
  151, 181,
  181, 212,
  212, 243,
  243, 273,
  273, 304,
  304, 334,
  334, 365 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 time = 15.5, 45, 74.5, 105, 135.5, 166, 196.5, 227.5, 258, 288.5, 319, 349.5 ;
}
