netcdf atmos_daily.00010101-00010701.ps.tile6 {
dimensions:
	time = UNLIMITED ; // (182 currently)
	phalf = 66 ;
	scalar_axis = 1 ;
	grid_yt = 10 ;
	grid_xt = 15 ;
	nv = 2 ;
	pfull = 65 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float bk(phalf) ;
		bk:_FillValue = 1.e+20f ;
		bk:missing_value = 1.e+20f ;
		bk:long_name = "vertical coordinate sigma value" ;
		bk:cell_methods = "time: point" ;
	float height10m(scalar_axis) ;
		height10m:_FillValue = 1.e+20f ;
		height10m:missing_value = 1.e+20f ;
		height10m:units = "m" ;
		height10m:long_name = "Height" ;
		height10m:cell_methods = "time: point" ;
		height10m:axis = "Z" ;
		height10m:positive = "up" ;
		height10m:standard_name = "height" ;
	float height2m(scalar_axis) ;
		height2m:_FillValue = 1.e+20f ;
		height2m:missing_value = 1.e+20f ;
		height2m:units = "m" ;
		height2m:long_name = "Height" ;
		height2m:cell_methods = "time: point" ;
		height2m:axis = "Z" ;
		height2m:positive = "up" ;
		height2m:standard_name = "height" ;
	float land_mask(grid_yt, grid_xt) ;
		land_mask:_FillValue = 1.e+20f ;
		land_mask:missing_value = 1.e+20f ;
		land_mask:valid_range = -0.01f, 1.01f ;
		land_mask:long_name = "fractional amount of land" ;
		land_mask:cell_methods = "time: point" ;
		land_mask:interp_method = "conserve_order1" ;
	float pk(phalf) ;
		pk:_FillValue = 1.e+20f ;
		pk:missing_value = 1.e+20f ;
		pk:units = "pascal" ;
		pk:long_name = "pressure part of the hybrid coordinate" ;
		pk:cell_methods = "time: point" ;
	float ps(time, grid_yt, grid_xt) ;
		ps:_FillValue = 1.e+20f ;
		ps:missing_value = 1.e+20f ;
		ps:units = "Pa" ;
		ps:long_name = "Surface Air Pressure" ;
		ps:cell_methods = "time: mean" ;
		ps:cell_measures = "area: area" ;
		ps:time_avg_info = "average_T1,average_T2,average_DT" ;
		ps:standard_name = "surface_air_pressure" ;
	float sftlf(grid_yt, grid_xt) ;
		sftlf:_FillValue = 1.e+20f ;
		sftlf:missing_value = 1.e+20f ;
		sftlf:units = "1.0" ;
		sftlf:long_name = "Fraction of the Grid Cell Occupied by Land" ;
		sftlf:cell_methods = "time: point" ;
		sftlf:cell_measures = "area: area" ;
		sftlf:standard_name = "land_area_fraction" ;
		sftlf:interp_method = "conserve_order1" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	float zsurf(grid_yt, grid_xt) ;
		zsurf:_FillValue = 1.e+20f ;
		zsurf:missing_value = 1.e+20f ;
		zsurf:units = "m" ;
		zsurf:long_name = "surface height" ;
		zsurf:cell_methods = "time: point" ;
		zsurf:interp_method = "conserve_order1" ;
	double grid_xt(grid_xt) ;
		grid_xt:units = "degrees_E" ;
		grid_xt:long_name = "T-cell longitude" ;
		grid_xt:axis = "X" ;
	double grid_yt(grid_yt) ;
		grid_yt:units = "degrees_N" ;
		grid_yt:long_name = "T-cell latitude" ;
		grid_yt:axis = "Y" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double pfull(pfull) ;
		pfull:units = "mb" ;
		pfull:long_name = "ref full pressure level" ;
		pfull:axis = "Z" ;
		pfull:positive = "down" ;
	double phalf(phalf) ;
		phalf:units = "mb" ;
		phalf:long_name = "ref half pressure level" ;
		phalf:axis = "Z" ;
		phalf:positive = "down" ;
	double scalar_axis(scalar_axis) ;
		scalar_axis:long_name = "none" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "area: 00010101.grid_spec.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Sat Aug 23 13:54:11 2025: ncks -d grid_xt,0,14 -d grid_yt,0,9 -d time,0,181 /work/cew/scratch//00010101.atmos_daily.tile6.nc -O /work/cew/scratch/atmos_subset/raw//00010101.atmos_daily.tile6.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 average_T1 = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 
    36, 37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 
    54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 
    72, 73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 
    90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 
    106, 107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 
    120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 
    134, 135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 
    148, 149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 
    162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 
    176, 177, 178, 179, 180, 181 ;

 average_T2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 
    37, 38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 
    55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 
    73, 74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 
    91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 
    107, 108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 
    121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 
    135, 136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 
    149, 150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 
    163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 
    177, 178, 179, 180, 181, 182 ;

 bk = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.00193294, 0.00749994, 0.01640714, 0.02841953, 
    0.04334756, 0.06103661, 0.0813586, 0.1042054, 0.1294836, 0.1571101, 
    0.1870091, 0.2191095, 0.2533426, 0.2896406, 0.3279357, 0.3681587, 
    0.4102391, 0.454293, 0.5001689, 0.5468886, 0.5935643, 0.6397641, 
    0.6851825, 0.729505, 0.7723162, 0.8125153, 0.8492141, 0.8817441, 
    0.909788, 0.9332725, 0.9524949, 0.9678352, 0.9798011, 0.9889621, 0.99575, 1 ;

 height10m = 10 ;

 height2m = 2 ;

 land_mask =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 pk = 1, 5.134703, 14.0424, 30.72784, 53.79506, 82.4549, 117.056, 158.6284, 
    208.79, 270.0273, 345.5085, 438.4194, 551.8527, 689.2505, 854.4094, 
    1051.478, 1284.95, 1559.651, 1880.717, 2253.565, 2683.865, 3177.496, 
    3740.5, 4379.036, 5099.326, 5907.593, 6810.008, 7812.624, 8921.319, 
    10141.74, 11285.93, 12188.79, 12884.3, 13400.12, 13758.85, 13979.1, 
    14076.26, 14063.13, 13950.46, 13747.31, 13461.45, 13099.54, 12667.38, 
    12170.08, 11612.19, 10997.8, 10330.65, 9611.055, 8843.304, 8045.85, 
    7236.312, 6424.557, 5606.509, 4778.059, 3944.972, 3146.775, 2416.634, 
    1778.226, 1246.215, 826.5195, 511.2139, 290.7407, 150, 68.893, 14.999, 0 ;

 ps =
  101712.3, 101782.5, 101844.1, 101902.7, 101954.6, 101997.3, 102033.4, 
    102064.2, 102088.4, 102100.8, 102097.9, 102077.7, 102040.9, 101990.5, 
    101917.2,
  101679.3, 101752.2, 101820.3, 101887, 101945.6, 101998.8, 102039.5, 
    102074.9, 102103.7, 102119.1, 102120.9, 102107.6, 102068.4, 102013.2, 
    101941.8,
  101629, 101709.6, 101785.1, 101861.3, 101927.7, 101987, 102036.5, 102078.9, 
    102111.5, 102131.3, 102139.4, 102129, 102096, 102041.5, 101969.9,
  101569.7, 101657, 101740.7, 101824.3, 101900.6, 101971.5, 102031.1, 
    102078.4, 102113.4, 102141.8, 102152.2, 102145.2, 102120.6, 102065.1, 
    101997.3,
  101494.6, 101592.5, 101680.7, 101774.9, 101861.2, 101942.5, 102012.7, 
    102069.5, 102112.2, 102144, 102159, 102158.9, 102137.1, 102089.4, 102020.8,
  101405, 101513.7, 101608.9, 101713.5, 101808.9, 101903.7, 101985, 102054.5, 
    102107.5, 102144.3, 102169.1, 102170, 102151.1, 102106.7, 102041.5,
  101299.4, 101418.4, 101520.1, 101638.4, 101742.8, 101848.6, 101944, 
    102027.2, 102093.3, 102138.2, 102168.9, 102178.4, 102164.1, 102126.6, 
    102063.5,
  101179.1, 101306.8, 101417.2, 101549.4, 101664.2, 101786.1, 101891.2, 
    101989.7, 102067.6, 102131.3, 102165.5, 102185.4, 102176.4, 102142.6, 
    102083,
  101039.4, 101171.3, 101295.1, 101440.9, 101571.1, 101706.7, 101826.7, 
    101942.4, 102030.8, 102110, 102158.2, 102186.3, 102185.5, 102157.6, 
    102103.2,
  100882.1, 101020.7, 101157.8, 101315.3, 101464.5, 101615.8, 101752.6, 
    101881, 101986.5, 102075.1, 102138.7, 102175.5, 102189, 102170.8, 102120.8,
  101731.4, 101778.5, 101818.3, 101845.3, 101861.6, 101868, 101863.8, 
    101855.9, 101843.2, 101818.8, 101781.2, 101731.8, 101671.7, 101602.9, 
    101525.8,
  101711.8, 101763.9, 101811.5, 101846, 101871.6, 101889.4, 101892.3, 
    101894.7, 101882.2, 101860.9, 101829.6, 101789.8, 101734.9, 101664, 
    101587.3,
  101679.8, 101737.5, 101792.8, 101844.3, 101881.7, 101907.3, 101921, 
    101923.8, 101918.3, 101900.5, 101873.8, 101834, 101780.6, 101716.8, 
    101636.5,
  101635.2, 101700.3, 101764.8, 101825, 101876.3, 101915.5, 101939.9, 
    101951.1, 101955.3, 101944.4, 101918.1, 101880.9, 101828.4, 101762.7, 
    101681.5,
  101577.1, 101658.3, 101730.6, 101798.2, 101862, 101914.9, 101956.4, 
    101978.9, 101985.4, 101978.5, 101956.9, 101921.2, 101870.5, 101803.7, 
    101719.1,
  101507.4, 101598.2, 101680.6, 101763.1, 101835.3, 101898.1, 101951.2, 
    101986, 102001.6, 102009.9, 101990.9, 101959.4, 101905.7, 101843, 101755.8,
  101424.2, 101528.6, 101622, 101716.7, 101797.6, 101874, 101936, 101986.6, 
    102012, 102027.9, 102016.8, 101986.5, 101935.9, 101875.1, 101791.1,
  101320, 101444.2, 101548.2, 101658.8, 101753, 101842.5, 101914.2, 101978.1, 
    102020.3, 102045.3, 102034.6, 102008.9, 101962.4, 101904.4, 101819.2,
  101199.7, 101341.5, 101462.1, 101591, 101695.8, 101799.7, 101884.7, 
    101960.4, 102013.8, 102051.5, 102050.8, 102029.9, 101979, 101921.3, 
    101848.3,
  101053.7, 101219.8, 101357.8, 101508.5, 101631.3, 101748.5, 101844.4, 
    101934.8, 101996.4, 102045.5, 102056.6, 102043.3, 102000.2, 101937.9, 
    101869.2,
  101710.1, 101719.9, 101705.1, 101677.2, 101630.8, 101564.5, 101477.3, 
    101369.9, 101238.4, 101072.6, 100877.9, 100657.2, 100413, 100171.1, 
    99942.59,
  101711.6, 101720.4, 101725.2, 101714.2, 101681.2, 101629.6, 101561.1, 
    101464.3, 101343, 101193.3, 101014.8, 100808.7, 100578.4, 100330.7, 100110,
  101700.2, 101725, 101736.9, 101743, 101728.8, 101696.8, 101644, 101566.8, 
    101462, 101324.7, 101157.7, 100963.3, 100744.2, 100501.9, 100275.3,
  101674.8, 101711.4, 101736.9, 101756.8, 101757.5, 101743.4, 101708.2, 
    101650, 101565.8, 101450.3, 101300.1, 101118.8, 100914.8, 100683.3, 
    100469.9,
  101640.3, 101688.6, 101725.3, 101758.1, 101774.7, 101784.4, 101768.9, 
    101728.7, 101665.2, 101573.6, 101448.5, 101282.7, 101102, 100892.3, 100685,
  101595.8, 101652, 101702.7, 101745.4, 101773.7, 101798.6, 101805.3, 
    101791.3, 101749.3, 101675, 101575.6, 101443.4, 101281.7, 101102.1, 
    100907.6,
  101539.4, 101603.6, 101668.2, 101719.6, 101770.6, 101803.6, 101830.4, 
    101836, 101817.2, 101768.4, 101693.2, 101588.4, 101459.4, 101304, 101128.5,
  101468.1, 101544, 101616, 101684.7, 101748.7, 101803.9, 101841.2, 101869.4, 
    101873.4, 101847.9, 101795.8, 101712.2, 101611.2, 101486.6, 101331.4,
  101391.7, 101477.8, 101557.3, 101638.5, 101714.5, 101786.6, 101840.3, 
    101879.7, 101906.3, 101906.3, 101876, 101814.4, 101741.3, 101635.9, 
    101505.9,
  101303.1, 101396.1, 101487.8, 101582.9, 101668.6, 101752.9, 101827.9, 
    101884.5, 101924.9, 101942, 101928.2, 101884.7, 101825.6, 101742.8, 
    101640.7,
  101665.6, 101604.3, 101512.2, 101389.9, 101232.2, 101054.9, 100859.9, 
    100668.4, 100471.3, 100268.2, 100135.8, 100036.7, 99970.12, 100010, 
    99987.55,
  101715.8, 101673.2, 101595.1, 101493.5, 101353.4, 101186.2, 100985.8, 
    100782, 100574.8, 100367.4, 100167.3, 100060.5, 99953.3, 99948.8, 99933.7,
  101750.3, 101722.5, 101664.5, 101590.1, 101471, 101324, 101143.2, 100935.2, 
    100713.3, 100487.6, 100269.1, 100098.7, 99971.12, 99898.38, 99896.64,
  101766.8, 101758.6, 101719.8, 101666.9, 101574.3, 101449.6, 101287.3, 
    101095.7, 100874.2, 100633.6, 100386.4, 100165.4, 100010.6, 99868.82, 
    99833.92,
  101768.6, 101772.4, 101755.7, 101720.8, 101658, 101563.2, 101432.2, 
    101263.9, 101065.8, 100825.4, 100562.1, 100311.1, 100094.4, 99925.64, 
    99794.02,
  101768.1, 101779.1, 101786.6, 101768.9, 101724.7, 101655.5, 101553.4, 
    101416, 101243.3, 101027.9, 100777.7, 100501.4, 100239, 100031.8, 99848.59,
  101762.6, 101784.2, 101792.6, 101800.1, 101776.7, 101732, 101657.2, 
    101548.7, 101407, 101228.6, 100998.2, 100749.9, 100457, 100192.7, 99977.5,
  101748.4, 101782.6, 101803.9, 101822.5, 101814.5, 101792.8, 101742.6, 
    101665.8, 101550.2, 101404.6, 101214.4, 100983.3, 100728.3, 100431.8, 
    100162.6,
  101718.9, 101770.8, 101807.7, 101839.6, 101851.8, 101850.4, 101821, 101765, 
    101681.8, 101563.9, 101408.3, 101214, 100982.9, 100720.9, 100424.9,
  101675.1, 101743.4, 101796.6, 101837.9, 101863.3, 101882.5, 101876.2, 
    101848.8, 101791.4, 101699.6, 101579.5, 101419, 101221.1, 100990.3, 
    100721.9,
  101061, 100928.6, 100839.1, 100777, 100745.7, 100767.4, 100794.9, 100785.1, 
    100760.2, 100729, 100667.4, 100573, 100454.6, 100320.2, 100180.4,
  101136.6, 101012.7, 100895.7, 100807.8, 100755.1, 100744.6, 100761.5, 
    100768.6, 100744.6, 100708.5, 100656.4, 100570.7, 100452.6, 100316.9, 
    100168.6,
  101252.2, 101129.9, 100991.2, 100871.9, 100775.7, 100730.4, 100731.1, 
    100743.3, 100735.8, 100697.8, 100649.3, 100577.9, 100469.7, 100335.6, 
    100181.2,
  101359.9, 101258.9, 101111.6, 100964.8, 100845.7, 100754, 100708.8, 
    100706.6, 100707.3, 100690.7, 100642.5, 100577.5, 100485.3, 100359.7, 
    100204.6,
  101457.6, 101376.8, 101259.4, 101125.1, 100969.9, 100837.7, 100742.1, 
    100694.3, 100683, 100665.6, 100644, 100580.1, 100496.1, 100386, 100243.8,
  101534.2, 101476, 101381.9, 101269.1, 101131.9, 100988.9, 100852.4, 
    100741.6, 100681.3, 100661.5, 100625.1, 100586.4, 100510.4, 100408.2, 
    100280.1,
  101616.8, 101572.7, 101503, 101407.9, 101289.5, 101154.8, 101021.4, 
    100879.1, 100761.2, 100655.8, 100636.5, 100576.8, 100522.6, 100433.2, 
    100311.2,
  101686.5, 101657.6, 101609, 101535, 101438.1, 101323.6, 101195.1, 101058.6, 
    100915, 100781.5, 100658.4, 100604.2, 100525, 100452.1, 100350.8,
  101720.1, 101711.6, 101688.5, 101641.6, 101571.9, 101480.7, 101368, 
    101234.4, 101106.1, 100944.7, 100804.9, 100661.9, 100569.5, 100474.5, 
    100376.6,
  101735.3, 101743.9, 101735.9, 101706.1, 101658.5, 101592.6, 101513.9, 
    101402, 101273.4, 101140, 100983.7, 100826.4, 100662.7, 100541.7, 100426.8,
  100507.3, 100537.7, 100505.3, 100472, 100408, 100338.4, 100265.3, 100196.7, 
    100133.6, 100080.5, 100049, 100028.6, 100026.5, 100037.9, 100055.1,
  100495.6, 100521.8, 100495.9, 100469.8, 100417.1, 100343.9, 100266.3, 
    100183.9, 100106.2, 100043.4, 99994.35, 99962.12, 99946.73, 99943.41, 
    99951.76,
  100497.9, 100500.5, 100473.7, 100456.2, 100417.4, 100356.1, 100273.2, 
    100191.4, 100111.7, 100037.3, 99970.91, 99918.87, 99883.05, 99865.89, 
    99858.16,
  100527.9, 100492.2, 100451.1, 100445.8, 100401, 100362.1, 100292.3, 
    100204.4, 100112.2, 100031.4, 99953.42, 99892.02, 99834.98, 99801.33, 
    99781.21,
  100587.6, 100537.6, 100461.8, 100431.6, 100389.6, 100368.3, 100312.7, 
    100236.9, 100141.7, 100053.5, 99962.38, 99887.52, 99819.18, 99764.51, 
    99726.73,
  100669.6, 100595.7, 100509.9, 100455, 100393.4, 100360.7, 100314.6, 
    100269.3, 100186.1, 100080.3, 99982.55, 99902.29, 99824.04, 99759.59, 
    99690.21,
  100803.3, 100691.4, 100576.7, 100515.8, 100442.8, 100380.2, 100329.5, 
    100281.9, 100234.5, 100148.2, 100030.1, 99925.7, 99856.59, 99768.22, 
    99698.56,
  100979.6, 100860, 100718.6, 100614, 100536.1, 100452.2, 100379.1, 100307.5, 
    100254.9, 100205.1, 100115, 99996.88, 99883.3, 99803.27, 99717.73,
  101142.7, 101048.5, 100918.1, 100793, 100686, 100578.2, 100486.5, 100396.4, 
    100318, 100251, 100184.3, 100097.6, 99976.38, 99861.58, 99755.65,
  101255.5, 101178.9, 101067.7, 100967.8, 100863.2, 100752.9, 100640.7, 
    100535.3, 100434.8, 100348.9, 100269.7, 100188, 100085.9, 99971.09, 
    99842.99,
  100226, 100198.9, 100160, 100143.1, 100134, 100136.2, 100155, 100186.4, 
    100229.5, 100286, 100353.4, 100429.5, 100511.1, 100594, 100676.6,
  100206.1, 100168.1, 100119.4, 100080.8, 100058.7, 100054.5, 100056.2, 
    100073.6, 100109.1, 100159.6, 100223.4, 100302.1, 100389.6, 100479.5, 
    100572.5,
  100186, 100147.7, 100087.4, 100038.8, 100001.3, 99978.44, 99975.98, 
    99982.47, 100004.5, 100041.8, 100099.7, 100170.2, 100258.1, 100352.7, 
    100452,
  100185.8, 100131, 100067.1, 100016.8, 99961.12, 99925.88, 99908.05, 
    99902.72, 99918.58, 99940.37, 99985.48, 100048.2, 100130.5, 100228.6, 
    100333.9,
  100176.9, 100117.3, 100064.4, 100011.7, 99943.26, 99895.77, 99857.27, 
    99844.84, 99845.12, 99865.23, 99890.77, 99941.65, 100012.4, 100102.5, 
    100207.3,
  100164.1, 100147.4, 100055.9, 100001.6, 99944.73, 99880.58, 99833.09, 
    99792.67, 99777.06, 99782.58, 99805.19, 99840.66, 99907.83, 99999.57, 
    100096.6,
  100154.5, 100156.4, 100083, 100008.3, 99941.87, 99884.99, 99825.4, 
    99771.89, 99709.22, 99693.5, 99705.25, 99726.76, 99783.84, 99875.23, 
    100000.3,
  100201, 100141.6, 100093.4, 100035.4, 99959.5, 99898.27, 99835.28, 
    99771.34, 99708.82, 99653.87, 99604.39, 99600.24, 99642.06, 99748.67, 
    99894.12,
  100281.2, 100188.8, 100096.5, 100052, 99980.3, 99922.01, 99865.55, 
    99804.75, 99728.68, 99669.12, 99605.77, 99564.87, 99545.47, 99623.49, 
    99771.44,
  100404.1, 100299.9, 100159, 100065.3, 100012.4, 99950.84, 99901.3, 99851.8, 
    99789.52, 99730.34, 99671.41, 99636.62, 99613.73, 99654.73, 99720.95,
  100797, 100773.9, 100756.9, 100752.3, 100755.3, 100766.1, 100778.4, 
    100794.6, 100816.8, 100842.3, 100873.1, 100900.5, 100928.8, 100953.8, 
    100978,
  100774, 100739, 100707, 100692.4, 100688, 100686.8, 100695, 100705.5, 
    100723.1, 100746.3, 100779.8, 100819.1, 100860.9, 100900.5, 100932.8,
  100759.3, 100712.4, 100666.8, 100634.9, 100615.2, 100612.3, 100610.5, 
    100612.8, 100623.7, 100641.4, 100671.5, 100709, 100752, 100798.8, 100847.1,
  100746.7, 100692.9, 100633.2, 100590.8, 100564.3, 100550.9, 100537.4, 
    100532, 100521.9, 100532, 100554.5, 100595.9, 100643.9, 100701.8, 100755.4,
  100747.9, 100691.8, 100619.9, 100571.5, 100525.6, 100500.2, 100475.7, 
    100448.9, 100425.6, 100416.3, 100425.1, 100459.5, 100508.8, 100570.1, 
    100635.9,
  100742.5, 100699.4, 100622.6, 100563, 100509.8, 100471.1, 100430.4, 
    100384.6, 100335.7, 100286, 100267.6, 100301.4, 100367, 100433.2, 100503.3,
  100751.5, 100707, 100636.7, 100572.8, 100508.6, 100454.9, 100400.1, 
    100333.3, 100245.7, 100129, 100079.1, 100093.8, 100174, 100268.5, 100350.8,
  100747.3, 100729.7, 100655.6, 100596.9, 100525.1, 100465.1, 100397.4, 
    100304.8, 100192.7, 100032.6, 99921.7, 99910.23, 99986.13, 100089.4, 
    100179,
  100760.8, 100739.6, 100681.7, 100627, 100552.8, 100483.6, 100416.2, 
    100320.6, 100196.7, 100032.1, 99879.52, 99815.49, 99848.78, 99937.74, 
    100012.5,
  100830.1, 100762.9, 100703.8, 100662.7, 100590.5, 100523, 100441.3, 
    100358.7, 100237.7, 100093.5, 99932.63, 99829.07, 99813.39, 99832.11, 
    99870.77,
  101253.6, 101265.8, 101263.5, 101261.5, 101260.2, 101256.9, 101251.6, 
    101248.6, 101242.5, 101229.9, 101218.1, 101193.9, 101164.9, 101131.1, 
    101092.5,
  101217.3, 101229.4, 101231.4, 101237.3, 101234.9, 101236.2, 101236.7, 
    101234.4, 101235.1, 101228, 101211.1, 101185.8, 101156.1, 101118.3, 
    101072.7,
  101179, 101188.3, 101189.1, 101192.8, 101194.9, 101198.3, 101196.2, 
    101192.6, 101193.8, 101188.6, 101183.1, 101169.5, 101146.6, 101111.1, 
    101070,
  101138.6, 101148.7, 101148.8, 101160.4, 101160.2, 101163.2, 101160.1, 
    101160.4, 101154.6, 101154, 101147.4, 101142.2, 101127.8, 101103.6, 
    101059.1,
  101104.8, 101111, 101110.8, 101120.2, 101121.4, 101119.9, 101117.5, 
    101114.4, 101107.8, 101107.4, 101105.6, 101102.4, 101092.4, 101071.8, 
    101032.1,
  101080.2, 101086, 101081.5, 101087.2, 101086.3, 101088.2, 101080.1, 
    101070.3, 101059.4, 101052, 101047.1, 101043.3, 101036.8, 101026, 100999.2,
  101052.2, 101053.4, 101054.2, 101053.7, 101051.1, 101048.1, 101036.6, 
    101024.1, 101005.2, 100992.6, 100980.8, 100977.4, 100976, 100970.6, 
    100954.5,
  101037.5, 101037, 101028.2, 101030.3, 101029.1, 101011.7, 100994.2, 
    100974.6, 100944.9, 100927.2, 100910.3, 100901, 100897.9, 100894.5, 
    100891.3,
  101007.1, 101022, 101015.7, 101011.5, 101004.8, 100996.9, 100969, 100933.5, 
    100890, 100851.7, 100828.2, 100820.1, 100813.8, 100818.3, 100817,
  100974.6, 101000.5, 101004.6, 101002.7, 100988.7, 100979.9, 100952.7, 
    100903.4, 100850.1, 100791.8, 100748.2, 100729.5, 100715.7, 100715.9, 
    100721.7,
  101210.4, 101212.4, 101207.3, 101185.1, 101165.1, 101135.2, 101091, 
    101043.2, 100994.1, 100953.9, 100912.7, 100875.5, 100854, 100840.4, 100835,
  101207.1, 101205.7, 101197.2, 101184.7, 101164.1, 101128.7, 101079.5, 
    101028.5, 100968.9, 100906.3, 100853.4, 100804.4, 100767.7, 100739.9, 
    100726.2,
  101177.8, 101180.7, 101177, 101167.6, 101150.2, 101120.1, 101072.7, 
    101011.1, 100946, 100874, 100805, 100734.3, 100679.5, 100635.5, 100613.5,
  101148.4, 101153.7, 101157.4, 101154.4, 101136.6, 101112.3, 101066.8, 
    101002.5, 100931.8, 100846.9, 100760.5, 100677, 100602.7, 100543.7, 
    100507.4,
  101109.1, 101115.8, 101123.9, 101126.6, 101117, 101106.4, 101068.5, 
    101012.9, 100935.1, 100844.8, 100746.4, 100640.9, 100549, 100467.6, 
    100417.7,
  101061.9, 101081.5, 101087.2, 101096.2, 101099.4, 101089.8, 101065.4, 
    101020.6, 100949.3, 100856.9, 100754, 100638.8, 100518.5, 100410.8, 
    100344.3,
  101011.7, 101039.7, 101048.5, 101061.4, 101066.7, 101069.5, 101058.3, 
    101025.4, 100972.8, 100890.8, 100791.2, 100669.8, 100540.2, 100406.5, 
    100309.9,
  100963, 100991.9, 101001.6, 101018.9, 101029, 101038.2, 101038.6, 101024.6, 
    100988.2, 100924, 100840.9, 100729.9, 100600.2, 100445, 100307.8,
  100907.7, 100939.1, 100958.9, 100978, 100991.2, 100999.7, 101008.8, 
    101001.1, 100980.9, 100947.3, 100885.4, 100796.1, 100684.4, 100549.8, 
    100418.2,
  100861.7, 100889.1, 100914.6, 100936.5, 100957.3, 100971.9, 100979.2, 
    100977.9, 100972.4, 100934.2, 100910.3, 100851.3, 100768.9, 100655.1, 
    100551.9,
  101065, 101053.3, 101047.4, 101044.4, 101044.1, 101056, 101074.5, 101103.4, 
    101131.9, 101168.9, 101202, 101240.1, 101272.5, 101301.4, 101321.4,
  101058.1, 101033.4, 101012, 100998.1, 100988.4, 100989, 100996.5, 101012.2, 
    101034.4, 101065.4, 101103.4, 101147.2, 101193.1, 101235.7, 101272.2,
  101034.1, 101003.5, 100973.1, 100946.1, 100921.3, 100904.8, 100898.3, 
    100904.8, 100921.4, 100948.4, 100987.8, 101035.5, 101091.3, 101147.9, 
    101198.1,
  101024.3, 100982.6, 100941.5, 100901, 100862, 100827, 100800.3, 100786.6, 
    100785.5, 100800.3, 100833.6, 100883.7, 100952.2, 101026.3, 101099.8,
  101007.1, 100957, 100911.9, 100859.8, 100804.2, 100749.1, 100696.3, 
    100657.7, 100634.9, 100629.2, 100649.2, 100698.8, 100775.2, 100867.7, 
    100967.1,
  100995.1, 100939.3, 100889.2, 100828, 100759, 100684.3, 100602.8, 100527, 
    100467.8, 100432.6, 100427.9, 100462.5, 100541.9, 100653, 100783,
  100984.1, 100922, 100869.2, 100802.5, 100722.8, 100631.1, 100528.6, 100422, 
    100317.7, 100233.3, 100189.5, 100195.3, 100269.8, 100396.7, 100561,
  100970.4, 100911.7, 100853.2, 100787.9, 100704.9, 100605.1, 100484.9, 
    100343.3, 100194.8, 100060.8, 99967.59, 99934.23, 99965.34, 100093.2, 
    100302.1,
  100948.9, 100897.2, 100834.4, 100768.4, 100687, 100590.2, 100467.1, 
    100318.1, 100156.1, 99994.95, 99873.94, 99806.75, 99791.12, 99885.21, 
    100117.9,
  100931.3, 100887.5, 100826.8, 100764, 100686.9, 100595, 100478.9, 100330.3, 
    100169.5, 100016.2, 99899.98, 99836.05, 99796.23, 99852.23, 100063.9,
  101839.6, 101864.4, 101860.8, 101861.3, 101863.6, 101856, 101848.8, 
    101835.5, 101807.7, 101765.3, 101699.3, 101623.9, 101541.1, 101448.4, 
    101341.7,
  101852.4, 101868, 101866.8, 101863.8, 101856.5, 101857, 101843.3, 101829.4, 
    101806.6, 101771.9, 101718.1, 101651.3, 101578, 101490.3, 101385.5,
  101849.8, 101864.9, 101865.4, 101862.6, 101855.3, 101847.8, 101833.7, 
    101818.6, 101797.5, 101773.7, 101737.5, 101683, 101609.7, 101527.5, 
    101431.2,
  101841.2, 101852.8, 101848.6, 101835.3, 101815.2, 101800.6, 101790.1, 
    101777.8, 101762.6, 101743.9, 101718.6, 101682, 101629, 101558.1, 101470.4,
  101830.7, 101831.4, 101817.9, 101790.1, 101769, 101750.6, 101736.5, 
    101724.6, 101715.6, 101705.8, 101693.5, 101670.9, 101631.8, 101575.4, 
    101498,
  101816.7, 101812.1, 101785.9, 101750, 101722, 101692.7, 101675.3, 101659.1, 
    101650.5, 101643, 101634.3, 101626.3, 101605, 101572.4, 101514.9,
  101802.5, 101786.3, 101747.9, 101705.6, 101665.3, 101628.5, 101599.9, 
    101579.6, 101567.4, 101567.1, 101569.3, 101569.3, 101559.8, 101537.4, 
    101505.4,
  101786.8, 101759.4, 101712.1, 101658.1, 101606.1, 101553.2, 101510.8, 
    101483.1, 101468.3, 101470.1, 101477.7, 101485.3, 101487.7, 101487, 
    101470.1,
  101772, 101731.9, 101678.3, 101610.6, 101541.4, 101471.8, 101413.1, 
    101372.1, 101350.1, 101349.8, 101365.3, 101389, 101411.7, 101427.8, 
    101424.1,
  101758.6, 101708, 101645.5, 101566.1, 101480.9, 101393.6, 101316.9, 
    101260.6, 101230.7, 101231.2, 101253.3, 101285.8, 101324.3, 101352.5, 
    101359,
  102585, 102628.2, 102636, 102631.2, 102611.7, 102583.5, 102558.6, 102523.8, 
    102474.1, 102395.3, 102310.2, 102213.1, 102098.8, 101983.5, 101873.8,
  102607.4, 102651.9, 102673.1, 102679.9, 102666.4, 102642.2, 102610.8, 
    102581.5, 102528.2, 102454.7, 102365.7, 102266.7, 102149, 102022.3, 
    101904.1,
  102627.2, 102680.8, 102704.7, 102724.3, 102722, 102712.6, 102677.8, 
    102628.9, 102572.9, 102509.7, 102423.5, 102319.2, 102196.4, 102064.1, 
    101936.1,
  102652.7, 102694.7, 102721.4, 102742.8, 102751.4, 102746.4, 102730.1, 
    102693.3, 102629.8, 102557.3, 102474.9, 102369.2, 102245.7, 102103.4, 
    101968,
  102682.3, 102709.6, 102748.3, 102763, 102765, 102759.8, 102760.5, 102732.6, 
    102685, 102606, 102520.5, 102417.7, 102291.6, 102146.2, 102007.5,
  102704.1, 102730.1, 102764.1, 102768.7, 102782.9, 102780.1, 102773.6, 
    102751.3, 102716.3, 102653.3, 102564.1, 102462.6, 102333.7, 102185.8, 
    102038.1,
  102717.1, 102750, 102766.6, 102791.4, 102794.6, 102796.6, 102788.5, 
    102766.5, 102733.5, 102678.7, 102600.1, 102506.5, 102375.6, 102228.6, 
    102077,
  102720, 102762.8, 102769.6, 102797.2, 102804.3, 102796.7, 102794, 102776.8, 
    102749.7, 102700.7, 102628.9, 102545.3, 102420.3, 102270.8, 102113.1,
  102721.1, 102749.7, 102757.9, 102786.7, 102799, 102794.5, 102794.8, 
    102777.4, 102752.4, 102709.7, 102647.6, 102569.5, 102457, 102313.1, 
    102155.7,
  102711.3, 102730, 102747.8, 102764.8, 102774, 102784.9, 102789.2, 102768.7, 
    102747.2, 102709.5, 102655.4, 102586.5, 102484.2, 102352.3, 102197.4,
  102593.7, 102623.4, 102658, 102687.2, 102702.3, 102695.2, 102672.2, 
    102632.8, 102577.7, 102500.5, 102421.5, 102339.8, 102250.4, 102150, 
    102053.6,
  102612.5, 102650.5, 102678.4, 102714.4, 102747.4, 102755.2, 102732.8, 
    102679.7, 102619.9, 102547.4, 102469.2, 102387.7, 102293.1, 102189.1, 
    102084.3,
  102662.6, 102701.8, 102723.6, 102756.5, 102768.6, 102783.6, 102771.6, 
    102730.4, 102677.5, 102606.4, 102516.6, 102429.4, 102334.4, 102225.5, 
    102112.4,
  102723.9, 102749.8, 102771.4, 102796, 102815.5, 102813, 102808.6, 102781, 
    102717.8, 102648, 102564, 102472, 102370.3, 102257.2, 102139.6,
  102777.9, 102794.7, 102828.5, 102841.3, 102848.1, 102848.4, 102846, 
    102823.1, 102762.5, 102689.7, 102607.9, 102508.7, 102401, 102283.6, 
    102164.9,
  102799.3, 102828.6, 102860.1, 102880, 102893.3, 102894.1, 102877.7, 102855, 
    102811.9, 102731.3, 102643.8, 102540.4, 102429.6, 102301.1, 102190.6,
  102810.7, 102857.8, 102880.3, 102894.8, 102912.3, 102925.2, 102912.6, 
    102882.6, 102832.2, 102759.2, 102673.2, 102564.3, 102451.4, 102314.9, 
    102212,
  102820.7, 102862.9, 102894.3, 102920, 102933, 102937.4, 102934.1, 102911.1, 
    102858.9, 102784.5, 102695.4, 102580.3, 102467, 102327, 102217.3,
  102826.3, 102870.9, 102908.7, 102936.5, 102957.1, 102950.9, 102953.8, 
    102925, 102875.8, 102800.3, 102708.8, 102591.6, 102472.9, 102330.7, 
    102215.2,
  102821.2, 102874.8, 102920.5, 102952.4, 102957.1, 102959.6, 102961, 
    102930.5, 102879.3, 102808.8, 102715.5, 102598.3, 102470.6, 102335.4, 
    102212.9,
  102264.8, 102265.9, 102237.1, 102210.1, 102201, 102179.4, 102152.9, 
    102105.6, 102030.4, 101941.4, 101851.3, 101775.3, 101709.3, 101661.8, 
    101631.9,
  102305.8, 102306.6, 102262.6, 102225.1, 102201.5, 102199.4, 102179.6, 
    102146, 102055.3, 101947.3, 101843.9, 101760.4, 101693.7, 101644, 101616.4,
  102345.5, 102347.3, 102328.2, 102272.7, 102227.4, 102204.4, 102184.7, 
    102158.8, 102088.1, 101978.2, 101859.4, 101753, 101678.9, 101635.2, 
    101602.5,
  102372, 102376.1, 102365, 102330.6, 102281.5, 102240.8, 102208, 102170.7, 
    102117.1, 102010.4, 101878.7, 101756.8, 101669.4, 101624.9, 101588.3,
  102395.8, 102401.4, 102407.6, 102384.1, 102330.9, 102276.4, 102234.7, 
    102187.9, 102130.6, 102053.2, 101919.5, 101775, 101670.2, 101619.9, 
    101579.6,
  102406.4, 102435.2, 102440.5, 102425.4, 102394.8, 102334.6, 102278.1, 
    102225, 102150.4, 102072.1, 101962.4, 101821.3, 101688.8, 101621.6, 
    101568.1,
  102437.6, 102462, 102463.8, 102451.5, 102428.2, 102380.9, 102321.7, 
    102263.2, 102190.2, 102106.9, 101994.9, 101870.4, 101719.6, 101626.1, 
    101564.9,
  102455.8, 102488.5, 102495.8, 102484.2, 102450.6, 102408, 102361, 102299.3, 
    102222.7, 102137.8, 102025.5, 101910.4, 101760.9, 101642.1, 101564.8,
  102474.6, 102511.7, 102522, 102508.1, 102478.2, 102431, 102388.3, 102331.5, 
    102254.1, 102167.6, 102055.5, 101934.3, 101794.5, 101656.1, 101566.8,
  102496.3, 102531.1, 102541.3, 102540.4, 102511.6, 102456.6, 102409.5, 
    102355.1, 102276.2, 102186.7, 102076.6, 101953.8, 101820.3, 101668.7, 
    101570.9,
  102089.2, 102098.9, 102093.1, 102069.6, 102026.4, 101987.9, 101958.4, 
    101884.5, 101842.8, 101777.9, 101705.2, 101633.5, 101554.1, 101481.5, 
    101414,
  102138.1, 102141.4, 102135.9, 102105.8, 102060, 102015, 101967.2, 101911.5, 
    101840.8, 101776.4, 101716.5, 101648.6, 101585.3, 101511.4, 101447.2,
  102157.9, 102171.8, 102163.9, 102138.7, 102076.7, 102030.4, 101978.4, 
    101914.2, 101847.1, 101793.1, 101737.4, 101669.6, 101601.1, 101533.3, 
    101483.5,
  102187.9, 102204.3, 102196.9, 102180.8, 102117.3, 102057, 101991.8, 
    101924.7, 101850.2, 101797.7, 101740.1, 101683, 101616, 101558.1, 101512.9,
  102226.7, 102238.4, 102228.3, 102202.9, 102150.3, 102075.6, 102007.7, 
    101939.5, 101859.2, 101798.3, 101743.7, 101695.6, 101632.1, 101576, 
    101532.3,
  102258.4, 102267.8, 102263.8, 102234.3, 102186.1, 102100.3, 102022, 
    101945.3, 101864.9, 101800.9, 101738.4, 101696.3, 101638.2, 101597, 
    101542.5,
  102285.1, 102287, 102289.1, 102262.1, 102220.9, 102130.8, 102044.8, 
    101956.7, 101873.9, 101803.2, 101739.9, 101700, 101641.6, 101623.1, 
    101552.3,
  102324.1, 102330.4, 102323.3, 102292.4, 102249.8, 102162.6, 102066.7, 
    101966.4, 101879.6, 101807.2, 101747.2, 101687.9, 101647.7, 101622.9, 
    101562.7,
  102353, 102358.3, 102353.1, 102323.7, 102272.1, 102196.2, 102093, 101985.4, 
    101890.2, 101809.8, 101739.1, 101682.9, 101641.3, 101608.8, 101571.3,
  102389.3, 102395.9, 102386.7, 102357, 102298.5, 102223.8, 102123.5, 
    102009.1, 101901.8, 101807.4, 101729.1, 101673.1, 101615.6, 101599.3, 
    101567.6,
  102291.9, 102317.8, 102353.6, 102368.2, 102361.4, 102344.1, 102310.4, 
    102266.7, 102205.4, 102127.2, 102043.4, 101925.4, 101830.8, 101745.3, 
    101704.2,
  102349, 102371.5, 102403.7, 102409.5, 102406, 102389.9, 102356.1, 102313.3, 
    102254.3, 102162.2, 102075.6, 101955, 101860.1, 101749.7, 101692.2,
  102386.2, 102415, 102449.4, 102460.3, 102461.4, 102438.3, 102404.7, 
    102353.9, 102297.5, 102216.3, 102118.7, 101992, 101886.8, 101752.6, 
    101687.4,
  102438.2, 102469.4, 102498.8, 102518.3, 102512.8, 102485.6, 102447.8, 
    102394.7, 102333.7, 102259.8, 102163.9, 102037.5, 101918.5, 101776, 
    101692.9,
  102475, 102510.7, 102551.3, 102562.5, 102558, 102524.4, 102485.8, 102430.6, 
    102367.3, 102291.6, 102203.1, 102082.3, 101961.7, 101810.7, 101698.8,
  102519.9, 102565.3, 102596, 102606.1, 102597.7, 102562.9, 102514.4, 
    102462.4, 102393.7, 102320.2, 102233.4, 102112.9, 101991.6, 101840.4, 
    101710,
  102564.5, 102602.7, 102630.1, 102639.2, 102629.3, 102595.2, 102542.8, 
    102487.4, 102419.2, 102345.3, 102257.9, 102141.2, 102017.3, 101868.6, 
    101724.2,
  102599.7, 102640.4, 102670.6, 102675.5, 102658.1, 102620.9, 102568.1, 
    102507.1, 102437.4, 102363.2, 102281.3, 102171.3, 102044, 101906.1, 
    101752.5,
  102633.1, 102674.9, 102691.3, 102697.4, 102679.7, 102639.2, 102584.4, 
    102520.5, 102450.5, 102385.5, 102309.3, 102204.7, 102086.3, 101949.8, 
    101799.2,
  102655.6, 102704, 102718.4, 102723, 102692.4, 102649.3, 102590.2, 102527.6, 
    102459.9, 102396.9, 102324.9, 102239, 102129.2, 101999.7, 101858.1,
  102482.8, 102519.1, 102548.9, 102571.2, 102589.1, 102601.6, 102605.4, 
    102597, 102577.5, 102546.1, 102506.9, 102458.6, 102405.4, 102350.6, 
    102279.5,
  102556.6, 102588.4, 102616, 102639.4, 102656.7, 102667.8, 102669.1, 102659, 
    102641.2, 102606.1, 102560.8, 102505.3, 102443.4, 102385.8, 102314,
  102624.6, 102655, 102684, 102709.5, 102724.8, 102736.9, 102733.2, 102720.2, 
    102695.9, 102659.8, 102612.9, 102551.3, 102484.9, 102416.6, 102340.5,
  102693.4, 102721, 102749.1, 102772.7, 102791.9, 102799.9, 102799.1, 
    102785.5, 102757.8, 102715.8, 102661.8, 102592.5, 102525.4, 102448.6, 
    102364.9,
  102755.2, 102782.9, 102816.4, 102841.2, 102855.1, 102866, 102863.5, 
    102844.4, 102812.5, 102764.4, 102708.9, 102634.4, 102561.8, 102478.7, 
    102389.5,
  102813.8, 102850, 102881.2, 102901.5, 102916.4, 102921.6, 102919.6, 
    102899.5, 102865.1, 102814.5, 102752.9, 102673.5, 102591.5, 102505.7, 
    102412,
  102874.1, 102911.3, 102944.5, 102965.3, 102980.2, 102983.9, 102974.8, 
    102950, 102910.9, 102858.5, 102791.5, 102711.1, 102619.2, 102526.5, 102426,
  102928, 102977.1, 102998.2, 103020.2, 103029.6, 103031.6, 103020.6, 
    102995.3, 102953.2, 102896.4, 102827.3, 102741.7, 102642.1, 102538.1, 
    102435.5,
  102978.6, 103025.1, 103042.7, 103058.5, 103065.5, 103065.8, 103057.1, 
    103034.2, 102988.6, 102928.8, 102857.3, 102768.6, 102661.8, 102546.1, 
    102433.5,
  103022.4, 103053.1, 103070, 103085.6, 103093.7, 103094.8, 103079.8, 
    103058.8, 103016.7, 102958.3, 102881.1, 102793.1, 102680.5, 102552.6, 
    102427.9,
  102038.8, 102111.7, 102171.4, 102213.6, 102246.1, 102266.5, 102271.9, 
    102264.5, 102254.9, 102236.2, 102206.3, 102174, 102128.4, 102072.1, 
    102005.8,
  102124.8, 102179.7, 102231.1, 102273.4, 102303.4, 102319.4, 102325.5, 
    102320.3, 102305.4, 102280.8, 102242.5, 102201.6, 102149.6, 102087.3, 
    102014.6,
  102201.9, 102254.3, 102305.9, 102337.5, 102363.8, 102376.9, 102379.9, 
    102370, 102350.5, 102322.3, 102278.9, 102226.2, 102161.2, 102084.8, 
    101996.6,
  102291.4, 102331.4, 102375.2, 102398, 102423.2, 102431.2, 102433.9, 102422, 
    102398, 102364.6, 102317.8, 102252.7, 102174.3, 102085.6, 101982.5,
  102380, 102407.8, 102448.2, 102463.5, 102484.9, 102491.5, 102493, 102476.5, 
    102448.9, 102404.7, 102348.3, 102276.9, 102184.8, 102079.7, 101958.8,
  102468.2, 102486, 102521.6, 102529, 102549.1, 102548.3, 102545.6, 102527, 
    102495.8, 102451, 102385.2, 102297.7, 102195, 102073.4, 101936.5,
  102549.1, 102561.6, 102589.8, 102594.6, 102610.1, 102606, 102601.7, 
    102580.5, 102542.6, 102489.9, 102414.8, 102322.1, 102203, 102069.5, 
    101913.2,
  102622.6, 102629.4, 102653.3, 102654.8, 102666.7, 102662.2, 102652.8, 
    102633.6, 102593.4, 102531.2, 102445.9, 102343.6, 102212.2, 102064.8, 
    101893,
  102689.4, 102692.2, 102707, 102701, 102706.4, 102699.6, 102691, 102670.9, 
    102634.1, 102574, 102481.9, 102363.5, 102223.5, 102061, 101882,
  102743.5, 102742.1, 102755, 102749.6, 102752.1, 102741.5, 102731.3, 
    102705.4, 102666.8, 102606, 102514.2, 102389.4, 102238.5, 102058.5, 
    101874.2,
  101073.3, 101112.8, 101184.6, 101275.3, 101372.3, 101468, 101541.2, 
    101600.4, 101629.2, 101639.6, 101632.1, 101650.4, 101664, 101680.9, 
    101719.4,
  101142.6, 101183.4, 101235.7, 101315.3, 101405.6, 101488.6, 101558.8, 
    101620.4, 101639.7, 101648.5, 101631.9, 101642.5, 101664.3, 101691.9, 
    101719,
  101238.1, 101267, 101303, 101369.3, 101450.7, 101523.1, 101576.1, 101639.3, 
    101657.2, 101648.2, 101629.6, 101639.2, 101651.9, 101677, 101706.3,
  101336.1, 101360.6, 101386.6, 101439.7, 101504.4, 101559.9, 101599.1, 
    101657.5, 101668.9, 101647.6, 101622.1, 101629.4, 101633.7, 101653.4, 
    101679.7,
  101433.4, 101456.7, 101475.8, 101512.9, 101555.7, 101599.1, 101627.6, 
    101668.6, 101674.7, 101646, 101615.5, 101613.9, 101609.7, 101629.4, 
    101654.1,
  101530.5, 101552.4, 101564.2, 101591.9, 101623.4, 101652.1, 101659.9, 
    101688.3, 101678.4, 101640.4, 101605.3, 101588.8, 101577.5, 101590.4, 
    101614.6,
  101624.1, 101638.7, 101652.8, 101673.9, 101687.6, 101700.4, 101696.4, 
    101707.1, 101690.9, 101638.7, 101593.5, 101564.1, 101546.2, 101549.1, 
    101565,
  101726.9, 101733, 101739.1, 101749, 101751.7, 101747.8, 101733.8, 101727.6, 
    101694.8, 101633.8, 101577, 101533.9, 101509.4, 101499.9, 101509.7,
  101832.8, 101826.7, 101829.9, 101822.4, 101811.3, 101791.2, 101766.7, 
    101744.9, 101701, 101631.5, 101562.4, 101503.3, 101469.6, 101447.4, 
    101440.7,
  101936.2, 101915.4, 101910.2, 101892.6, 101868.5, 101835, 101797.2, 
    101760.6, 101707.3, 101626.4, 101546.9, 101470.3, 101425.4, 101390, 
    101370.6,
  100830.1, 100895.9, 100997.3, 101120.2, 101252.2, 101370.8, 101480.9, 
    101584.9, 101678.8, 101776.4, 101866.8, 101948, 102020.8, 102095.5, 102158,
  100805.8, 100877.8, 100979.1, 101102.5, 101233.4, 101352.1, 101464.8, 
    101569.6, 101667.1, 101769.9, 101864.9, 101954.1, 102026.8, 102107, 
    102176.6,
  100800.9, 100871.1, 100955.6, 101082, 101216.8, 101332.8, 101444.1, 
    101557.8, 101653.3, 101758.2, 101853.5, 101941.6, 102016.2, 102096.2, 
    102170.7,
  100798.2, 100863.5, 100943.3, 101064.6, 101200, 101315.5, 101421.6, 
    101536.2, 101629.6, 101737.5, 101833.3, 101922.5, 102002.4, 102084, 
    102161.9,
  100782.6, 100847.8, 100932.7, 101047.6, 101175.8, 101299.3, 101395.9, 
    101512.8, 101603.2, 101708.8, 101807.1, 101895.2, 101974.4, 102055.6, 
    102135,
  100761.4, 100837.1, 100918, 101039.9, 101155.1, 101279.2, 101366.6, 
    101481.5, 101568.8, 101673.9, 101770.7, 101858.9, 101938.9, 102020.2, 
    102099.3,
  100731.4, 100819.4, 100890.8, 101025.9, 101129.4, 101258.2, 101334.1, 
    101449, 101530.7, 101631.4, 101725.5, 101813.3, 101893, 101972.8, 102049.6,
  100702.4, 100804.2, 100858, 101003.8, 101103, 101235, 101300.8, 101411, 
    101483.6, 101580.5, 101671.1, 101756.8, 101834.1, 101913.1, 101990.8,
  100703.8, 100798, 100829.1, 100975.5, 101073.7, 101203, 101263.8, 101366.3, 
    101436.5, 101524.5, 101610.7, 101691.2, 101765.8, 101841.4, 101914.6,
  100750.1, 100803.9, 100816.7, 100945.9, 101052, 101169.9, 101228.4, 
    101315.2, 101383.6, 101459.5, 101542.1, 101617.5, 101686.5, 101759.4, 
    101829.4,
  101414, 101540.4, 101668.3, 101792.9, 101902.4, 102006.6, 102104.4, 
    102197.9, 102284, 102368.6, 102444.3, 102518.9, 102585.6, 102650.3, 
    102705.5,
  101418, 101544.9, 101678.1, 101799.1, 101910.2, 102014.6, 102112.3, 
    102206.8, 102294.8, 102381, 102463.6, 102543.2, 102613.5, 102681.1, 
    102742.8,
  101433.7, 101552.6, 101683, 101802, 101912.5, 102017.1, 102117.2, 102211.5, 
    102301.1, 102388.7, 102476.6, 102557.1, 102634.3, 102706, 102770.1,
  101449.1, 101561.8, 101686.8, 101802.6, 101913.7, 102016, 102115.5, 
    102210.5, 102299.2, 102390.7, 102478.3, 102562.3, 102643.3, 102718.3, 
    102786,
  101464.6, 101565.4, 101687.2, 101798.4, 101911.5, 102012.4, 102109.2, 
    102204.2, 102293.8, 102383.3, 102473.5, 102558.4, 102640.1, 102719, 
    102792.6,
  101469.7, 101568.1, 101684.2, 101790.5, 101900.9, 102002.3, 102097, 
    102191.8, 102282.2, 102374.6, 102460.8, 102546.3, 102630.2, 102710.1, 
    102787.2,
  101463.7, 101563, 101672.4, 101777.4, 101885.2, 101985.5, 102076.1, 
    102171.3, 102261.5, 102353.7, 102441.9, 102525.3, 102606.4, 102687.8, 
    102765.9,
  101443.1, 101548.1, 101652.4, 101757.9, 101860.4, 101963.6, 102050.9, 
    102144, 102234.4, 102326.2, 102412.6, 102494.1, 102574.3, 102653, 102730.3,
  101403.2, 101522.8, 101621.8, 101732.7, 101826.9, 101934.5, 102018.6, 
    102110.6, 102198.1, 102287.7, 102372.4, 102452.7, 102528.3, 102604.9, 
    102679.3,
  101346.7, 101487.4, 101580.1, 101700, 101786.7, 101898.1, 101980.5, 
    102074.2, 102156.1, 102242.7, 102320.2, 102399.1, 102473.4, 102547.4, 
    102619.2,
  101499.7, 101625.4, 101749.4, 101861.6, 101967.2, 102061.5, 102154.3, 
    102244.8, 102330.8, 102412, 102489.2, 102561.9, 102629.3, 102691.1, 
    102747.8,
  101535.8, 101638.4, 101767.8, 101873.5, 101980.6, 102075.2, 102169.2, 
    102258.2, 102346.4, 102428.7, 102509.9, 102584.3, 102654.3, 102719.3, 
    102781.5,
  101538.5, 101640.5, 101772.1, 101875.5, 101985.4, 102080.5, 102174.2, 
    102262.8, 102352.8, 102436.1, 102519, 102596.3, 102669.1, 102737.9, 
    102805.7,
  101566.4, 101656.8, 101778.8, 101884.9, 101988.8, 102082.9, 102174.9, 
    102263.9, 102353.2, 102436.6, 102519.9, 102597, 102672.5, 102745.1, 
    102817.3,
  101574.9, 101669.4, 101777.4, 101885.3, 101984.4, 102079.6, 102168.2, 
    102256.3, 102343.5, 102426.6, 102507.3, 102586.6, 102663, 102738.6, 
    102811.7,
  101575.4, 101686.3, 101775.5, 101885.8, 101973.8, 102070.2, 102152.4, 
    102239.9, 102322.6, 102406.6, 102484, 102563.5, 102638.6, 102716.6, 
    102789.9,
  101580.1, 101690.6, 101767.1, 101879.3, 101957, 102055.8, 102129.2, 
    102214.8, 102292.3, 102373.7, 102448.1, 102524.3, 102599.5, 102676.3, 
    102748.4,
  101575.2, 101683.4, 101757.5, 101866.4, 101933.4, 102033, 102098.6, 
    102182.4, 102252, 102329, 102398.8, 102471.1, 102542.7, 102616.9, 102688.5,
  101565.2, 101670.8, 101744.4, 101845.9, 101908.3, 102004.2, 102063.2, 
    102142.1, 102204.8, 102273.1, 102336.2, 102404.6, 102472.1, 102542.8, 
    102609.1,
  101546.4, 101653.8, 101728.9, 101821.7, 101879.7, 101965.1, 102024.2, 
    102095, 102147.4, 102208.9, 102264.4, 102325.6, 102387.1, 102452.2, 
    102517.9,
  101328.9, 101441.1, 101544.4, 101640.5, 101730.6, 101826.6, 101919.1, 
    102013.2, 102104.4, 102194.3, 102283.2, 102367.5, 102447.5, 102525.1, 
    102597.1,
  101306.9, 101411.4, 101514.1, 101609, 101700, 101793.2, 101886.3, 101979.8, 
    102073.1, 102164.9, 102255.2, 102345.2, 102430.9, 102514, 102592.4,
  101264.1, 101370.5, 101480.5, 101568.9, 101661.1, 101750.2, 101845.3, 
    101939.9, 102036, 102130.5, 102222.9, 102314.7, 102406.3, 102495.7, 
    102579.6,
  101238.3, 101336.8, 101449.7, 101531.2, 101624.3, 101708.2, 101800.7, 
    101895.6, 101989.8, 102084.8, 102180.4, 102273.7, 102368.8, 102463, 
    102553.3,
  101212.1, 101301.3, 101413, 101493, 101580.5, 101661.9, 101749.5, 101842.1, 
    101939.3, 102034.7, 102132.2, 102228.6, 102325.1, 102421.6, 102518,
  101184.7, 101278, 101378.7, 101457.3, 101536.7, 101613.3, 101697.3, 
    101787.3, 101881.8, 101978.5, 102077.1, 102177.4, 102276.4, 102374.9, 
    102471.6,
  101159, 101255.2, 101343.8, 101420.6, 101493, 101563.7, 101641, 101728.5, 
    101823.3, 101917.4, 102017.4, 102117.4, 102219, 102322.5, 102423.7,
  101147.6, 101232.1, 101312, 101384.8, 101450.6, 101515.6, 101586.7, 
    101667.9, 101761.2, 101855.8, 101955.3, 102055.5, 102157.9, 102262.9, 
    102367.2,
  101137, 101208.5, 101281, 101347.9, 101406.7, 101467.8, 101533.1, 101609.4, 
    101698.1, 101791.8, 101890.8, 101989.9, 102092.9, 102196.9, 102305.7,
  101125.3, 101190.5, 101253.1, 101315.7, 101366.4, 101421.8, 101482.1, 
    101553, 101635.3, 101728.5, 101825.9, 101925.2, 102026.7, 102129.4, 
    102237.5,
  101246.7, 101340.7, 101434.9, 101534.8, 101633.8, 101735.5, 101830.8, 
    101920.8, 102008.2, 102091.8, 102172.1, 102251, 102327.1, 102403.3, 
    102469.6,
  101189.8, 101288.7, 101386.6, 101489.9, 101590.1, 101694.7, 101796.9, 
    101892.2, 101985.3, 102072, 102154.8, 102236.7, 102314.8, 102394.4, 
    102466.1,
  101125.3, 101224.9, 101326, 101429, 101536.4, 101644.7, 101756, 101855.9, 
    101956.4, 102046.9, 102132.6, 102218.5, 102297.7, 102379, 102454.1,
  101068.3, 101169.7, 101272.3, 101376.7, 101487.7, 101597.4, 101713.9, 
    101819.6, 101922.9, 102021.8, 102107.8, 102195.5, 102276.1, 102360, 
    102439.6,
  101010, 101112.5, 101216.3, 101320.1, 101431.7, 101545.6, 101661.6, 
    101780.4, 101884, 101988.4, 102077.4, 102167.8, 102252, 102337.3, 102419.2,
  100954, 101061.3, 101165.2, 101269.3, 101380.1, 101498.8, 101612.4, 
    101735.3, 101843.5, 101951.6, 102044.8, 102135.8, 102223, 102310.8, 
    102394.5,
  100896.8, 101007.6, 101118.7, 101220.7, 101332.1, 101449.1, 101564.9, 
    101686.2, 101798.6, 101911, 102006.9, 102099.8, 102189.3, 102279.9, 
    102365.4,
  100840, 100955.1, 101074.5, 101178.6, 101286.9, 101405, 101520.4, 101640.6, 
    101753.9, 101865.4, 101967.5, 102060.5, 102151.1, 102243.1, 102331.6,
  100782.5, 100905.5, 101031.5, 101139, 101246.8, 101362.6, 101477.4, 
    101596.2, 101708.4, 101820.8, 101923.5, 102019, 102110.7, 102201.9, 
    102291.3,
  100728.4, 100862, 100990.7, 101102.5, 101211.8, 101325.9, 101437.8, 
    101554.9, 101666.6, 101774.4, 101879.5, 101974.1, 102064.8, 102154, 
    102244.8,
  101384.1, 101464.7, 101543.6, 101620.7, 101700, 101775.8, 101851.8, 
    101923.4, 101996.8, 102069.1, 102140.5, 102206.4, 102269.6, 102331.4, 
    102388.6,
  101309.3, 101387, 101466.6, 101547.7, 101629.7, 101708.6, 101789.2, 
    101865.2, 101942, 102018.7, 102092.9, 102164.3, 102231.9, 102298.2, 
    102360.4,
  101213.1, 101293.8, 101377.5, 101460.8, 101546, 101630.7, 101713.9, 
    101795.9, 101877.5, 101960.8, 102037.8, 102113.8, 102186.6, 102255.7, 
    102319.2,
  101118.6, 101199.8, 101284.5, 101370.6, 101453.6, 101543.3, 101626.4, 
    101714.7, 101800.4, 101887.6, 101968.6, 102049.8, 102127.5, 102200.3, 
    102267.6,
  101020.7, 101099.2, 101184, 101268.6, 101353.7, 101441.9, 101530.2, 
    101619.6, 101709.5, 101799.7, 101887.6, 101973.2, 102057, 102135.1, 
    102206.8,
  100920.2, 101000.4, 101085.6, 101166.9, 101250.7, 101334.6, 101421.5, 
    101511, 101604.2, 101699.1, 101793.2, 101887.6, 101976.7, 102060.8, 
    102135.9,
  100814.1, 100899.4, 100984.1, 101064.6, 101143.9, 101224, 101307.9, 
    101394.2, 101486.7, 101585.5, 101681.8, 101783.6, 101878.2, 101968.5, 
    102050.4,
  100704.6, 100796.1, 100881.6, 100963.6, 101041.3, 101116.1, 101191.1, 
    101276.5, 101360.9, 101458.8, 101559.2, 101663.8, 101765.7, 101863.3, 
    101952.5,
  100586.1, 100688, 100779.9, 100862.3, 100939.9, 101008.6, 101078.8, 
    101151.5, 101235.4, 101324.8, 101423.4, 101526.9, 101633.8, 101739, 
    101836.2,
  100479.9, 100580.5, 100682.5, 100767, 100845.2, 100909.1, 100973.8, 
    101038.8, 101108.3, 101190.1, 101286.6, 101382.1, 101491, 101599.3, 
    101705.8,
  101221.4, 101270.8, 101316, 101368.3, 101419.8, 101472, 101522.3, 101573.1, 
    101621.3, 101664, 101703.3, 101741.8, 101791.3, 101854.2, 101923.7,
  101128.6, 101176.9, 101223.3, 101279.1, 101332.8, 101388.9, 101443.9, 
    101498.8, 101551, 101596, 101636.8, 101674, 101720.6, 101783.2, 101854.7,
  101012.2, 101064.9, 101111.5, 101175.4, 101237, 101301.1, 101360.6, 
    101420.1, 101475.5, 101524.9, 101564.7, 101599.7, 101641.7, 101696.7, 
    101770.5,
  100897, 100947.5, 100995.8, 101057, 101121.6, 101193.3, 101262.1, 101331.3, 
    101394.4, 101453.7, 101499.6, 101535.2, 101572.6, 101619, 101691.3,
  100778.5, 100820.9, 100869.1, 100930.9, 100999, 101075, 101152, 101229.8, 
    101303.3, 101369.1, 101427.2, 101473, 101509.4, 101548.4, 101613.1,
  100672, 100708.6, 100750.2, 100804.9, 100868.8, 100945.5, 101028, 101115.4, 
    101201.2, 101280.8, 101351.8, 101411.6, 101459.3, 101501.5, 101550.4,
  100566.9, 100606.6, 100645.5, 100700.1, 100755.5, 100826.3, 100903.1, 
    100992, 101087.8, 101182.8, 101267.9, 101344.1, 101408.4, 101460.5, 
    101507.3,
  100475.7, 100514, 100547.5, 100599, 100656.1, 100725.7, 100797.8, 100879.4, 
    100967.6, 101070.9, 101175, 101267.3, 101347.3, 101423.2, 101483,
  100411.1, 100440.3, 100468.5, 100518.2, 100570.8, 100641.6, 100715.3, 
    100787.8, 100867.1, 100958.7, 101065.7, 101176.7, 101274.1, 101359.9, 
    101436.4,
  100356.3, 100383.8, 100408.9, 100453.6, 100506.1, 100568.3, 100644.9, 
    100726.1, 100797.7, 100867.1, 100956.5, 101068.5, 101184.4, 101288.5, 
    101381.6,
  101275.6, 101291.1, 101308.7, 101327.7, 101343.1, 101364.5, 101385.7, 
    101412, 101422.4, 101444.6, 101478.4, 101545.7, 101646.5, 101780.1, 
    101914.6,
  101252.3, 101269.6, 101285.6, 101302.6, 101321.2, 101350, 101383.2, 
    101412.2, 101432, 101460.3, 101491.8, 101551.6, 101645.5, 101760.8, 
    101890.1,
  101228.8, 101244.5, 101259.3, 101278, 101305.5, 101340.3, 101379.6, 
    101422.3, 101462.2, 101494.8, 101527.3, 101569.6, 101641.8, 101747.1, 
    101866.3,
  101211.8, 101218.6, 101235.1, 101252.6, 101278.4, 101315.3, 101363.4, 
    101411.5, 101461.2, 101508.5, 101553, 101599.6, 101657.3, 101749.8, 
    101852.1,
  101215.2, 101209.3, 101213, 101229.9, 101257.4, 101285.4, 101335.7, 
    101389.8, 101450.2, 101504.8, 101558.9, 101611.2, 101668.3, 101743.5, 
    101840.4,
  101212.6, 101219.7, 101221, 101224.5, 101234.6, 101250.9, 101291.8, 
    101343.5, 101406, 101472.4, 101537.6, 101599.7, 101662.3, 101739.7, 
    101825.5,
  101192.9, 101212.7, 101213.9, 101226.7, 101231.3, 101239.1, 101254.9, 
    101289.6, 101347.1, 101414.2, 101488.5, 101562.6, 101635.6, 101712, 
    101797.9,
  101173.8, 101184.2, 101187.2, 101204, 101212.9, 101232, 101236.8, 101250.9, 
    101284.7, 101345, 101422.5, 101506.2, 101590.2, 101673.8, 101760.2,
  101157.4, 101163.4, 101170.4, 101182.5, 101199.2, 101217.6, 101233.5, 
    101235.8, 101242.6, 101279.8, 101350, 101439, 101535.1, 101622.9, 101714.9,
  101140.5, 101143, 101151.5, 101162.2, 101179.2, 101199.4, 101216, 101235.2, 
    101234.8, 101242.6, 101284.9, 101366.7, 101472.6, 101571.3, 101667.1,
  101342.7, 101398.6, 101454.9, 101513.5, 101577.2, 101641.8, 101704.5, 
    101772.9, 101841.3, 101911.8, 101983.6, 102061.5, 102138.7, 102211.7, 
    102284.2,
  101335.2, 101381.2, 101435.4, 101497.5, 101556.9, 101618.1, 101679.9, 
    101746.1, 101813.8, 101888.6, 101961.4, 102035.5, 102108.6, 102183.1, 
    102255,
  101329.2, 101379.8, 101416.3, 101469.8, 101522.4, 101579.4, 101642.6, 
    101709, 101777.8, 101851.9, 101923.8, 101997.8, 102071.8, 102143, 102212.1,
  101341.9, 101377.6, 101403.6, 101453.4, 101492.8, 101540.3, 101599.2, 
    101665.8, 101736.8, 101810.6, 101885.5, 101958.2, 102029.4, 102097.1, 
    102165,
  101364.1, 101377, 101388.6, 101439.1, 101455.1, 101500.5, 101550.3, 
    101616.3, 101691.1, 101765, 101838.3, 101908.9, 101978, 102043.2, 102108.5,
  101378.6, 101417.5, 101399.4, 101418, 101430, 101460.8, 101504, 101562, 
    101639.8, 101714.8, 101789, 101858.6, 101925.6, 101985.6, 102046.6,
  101384.4, 101410.4, 101401.5, 101410.3, 101406.5, 101426.4, 101459.8, 
    101511.9, 101582.3, 101658.8, 101732.7, 101798.4, 101862.1, 101920.8, 
    101976.5,
  101397, 101411.1, 101400.7, 101408.9, 101395.1, 101406.3, 101420.7, 
    101464.4, 101528, 101600.3, 101672.4, 101736.7, 101795.1, 101851.3, 
    101903.8,
  101409.1, 101412.3, 101404.6, 101401.2, 101393.5, 101394.8, 101398.8, 
    101426.5, 101472.8, 101538.7, 101609.4, 101670.7, 101725.3, 101776.7, 
    101825.5,
  101424.1, 101417.5, 101407.8, 101400.5, 101394.7, 101392.9, 101380, 101398, 
    101429.3, 101480.6, 101543.7, 101602.8, 101653.1, 101698.5, 101740,
  101678.4, 101737.6, 101795.1, 101855, 101914.5, 101975.8, 102033, 102087.3, 
    102142.9, 102193.4, 102243.8, 102293.8, 102338.2, 102380.8, 102419,
  101617.3, 101677.3, 101737.5, 101799.3, 101863.3, 101925, 101981.2, 
    102035.6, 102088.7, 102140.8, 102188.2, 102236.9, 102279.7, 102320.6, 
    102356.3,
  101549, 101609.6, 101671.5, 101733.8, 101799.6, 101863.2, 101920.6, 
    101977.3, 102029.3, 102079.2, 102124.3, 102170, 102213.3, 102252.9, 
    102286.6,
  101474.2, 101532.7, 101599.2, 101666.4, 101732.2, 101799.2, 101859, 
    101913.7, 101965.9, 102012.8, 102059.5, 102101.2, 102141.8, 102180.2, 
    102212.5,
  101396.4, 101452.3, 101515.4, 101585.8, 101655.5, 101725.1, 101787.5, 
    101842.6, 101896.7, 101942.8, 101987.6, 102027.8, 102065.5, 102100.2, 
    102130.4,
  101310.9, 101368, 101427.9, 101501, 101575.3, 101646.6, 101713.1, 101769, 
    101822, 101868.7, 101913.4, 101953.4, 101987, 102018.5, 102044,
  101223.1, 101278.8, 101340.3, 101409.6, 101486.7, 101561.8, 101631.5, 
    101690.4, 101743.3, 101788.8, 101832.9, 101871.5, 101904, 101931.1, 
    101950.9,
  101138.9, 101196.4, 101254, 101318.7, 101393.8, 101472.6, 101543.8, 
    101607.9, 101658.7, 101704.9, 101745.8, 101785.5, 101814.4, 101836.5, 
    101848,
  101053.5, 101114.9, 101171.6, 101231.9, 101302.6, 101377.5, 101453.5, 
    101519.5, 101572.7, 101618, 101656.2, 101690.5, 101718, 101735.6, 101743.1,
  100966.4, 101031.7, 101097.1, 101151.1, 101213.1, 101285.5, 101358.7, 
    101429.4, 101482.8, 101528.1, 101563.9, 101595.6, 101619.3, 101631.7, 
    101638.3,
  101919, 101917, 101921.4, 101919.7, 101920, 101924.1, 101929, 101930.4, 
    101931.9, 101935.9, 101941.4, 101952.1, 101964.5, 101981.3, 101999.8,
  101872.9, 101871.8, 101873.8, 101873.1, 101871.2, 101868.7, 101861.3, 
    101853.5, 101848.9, 101847.2, 101845.2, 101853.3, 101864.7, 101881, 
    101900.4,
  101829.7, 101825.7, 101820.3, 101813.5, 101804.5, 101793.6, 101778.4, 
    101763.6, 101751.1, 101743, 101743.6, 101750.6, 101759.2, 101774.5, 
    101796.4,
  101776.8, 101769.3, 101766.3, 101754.3, 101739.7, 101718.4, 101696.6, 
    101673.9, 101654.2, 101643.9, 101640.2, 101639.5, 101648.6, 101662.7, 
    101681.6,
  101722.1, 101712.5, 101703.4, 101686.3, 101663.2, 101635.7, 101607.8, 
    101578.4, 101555, 101541.5, 101531.1, 101533, 101538.9, 101551, 101567.2,
  101662.3, 101650.2, 101636.3, 101613.8, 101584.2, 101552.2, 101517.4, 
    101483, 101456.3, 101437.7, 101427.1, 101424.1, 101425.5, 101432.2, 
    101444.2,
  101599.3, 101583.1, 101565, 101536, 101502, 101465.6, 101424.1, 101385.9, 
    101357.2, 101334, 101319.2, 101308.4, 101303.9, 101304.5, 101313.6,
  101532.2, 101511.6, 101486.8, 101456.8, 101417.6, 101375.4, 101329.8, 
    101289.4, 101256.6, 101230.1, 101207.4, 101190.4, 101178.7, 101174.8, 
    101177.6,
  101461.7, 101436.7, 101410.8, 101373.8, 101331.4, 101282.3, 101234.2, 
    101189.1, 101150.2, 101118.7, 101090.1, 101066.7, 101049.9, 101037.5, 
    101033.3,
  101384.5, 101358.7, 101325.1, 101288.7, 101242, 101190.6, 101135.3, 
    101085.3, 101044.1, 101006.9, 100975.7, 100944.5, 100920.2, 100900.5, 
    100885.9,
  101332.5, 101306.6, 101287.8, 101268.8, 101262.3, 101260.9, 101261.9, 
    101279.9, 101305.1, 101335.4, 101370.5, 101410.7, 101456.8, 101507.1, 
    101562.2,
  101290.6, 101249.4, 101222, 101193.5, 101180.3, 101167.4, 101164.8, 
    101178.6, 101198.3, 101223.9, 101255.7, 101290.6, 101330.6, 101377, 
    101430.1,
  101240.4, 101190.2, 101154, 101114.1, 101090.8, 101066.5, 101063.9, 
    101069.9, 101082.5, 101101.7, 101122.8, 101150, 101187.1, 101230.9, 
    101281.1,
  101191.3, 101131.9, 101085.5, 101033.8, 100996.7, 100961.1, 100954.4, 
    100952.5, 100959.9, 100968.5, 100979.8, 100999.4, 101029.6, 101065.4, 
    101111.2,
  101140.5, 101070.2, 101009.7, 100946.9, 100898.1, 100859.5, 100844, 
    100832.4, 100829.3, 100822.8, 100824.5, 100834.3, 100854.1, 100883.2, 
    100922.5,
  101089.8, 101007.5, 100935, 100861.8, 100801.5, 100752.1, 100726, 100705.9, 
    100689.6, 100671.1, 100662.1, 100659.8, 100668.6, 100688.2, 100718.7,
  101039.5, 100945.2, 100859.5, 100774.4, 100701.5, 100642, 100604.9, 
    100573.9, 100542.1, 100512, 100489, 100476.1, 100473.4, 100483, 100504.8,
  100990.7, 100882.4, 100784.5, 100687.9, 100600.9, 100534.4, 100485.3, 
    100442.3, 100397.3, 100355.7, 100321.4, 100292.9, 100279.9, 100278, 100289,
  100945.4, 100821.6, 100711.3, 100599.8, 100502.3, 100427.9, 100364.4, 
    100308.7, 100248.6, 100197.4, 100145.4, 100108.1, 100081.3, 100069.8, 
    100072.4,
  100902, 100763.5, 100639.3, 100515.2, 100409.6, 100323.9, 100250, 100182.3, 
    100109.3, 100039.7, 99979.41, 99925.99, 99887.69, 99864.34, 99858.17,
  100819.9, 100784.4, 100746, 100719.1, 100702.2, 100699.7, 100705.2, 
    100721.9, 100750.8, 100791.5, 100839.5, 100899.5, 100963.8, 101038.3, 
    101116.4,
  100756.9, 100705.9, 100663.1, 100628, 100602.6, 100591.2, 100593.9, 
    100612.3, 100639.2, 100678.9, 100725.7, 100784.7, 100850.9, 100925.2, 
    101004.8,
  100682.7, 100622.6, 100577.7, 100533.8, 100508, 100492.4, 100490, 100500.7, 
    100525.2, 100562.6, 100610.3, 100668.3, 100731.6, 100808.5, 100885.4,
  100611.6, 100544.8, 100492.9, 100438.1, 100408.1, 100384, 100381.3, 
    100393.7, 100415.1, 100451.7, 100497.6, 100554.4, 100616.7, 100690.8, 
    100772.6,
  100543.3, 100467.7, 100402.7, 100345.1, 100310.1, 100285.4, 100277.3, 
    100283.2, 100304.2, 100336.1, 100380.6, 100435.4, 100500.6, 100573.3, 
    100654.2,
  100477.8, 100395.1, 100319, 100254.1, 100209.7, 100184.3, 100173.5, 100173, 
    100187.8, 100217.8, 100262.2, 100317.7, 100381.8, 100453.9, 100537.5,
  100416.7, 100325.9, 100239.5, 100167.9, 100119.4, 100088, 100066.3, 100062, 
    100076.6, 100101.9, 100142.2, 100193.2, 100259.4, 100336.7, 100418.7,
  100362.4, 100264.9, 100168.5, 100089.4, 100032.3, 99990.2, 99964.72, 
    99950.45, 99958.17, 99977.55, 100017.5, 100068.9, 100134.3, 100209.8, 
    100295.1,
  100315.1, 100210.4, 100103.1, 100016.8, 99946.7, 99900.05, 99866.58, 
    99846.87, 99844.97, 99862.7, 99890.06, 99938.88, 100001.4, 100079.3, 
    100165,
  100276.4, 100162.1, 100046.6, 99949.67, 99869.29, 99816.8, 99769.66, 
    99742.07, 99731.05, 99736.03, 99761.3, 99805.59, 99865.55, 99944.04, 
    100031.9,
  101133.5, 101171.7, 101212.5, 101262.3, 101312.3, 101366.9, 101423, 
    101478.4, 101534, 101589.7, 101648.7, 101705.9, 101765.3, 101827.1, 
    101885.9,
  101087.9, 101128.4, 101171.1, 101220.8, 101271.1, 101320.8, 101368.7, 
    101419.6, 101471.4, 101524.5, 101581.2, 101637.3, 101694.8, 101755.2, 
    101815.2,
  101043.5, 101079.3, 101117.3, 101164.1, 101206, 101251.1, 101297.9, 
    101344.2, 101394.1, 101444.4, 101497, 101553.1, 101612.3, 101670.5, 
    101733.7,
  101001.5, 101033.2, 101072.3, 101110.8, 101154.9, 101191.9, 101231.3, 
    101271, 101315.2, 101363.1, 101413.8, 101466, 101522.3, 101578.8, 101641,
  100952.6, 100983.8, 101015.1, 101051, 101085.6, 101119, 101152.2, 101188.2, 
    101227.7, 101271.3, 101316.2, 101367.3, 101420.8, 101477.3, 101536.4,
  100902.6, 100930.3, 100958.1, 100993.9, 101022.9, 101051.8, 101077.7, 
    101107.2, 101140.2, 101176.2, 101218.7, 101263.6, 101312.4, 101367.5, 
    101425.1,
  100853.9, 100875.5, 100898.7, 100929.8, 100951.1, 100975.2, 100995.8, 
    101016.7, 101043.5, 101075.7, 101110.7, 101153.6, 101198.8, 101250.8, 
    101305,
  100802.6, 100820, 100835.4, 100861.9, 100879.2, 100898.3, 100913.4, 
    100929.7, 100950.6, 100977.4, 101005.3, 101040.8, 101082.4, 101129.9, 
    101180.4,
  100750.1, 100763.5, 100772.2, 100794.8, 100805.5, 100818, 100828.6, 
    100839.7, 100854.5, 100874.5, 100899.5, 100929.2, 100963.5, 101005.2, 
    101052.5,
  100698.3, 100703.4, 100705.8, 100723.1, 100727.1, 100737.8, 100741.1, 
    100748.5, 100757, 100773, 100792.3, 100817.1, 100846.2, 100881.6, 100924.3,
  101840.2, 101873.6, 101906.6, 101935.5, 101971.3, 102006.6, 102047.7, 
    102087.1, 102129.2, 102173.9, 102218.2, 102262.4, 102307.4, 102350.8, 
    102393,
  101793, 101816.4, 101843.7, 101872.8, 101906.9, 101940.6, 101981, 102023, 
    102066.3, 102111.4, 102159.7, 102207.9, 102257.4, 102303.6, 102349.7,
  101731, 101750.2, 101776.9, 101802.9, 101835.4, 101872, 101911.8, 101956.2, 
    102003.5, 102052.2, 102102.5, 102154.2, 102206, 102259.9, 102308.6,
  101671.2, 101686.4, 101707.9, 101731.2, 101761.3, 101797.8, 101840.4, 
    101887.2, 101935.4, 101987.8, 102042.2, 102097.6, 102154.3, 102211.8, 
    102265.5,
  101610.7, 101619.5, 101636.2, 101656, 101684.3, 101720.1, 101762.6, 
    101810.4, 101863.4, 101916.4, 101973.5, 102033.9, 102094.9, 102157.1, 
    102217.2,
  101547, 101551.6, 101563.1, 101579, 101605.1, 101638.1, 101680.2, 101727, 
    101780.4, 101837.1, 101896.2, 101959.4, 102024.4, 102090.4, 102155,
  101485.7, 101484.7, 101490.4, 101501, 101521.2, 101550.1, 101587, 101634, 
    101686.3, 101745.5, 101806.5, 101873, 101941.1, 102011.5, 102082.9,
  101426.2, 101417.2, 101416.7, 101420.3, 101433.7, 101456.6, 101490.9, 
    101535, 101585.7, 101642.8, 101705.8, 101772.7, 101845, 101919.3, 101994.3,
  101366.8, 101352.6, 101343.4, 101340.9, 101347.4, 101361.2, 101388.3, 
    101426.2, 101475.2, 101531.5, 101593.7, 101662.2, 101735.7, 101814.2, 
    101894.8,
  101309.5, 101287.4, 101270.5, 101260.8, 101255.3, 101262.5, 101281.6, 
    101313.5, 101357.6, 101410.7, 101471.4, 101538.4, 101612.4, 101691, 
    101776.5,
  102225.1, 102264.3, 102297.1, 102326, 102348.1, 102365.2, 102380.1, 
    102381.5, 102383, 102375.6, 102371.3, 102367.1, 102361.8, 102357, 102351.5,
  102217.8, 102257.5, 102287.2, 102319, 102341.5, 102359.1, 102373.3, 
    102381.8, 102376.9, 102367.6, 102359.8, 102350.5, 102341.8, 102327.8, 
    102312.1,
  102206.9, 102247.3, 102281.9, 102312.4, 102334.3, 102353, 102364.3, 
    102371.2, 102370.4, 102363.1, 102350.7, 102333.4, 102314.4, 102295.2, 
    102271,
  102185, 102227.6, 102265.3, 102295.5, 102318.2, 102336.9, 102346.6, 
    102354.4, 102349.6, 102340.6, 102325, 102306.1, 102284.8, 102259.1, 
    102229.1,
  102158.5, 102200.7, 102241.1, 102275.6, 102301.5, 102316.8, 102322.7, 
    102325.1, 102321.7, 102313.1, 102293.3, 102269, 102238.6, 102208, 102172.6,
  102124.9, 102169.1, 102208.3, 102242.4, 102270.8, 102285.8, 102292.6, 
    102288.6, 102281.4, 102268.4, 102248, 102219.1, 102185, 102146.5, 102108.5,
  102086, 102131.4, 102170.8, 102201.2, 102224.1, 102240.5, 102245.9, 
    102242.3, 102230.8, 102214.1, 102191.7, 102157.7, 102120.2, 102075.9, 
    102027.6,
  102037.5, 102080.4, 102117.8, 102144.4, 102164.8, 102181.7, 102187.2, 
    102183.6, 102171.3, 102152.3, 102122.2, 102085.9, 102042.7, 101992, 
    101937.8,
  101981.2, 102020.4, 102056.1, 102080.8, 102098.1, 102109.3, 102114.8, 
    102109.6, 102098.8, 102076.2, 102043.1, 102002, 101955, 101898.4, 101838.2,
  101919, 101953.5, 101983.7, 102005.7, 102022, 102030.6, 102032.6, 102026.9, 
    102014.6, 101990.4, 101955.4, 101909.9, 101853.9, 101792.1, 101725.2,
  102298.4, 102285.6, 102272.2, 102247.1, 102222.9, 102205, 102179.6, 102161, 
    102152.5, 102143.4, 102139.2, 102133, 102123.1, 102114.1, 102103.5,
  102306.3, 102284.9, 102261.5, 102234, 102207.3, 102176.1, 102147.2, 
    102123.4, 102104.7, 102091.3, 102081.7, 102070.1, 102058.6, 102047, 
    102032.1,
  102302.5, 102271.5, 102245.1, 102205.8, 102170.9, 102135.1, 102103.9, 
    102070.2, 102047.8, 102030.4, 102014.5, 101999.7, 101987.7, 101974.4, 
    101961.2,
  102297.1, 102255.6, 102224.7, 102177.4, 102136.9, 102096.5, 102057.3, 
    102020.3, 101990.4, 101967.2, 101947.4, 101927.9, 101910.9, 101892.7, 
    101873.4,
  102278.3, 102231.1, 102195.1, 102137.5, 102091, 102044.2, 101999.7, 
    101957.6, 101922.7, 101895.3, 101869.7, 101846.9, 101825.8, 101803.6, 
    101781.7,
  102258.2, 102204.1, 102158.1, 102098.9, 102042.3, 101988, 101936.8, 
    101890.6, 101851.9, 101818.9, 101789.3, 101765.1, 101742.2, 101717.8, 
    101694.4,
  102237.3, 102172.6, 102119.3, 102051.7, 101988.7, 101926.7, 101867.6, 
    101814.9, 101772, 101732.6, 101699.9, 101678.3, 101656.9, 101642.3, 101629,
  102210.2, 102140.7, 102077.1, 102003.1, 101931.7, 101859.2, 101790.4, 
    101731.7, 101678.8, 101642, 101615.8, 101601.4, 101595.4, 101593.1, 
    101593.6,
  102177.1, 102101.3, 102026.4, 101945.1, 101864.3, 101783.2, 101709.8, 
    101644.3, 101593.8, 101558, 101537, 101525.4, 101525.2, 101533.5, 101549.9,
  102137.1, 102058.2, 101978.9, 101889.3, 101799, 101710, 101629.2, 101555.1, 
    101505.5, 101470.4, 101454.1, 101452.8, 101462.2, 101482.8, 101508.1,
  102406.5, 102400.7, 102392.9, 102387.2, 102395.5, 102403.8, 102408.5, 
    102407.1, 102414.7, 102418.5, 102419.9, 102413.5, 102408.8, 102402.6, 
    102392.2,
  102405.9, 102386.5, 102375.7, 102378.5, 102386, 102384.5, 102390.1, 
    102393.2, 102393, 102389.3, 102387.6, 102380.9, 102376.2, 102366, 102352.9,
  102386.7, 102369.6, 102366.9, 102364.1, 102365.6, 102365.4, 102366.2, 
    102361.2, 102358, 102355.5, 102350.4, 102346, 102336.9, 102324.7, 102310.5,
  102364.7, 102352.7, 102350, 102345.6, 102347.1, 102346.3, 102345.1, 
    102344.3, 102335.6, 102325.6, 102317.6, 102307.7, 102292.1, 102273.2, 
    102253.4,
  102340.7, 102331.9, 102326.9, 102324.2, 102326, 102327.9, 102325, 102321.6, 
    102312.5, 102299.3, 102285.9, 102267.8, 102241.9, 102212.5, 102193.1,
  102323.3, 102312.6, 102304.5, 102297.7, 102296.3, 102303.2, 102308.2, 
    102311.8, 102305, 102288.1, 102264, 102238.7, 102210.5, 102183, 102167.6,
  102298.8, 102285.1, 102273.4, 102272.1, 102277.4, 102293.8, 102304.6, 
    102315.9, 102324.3, 102321.2, 102304.9, 102280.9, 102254, 102226.6, 102220,
  102280.5, 102260.3, 102248.6, 102248.2, 102257.6, 102287.1, 102317.7, 
    102347.6, 102371.8, 102379.7, 102378.7, 102360.8, 102351.5, 102333.8, 
    102325.6,
  102251.5, 102233.7, 102225.2, 102230.9, 102261.2, 102293.4, 102336.9, 
    102378.5, 102402, 102418.4, 102427.5, 102425, 102421.4, 102412.3, 102405.1,
  102226.8, 102212, 102218.8, 102229.5, 102256.7, 102302.5, 102352, 102394, 
    102421.2, 102444.6, 102456.9, 102466.2, 102463.2, 102458.9, 102448.8,
  102439.1, 102455, 102484.1, 102495.1, 102521, 102525.1, 102538.5, 102557.4, 
    102572.4, 102586, 102593.3, 102599.6, 102600.8, 102599.2, 102592.9,
  102460.8, 102474.4, 102499, 102509.4, 102534.8, 102536.9, 102551.9, 
    102561.7, 102562.4, 102568.7, 102581.1, 102585.4, 102584.1, 102581, 102578,
  102477.3, 102504.3, 102518, 102519.2, 102538.2, 102538.6, 102548, 102540.9, 
    102542.5, 102550, 102550, 102556, 102555.3, 102555, 102553.7,
  102484.1, 102518.6, 102523.8, 102526.2, 102549.9, 102549.4, 102544.2, 
    102535.3, 102527.9, 102525.5, 102521, 102517, 102514.9, 102517.5, 102520.2,
  102497.6, 102521.5, 102519, 102526.3, 102553.8, 102565, 102544, 102524, 
    102511, 102501.3, 102491.1, 102484.2, 102483.4, 102482.3, 102481.9,
  102495.2, 102501.9, 102520.8, 102520.1, 102537.8, 102549.2, 102544.1, 
    102526.6, 102499.4, 102481.8, 102461.7, 102447.4, 102446.5, 102460, 
    102479.9,
  102497.5, 102506.9, 102503.5, 102521.8, 102557.4, 102578.5, 102570.2, 
    102538.8, 102499.2, 102463.1, 102426.2, 102397.7, 102392.1, 102410.7, 
    102455.2,
  102503.4, 102515.2, 102514.6, 102545.9, 102576.5, 102604.6, 102586.3, 
    102576.1, 102532.6, 102477.7, 102429.7, 102392.6, 102382.7, 102407.1, 
    102455.7,
  102549.6, 102557.1, 102572.4, 102590.1, 102607.9, 102629.4, 102633.7, 
    102622.2, 102581, 102525.9, 102478.6, 102440.6, 102434.1, 102453.8, 
    102490.9,
  102580.2, 102593.8, 102621, 102618.6, 102631.4, 102648, 102649.7, 102650.7, 
    102623.2, 102581.7, 102536.2, 102511.4, 102501.6, 102506.2, 102525.9,
  102071.4, 102118.4, 102173.5, 102204.6, 102243.1, 102269.4, 102289.3, 
    102305.8, 102319.4, 102334.7, 102348, 102358.2, 102361.8, 102355, 102347,
  102120.4, 102159.3, 102200.8, 102219.3, 102259, 102283.3, 102298.7, 
    102301.8, 102317.1, 102332.6, 102345.9, 102355.8, 102362.9, 102354.1, 
    102342.2,
  102142.5, 102183.7, 102213.6, 102240.9, 102275.9, 102286.4, 102278.6, 
    102283.6, 102296.4, 102315.9, 102327.2, 102335, 102347.2, 102352.4, 
    102343.9,
  102171.9, 102201.2, 102216.3, 102244.7, 102275.6, 102276.2, 102263.5, 
    102268.6, 102284.4, 102303.7, 102318.3, 102324.7, 102327.4, 102334.8, 
    102334.5,
  102189.7, 102205.1, 102214.1, 102235.1, 102251.3, 102265.7, 102251.3, 
    102256.7, 102271.5, 102283.5, 102300, 102311.4, 102321, 102326.2, 102325.7,
  102174.4, 102206.9, 102204.4, 102231.4, 102249.2, 102232.4, 102227.5, 
    102228.5, 102242.9, 102261.9, 102279.3, 102304.2, 102324.8, 102330, 
    102322.4,
  102175, 102198.5, 102192.2, 102220.9, 102254.2, 102221.3, 102208.6, 
    102194.6, 102195.1, 102199.5, 102216.9, 102249.6, 102291.7, 102321.5, 
    102331.3,
  102200.6, 102203, 102200.8, 102217.2, 102247.7, 102211.1, 102189.9, 
    102163.7, 102154.3, 102153.1, 102171.4, 102207, 102255.6, 102298.5, 
    102318.2,
  102265.1, 102250.2, 102243, 102246.8, 102249, 102223.4, 102181.9, 102146.5, 
    102120.3, 102114.6, 102137, 102185.3, 102242.1, 102288.6, 102317.3,
  102285, 102287.7, 102283.9, 102261.9, 102253, 102226.4, 102176.9, 102134.4, 
    102100.1, 102094.3, 102120, 102189.6, 102239.2, 102275, 102298.9,
  101795.3, 101852.3, 101885.8, 101928, 101974.4, 101999.1, 102016.2, 
    102040.8, 102052.7, 102065.7, 102067.1, 102055, 102025.6, 101979.4, 
    101927.5,
  101810.1, 101865.6, 101905.2, 101944.1, 101978.9, 102001.8, 102028, 102062, 
    102069.6, 102082.2, 102078.1, 102071.7, 102054.4, 102004.4, 101944.1,
  101827.1, 101874.7, 101902.6, 101933.4, 101971.2, 102000.1, 102027.4, 
    102065, 102087.7, 102108.4, 102110.1, 102090.8, 102070.5, 102035.8, 
    101973.2,
  101845.1, 101875.7, 101913.7, 101938.5, 101964.9, 101997.6, 102024.5, 
    102063, 102097, 102120.6, 102133.3, 102126.9, 102097.1, 102058, 102006.7,
  101845.2, 101868.3, 101911.6, 101931.5, 101950.7, 101989.7, 102024.7, 
    102054.3, 102090.5, 102117.5, 102144.8, 102146.1, 102125.3, 102075, 102035,
  101841.4, 101862.1, 101900.8, 101920, 101940.3, 101980.9, 102023, 102064.7, 
    102108.4, 102140.8, 102157, 102160.9, 102148.3, 102110.6, 102055,
  101848.1, 101859.7, 101895.2, 101921.6, 101934.2, 101974.4, 102023.2, 
    102067.1, 102124.8, 102149.8, 102169, 102175.1, 102177.7, 102167.4, 
    102104.3,
  101861.8, 101871.8, 101903.6, 101920.1, 101939, 101968.2, 102026.3, 
    102076.4, 102128.2, 102164.5, 102186.3, 102202.1, 102201.9, 102194.5, 
    102154.9,
  101896.5, 101903.1, 101913.6, 101908.8, 101931, 101968.4, 102028.5, 
    102078.3, 102128.2, 102167.7, 102193.7, 102214.9, 102225.4, 102217.9, 
    102196.3,
  101915.4, 101911.4, 101915.7, 101913, 101929.7, 101966.2, 102023.3, 
    102073.5, 102127.2, 102163.2, 102195.8, 102220.1, 102233.4, 102231.3, 
    102215.4,
  101933, 101960.9, 101977.4, 101985.7, 102016.9, 102045.3, 102057.8, 
    102046.1, 102039.3, 102018.9, 101979.7, 101935.2, 101868.4, 101797.7, 
    101710.4,
  101976.4, 101988.8, 102012.4, 102033, 102048.1, 102062, 102064.8, 102077.2, 
    102072.9, 102052, 102005.5, 101950.7, 101887, 101808.3, 101715.2,
  102023.6, 102022.3, 102049.1, 102052.2, 102061.3, 102077.2, 102082.7, 
    102092.9, 102093.1, 102085.1, 102063.3, 101986.7, 101912.3, 101826.4, 
    101718.9,
  102049.4, 102046.2, 102082.5, 102086.5, 102088.6, 102093.7, 102104.6, 
    102110.7, 102117.2, 102110, 102082.1, 102033.5, 101944.6, 101853.9, 
    101731.1,
  102072.1, 102078.6, 102097.4, 102106.4, 102118.3, 102124.5, 102142, 102154, 
    102164.4, 102148.6, 102114.8, 102065.4, 101991.8, 101880.5, 101752.5,
  102098.3, 102114.5, 102135.8, 102147, 102157.4, 102167.8, 102194.2, 
    102201.7, 102224, 102209.4, 102163.5, 102100.7, 102032.4, 101918.4, 
    101778.4,
  102123.5, 102145.2, 102177.8, 102193.6, 102206.5, 102224.2, 102247.4, 
    102257.2, 102267.1, 102266.6, 102230.4, 102159.3, 102073.4, 101967.9, 
    101817,
  102140.7, 102172.3, 102215.5, 102235, 102258.7, 102294, 102307.7, 102312.9, 
    102314.4, 102304.6, 102277.4, 102221.9, 102129.2, 102021.9, 101876.6,
  102154.9, 102191, 102236, 102291, 102333.7, 102352.3, 102371, 102380.8, 
    102376.5, 102361.2, 102331.7, 102279.2, 102199.2, 102098.3, 101950.1,
  102168.8, 102216.9, 102284.9, 102337.4, 102373.7, 102397.1, 102428.7, 
    102434, 102425, 102407.4, 102377.8, 102331.6, 102258.1, 102167.7, 102035.3,
  102234.4, 102230.1, 102221.7, 102202.1, 102182.3, 102152, 102137.5, 
    102117.9, 102112, 102082.2, 102081.8, 102043.6, 101979, 101903, 101834.2,
  102299.9, 102298.7, 102292.2, 102276.2, 102256.9, 102236.3, 102211.1, 
    102179.1, 102170.3, 102139, 102112.8, 102077.8, 102022.5, 101904.7, 
    101832.4,
  102358.6, 102360, 102358.5, 102340.9, 102321.2, 102294.8, 102268.8, 102234, 
    102211.1, 102184, 102158.8, 102112.6, 102054.6, 101932, 101844.8,
  102411.2, 102417.8, 102419.6, 102406.2, 102386.3, 102359.6, 102331, 
    102292.9, 102257.5, 102224.6, 102190.4, 102149.6, 102077.3, 101957.7, 
    101849.7,
  102461.5, 102476.3, 102481.5, 102472.8, 102454.3, 102427.4, 102391.7, 
    102352.2, 102305.8, 102265, 102220.3, 102174.8, 102107.9, 101986.5, 
    101864.5,
  102517.5, 102538.8, 102547.7, 102546, 102532.4, 102505.8, 102469.9, 
    102422.3, 102367.8, 102318, 102263.2, 102201.5, 102142.2, 102011.2, 
    101876.8,
  102575.6, 102604.7, 102620.5, 102624.9, 102617.4, 102594.1, 102553.9, 
    102506.4, 102442.5, 102380.4, 102315.5, 102238.6, 102175.6, 102042.4, 
    101896.2,
  102635.8, 102670.2, 102689.8, 102699.1, 102698.8, 102686.8, 102654.6, 
    102601.5, 102532.2, 102454.3, 102381.4, 102287.7, 102211.3, 102089.2, 
    101925.9,
  102689.5, 102728.6, 102752.5, 102769.7, 102775.5, 102763.3, 102737.4, 
    102693.5, 102633.3, 102543.7, 102452.3, 102351.4, 102249.1, 102137.3, 
    101965.4,
  102740.6, 102787, 102818, 102842.8, 102850.1, 102845.8, 102825, 102784.4, 
    102723, 102636.8, 102531, 102422.2, 102297, 102182.6, 102013.8,
  102376.7, 102366.8, 102353.7, 102321.7, 102293.5, 102246, 102230, 102169.9, 
    102166.3, 102091.3, 102071.8, 102081.5, 102050.2, 102063.4, 102068.9,
  102468.8, 102456.2, 102444.5, 102422.3, 102402.6, 102359.6, 102339.5, 
    102283.2, 102275.5, 102201.2, 102205.8, 102170.4, 102125.7, 102111.4, 
    102110.1,
  102554.7, 102544.6, 102536.8, 102511.4, 102488.8, 102447.2, 102417.3, 
    102365, 102348.6, 102281.9, 102281.3, 102232.3, 102209.2, 102173.4, 
    102150.8,
  102644.6, 102637.2, 102627.7, 102608.4, 102586.6, 102550.2, 102518.2, 
    102460, 102436.1, 102374.8, 102362.6, 102296.1, 102265.2, 102210.7, 
    102179.6,
  102733.4, 102727.8, 102717.4, 102697.8, 102675.3, 102637.7, 102602.5, 
    102548.9, 102512.8, 102450.9, 102433.5, 102356, 102315.9, 102250.7, 
    102215.2,
  102823, 102819, 102812, 102791.7, 102765.4, 102732, 102692.2, 102641.2, 
    102595, 102523.5, 102488.8, 102408.7, 102358.7, 102288.4, 102220.6,
  102904.4, 102906.1, 102902.4, 102885.8, 102857.4, 102819.2, 102776.8, 
    102721.1, 102670.4, 102595.3, 102543.4, 102459.2, 102395.3, 102322.2, 
    102228.2,
  102991.4, 102993.1, 102987.5, 102968.9, 102945.6, 102910.9, 102867.5, 
    102805.2, 102747.8, 102663.2, 102595.2, 102501.5, 102429.8, 102351.1, 
    102229.5,
  103072.9, 103076, 103075.2, 103058.1, 103032.9, 102991.1, 102948.8, 
    102885.2, 102820.4, 102729.2, 102644.9, 102542.6, 102456.7, 102368.3, 
    102239.3,
  103151.8, 103161, 103163.8, 103146.5, 103121.2, 103075.9, 103027, 102963.8, 
    102892.1, 102797.5, 102695, 102578.8, 102475.4, 102379.5, 102243.5,
  102512.6, 102524.3, 102530.8, 102524.6, 102519.2, 102494.9, 102467.7, 
    102424.8, 102388.1, 102324.1, 102277.3, 102205.6, 102139.7, 102080.2, 
    102035,
  102612, 102617, 102627.5, 102621.8, 102615.5, 102600.7, 102578.1, 102544.4, 
    102503.5, 102452.9, 102406.3, 102339.9, 102288.1, 102237.5, 102187.1,
  102695.8, 102704.2, 102715.3, 102713.3, 102708, 102694, 102673.8, 102644.4, 
    102609.7, 102565.2, 102516.9, 102460.6, 102412.4, 102363.6, 102315.6,
  102788.9, 102799, 102809.9, 102808.8, 102803.5, 102789.6, 102769.3, 102742, 
    102710.3, 102672.3, 102632.8, 102588.1, 102542.7, 102497, 102449.2,
  102877.5, 102886.6, 102900.1, 102897.6, 102892, 102875.2, 102855.8, 
    102828.3, 102801.6, 102765.1, 102731, 102692.5, 102650.6, 102605.9, 
    102558.7,
  102970.2, 102979.1, 102991.9, 102989.1, 102983.2, 102966, 102944.1, 
    102915.8, 102887, 102852.2, 102822.1, 102785.2, 102750, 102704.1, 102659.6,
  103051.2, 103064.9, 103077.3, 103074.9, 103067.4, 103050.4, 103029.2, 
    102998.4, 102968.7, 102933.6, 102902.7, 102865.6, 102836.1, 102800.5, 
    102750,
  103135.9, 103149.2, 103159.8, 103159.3, 103151.4, 103134.2, 103110.2, 
    103081.7, 103046.2, 103009.4, 102976.4, 102937.9, 102902.3, 102866.4, 
    102820.1,
  103211.1, 103227.6, 103237.4, 103237.1, 103229.8, 103212.8, 103186, 103155, 
    103118.9, 103076.2, 103040.9, 103000.3, 102960, 102920.6, 102870.5,
  103285, 103297.4, 103306.8, 103308.3, 103302.8, 103284, 103259.6, 103224.4, 
    103184.8, 103139, 103098.2, 103048.9, 103008.8, 102956.6, 102906.3,
  102577.4, 102602.5, 102621.8, 102634.5, 102640.1, 102641.5, 102639.7, 
    102630.1, 102615.7, 102591.2, 102559.5, 102517.5, 102468.9, 102406.7, 
    102341.7,
  102679.1, 102697.1, 102720.1, 102731.1, 102741.8, 102742.9, 102740.3, 
    102733.6, 102720.8, 102699.5, 102669.6, 102632.2, 102590, 102532.9, 
    102470.3,
  102766, 102787.8, 102815.5, 102829, 102841.2, 102846.1, 102847.8, 102842.5, 
    102830.1, 102810, 102783.3, 102745.7, 102704.7, 102651.2, 102590.7,
  102858.2, 102883, 102909.4, 102925.1, 102940.2, 102945.4, 102949.5, 
    102945.8, 102935.5, 102917.7, 102892, 102857.5, 102817.1, 102768.2, 
    102710.4,
  102946.5, 102973.3, 103003.3, 103021.2, 103041.4, 103049.4, 103055.5, 
    103051.1, 103040.9, 103022.4, 102998.4, 102965.8, 102927, 102878.4, 
    102826.5,
  103038.3, 103065.1, 103096.4, 103116.5, 103136.3, 103145.9, 103154.4, 
    103152, 103144, 103124.3, 103100.5, 103068.4, 103031.4, 102985.6, 102930.3,
  103125.1, 103153, 103183.3, 103206, 103226.9, 103240.1, 103249.1, 103250.7, 
    103242.8, 103227.6, 103202.2, 103171.2, 103133, 103088.7, 103038,
  103206.7, 103240.6, 103274.7, 103298.7, 103318.3, 103329.9, 103337.1, 
    103338.3, 103329.1, 103314.4, 103293.6, 103263.2, 103229.5, 103193.8, 
    103142.9,
  103284.2, 103317.8, 103352.9, 103374.7, 103395.1, 103405.8, 103419.8, 
    103418.9, 103415, 103398.7, 103377.5, 103347, 103308.3, 103273.7, 103229.2,
  103349.1, 103383.4, 103419.9, 103443.1, 103468.7, 103480.2, 103491.9, 
    103486.2, 103482.4, 103467.1, 103448, 103422.5, 103386.5, 103347.4, 
    103305.7,
  102585.3, 102613.1, 102643.6, 102660.9, 102675, 102682.1, 102683.1, 
    102678.9, 102671.2, 102658.7, 102644.9, 102621.9, 102597.3, 102555.4, 
    102507,
  102693.2, 102714.3, 102742.5, 102759.2, 102776.1, 102784.4, 102788.1, 
    102782.3, 102772.6, 102758.4, 102742.4, 102723, 102696.2, 102659.2, 
    102617.1,
  102779.7, 102814.5, 102845.3, 102864.8, 102879, 102888.7, 102891.5, 
    102887.4, 102878.3, 102861.9, 102844.1, 102819.7, 102794.1, 102761.1, 
    102717.8,
  102876.9, 102911, 102938.5, 102963.1, 102981.8, 102988.7, 102993, 102988.7, 
    102980.8, 102964.4, 102945.1, 102919.9, 102891.5, 102857.7, 102815,
  102960, 102998, 103030.3, 103054.8, 103074.8, 103086.3, 103091.4, 103088, 
    103079.2, 103065.7, 103045.1, 103020.9, 102986.8, 102951.1, 102907.7,
  103037.8, 103077.5, 103114.2, 103142.1, 103166.9, 103178.8, 103184.2, 
    103183.2, 103176.4, 103163.5, 103144.2, 103117.4, 103088.5, 103050.3, 
    103002.7,
  103103.8, 103145.6, 103187.9, 103218, 103245.1, 103264.4, 103275.4, 
    103277.7, 103273.4, 103256.5, 103241.1, 103211.4, 103178.6, 103137.1, 
    103091.6,
  103159.9, 103204.6, 103249.6, 103286.4, 103318, 103340.2, 103355.9, 
    103361.6, 103358.2, 103345.6, 103330.3, 103304.9, 103272, 103228, 103178.4,
  103202.9, 103252.1, 103302.9, 103343.2, 103378, 103405.6, 103423.7, 
    103433.7, 103431.6, 103419.8, 103403.3, 103376.2, 103345.8, 103306.4, 
    103257.6,
  103238, 103290.1, 103341.9, 103385, 103424.5, 103454.9, 103480.5, 103495.3, 
    103494.7, 103487.9, 103473, 103445.6, 103409.8, 103368.6, 103324.5,
  102585.7, 102607.7, 102627.4, 102638.9, 102648.9, 102656.7, 102660.7, 
    102661.1, 102657.6, 102649.8, 102639.3, 102619.8, 102602.7, 102566.4, 
    102540.2,
  102674.3, 102696.7, 102717.8, 102733.7, 102747.8, 102757.4, 102761.2, 
    102760.6, 102756.3, 102747.8, 102734.1, 102713.5, 102690.4, 102655.1, 
    102620.3,
  102742.8, 102772.2, 102799.8, 102819.8, 102838.9, 102851.6, 102857.9, 
    102858.2, 102853.7, 102842.6, 102826.3, 102804.2, 102777.1, 102741.1, 
    102698.6,
  102811.8, 102844.1, 102871.4, 102897.8, 102916.5, 102929.3, 102940.7, 
    102944.3, 102939.8, 102930.2, 102915, 102889.6, 102859.1, 102821.9, 
    102778.5,
  102870.4, 102905.9, 102938.3, 102967.2, 102988, 103007.9, 103024.9, 103032, 
    103029.2, 103016.2, 102997.4, 102970.4, 102939, 102896.5, 102851,
  102924.9, 102966, 102998.5, 103030.6, 103054.5, 103077.4, 103093.8, 
    103106.4, 103106.9, 103094.3, 103072.9, 103043.7, 103009, 102970.5, 
    102922.2,
  102967.4, 103013.6, 103051.5, 103087.8, 103115.5, 103142, 103159.9, 103173, 
    103175.6, 103169.6, 103151.7, 103123, 103083.8, 103035.6, 102991.6,
  103004.9, 103055, 103100.7, 103136.8, 103166.5, 103194.1, 103211.4, 
    103225.1, 103233, 103229, 103214.3, 103183.4, 103144.1, 103099.5, 103050.3,
  103034.1, 103087, 103137.3, 103175.4, 103208.4, 103240.3, 103260.5, 
    103272.8, 103278.3, 103280, 103266.1, 103244, 103205.5, 103156.4, 103100.1,
  103052.3, 103109.8, 103160.9, 103204, 103246.1, 103280.3, 103297.8, 
    103304.4, 103311.8, 103311.7, 103307.1, 103280.1, 103245.9, 103195.2, 
    103139.2,
  102548.3, 102568.9, 102573, 102576.5, 102572, 102561.4, 102546.4, 102522.8, 
    102501.9, 102468.7, 102435.8, 102401.5, 102360.5, 102319.1, 102272.2,
  102634.1, 102651.8, 102660, 102666.1, 102667.3, 102661.1, 102649.4, 
    102629.6, 102605.3, 102572.1, 102540.5, 102503.2, 102463.4, 102417.1, 
    102363.5,
  102702.7, 102722.7, 102736.2, 102747.6, 102749.8, 102746.8, 102736.4, 
    102719.4, 102696.5, 102664.4, 102633.7, 102597.2, 102556, 102504.7, 102448,
  102771.1, 102796.1, 102813.3, 102829, 102834.9, 102835.5, 102826.4, 
    102808.5, 102784.5, 102755, 102720.5, 102681.8, 102639.5, 102588.8, 
    102530.3,
  102828.5, 102858.9, 102882.6, 102901.4, 102913.1, 102915.5, 102908.4, 
    102894.9, 102870.7, 102840.4, 102805, 102765, 102722, 102666.1, 102602.3,
  102882, 102913.3, 102943.5, 102967, 102987.8, 102993, 102987, 102974.3, 
    102952.5, 102924, 102885.9, 102843, 102796.3, 102741.7, 102673.1,
  102926.3, 102962.4, 103001, 103030.5, 103051.5, 103060.8, 103063.9, 
    103050.2, 103030.6, 102999.7, 102963.3, 102919.2, 102867.8, 102807, 
    102737.6,
  102967.5, 103009.9, 103048, 103084, 103107.8, 103121.9, 103127, 103119.2, 
    103099.6, 103070.8, 103031.6, 102985.3, 102936.2, 102873.2, 102797.7,
  103009, 103050.1, 103097, 103131.4, 103154.8, 103170.3, 103179.4, 103172.4, 
    103154.1, 103123, 103087.4, 103043.1, 102991.7, 102924.8, 102846.1,
  103043.6, 103094.1, 103141.3, 103172, 103198.6, 103215.1, 103227.4, 
    103225.5, 103203.6, 103170.3, 103130.9, 103090.7, 103038.2, 102972, 
    102888.5,
  102503.4, 102503.4, 102498.6, 102485.8, 102468.9, 102440.7, 102408.8, 
    102375.5, 102343.6, 102308.7, 102271.1, 102230.1, 102192.6, 102151.3, 
    102109.7,
  102588.2, 102585.3, 102583.8, 102576.4, 102564.5, 102547.5, 102524.4, 
    102496.7, 102460.6, 102425, 102389.6, 102354.4, 102319.3, 102277.4, 
    102230.4,
  102663.1, 102668.5, 102668.8, 102664.1, 102653.4, 102642.1, 102621.5, 
    102597, 102574.2, 102546.9, 102513.9, 102477.5, 102434.2, 102384.1, 
    102328.1,
  102734.7, 102744.7, 102746.6, 102745.4, 102740.4, 102730.4, 102717.6, 
    102700.1, 102675.2, 102643.9, 102613.5, 102576.1, 102532.4, 102480.6, 
    102422,
  102810.2, 102820.1, 102825.7, 102826.6, 102822.2, 102812.7, 102798.1, 
    102780.2, 102758.9, 102730.8, 102701.1, 102660.1, 102615.4, 102559.2, 
    102501.8,
  102876, 102888.5, 102896.7, 102899.2, 102897.5, 102892, 102882.7, 102866, 
    102841.2, 102813.3, 102780.9, 102741.9, 102694, 102637.1, 102576.8,
  102939.6, 102957.7, 102971.4, 102976.3, 102981, 102972.2, 102964.3, 
    102947.1, 102927.4, 102897.3, 102860.6, 102818.3, 102765.3, 102706.3, 
    102640.4,
  102989.5, 103011.9, 103028.2, 103046.2, 103059.1, 103055.9, 103049.2, 
    103033.8, 103009.6, 102978.6, 102940.8, 102896.5, 102840.9, 102777.6, 
    102704.4,
  103042.3, 103071.7, 103090, 103113.4, 103122.7, 103125.2, 103115.2, 
    103100.2, 103080.3, 103047.7, 103007, 102959.1, 102898, 102837.5, 102754.3,
  103087.4, 103116.6, 103142.5, 103168.2, 103179, 103184.2, 103185.8, 
    103169.1, 103147.8, 103120.3, 103077.9, 103025.1, 102955.5, 102884.5, 
    102795.9,
  102435.2, 102420.6, 102398.3, 102354.3, 102304.8, 102249.1, 102190, 
    102122.7, 102023.8, 101969.9, 101903.1, 101846.6, 101777.7, 101715.5, 
    101648.9,
  102512.9, 102500.4, 102488.7, 102459.4, 102420, 102366.3, 102306.2, 
    102249.4, 102194.2, 102133.6, 102057, 101999.8, 101934.3, 101879.2, 
    101818.8,
  102575.9, 102572.8, 102576.8, 102558.4, 102529.7, 102492.2, 102447.5, 
    102390.3, 102327.5, 102266.9, 102211.4, 102159, 102100.7, 102046.8, 
    101983.9,
  102635.6, 102642.4, 102645.1, 102636.8, 102624.8, 102598.7, 102564.1, 
    102524, 102481.7, 102427, 102368.6, 102310.1, 102250, 102194.1, 102132.2,
  102686.1, 102697, 102704.8, 102708.4, 102699, 102685.5, 102664.6, 102630.2, 
    102590.5, 102542.3, 102493.5, 102440.7, 102384.7, 102326.9, 102266,
  102735.3, 102753.5, 102761.6, 102769.3, 102768.2, 102761.3, 102745.6, 
    102723, 102693.4, 102653.6, 102605.7, 102551.8, 102494.8, 102438.4, 
    102380.2,
  102782.7, 102800.6, 102816, 102825, 102825.4, 102821.2, 102809.6, 102792.8, 
    102766.8, 102734.1, 102692.4, 102643.6, 102590.7, 102534.9, 102477.5,
  102814.6, 102840.1, 102864.2, 102878.7, 102887.9, 102886, 102879.2, 102865, 
    102840.4, 102808.1, 102769.8, 102725.8, 102672.9, 102619, 102564.5,
  102846.8, 102881.8, 102913.1, 102927.9, 102937.3, 102936.6, 102930.4, 
    102918.2, 102903.3, 102874.3, 102830.9, 102788.4, 102740.9, 102691.4, 
    102633.4,
  102867.2, 102906.9, 102939.7, 102964.5, 102978.6, 102984.1, 102987.3, 
    102975.7, 102956.3, 102933.9, 102898.7, 102846.4, 102792.6, 102747.7, 
    102684.6,
  102491.1, 102469.3, 102426, 102390.3, 102334.6, 102270.1, 102177.6, 
    102075.8, 101978.1, 101867.7, 101769.6, 101697.8, 101637.7, 101589.2, 
    101537,
  102557.5, 102548.6, 102520, 102471.1, 102419.4, 102361.4, 102284.9, 
    102189.3, 102080.3, 101973.9, 101874.6, 101792.1, 101728.3, 101677, 
    101626.8,
  102602, 102587.5, 102572.2, 102542, 102497.3, 102449, 102391.7, 102305.2, 
    102203.8, 102093.3, 101985.8, 101895.5, 101827.3, 101773.1, 101724.1,
  102642, 102651.3, 102647.1, 102624.4, 102588.6, 102535.6, 102476.5, 
    102403.1, 102319.4, 102223.3, 102120.3, 102023.8, 101946.3, 101888.1, 
    101836.5,
  102665.1, 102676.8, 102677.8, 102668.1, 102644, 102611.8, 102567.3, 
    102514.1, 102441.6, 102353.9, 102262.2, 102163.4, 102084, 102020.2, 
    101962.2,
  102686.5, 102708.5, 102719.9, 102721.3, 102710, 102684.9, 102644.7, 
    102594.1, 102537.1, 102471.3, 102398, 102310.9, 102234.2, 102164.6, 
    102102.7,
  102682.8, 102710.4, 102734.2, 102744.3, 102746.7, 102732, 102709.7, 
    102675.2, 102628.3, 102574.2, 102512.7, 102443.5, 102375.7, 102303.7, 
    102239.1,
  102674.7, 102714.5, 102744.5, 102763.3, 102778.2, 102778.8, 102757.9, 
    102733.5, 102697.7, 102646.9, 102599.4, 102545.1, 102489, 102431.6, 
    102369.6,
  102651.1, 102695.4, 102735.7, 102760.9, 102781.1, 102787.2, 102780.4, 
    102770.2, 102756.6, 102724.8, 102679, 102631, 102575.5, 102521.7, 102469.9,
  102620.7, 102669.6, 102718.1, 102749.2, 102773.1, 102786.4, 102792.5, 
    102787, 102777.3, 102755.5, 102726, 102684.6, 102647.8, 102594.5, 102541.3,
  102677.6, 102668.8, 102636, 102591.1, 102538.7, 102462.5, 102384.1, 
    102308.2, 102220.6, 102124.3, 102025.4, 101940.4, 101879.3, 101830.9, 
    101784.8,
  102727.8, 102712.7, 102691.7, 102652.3, 102601.6, 102541.4, 102466.2, 
    102387.5, 102294.8, 102198.7, 102102.1, 102016.7, 101943.2, 101882.1, 
    101823.9,
  102766.5, 102752.2, 102735.9, 102702.4, 102658.1, 102603.6, 102534.7, 
    102459.6, 102368.8, 102279.5, 102185.2, 102090.4, 102007.1, 101928.8, 
    101855.5,
  102789.1, 102790.7, 102784, 102757.7, 102710.9, 102663.9, 102599.9, 
    102526.5, 102433.7, 102332.7, 102237.2, 102143.8, 102056.1, 101969.4, 
    101890,
  102794.6, 102807.6, 102806.4, 102789.4, 102756.8, 102704.6, 102644.3, 
    102572, 102487.7, 102385.6, 102279.1, 102182.8, 102082.9, 101993.7, 
    101914.2,
  102801.5, 102821.9, 102826.9, 102825, 102800.1, 102754.6, 102690.2, 
    102618.7, 102530.5, 102431, 102309.1, 102200.5, 102096.6, 102009.9, 
    101932.3,
  102796.6, 102825.6, 102847.1, 102844.4, 102829, 102796.2, 102734.3, 
    102661.4, 102585.9, 102477.5, 102349.9, 102228.5, 102115.3, 102027.8, 
    101956.4,
  102780.9, 102817.9, 102848.6, 102854.2, 102847.9, 102828.3, 102786.8, 
    102706.4, 102620, 102519.3, 102393.9, 102268.9, 102150.2, 102057.3, 
    101988.2,
  102754.9, 102798, 102833.2, 102854.5, 102850, 102840.4, 102809, 102749.3, 
    102658.8, 102554.3, 102433, 102311.5, 102191.5, 102097.3, 102025.6,
  102722, 102765.9, 102805.1, 102834.6, 102844.1, 102843.7, 102811.3, 
    102768.2, 102693, 102591.7, 102472.4, 102353.3, 102237.6, 102142.5, 
    102072.1,
  102791.9, 102778.3, 102756.2, 102725.8, 102674.5, 102612.4, 102549.9, 
    102475.9, 102404.7, 102348, 102313.4, 102278, 102244, 102201.7, 102175.5,
  102825.6, 102804.4, 102777.4, 102747.5, 102696.5, 102633.1, 102557.6, 
    102485.3, 102415.7, 102350.6, 102300.1, 102255.1, 102212.3, 102175, 102157,
  102838.8, 102820.5, 102791.2, 102759.7, 102714.9, 102650.4, 102573.7, 
    102494.3, 102415.1, 102340.8, 102278.6, 102225.5, 102180.5, 102154.9, 
    102135.5,
  102843.4, 102835.1, 102812.2, 102775.6, 102726.6, 102659.2, 102580.2, 
    102497.6, 102416.9, 102339.7, 102266.1, 102200.7, 102154.1, 102132.9, 
    102103.3,
  102842.6, 102834.9, 102809.5, 102777.4, 102727.6, 102657.5, 102578.3, 
    102494.4, 102412.2, 102329.4, 102248.3, 102180.9, 102140.5, 102108.4, 
    102060,
  102842.1, 102838.4, 102808.7, 102774.6, 102727, 102655.5, 102572, 102484.2, 
    102394.4, 102313.4, 102232.6, 102166.5, 102114.8, 102064.2, 102025.1,
  102835.5, 102823.6, 102807.4, 102764.9, 102705.2, 102633.4, 102552.5, 
    102464.3, 102373, 102285.8, 102207.5, 102140.6, 102078.6, 102026.8, 
    101985.8,
  102822.1, 102807.2, 102793.6, 102746.5, 102687.2, 102616.5, 102531.3, 
    102440.4, 102343.1, 102254.5, 102178.1, 102107.2, 102036.4, 101980.1, 
    101939.7,
  102803.4, 102782.7, 102764.6, 102722.1, 102656.4, 102580.7, 102495.7, 
    102399.8, 102301.6, 102214.5, 102135.9, 102056.1, 101986, 101930.8, 
    101882.3,
  102781.6, 102764.9, 102737.9, 102695.7, 102623.1, 102541.5, 102455.9, 
    102353.4, 102255.3, 102162.7, 102073.7, 101995, 101929.3, 101866.3, 
    101814.8,
  102572.8, 102572.1, 102566.7, 102565.4, 102560.6, 102559.6, 102557.4, 
    102561.8, 102573.7, 102586.8, 102600.7, 102613.2, 102621.9, 102622.6, 
    102634.2,
  102538.1, 102528.1, 102520, 102519.4, 102514.6, 102512.9, 102515.2, 
    102526.5, 102540.5, 102551.9, 102565.2, 102580.6, 102604.2, 102630.1, 
    102651,
  102488.9, 102481.2, 102474.7, 102473.4, 102471.4, 102473.8, 102480.2, 
    102493.9, 102512.2, 102529.9, 102550.3, 102575, 102601, 102620.4, 102630.6,
  102435.2, 102427.8, 102420, 102418.4, 102416.9, 102421, 102432.3, 102448.6, 
    102468.6, 102488.7, 102511.6, 102540.2, 102573.1, 102597.5, 102612.8,
  102371.6, 102366.7, 102359.3, 102359, 102362.6, 102368.1, 102382.9, 
    102402.9, 102426.2, 102450.4, 102476.9, 102506.3, 102535.5, 102558.5, 
    102580.5,
  102302.9, 102297.4, 102292, 102293.2, 102296.7, 102305.8, 102323.3, 
    102347.3, 102373.1, 102401, 102432.6, 102466, 102496.6, 102524.8, 102547,
  102232.7, 102222.5, 102218.5, 102219.4, 102225.4, 102237.7, 102257.6, 
    102285, 102315.6, 102349.5, 102384.4, 102414.2, 102443.5, 102474.5, 
    102496.1,
  102159.2, 102146.5, 102140.3, 102139.4, 102147, 102162.2, 102185.1, 
    102215.6, 102251.2, 102289.7, 102324.2, 102353.4, 102384.9, 102415.5, 
    102439.2,
  102083.8, 102065.9, 102057, 102053.8, 102063.6, 102079.1, 102105.2, 
    102139.9, 102179.8, 102214.8, 102245.7, 102275.2, 102309.1, 102338, 
    102362.2,
  102003.2, 101984.2, 101972.6, 101968.9, 101975.3, 101992.2, 102017.5, 
    102051.1, 102090.6, 102124.8, 102157.6, 102193.2, 102222.6, 102244.2, 
    102262.8,
  102228.4, 102283.2, 102329.8, 102374.1, 102418.1, 102458.6, 102492.2, 
    102522.3, 102547.6, 102570.3, 102584.7, 102596.9, 102604, 102591.8, 
    102562.2,
  102198.5, 102251.9, 102302.2, 102352.4, 102396.6, 102437.2, 102473.3, 
    102507.6, 102534, 102557, 102575.9, 102586.5, 102589.9, 102587.8, 102578.5,
  102161.3, 102208.7, 102262, 102315.9, 102362.4, 102409.1, 102447.2, 
    102484.1, 102515.8, 102542, 102566.1, 102581.5, 102588.9, 102587.7, 
    102573.1,
  102109.8, 102161.5, 102221.3, 102272.1, 102320.7, 102367.9, 102410.6, 
    102451.1, 102484.6, 102517.5, 102539.1, 102555.9, 102565.5, 102570.9, 
    102570.6,
  102050.4, 102101.8, 102162, 102213.6, 102266.4, 102314.3, 102362.5, 
    102405.3, 102444.3, 102479, 102512.1, 102530.5, 102542.9, 102544, 102544.1,
  101985, 102037.4, 102093.1, 102146.5, 102201.3, 102252.5, 102301, 102346.8, 
    102389.9, 102426.9, 102461.1, 102487.1, 102506.5, 102519, 102518,
  101911.2, 101963, 102014.6, 102067.1, 102120.2, 102172.1, 102224, 102272.1, 
    102318, 102360.2, 102397.7, 102426.8, 102452.7, 102469, 102479.1,
  101830, 101879, 101928, 101979.4, 102031, 102082.7, 102133.3, 102181.1, 
    102227.8, 102273.9, 102312.2, 102349.3, 102378.8, 102403.9, 102419.8,
  101742.8, 101787.1, 101833.2, 101882.5, 101931, 101982.2, 102032.6, 
    102081.9, 102128.6, 102173.2, 102216.2, 102254.9, 102290.3, 102319.9, 
    102343.1,
  101649.6, 101691.6, 101734, 101777.7, 101823.6, 101870.6, 101917.9, 
    101966.4, 102014.2, 102060.2, 102103.3, 102142.6, 102179.6, 102213.7, 
    102242.1,
  102305.8, 102352.4, 102395.5, 102438.1, 102469.5, 102494.6, 102504.2, 
    102500.2, 102489.8, 102473.6, 102451.4, 102418.6, 102363.1, 102320.2, 
    102277.6,
  102287.1, 102333.8, 102383.2, 102428, 102460.1, 102480.9, 102503.3, 102507, 
    102501.1, 102484.6, 102461.9, 102428.9, 102377.5, 102332.2, 102288.5,
  102256.2, 102297.8, 102349.8, 102392.4, 102435.9, 102474.2, 102497.2, 
    102506, 102504.8, 102491.8, 102465.3, 102440.7, 102386.9, 102331.3, 
    102284.5,
  102222.8, 102272, 102322.2, 102363.3, 102408.4, 102442.5, 102473.7, 
    102489.4, 102492.5, 102483.7, 102463.7, 102429.7, 102386.5, 102327.7, 
    102276.8,
  102191, 102241.4, 102284.1, 102330.3, 102374.3, 102410.9, 102444.9, 
    102468.4, 102475.4, 102473, 102452, 102417.3, 102378.8, 102318.4, 102259.4,
  102156.6, 102209, 102252.4, 102297.6, 102340.4, 102377.6, 102409.9, 
    102431.5, 102446.4, 102445.3, 102427.1, 102395.6, 102360.3, 102300.1, 
    102232.9,
  102126.2, 102175.2, 102222.3, 102262.8, 102302.6, 102341.7, 102373.1, 
    102395.3, 102411.3, 102417, 102400, 102373.6, 102329.8, 102276.1, 102208.2,
  102097.2, 102146.3, 102192, 102233.3, 102268.8, 102303.4, 102334.9, 
    102359.4, 102374.4, 102378.1, 102369.1, 102337.5, 102296.8, 102238.2, 
    102173.6,
  102069.3, 102119, 102162.4, 102204.3, 102240.3, 102272.6, 102294.4, 
    102316.5, 102333.9, 102337.9, 102328.8, 102296.2, 102253.2, 102199, 102136,
  102043.7, 102093.6, 102137.6, 102178.4, 102219.5, 102249.5, 102263.9, 
    102274.7, 102287, 102289.6, 102281.7, 102250.2, 102211.3, 102154.5, 
    102092.2,
  102550.6, 102580.5, 102592.9, 102593.3, 102590, 102587.1, 102565, 102522, 
    102465.4, 102391.6, 102305.7, 102198.3, 102080, 101952.9, 101817.8,
  102583, 102604.4, 102621.3, 102628.6, 102618.2, 102611.1, 102591.3, 
    102551.3, 102496.1, 102420.6, 102336.7, 102237.1, 102122.6, 102004.4, 
    101875.1,
  102606.5, 102623, 102637.1, 102646.5, 102640.1, 102639.2, 102620.4, 
    102577.7, 102524.2, 102451.1, 102366.8, 102274.1, 102164.8, 102047.2, 
    101927.5,
  102632.9, 102656.8, 102666, 102660.5, 102655.2, 102648.3, 102636.2, 
    102602.1, 102548.1, 102475, 102388.8, 102299.8, 102195.5, 102081.7, 
    101966.7,
  102660.2, 102680.8, 102690.3, 102689.2, 102678.8, 102664.8, 102648.7, 
    102617.2, 102564.8, 102496.2, 102410.1, 102320.1, 102222.6, 102107.3, 
    101997.2,
  102684, 102702.9, 102718.4, 102713.3, 102698.5, 102677.4, 102661.5, 
    102626.7, 102573.7, 102506.3, 102422.3, 102334.5, 102235.9, 102122.3, 
    102016.1,
  102710.3, 102731, 102744.1, 102739.8, 102726.4, 102700.1, 102667.7, 
    102632.7, 102579.5, 102508.8, 102427.1, 102339.4, 102238.8, 102132.4, 
    102023.6,
  102729.9, 102754.5, 102760.5, 102757.3, 102745.9, 102710.2, 102681.4, 
    102635.6, 102575, 102506.2, 102426.3, 102332.4, 102234.9, 102127.2, 
    102014.3,
  102752.6, 102768.6, 102778.3, 102779.9, 102762.9, 102715.9, 102677.8, 
    102631.8, 102567.6, 102497.5, 102411.2, 102317.3, 102219, 102111.9, 
    101997.4,
  102770.8, 102791, 102795.4, 102790.4, 102771.3, 102727.8, 102669.4, 
    102619.7, 102552.3, 102477.9, 102386.2, 102292.1, 102191.3, 102082.7, 
    101968.9,
  102597, 102603.3, 102585.7, 102546.8, 102497.7, 102439.1, 102370.7, 
    102283.5, 102178, 102055.3, 101922, 101785, 101651.1, 101516.4, 101389.2,
  102643, 102638.9, 102620.6, 102585.3, 102536.2, 102463.8, 102389, 102295.7, 
    102186.8, 102056.3, 101916, 101771.4, 101625.6, 101480, 101337,
  102680.8, 102669.6, 102646.8, 102616.7, 102568.6, 102495.2, 102411.3, 
    102315.3, 102203.4, 102069.8, 101920.9, 101766, 101603.7, 101442.9, 
    101292.6,
  102713.8, 102706.2, 102685.6, 102652.8, 102599.7, 102526.9, 102439.6, 
    102336.3, 102218.7, 102083.2, 101925.9, 101758.2, 101584.4, 101411.9, 
    101249.1,
  102748.7, 102740.5, 102719.7, 102684.1, 102629.9, 102555.8, 102464.5, 
    102359.8, 102238.2, 102096.9, 101935.9, 101760.1, 101571.2, 101387.2, 
    101217.2,
  102793, 102777.3, 102752.9, 102716.4, 102662.9, 102584.6, 102492.6, 
    102383.3, 102255, 102110.3, 101939.9, 101753.7, 101558.7, 101363, 101184.5,
  102831.3, 102818.9, 102794.8, 102753.6, 102695.6, 102614.5, 102515.3, 
    102403.8, 102273.8, 102122.2, 101948.6, 101754.4, 101551.3, 101343.5, 
    101164.8,
  102874.6, 102862.2, 102832.1, 102790.2, 102727.4, 102644.8, 102544, 
    102426.2, 102289.9, 102134.4, 101955.1, 101753.5, 101544.9, 101328.1, 
    101145.6,
  102912.4, 102902.1, 102868.4, 102824.5, 102758.3, 102670.9, 102564.6, 
    102447, 102305.8, 102145.7, 101964.8, 101756.9, 101542.5, 101321.5, 
    101139.1,
  102948.5, 102936.5, 102900.7, 102856.1, 102786.1, 102698, 102584.7, 
    102465.9, 102320.7, 102158.3, 101975.9, 101766.3, 101548.1, 101322.3, 
    101133,
  102517.5, 102511.8, 102495.3, 102464.6, 102424.7, 102375.3, 102307.4, 
    102235.5, 102168.2, 102104.8, 102035.6, 102015.6, 101976.7, 101954.7, 
    101913,
  102549.7, 102534.8, 102516.2, 102479.9, 102435.5, 102377.6, 102310.8, 
    102241, 102161.5, 102074.9, 102033, 102033.3, 102014.5, 101979.7, 101911.6,
  102576.5, 102552.8, 102532.5, 102494.8, 102445.4, 102379.3, 102306.6, 
    102230.4, 102141.1, 102069.6, 102078.4, 102036.7, 102009.2, 101957.3, 
    101916.5,
  102601.6, 102573.9, 102549.9, 102506.1, 102449.9, 102379.3, 102300.9, 
    102212.6, 102116.4, 102086.2, 102067.1, 102023.3, 102003.8, 101963.6, 
    101939.4,
  102622.4, 102591.9, 102561.5, 102513.4, 102452.9, 102374.2, 102288.1, 
    102198.5, 102117, 102088.9, 102046.2, 102024.3, 102008.1, 101986.4, 
    101979.3,
  102642.5, 102607.1, 102572.8, 102518.4, 102452.2, 102367.6, 102273.1, 
    102173.9, 102107.8, 102068.3, 102028.1, 102015.5, 101994.3, 101986.1, 
    101984.5,
  102661.5, 102618.7, 102579.6, 102518.9, 102447.3, 102355.1, 102254.4, 
    102154.5, 102090.6, 102038.3, 102002.6, 101986, 101970.2, 101974.8, 
    101979.9,
  102680.1, 102631.6, 102584.5, 102519.2, 102438.5, 102340.7, 102232.7, 
    102132.5, 102063.3, 102003.3, 101960, 101939, 101932.4, 101936.5, 101951.3,
  102695.4, 102643.7, 102587.7, 102515.3, 102427.3, 102322.8, 102208.6, 
    102109.4, 102028, 101961.6, 101914.7, 101888.2, 101883.6, 101893.1, 
    101912.1,
  102713.4, 102653.4, 102590, 102509.6, 102414.8, 102303.2, 102182.2, 
    102079.6, 101987.4, 101910.8, 101856.5, 101824.3, 101820.5, 101828, 
    101856.9,
  102381.1, 102374.3, 102359.2, 102333.4, 102294.7, 102246.9, 102191.4, 
    102119, 102041, 101943.7, 101841.5, 101714.3, 101628.2, 101525.6, 101547.1,
  102434.9, 102427.4, 102410.3, 102381.9, 102341, 102288.6, 102229.7, 102156, 
    102077.2, 101977.8, 101877.1, 101742.1, 101659.3, 101518.9, 101592.9,
  102488, 102476.6, 102454.6, 102426, 102384.7, 102331.9, 102271.2, 102191, 
    102111.2, 102008.9, 101911.5, 101786.1, 101702.2, 101576.6, 101596.4,
  102544.4, 102529, 102503.5, 102470.2, 102425.5, 102369.7, 102307.6, 
    102228.6, 102140.1, 102041.1, 101944.4, 101836.2, 101730.4, 101619.9, 
    101584,
  102594.9, 102575.7, 102549.2, 102513.1, 102463.5, 102408, 102342.2, 
    102259.1, 102172, 102082.1, 101988.1, 101894.9, 101791.4, 101687.3, 
    101597.2,
  102644.3, 102619.7, 102587.9, 102548.6, 102497, 102439.4, 102365.3, 
    102286.2, 102210.1, 102123.4, 102036.5, 101951.6, 101850.2, 101750, 
    101654.1,
  102697.9, 102668.5, 102630.9, 102582.8, 102527.9, 102465, 102389.1, 
    102313.7, 102248.9, 102171.2, 102091.4, 102016.6, 101916.4, 101823.9, 
    101722.4,
  102739.9, 102701.9, 102660, 102611.6, 102552.2, 102484.9, 102408, 102349.3, 
    102288.4, 102216.7, 102141.9, 102067.8, 101981.9, 101896.6, 101802.4,
  102774.7, 102728.8, 102681.4, 102631.3, 102567.8, 102501.7, 102429.2, 
    102384.8, 102326.9, 102267.9, 102199.8, 102127, 102048.8, 101971.8, 101885,
  102794.7, 102745.6, 102699.6, 102638.9, 102577.9, 102509.8, 102457, 
    102419.1, 102362.6, 102308.8, 102245.6, 102183.9, 102114.7, 102045.5, 
    101970.7,
  101946.2, 101899, 101875.2, 101921.1, 101946.9, 101926.8, 101895.9, 
    101827.6, 101747.3, 101658.6, 101583.7, 101531.7, 101500.9, 101483.8, 
    101479.8,
  102004.8, 101964.1, 101951.6, 101941.7, 101975.6, 101954.8, 101927.1, 
    101856.2, 101769.7, 101669.8, 101592, 101524, 101483.8, 101446.7, 101440.1,
  102101.6, 102054.5, 102016.8, 101976.9, 101981.8, 101986.3, 101942.6, 
    101879.3, 101792.4, 101679.8, 101595.5, 101519.1, 101461.9, 101413.2, 
    101405,
  102206.1, 102150, 102094.2, 102049, 102015.7, 102022.4, 101973, 101907.8, 
    101816.9, 101691.9, 101592.4, 101499.6, 101429.7, 101369.4, 101349.7,
  102310.3, 102249.8, 102183.4, 102127.7, 102068.6, 102039.7, 102011, 
    101935.3, 101849.8, 101721.3, 101603.7, 101494.5, 101414.1, 101341, 
    101300.5,
  102420.9, 102356.2, 102279.6, 102208, 102142.1, 102076.3, 102056, 101966.8, 
    101876.9, 101744.3, 101612.9, 101486.5, 101392.7, 101307, 101255.5,
  102527.2, 102460.8, 102378.9, 102292.6, 102215.1, 102130.8, 102090.6, 
    102009.9, 101909.6, 101773.8, 101630.9, 101485.6, 101382.3, 101279.3, 
    101212,
  102630.5, 102558.7, 102476.2, 102389.4, 102295.4, 102203.6, 102122.1, 
    102053.4, 101944.5, 101802.5, 101652.2, 101486.5, 101370.9, 101252.9, 
    101170.5,
  102723.2, 102652.5, 102568.6, 102472.5, 102373.1, 102276, 102171.5, 
    102097.4, 101980.9, 101836.7, 101680.3, 101496.2, 101366.5, 101229.4, 
    101130.6,
  102807.9, 102738.6, 102657.4, 102555.1, 102449, 102343.3, 102233.9, 
    102136.9, 102021.7, 101869.7, 101710.3, 101512, 101363.8, 101207.2, 
    101091.8,
  101997.4, 101934.2, 101915.8, 101952.7, 101973.2, 101984.3, 102000.1, 
    101991, 102004, 102050.1, 102097, 102142.3, 102191.4, 102238.2, 102285.5,
  102022.9, 101961.9, 101938.5, 101954.8, 101975.3, 101973.2, 101971.4, 
    101974.6, 102007.6, 102038.3, 102076.4, 102108.1, 102140.8, 102184.9, 
    102227.7,
  102077.5, 102003.6, 101953.4, 101927.8, 101969.7, 101961.3, 101958.4, 
    101962.9, 101981.5, 102002.3, 102041.4, 102061.2, 102090, 102129.2, 
    102162.4,
  102133.4, 102051.5, 101983.2, 101934.1, 101944.4, 101956.3, 101938.4, 
    101946.2, 101950.5, 101966.2, 101998.4, 102004.4, 102026.9, 102056.5, 
    102081.8,
  102190.6, 102103.3, 102012.7, 101955.1, 101910.4, 101938.4, 101923.3, 
    101921.6, 101921.9, 101923.2, 101949.2, 101948.1, 101961, 101977.9, 
    101998.3,
  102251, 102159.3, 102048.7, 101977.3, 101913.7, 101908.5, 101909.4, 
    101885.4, 101885.2, 101875.4, 101891.7, 101881.9, 101881.9, 101888.2, 
    101897,
  102308.2, 102211.6, 102092.4, 101995.5, 101925.3, 101874.2, 101891.9, 
    101852.3, 101848.4, 101828.2, 101831.5, 101810.5, 101799.6, 101792.5, 
    101790.8,
  102371, 102264.5, 102138.9, 102019.7, 101937.2, 101857.2, 101863.8, 
    101820.9, 101806.7, 101775, 101765.7, 101736.1, 101713, 101692.3, 101677.2,
  102436.6, 102316.9, 102188.1, 102049.7, 101947.8, 101858.9, 101822.9, 
    101799.2, 101763.8, 101725.4, 101701.5, 101660.6, 101622.8, 101587.6, 
    101557.6,
  102499.2, 102373.3, 102236.6, 102085.9, 101961.6, 101866.5, 101787.9, 
    101780.7, 101718.4, 101678.7, 101633.8, 101587.1, 101534.8, 101482.2, 
    101437.1,
  102241.4, 102309.2, 102413.8, 102500.2, 102594.6, 102688.5, 102786.6, 
    102874.1, 102953, 103034.9, 103099.6, 103172.2, 103240.2, 103313.6, 
    103386.8,
  102257, 102320.2, 102416.4, 102523.2, 102610.3, 102710.4, 102801.7, 
    102892.6, 102969.7, 103052.1, 103117.3, 103189.8, 103260, 103337.8, 103414,
  102264.8, 102337.8, 102416.1, 102540.1, 102609.4, 102721.7, 102803.9, 
    102896.5, 102971.3, 103053.8, 103123.9, 103205.2, 103284.8, 103362.3, 
    103433.4,
  102272.9, 102356.5, 102412.5, 102542.6, 102608.1, 102722.3, 102797.4, 
    102890.4, 102964, 103048, 103123.3, 103206.7, 103284.8, 103353.1, 103423.5,
  102280.1, 102370.5, 102411.3, 102540.1, 102601.2, 102707.2, 102779.5, 
    102869.8, 102942.3, 103028, 103103.5, 103187.5, 103260, 103333.1, 103399.8,
  102290, 102376.2, 102406.1, 102530.9, 102587.5, 102681.8, 102754.4, 102837, 
    102909.7, 102992.5, 103067.4, 103145.3, 103216, 103283.3, 103349.6,
  102299, 102377.2, 102396.3, 102510, 102560, 102648.1, 102713, 102792.2, 
    102862.2, 102939.3, 103011.4, 103085.7, 103152.7, 103217.7, 103281.7,
  102306.2, 102370.6, 102379.8, 102480.2, 102523.5, 102601.5, 102663.4, 
    102738.2, 102801.6, 102871.2, 102939.6, 103006.4, 103068, 103132.1, 
    103191.2,
  102311.6, 102354.7, 102359.5, 102440.3, 102480.1, 102545.5, 102602.7, 
    102668.4, 102726.4, 102790.6, 102849.8, 102910.5, 102967.1, 103024.1, 
    103083.6,
  102309.6, 102334, 102335.2, 102390.2, 102434.1, 102480.4, 102534.5, 
    102592.1, 102638.6, 102694.4, 102744.5, 102796.9, 102848.9, 102898.8, 
    102954,
  102764.3, 102830.3, 102878.9, 102935, 102990.6, 103066.2, 103123.4, 
    103185.9, 103252.2, 103316.8, 103376.8, 103437.6, 103495.8, 103555.8, 
    103612.3,
  102815.4, 102889.1, 102941.1, 103016.8, 103086.1, 103159.3, 103214.5, 
    103280.1, 103338, 103395.5, 103450.8, 103507.6, 103562.5, 103619.5, 
    103676.3,
  102854.6, 102958.2, 103020.8, 103098.2, 103158.6, 103224.4, 103279.2, 
    103340.8, 103397.4, 103455.6, 103509.6, 103564.8, 103617, 103671.1, 
    103721.6,
  102886.2, 102987.7, 103061.3, 103139.9, 103208.3, 103273.3, 103335.1, 
    103397.4, 103451.2, 103504.5, 103558.4, 103611.8, 103659.4, 103705.9, 
    103753.8,
  102899.5, 103010.1, 103093.1, 103170.9, 103242.6, 103308.1, 103370.5, 
    103429.9, 103486, 103535.8, 103588, 103638.2, 103679.7, 103719.9, 103760.2,
  102909.3, 103017.1, 103104.3, 103185.5, 103261.5, 103329.7, 103396.9, 
    103454.7, 103506, 103555.2, 103600.4, 103645.6, 103682.9, 103716.2, 
    103748.8,
  102913.1, 103020.5, 103112.2, 103196.6, 103272.7, 103344.3, 103406.5, 
    103462.5, 103511.4, 103557, 103596.2, 103633, 103666, 103693.3, 103717.8,
  102914.1, 103021.1, 103114.9, 103199.1, 103276.9, 103346.7, 103407.1, 
    103458.1, 103501.7, 103542.2, 103572.7, 103602.6, 103629.5, 103650.6, 
    103666.4,
  102913.7, 103019, 103116.6, 103198.2, 103273.6, 103342.2, 103392.1, 
    103438.9, 103476.2, 103507.1, 103533.5, 103555.9, 103574.9, 103590.6, 
    103603.6,
  102911.7, 103013.3, 103113.1, 103190.1, 103265.4, 103322, 103365.9, 
    103403.3, 103435.5, 103460.4, 103479.6, 103495.1, 103506.2, 103515.1, 
    103523.4,
  102087.7, 102114, 102080.5, 102106.2, 102141.3, 102196.4, 102264.3, 
    102324.9, 102395.7, 102490.8, 102588.2, 102699.7, 102795.6, 102890.6, 
    102985.7,
  102281.1, 102277.5, 102294, 102300.8, 102324.6, 102360.8, 102416.9, 
    102475.8, 102547.4, 102627.1, 102705.5, 102793.7, 102875.1, 102963.2, 
    103047.3,
  102381.6, 102396, 102422.8, 102427.6, 102443.7, 102483.6, 102537.4, 
    102592.8, 102656.2, 102721.8, 102790.2, 102872.1, 102951.6, 103032.8, 
    103104.3,
  102468.3, 102529.4, 102543.4, 102564, 102572.3, 102619.9, 102662.6, 
    102715.3, 102768.8, 102821.6, 102882.3, 102953, 103018.7, 103084.4, 103148,
  102560, 102620.1, 102629.2, 102669.8, 102683.4, 102731, 102764.2, 102810, 
    102852.5, 102902.3, 102956, 103017, 103077.3, 103133.4, 103191.7,
  102634.5, 102686.2, 102713.2, 102755.8, 102783.5, 102819, 102849.2, 
    102889.5, 102931.5, 102977.8, 103024.4, 103073.6, 103126.2, 103170.1, 
    103224.6,
  102698.2, 102730.9, 102786.7, 102819, 102849.9, 102879.2, 102912.9, 
    102949.1, 102990.2, 103029.5, 103073.4, 103114.8, 103157.7, 103200.6, 
    103247.1,
  102742.6, 102771.3, 102835.5, 102860.2, 102898.8, 102923.3, 102958.7, 
    102993.4, 103033.1, 103068.7, 103103.7, 103138.4, 103179.8, 103220.1, 
    103260.9,
  102765.4, 102799.9, 102857, 102882.9, 102923.1, 102949.1, 102985.2, 
    103015.2, 103051.9, 103086.1, 103119.1, 103149.2, 103184.5, 103224.3, 
    103259.3,
  102774.7, 102813.4, 102862.7, 102892.4, 102929.9, 102959, 102995.2, 
    103020.3, 103055.9, 103087.9, 103118.6, 103147.6, 103180.2, 103211.1, 
    103234.9,
  101181.4, 101095.4, 101004.4, 100927.3, 100851, 100824.1, 100861, 101013.2, 
    101202.4, 101418.7, 101598.9, 101824.6, 102000.1, 102116.7, 102272.4,
  101236.6, 101159.5, 101083.3, 101031.8, 100981.8, 100965.5, 100997.5, 
    101169.1, 101397, 101570.4, 101706.1, 101895.4, 102030.7, 102155.5, 
    102295.6,
  101369.4, 101300.2, 101216.4, 101152.7, 101112.4, 101103.7, 101138.8, 
    101285.5, 101459.5, 101612.7, 101762.6, 101954.9, 102074.2, 102193.1, 
    102315,
  101474.7, 101405.7, 101329.6, 101268.1, 101244.9, 101241.6, 101291, 
    101428.5, 101596.3, 101752.7, 101859.7, 102022.5, 102121, 102241.2, 
    102339.3,
  101587.6, 101531.7, 101474.1, 101420.9, 101397.7, 101398.2, 101459.7, 
    101571.2, 101706.1, 101840.2, 101934.8, 102085.4, 102161.6, 102289.6, 
    102370.7,
  101697.9, 101660.8, 101606.5, 101563.5, 101546.7, 101564.1, 101635, 
    101733.4, 101845.9, 101953.2, 102029.4, 102148.3, 102212.7, 102329, 
    102393.7,
  101821.9, 101791.1, 101744.5, 101718.3, 101713.7, 101744.4, 101803.2, 
    101869, 101961.6, 102047.7, 102111.1, 102199.4, 102260.9, 102363.9, 
    102413.7,
  101952.1, 101926.2, 101893.4, 101873, 101875, 101903.7, 101949.2, 101996.2, 
    102085.1, 102139.6, 102186, 102253.9, 102311.6, 102385.9, 102426.2,
  102091.8, 102063.4, 102035.2, 102016.7, 102017.3, 102040.5, 102066.9, 
    102110.8, 102167.6, 102208.3, 102243.6, 102300.6, 102351.7, 102402.4, 
    102426.7,
  102210.4, 102188, 102161.3, 102145.8, 102141.1, 102156.4, 102174.8, 
    102208.5, 102243.9, 102269.5, 102301.6, 102346.7, 102378.4, 102407.2, 
    102414.4,
  100664.2, 100622.7, 100616, 100668.8, 100769.4, 100921, 101132.5, 101333, 
    101504.3, 101665.8, 101804.3, 101936.2, 102051.1, 102153.2, 102250.8,
  100628.1, 100561.6, 100544.3, 100563.6, 100645.7, 100782.4, 100993.7, 
    101226.5, 101418.1, 101594.6, 101739.8, 101874.9, 101994.7, 102102.6, 
    102200.5,
  100600.4, 100512.2, 100467.3, 100453.8, 100519.5, 100652.5, 100881.1, 
    101145.6, 101327.3, 101516.8, 101668, 101811.8, 101935.2, 102043.9, 
    102143.7,
  100587.3, 100474.1, 100400.6, 100360, 100397.9, 100524.3, 100753.1, 
    101049.5, 101243.7, 101448.3, 101606.6, 101754.5, 101881.7, 101992.5, 
    102089.1,
  100591.8, 100460.6, 100353.9, 100283.4, 100287, 100396.5, 100634.2, 
    100959.9, 101167.1, 101379.4, 101546.2, 101697.8, 101828.3, 101938.4, 
    102032.7,
  100612.1, 100466.7, 100337.4, 100224.7, 100198.8, 100265.9, 100550.3, 
    100885.1, 101118.1, 101317.2, 101495.8, 101646.7, 101779.1, 101890.2, 
    101980.9,
  100644.3, 100491.1, 100347.2, 100202.4, 100143.4, 100155.9, 100471.7, 
    100820.4, 101072.7, 101265.2, 101451.4, 101600.9, 101731.6, 101843.4, 
    101928.7,
  100683.1, 100528.3, 100381.2, 100222.7, 100131.9, 100107.2, 100431.1, 
    100802.1, 101053.3, 101230.8, 101412.5, 101567.5, 101686.2, 101799.5, 
    101878.9,
  100729, 100575.2, 100431.8, 100274.6, 100180.2, 100152.2, 100426.6, 
    100801.2, 101048.6, 101220.4, 101381.5, 101545.1, 101647, 101758.4, 
    101828.3,
  100781.3, 100630.6, 100492.5, 100352.8, 100271.9, 100260.4, 100474.6, 
    100841.2, 101055.7, 101232.2, 101366.5, 101530.7, 101615.7, 101720.9, 
    101780.2,
  101637, 101717, 101772, 101838.6, 101897.1, 101956.6, 102010.4, 102061.7, 
    102110.2, 102154.5, 102195.9, 102235.3, 102273.3, 102310.2, 102344.9,
  101543, 101612.9, 101671.5, 101742.5, 101808.1, 101874.3, 101935, 101990.5, 
    102043.9, 102092.9, 102138.6, 102180.4, 102220.3, 102259.2, 102295.1,
  101424.1, 101496.4, 101560.7, 101639.1, 101709.5, 101779.5, 101847, 
    101907.5, 101963.7, 102015.1, 102063.8, 102108.6, 102152, 102192.9, 
    102231.1,
  101287.7, 101359.7, 101430.3, 101514.5, 101594.2, 101672.2, 101746.4, 
    101813.5, 101875.8, 101933.5, 101986.6, 102033.5, 102077.6, 102119.1, 
    102158.4,
  101141.6, 101207.6, 101283.9, 101374.1, 101466.4, 101551.9, 101633.7, 
    101705.9, 101775.6, 101837.4, 101896.7, 101947.7, 101994.5, 102036.6, 
    102077.8,
  100982.9, 101036.4, 101112.4, 101211.4, 101315.8, 101415.1, 101510.6, 
    101591.8, 101667.6, 101735.2, 101798.3, 101854.9, 101906.2, 101952.3, 
    101995.8,
  100817.4, 100856.5, 100922.5, 101026.4, 101144.8, 101262.4, 101369.7, 
    101465.9, 101551.5, 101625.8, 101693.6, 101756, 101811.6, 101862.2, 
    101909.4,
  100655.3, 100678, 100725, 100824.9, 100952.4, 101097.6, 101223.6, 101332.5, 
    101427, 101513.5, 101586.8, 101654.8, 101714.3, 101766.4, 101813.1,
  100508.3, 100513.4, 100537.8, 100621.9, 100745.3, 100908.1, 101062.3, 
    101192.2, 101298.8, 101393.3, 101475.2, 101545.8, 101608.6, 101663.7, 
    101712.6,
  100381.4, 100367.7, 100377.2, 100442.7, 100555, 100713.8, 100892.6, 
    101044.5, 101164.4, 101273.3, 101360, 101437.9, 101500.3, 101557.6, 101605,
  102344.1, 102367.7, 102380.4, 102388.2, 102392.4, 102388, 102375.3, 102359, 
    102337.6, 102312.6, 102283.2, 102247.8, 102210, 102166.7, 102121.3,
  102331.5, 102345.7, 102361.2, 102374.5, 102372.2, 102374.8, 102372.9, 
    102365, 102351.9, 102335.4, 102313, 102284.9, 102253.4, 102218.1, 102181.5,
  102299.6, 102318, 102334.8, 102349, 102360.1, 102362.9, 102365.1, 102361.7, 
    102352.2, 102339.9, 102320.4, 102298.7, 102270.8, 102241.2, 102208.7,
  102264.7, 102283.3, 102301.7, 102317, 102329.1, 102339.7, 102345.4, 
    102355.3, 102351.3, 102342.9, 102331.9, 102312.4, 102297.3, 102268, 
    102242.9,
  102228, 102247.5, 102267.5, 102288.5, 102304.7, 102319.1, 102331.7, 
    102337.7, 102342.2, 102341.5, 102339.8, 102330.1, 102318.1, 102299.7, 
    102280.9,
  102182.7, 102203.8, 102229, 102252, 102275.3, 102295.3, 102312.7, 102328.6, 
    102344.7, 102355.9, 102357.1, 102353, 102348.7, 102328.8, 102312.8,
  102135, 102161.3, 102188.7, 102217.1, 102242.4, 102266.8, 102290, 102307.6, 
    102322.9, 102344.9, 102348.3, 102351.2, 102348.9, 102340.3, 102327.7,
  102084, 102112, 102142.1, 102171.8, 102203.4, 102229.8, 102255.3, 102280.6, 
    102298.5, 102320.7, 102333.6, 102335.9, 102335.3, 102329.7, 102326.6,
  102029.6, 102058.8, 102091.9, 102127.2, 102162.8, 102197.6, 102226.1, 
    102248.6, 102269.8, 102291.4, 102307.2, 102313.4, 102320.3, 102313.5, 
    102303.4,
  101968.5, 102002.1, 102036.6, 102073.1, 102107.2, 102145.1, 102178.9, 
    102207.4, 102232.5, 102253.9, 102267.7, 102275.4, 102279.4, 102275, 
    102263.4,
  102349.1, 102307, 102253.7, 102185.6, 102103, 102015.7, 101891.3, 101794.1, 
    101670.5, 101537.1, 101376.8, 101239.8, 101093.5, 100937.9, 100812.7,
  102402.3, 102369.5, 102331.5, 102281.3, 102216, 102139.8, 102047.6, 
    101953.7, 101826, 101710.2, 101576.8, 101456.5, 101326, 101180.8, 101055.6,
  102454.7, 102428.8, 102397.2, 102353.3, 102300.1, 102231.5, 102152.3, 
    102068.2, 101965.8, 101865.4, 101754.5, 101645.3, 101524.7, 101409.2, 
    101289.4,
  102500.9, 102482, 102455.1, 102422, 102379, 102328.9, 102265, 102196.5, 
    102110.4, 102017.9, 101914.5, 101818.9, 101713.9, 101611.2, 101508.2,
  102553.9, 102536.9, 102515.7, 102487.8, 102449.4, 102406, 102355.9, 
    102297.2, 102222.2, 102142.6, 102053.2, 101966.2, 101877.5, 101792.1, 
    101707.1,
  102604.3, 102592.3, 102576.9, 102555.7, 102525.8, 102490.2, 102445.5, 
    102395, 102338.6, 102267, 102185, 102100.9, 102023.4, 101945, 101867.7,
  102656, 102648.6, 102636.4, 102616.4, 102592, 102562.4, 102528.5, 102485.1, 
    102428.6, 102376.7, 102309.3, 102233.3, 102160.6, 102087.8, 102012.8,
  102697.6, 102697.7, 102691.6, 102674.8, 102654.3, 102624.9, 102591.8, 
    102563.1, 102517.5, 102465.7, 102405.4, 102345.7, 102278.2, 102215, 
    102147.5,
  102734.1, 102745.1, 102750.7, 102746.4, 102731.6, 102709.5, 102682.1, 
    102638.2, 102592.2, 102540.5, 102484.8, 102432.8, 102369.6, 102313.1, 
    102249.7,
  102751.4, 102771.4, 102783.1, 102780.9, 102770.6, 102754.1, 102733.5, 
    102692.6, 102652.5, 102606.3, 102552.5, 102503.4, 102443.1, 102384.2, 
    102323.7,
  101860.1, 101659, 101500.9, 101337.7, 101176, 101050.1, 100939.5, 100887.5, 
    100837.7, 100792.1, 100740.2, 100663.1, 100571.5, 100485.9, 100413.6,
  101974.4, 101822.2, 101677.2, 101453.6, 101315, 101180.7, 101056.5, 
    100982.1, 100916.5, 100855.8, 100793.6, 100725.4, 100641.4, 100550.1, 
    100471.1,
  102132.8, 101992.8, 101856.7, 101640.3, 101496.8, 101297.2, 101185.9, 
    101094.4, 101012.5, 100945.7, 100871.3, 100797, 100709.4, 100616.3, 
    100530.7,
  102267.1, 102154.3, 102026.5, 101834.7, 101681.6, 101483.7, 101363, 101250, 
    101152.1, 101067.3, 100982, 100897.4, 100808.2, 100718.6, 100634.1,
  102386, 102286.2, 102177.6, 102044.6, 101885, 101716.2, 101582.9, 101452.4, 
    101340.2, 101239.7, 101141.5, 101045.2, 100945.9, 100854.6, 100770.1,
  102504.5, 102421.5, 102316.2, 102212.5, 102082.8, 101938, 101801.7, 
    101676.5, 101561.8, 101446.1, 101332.3, 101227.4, 101129.4, 101037.7, 
    100960.7,
  102617, 102541, 102457.9, 102359.2, 102253.2, 102137.3, 102016.4, 101896.3, 
    101783.8, 101672.1, 101556.1, 101441.4, 101337.4, 101246.8, 101171.5,
  102732.2, 102667.8, 102596.2, 102508.9, 102416.1, 102315.2, 102212.2, 
    102107.3, 101995.1, 101887.8, 101775.5, 101662.1, 101554.4, 101462.5, 
    101387.5,
  102833.2, 102784.5, 102729.4, 102658.2, 102576.5, 102487.4, 102393.5, 
    102299.7, 102201.3, 102097.6, 101989.2, 101882, 101777.1, 101685.3, 
    101604.5,
  102920.2, 102884.5, 102840.5, 102784.4, 102719.3, 102641.3, 102560.8, 
    102472.9, 102385.2, 102289.4, 102187.4, 102085.2, 101986.8, 101897.2, 
    101816.6,
  101410.8, 101327.8, 101293.4, 101279.8, 101235.7, 101217.6, 101183.3, 
    101144.1, 101107.4, 101078.2, 101053.9, 101044.6, 101044.3, 101058.4, 
    101072,
  101417.2, 101296.7, 101269.2, 101240.6, 101217.6, 101209.9, 101180.8, 
    101140.6, 101101.4, 101070, 101044.3, 101029.2, 101025.3, 101027, 101037.4,
  101425.1, 101292.3, 101282.7, 101209.9, 101203.8, 101194.5, 101175.5, 
    101139.7, 101100.5, 101069.2, 101038.4, 101023.2, 101016.7, 101010.9, 
    101009.3,
  101438.5, 101362.7, 101270.9, 101171.2, 101175.3, 101164.3, 101163.8, 
    101138.6, 101107.8, 101078.1, 101046.6, 101024.6, 101008.2, 100996.9, 
    100989.4,
  101546.7, 101456.1, 101282.3, 101190, 101164.8, 101146.5, 101146.3, 
    101130.9, 101110, 101080.6, 101042.4, 101012.3, 100984.8, 100968.4, 
    100957.1,
  101680.7, 101564.9, 101384.7, 101273.9, 101202.8, 101164.6, 101154.6, 
    101136.5, 101107, 101071.8, 101030.3, 100989.6, 100953.7, 100931, 100922,
  101856.3, 101711.5, 101537.8, 101398.4, 101291.3, 101232.5, 101191.5, 
    101166.6, 101128.2, 101081.6, 101028.2, 100974.3, 100929, 100900.5, 
    100894.1,
  102041.9, 101874.6, 101706, 101552.1, 101431.6, 101337.4, 101274.7, 
    101226.4, 101182.1, 101124.5, 101059.2, 100991, 100935.3, 100896.9, 
    100885.3,
  102215.7, 102064.8, 101900.9, 101736.4, 101610.1, 101497.2, 101410.5, 
    101331.6, 101274.6, 101210, 101132.3, 101050.3, 100978.1, 100926.6, 
    100903.5,
  102377.4, 102248.9, 102106.2, 101946.6, 101825.5, 101698.3, 101599.2, 
    101500.8, 101412.6, 101339.5, 101251.1, 101157.1, 101066.4, 100995.9, 
    100951.2,
  101282.1, 101304.4, 101312.6, 101306.6, 101306.6, 101301.3, 101302.7, 
    101300.7, 101293.2, 101280.1, 101259.3, 101230.7, 101198.1, 101155.1, 
    101108.5,
  101266.1, 101287, 101290.1, 101285.3, 101279, 101265, 101258.1, 101252.4, 
    101246.5, 101235.2, 101211.2, 101180.2, 101135.9, 101089.3, 101037.2,
  101226.7, 101255.2, 101267.1, 101269.3, 101251.5, 101232, 101220.5, 101215, 
    101209.2, 101193.8, 101161.1, 101122.2, 101073, 101023, 100962.7,
  101173.6, 101231.7, 101242, 101256.3, 101241, 101222.5, 101199.9, 101185.6, 
    101167.6, 101149.7, 101116.1, 101071.6, 101013, 100953.8, 100883.2,
  101125.5, 101197.6, 101201.6, 101231, 101223.2, 101211.2, 101186.8, 
    101165.8, 101138.6, 101109.2, 101066.8, 101016.9, 100957.9, 100890.9, 
    100812.6,
  101073.9, 101169.2, 101161, 101201.3, 101191.7, 101190.3, 101163.8, 
    101141.2, 101107.4, 101071.1, 101021.9, 100967.8, 100903.6, 100829.5, 
    100744.8,
  101038.6, 101133.1, 101118.8, 101156.5, 101151.4, 101151.2, 101128, 
    101103.5, 101066.4, 101027.1, 100973.2, 100917.8, 100848.6, 100770, 
    100678.9,
  101087.5, 101093.2, 101092.9, 101113.9, 101106.8, 101105.4, 101081.6, 
    101059.2, 101022.4, 100980.9, 100925.6, 100866.1, 100796.2, 100713.9, 
    100615.5,
  101193.9, 101097, 101084.1, 101079.4, 101063.6, 101050.4, 101027.7, 
    101003.8, 100971.8, 100934.2, 100878.5, 100812.9, 100740.4, 100657.8, 
    100556.8,
  101340.9, 101184.8, 101107.9, 101071.6, 101039.2, 101004.5, 100973.1, 
    100945.4, 100920, 100881.7, 100829.4, 100763.3, 100686.3, 100603.9, 
    100502.2,
  101323.6, 101309.3, 101300.9, 101293.2, 101298.4, 101304.4, 101316.6, 
    101330.1, 101347.2, 101366.8, 101389.6, 101417.7, 101452, 101484.2, 
    101516.7,
  101305.1, 101284.1, 101266, 101253.4, 101254.1, 101255, 101259.3, 101266.4, 
    101278.1, 101290.6, 101308.2, 101333, 101360.7, 101388.6, 101419,
  101279.6, 101254.8, 101230.3, 101210.7, 101202.1, 101197, 101196.2, 
    101194.7, 101200.5, 101206.7, 101218.9, 101235.7, 101254.6, 101276.4, 
    101298.8,
  101261.4, 101230.1, 101199, 101173.1, 101153.8, 101141.6, 101132.3, 
    101125.5, 101120.5, 101119.8, 101122.5, 101130.9, 101139.5, 101150.9, 
    101165.7,
  101238.2, 101202.9, 101164.2, 101135.3, 101105.9, 101086.7, 101068.4, 
    101053.2, 101038.2, 101028.5, 101022.2, 101019.2, 101015.4, 101016.8, 
    101020.4,
  101214.3, 101174, 101132.1, 101095.6, 101059.5, 101028.8, 101003, 100977, 
    100953.3, 100934.2, 100916.7, 100901.1, 100882.8, 100870.1, 100863.2,
  101186.2, 101144.5, 101099.5, 101054.2, 101010.2, 100973.4, 100935.9, 
    100902.2, 100868.5, 100836.7, 100808.8, 100779.2, 100747.6, 100717.1, 
    100696.6,
  101148.4, 101116.1, 101061.9, 101016.3, 100964.8, 100919.4, 100870.9, 
    100827.1, 100782, 100738.5, 100696.9, 100654.4, 100603.6, 100557.4, 
    100521.8,
  101111, 101083.1, 101026.5, 100977.9, 100917.5, 100863.7, 100804.9, 
    100751.5, 100694.7, 100640, 100583.1, 100525.1, 100456.7, 100393, 100340,
  101087.5, 101041.2, 100990.6, 100938.5, 100873.2, 100810.5, 100742.6, 
    100677.5, 100608.7, 100540.2, 100468, 100392, 100306.5, 100225.6, 100153,
  101848.2, 101898.4, 101945.6, 101991.9, 102031.4, 102068.3, 102100.2, 
    102125.7, 102146.1, 102164.6, 102180.2, 102196.8, 102211.7, 102224.7, 
    102237.3,
  101839.5, 101885.1, 101930.3, 101974.4, 102009.5, 102038.4, 102063.5, 
    102084.9, 102098.6, 102110.3, 102119.3, 102132.2, 102139.9, 102149.2, 
    102156.3,
  101814.2, 101856.1, 101895.4, 101933.5, 101966.2, 101991.7, 102011.5, 
    102027.3, 102036.8, 102044, 102049.8, 102057.1, 102060.8, 102065.7, 102068,
  101794.1, 101829.8, 101866.7, 101899.4, 101925.5, 101945.3, 101960.3, 
    101966.8, 101969.8, 101968, 101970.5, 101967.9, 101966.3, 101964.1, 
    101962.5,
  101763.5, 101794.2, 101822.8, 101849.1, 101869.1, 101883.1, 101893, 101893, 
    101891.4, 101884, 101881, 101872.3, 101865.5, 101857, 101850,
  101729.1, 101755.6, 101779.9, 101801.8, 101813.6, 101821.7, 101823.4, 
    101816.1, 101805.8, 101790.8, 101780.1, 101763.4, 101750.2, 101734.6, 
    101721.6,
  101687.2, 101706.5, 101724.5, 101739.1, 101745.1, 101747, 101741.1, 
    101727.8, 101709.4, 101688.7, 101669, 101645.8, 101623.1, 101601.3, 
    101581.7,
  101648.9, 101656.5, 101672.2, 101677.9, 101678.7, 101671.3, 101658, 
    101634.8, 101607.5, 101576.1, 101545.4, 101511.5, 101481, 101452, 101425.5,
  101606.2, 101607.6, 101613.1, 101611.4, 101602.8, 101588.9, 101566.4, 
    101534.2, 101495.1, 101451.9, 101409.7, 101365.4, 101324.3, 101286.7, 
    101251.2,
  101563.1, 101557.8, 101553.1, 101543.4, 101526.2, 101504.2, 101471.1, 
    101429, 101375.7, 101319.4, 101263.3, 101206.3, 101154.6, 101106.2, 
    101062.7,
  102204.5, 102240.5, 102254.6, 102278.6, 102294.1, 102309.4, 102317.7, 
    102306.5, 102293, 102280.3, 102260.1, 102243.3, 102219.7, 102195.7, 
    102169.8,
  102256.9, 102277.7, 102298.8, 102308.5, 102318.4, 102323, 102323.5, 
    102307.1, 102284.9, 102265.7, 102241.6, 102212.1, 102180.3, 102146, 
    102109.5,
  102281.9, 102291.1, 102313.5, 102319.7, 102326.7, 102322.5, 102307.8, 
    102287.3, 102261.1, 102235, 102201.5, 102168.8, 102130.1, 102093.3, 
    102053.5,
  102310.1, 102314, 102330.5, 102331.2, 102325.5, 102310.6, 102290.8, 
    102262.4, 102233.5, 102198.9, 102162.5, 102118, 102071.2, 102026.1, 
    101981.9,
  102317.7, 102319.6, 102332.2, 102325.3, 102311.4, 102288.8, 102261.9, 
    102230.2, 102195.6, 102154.8, 102108, 102058.5, 102009.8, 101959.4, 
    101909.2,
  102322.1, 102322.8, 102326.1, 102307.2, 102292.8, 102261.9, 102230.9, 
    102195.1, 102149.9, 102101.6, 102050.3, 101996.4, 101940.9, 101882.2, 
    101827.7,
  102316.1, 102311.1, 102306.7, 102284.2, 102262.8, 102229.1, 102193, 
    102149.3, 102097.8, 102045.7, 101988.2, 101928.1, 101865.2, 101803.2, 
    101741.9,
  102309.2, 102297, 102284.4, 102261, 102237.1, 102191.3, 102149.9, 102097.7, 
    102041.5, 101981.9, 101917.6, 101850.8, 101783.6, 101716.2, 101650.5,
  102289.8, 102275.9, 102257.8, 102232.6, 102201, 102145.6, 102098.4, 
    102039.2, 101975.7, 101910.7, 101842, 101768.5, 101696.5, 101626.7, 
    101556.8,
  102273.7, 102255.4, 102233.7, 102197.9, 102152.4, 102095.6, 102040.4, 
    101973.9, 101906.5, 101833.3, 101758.5, 101682.6, 101608.1, 101533, 101455,
  101589.2, 101571.9, 101530.2, 101478, 101438.1, 101433.2, 101476, 101462.7, 
    101569.7, 101645.9, 101623.5, 101679.2, 101696, 101710.7, 101718.7,
  101668.1, 101650.9, 101618.3, 101584.3, 101568, 101545.5, 101601.9, 
    101656.7, 101706.9, 101681.9, 101654.8, 101679.6, 101681.9, 101680, 101674,
  101729.6, 101713.4, 101690.8, 101680.2, 101673.3, 101682.3, 101708.5, 
    101691.8, 101708.1, 101687.1, 101689.2, 101677.3, 101661.9, 101648, 
    101635.5,
  101802.5, 101789.5, 101768.3, 101771.7, 101764, 101773.1, 101770.9, 101759, 
    101764, 101720.5, 101702.2, 101666.3, 101637.9, 101608.7, 101582.3,
  101871.7, 101857.7, 101837.1, 101856.4, 101852.5, 101840.9, 101820.3, 
    101795.2, 101773.9, 101727.6, 101696.3, 101645.5, 101606.7, 101564.6, 
    101524.7,
  101944.1, 101929.1, 101904.3, 101930.6, 101917.7, 101887.9, 101857.8, 
    101832.1, 101787.2, 101737.2, 101680.4, 101618.2, 101562.8, 101507.6, 
    101451,
  102012.6, 101996, 101967.1, 101994.6, 101970.5, 101925.8, 101881.4, 
    101844.8, 101783.5, 101726.4, 101648.7, 101580.2, 101509.8, 101443.9, 
    101370.5,
  102087.7, 102060.3, 102034.4, 102047.2, 102010.5, 101957.7, 101900.2, 
    101852.5, 101778.5, 101703.9, 101613.2, 101530.6, 101446.9, 101364.2, 
    101276.2,
  102156.4, 102123, 102094.8, 102095.1, 102046, 101977.3, 101907.2, 101845.2, 
    101760.1, 101667, 101569.1, 101470.3, 101374, 101277, 101177.6,
  102218.9, 102182.1, 102152.5, 102129.1, 102067.2, 101985.2, 101909.5, 
    101830.7, 101730.3, 101625, 101514.2, 101399.6, 101292, 101177.8, 101076.1,
  100952.6, 100821.1, 100691.4, 100542.5, 100451.9, 100397.8, 100639.4, 
    101003.6, 101146, 101310.2, 101448.3, 101522.6, 101596.9, 101645, 101684.1,
  101009.1, 100883.2, 100759.1, 100595.1, 100491.7, 100412, 100596, 100978.8, 
    101164.8, 101272.7, 101401.8, 101476.8, 101550.3, 101594.2, 101628.8,
  101085.2, 100978.5, 100864.5, 100706.8, 100614.6, 100499.4, 100606.1, 
    100932.9, 101156.9, 101241.4, 101365.2, 101439.8, 101504.5, 101541, 101570,
  101146.5, 101042.3, 100934, 100815, 100722.4, 100651.9, 100746.3, 100971.4, 
    101188, 101249.6, 101353.3, 101411.8, 101467.8, 101492, 101516.2,
  101212.2, 101113.4, 101015, 100924.1, 100843.5, 100820.5, 100883.7, 
    101009.3, 101221.6, 101254.7, 101355, 101391.8, 101435.9, 101447.1, 
    101461.1,
  101260.2, 101178.2, 101077.6, 101007.7, 100937.3, 100943.6, 101018.8, 
    101120.5, 101278.4, 101278.4, 101360.6, 101380, 101407.3, 101409, 101410.5,
  101312.6, 101244, 101136.6, 101083.8, 101029.1, 101066.8, 101132.6, 
    101211.8, 101312.6, 101306.4, 101361.5, 101369.5, 101378.5, 101373.8, 
    101365.4,
  101372.5, 101282.4, 101192.5, 101140.5, 101101.5, 101160.8, 101226.2, 
    101304, 101344.8, 101341.5, 101359.6, 101359.8, 101352, 101337.9, 101320.4,
  101432.9, 101315.2, 101249.1, 101191.5, 101169, 101242.6, 101302.7, 
    101367.9, 101361.8, 101361.5, 101354.7, 101344.4, 101321.8, 101297.6, 
    101270.5,
  101492.6, 101357.8, 101293.4, 101240.8, 101227.2, 101307.4, 101359.3, 
    101410.4, 101385.1, 101376.7, 101347.5, 101324.5, 101285.1, 101254.3, 
    101224,
  100840.8, 100831, 100797.4, 100810, 100855.1, 100970.3, 101177.3, 101349.6, 
    101468.5, 101576.7, 101652.8, 101723.9, 101777.2, 101819.7, 101852.9,
  100796.1, 100789.1, 100800.1, 100835.9, 100889.3, 100958.2, 101128.6, 
    101312.2, 101435.9, 101551.6, 101629.9, 101705.1, 101759.2, 101806, 
    101842.6,
  100867.9, 100815, 100808, 100845.7, 100904, 100956.4, 101094.5, 101286.8, 
    101406.2, 101522.6, 101610.7, 101689.8, 101746.7, 101798.2, 101835.7,
  100938.5, 100887.8, 100856.7, 100874.1, 100942, 100991.5, 101101.6, 
    101278.6, 101392.6, 101506.9, 101593.5, 101669.4, 101727.6, 101779.4, 
    101815.4,
  101023.3, 100963.2, 100936.6, 100933.8, 100969.9, 101025.4, 101112.6, 
    101274.4, 101387, 101491.8, 101580.7, 101652.7, 101708.8, 101757.8, 
    101791.7,
  101054.2, 101047.6, 100988.3, 100983.1, 100996.2, 101058.5, 101142.1, 
    101290.2, 101402.9, 101482.9, 101567.6, 101634.4, 101685, 101730.1, 
    101761.2,
  101070.3, 101126.6, 101020.7, 101021.9, 101023.9, 101083.3, 101158.2, 
    101299.6, 101416, 101474.8, 101551.4, 101613.1, 101658.8, 101704.4, 
    101729.2,
  101127, 101174.7, 101049.8, 101054.4, 101046.4, 101111.3, 101179.6, 
    101330.1, 101427.8, 101470.2, 101527.9, 101584.8, 101623.4, 101665.9, 
    101687.6,
  101186.1, 101219.6, 101088.2, 101087.5, 101072.3, 101134.2, 101201.1, 
    101352.6, 101423.2, 101459.7, 101505.7, 101551.9, 101583.4, 101620.2, 
    101637.1,
  101238.7, 101229.3, 101152.2, 101108.4, 101103.2, 101157.8, 101236, 
    101372.6, 101418.1, 101448.2, 101478.6, 101512.3, 101538.9, 101569.4, 
    101578.4,
  101153.7, 101167.4, 101226.4, 101325.6, 101450.5, 101559, 101683.6, 
    101762.4, 101841.7, 101909.5, 101969.8, 102020.6, 102063.8, 102094.3, 
    102110.8,
  101177.1, 101207.4, 101286.9, 101379.3, 101494.4, 101597, 101730.3, 
    101809.5, 101897.3, 101969.6, 102033.4, 102084.1, 102123.5, 102149.6, 
    102170.1,
  101261, 101290.3, 101364.3, 101435, 101569.7, 101654.5, 101785.5, 101852.7, 
    101939.4, 102009.5, 102073.1, 102128.7, 102175.5, 102210.6, 102231.7,
  101322.8, 101358.8, 101436.4, 101506.2, 101647.7, 101722.8, 101843.5, 
    101909.1, 101998, 102067.6, 102129.6, 102183.1, 102228, 102261.7, 102285,
  101380.2, 101440.6, 101503.6, 101596.6, 101710.7, 101791.6, 101907, 
    101970.6, 102050.2, 102114.5, 102174.7, 102229.4, 102274.3, 102313.3, 
    102342.2,
  101443.1, 101506.1, 101578.8, 101661.5, 101784.2, 101856.7, 101965.1, 
    102031.8, 102114.4, 102173.6, 102230.3, 102282, 102325.9, 102366.2, 
    102391.2,
  101497.2, 101567.9, 101654, 101723.8, 101850.1, 101915, 102024, 102100.4, 
    102178, 102233.4, 102285.9, 102330.8, 102373.8, 102405, 102444.1,
  101550, 101628.7, 101711.1, 101787.7, 101903.6, 101982.3, 102084.2, 
    102168.1, 102239.8, 102294.8, 102346.2, 102392.4, 102428.4, 102462.4, 
    102493.6,
  101580.8, 101682.4, 101767, 101861.6, 101950, 102045.7, 102139.7, 102225.5, 
    102296.7, 102356.1, 102404.6, 102449.2, 102484.1, 102510.4, 102525.6,
  101604.5, 101727.9, 101801.9, 101918.6, 102000.6, 102102.9, 102192.2, 
    102277.8, 102351.9, 102409.3, 102460, 102508.5, 102541.9, 102559.5, 
    102562.4,
  101459.5, 101478.7, 101512.1, 101532.8, 101549.5, 101598.4, 101624.9, 
    101656.2, 101668.6, 101673.1, 101718.4, 101731.3, 101745.1, 101751.6, 
    101748.1,
  101555.1, 101591.7, 101632.8, 101661.8, 101683, 101710.1, 101723.1, 
    101774.6, 101804.8, 101813.9, 101854.1, 101860.1, 101872.5, 101874, 
    101866.3,
  101597.9, 101656.6, 101708.8, 101751.5, 101786.8, 101837.2, 101869.4, 
    101920, 101911.8, 101930.9, 101963.7, 101964.9, 101978, 101977.7, 101971,
  101659.2, 101736.7, 101805.4, 101861, 101897.8, 101944.8, 101970.2, 
    102013.8, 102020.9, 102063, 102081.7, 102089.5, 102099.7, 102092.6, 
    102084.2,
  101709.1, 101798.4, 101879.5, 101946.6, 102004.2, 102058.2, 102094.5, 
    102131.9, 102148.5, 102179.9, 102194, 102206.4, 102211.6, 102203.8, 
    102188.7,
  101742.7, 101849.4, 101954.6, 102038.7, 102105, 102156.9, 102203.7, 
    102233.3, 102255.9, 102288.5, 102311, 102323.3, 102325.9, 102315.9, 
    102296.3,
  101780.5, 101897.8, 102030.2, 102118.1, 102196, 102255.4, 102299, 102336, 
    102373.3, 102405.9, 102424, 102430.1, 102433.4, 102422.1, 102397.8,
  101818.1, 101950.7, 102092.6, 102190, 102281.9, 102349, 102402.1, 102450, 
    102483.9, 102506.2, 102526.4, 102533.1, 102533.8, 102516.4, 102488.1,
  101852.6, 102008.9, 102157.6, 102262.2, 102361.2, 102432.5, 102493.2, 
    102540.2, 102577.1, 102605.3, 102627, 102634.5, 102630.1, 102606.5, 
    102569.6,
  101939.4, 102077.9, 102222.4, 102336.4, 102439.6, 102519.3, 102586.5, 
    102641.5, 102683.8, 102710.8, 102726.2, 102724.9, 102714.8, 102691.8, 
    102654.3,
  101406, 101379.7, 101368.6, 101330.5, 101286.8, 101225.4, 101152.9, 
    101057.6, 100943.2, 100814.2, 100674.5, 100526.3, 100369.2, 100204, 100024,
  101439.6, 101433, 101433.1, 101410.6, 101377.5, 101327.4, 101261.8, 
    101177.5, 101070.6, 100947.2, 100810.9, 100668.5, 100516.2, 100351.5, 
    100171,
  101448.1, 101477.6, 101482.1, 101476.6, 101456.8, 101420.1, 101364.6, 
    101293.9, 101202.8, 101089, 100957.6, 100815, 100660.6, 100496.4, 100320.2,
  101440.6, 101494.3, 101516.8, 101537.2, 101527.7, 101509.1, 101467.5, 
    101406.4, 101325.9, 101225, 101103.1, 100966.5, 100818.9, 100656.9, 
    100480.3,
  101382.3, 101482.7, 101520.3, 101577.3, 101589.5, 101588.2, 101561.3, 
    101520.1, 101451.5, 101362.9, 101251.4, 101122.8, 100977.8, 100823.1, 
    100654.3,
  101271, 101444.7, 101505, 101601.6, 101627.4, 101660.4, 101646.5, 101621.4, 
    101569.1, 101494.2, 101395.6, 101277.2, 101141.1, 100990.6, 100828.2,
  101088.9, 101348.2, 101444.7, 101601.7, 101651.6, 101710.6, 101723.1, 
    101720.1, 101681.4, 101622.4, 101537.6, 101429.6, 101301.9, 101160.8, 
    101006.2,
  100899.9, 101231.2, 101377.1, 101572.5, 101669.9, 101758.1, 101785.7, 
    101804.3, 101784.4, 101742.8, 101671.9, 101580.2, 101464.4, 101332.3, 
    101185,
  100769.3, 101130.7, 101326.8, 101544.9, 101677.3, 101790.7, 101839.3, 
    101875.5, 101873.5, 101852.1, 101796.3, 101719.9, 101615.5, 101496.1, 
    101359.4,
  100866.8, 101133.5, 101336.7, 101550.2, 101699.3, 101827.1, 101902.2, 
    101946, 101961.5, 101951.6, 101914.6, 101850.5, 101762.4, 101652, 101525.8,
  100979.1, 100886.1, 100768.6, 100646.7, 100515.7, 100384.9, 100272.9, 
    100171.7, 100079.9, 99982.82, 99886.05, 99780.74, 99681.13, 99609.93, 
    99557.08,
  101004.3, 100904, 100782.7, 100659.8, 100532.4, 100399.7, 100285.2, 
    100171.4, 100066.5, 99955.22, 99849.88, 99745.88, 99656.93, 99576.54, 
    99508.94,
  101018.6, 100922.5, 100806.7, 100689.8, 100558.1, 100425.7, 100302.3, 
    100184.3, 100073.5, 99952.47, 99835.74, 99723.59, 99616.61, 99515.63, 
    99426.73,
  101027.6, 100939.1, 100830.4, 100719.9, 100584.9, 100450.3, 100320.8, 
    100195.5, 100070.3, 99937.09, 99805.61, 99685.05, 99567.09, 99455.04, 
    99353.32,
  101034, 100953.2, 100850.9, 100749.8, 100622.3, 100482.2, 100348.8, 
    100224.8, 100090.6, 99949.05, 99805.32, 99671.59, 99539.52, 99410.62, 
    99288.83,
  101011.9, 100950, 100859.7, 100766.6, 100651.5, 100515.8, 100384.5, 100256, 
    100115, 99969.52, 99813.87, 99662.94, 99516.41, 99375.27, 99234.21,
  100968.6, 100925.3, 100846.4, 100772.8, 100675.5, 100552.6, 100427.1, 
    100300.9, 100160.1, 100008, 99843.2, 99675.94, 99510.81, 99353.7, 99192.66,
  100909.3, 100882.2, 100813, 100766.9, 100681.4, 100585.5, 100474.1, 
    100354.9, 100215, 100058.2, 99884.86, 99704.28, 99522.07, 99348.46, 
    99169.97,
  100858.3, 100838.7, 100785, 100760.5, 100691, 100613.6, 100516.6, 100410.7, 
    100278, 100123.2, 99944.2, 99755.79, 99559.23, 99366.66, 99169.77,
  100842.6, 100813.2, 100765.4, 100754.6, 100713.6, 100654.9, 100565.2, 
    100470, 100344.2, 100192.8, 100014.2, 99819.62, 99614.32, 99406.32, 
    99191.43,
  101043.2, 101030.6, 101015, 101014, 101022.6, 101039.6, 101054.8, 101070.1, 
    101084, 101100.8, 101119.5, 101138.3, 101166.6, 101190.2, 101209.8,
  101005.5, 100981.6, 100967.4, 100968, 100973.3, 100985.7, 100997.5, 
    101011.5, 101023.2, 101038, 101053.3, 101072, 101085.5, 101100, 101110.1,
  100970.8, 100943.2, 100927.3, 100917.4, 100916.4, 100931, 100939.7, 
    100951.7, 100960.3, 100971.5, 100980.8, 100988.9, 100996.1, 101004, 
    101012.5,
  100937.1, 100901.4, 100879.2, 100867, 100864.9, 100873.1, 100878.1, 
    100886.8, 100892.2, 100899, 100905.7, 100907.9, 100912, 100914.7, 100914.6,
  100905.3, 100863.2, 100834.2, 100816.9, 100809.4, 100813.8, 100815.8, 
    100819.1, 100821.1, 100822.5, 100823.4, 100821, 100820.2, 100818, 100816.2,
  100872.1, 100824.8, 100789.9, 100767.1, 100751.7, 100748.6, 100750.5, 
    100746.4, 100745.2, 100742.1, 100738.7, 100732.9, 100731.9, 100727.4, 
    100720.2,
  100842.7, 100784.9, 100743.2, 100713.2, 100696.2, 100684.3, 100680.2, 
    100670.3, 100665.1, 100654.6, 100649.2, 100641.2, 100637.8, 100630.3, 
    100621.1,
  100814.6, 100750.1, 100701.1, 100658.3, 100637.4, 100611.7, 100606.9, 
    100592.3, 100581.9, 100567.2, 100556.4, 100545.6, 100539.2, 100525.5, 
    100509.4,
  100785.1, 100711.2, 100656, 100607.6, 100578.5, 100539.2, 100533.4, 
    100513.7, 100498.4, 100478.2, 100463.9, 100448.6, 100434.2, 100413.2, 
    100392.9,
  100759.2, 100674.7, 100614.9, 100561.3, 100519.2, 100471.1, 100462, 
    100434.5, 100413.9, 100389.2, 100371.4, 100347.3, 100324.8, 100297.2, 
    100265.3,
  102042.8, 102088, 102127, 102142.2, 102157.2, 102164.4, 102162.3, 102152.8, 
    102140.8, 102128.8, 102112.9, 102094.3, 102075.1, 102053, 102031.7,
  102049.6, 102082.4, 102117.3, 102128, 102135.4, 102133.1, 102126.8, 102115, 
    102099.8, 102081.1, 102057.4, 102030.9, 102006.2, 101983.6, 101963.8,
  102033.3, 102066.6, 102092.2, 102103, 102104.2, 102100, 102087.5, 102069.1, 
    102046.5, 102022.2, 101993.9, 101969.3, 101944.7, 101922.3, 101897.3,
  102018.7, 102060.4, 102078.9, 102079.5, 102078, 102064.6, 102047.8, 
    102024.3, 101995, 101963.3, 101932.8, 101902.5, 101876.3, 101847.1, 
    101817.5,
  101994.4, 102030.8, 102052.1, 102053.1, 102045.8, 102027.7, 102000.1, 
    101972.8, 101936.8, 101901.6, 101866.7, 101836.2, 101802.7, 101771.1, 
    101737.8,
  101975.9, 102006.2, 102020.9, 102023.6, 102007.7, 101987.9, 101951.8, 
    101920.3, 101877.6, 101837.4, 101800.6, 101766, 101728, 101689.5, 101645.3,
  101940.9, 101973.8, 101984.2, 101987, 101966.8, 101937.2, 101900.3, 
    101861.3, 101815.2, 101772.5, 101732.3, 101691.7, 101648.4, 101598.6, 
    101545.6,
  101911.2, 101944.4, 101950.4, 101944.5, 101915.6, 101888.2, 101848.3, 
    101801.5, 101752.3, 101705.5, 101662.5, 101615.3, 101559.1, 101500.2, 
    101435.6,
  101880.6, 101912.8, 101913.1, 101905, 101874.7, 101836.3, 101791.1, 
    101740.5, 101686.5, 101640.2, 101590.5, 101529.3, 101464.1, 101392.5, 
    101315.5,
  101849, 101877.3, 101872.8, 101857.4, 101825.8, 101786, 101735.8, 101679, 
    101623.7, 101570.3, 101508.4, 101439.9, 101359.9, 101275.3, 101182.3,
  102368.8, 102385.9, 102386.3, 102386.3, 102383.5, 102365.8, 102338.7, 
    102307.2, 102272.1, 102226.3, 102176, 102119.2, 102058.8, 101994.1, 
    101923.5,
  102423.4, 102430.7, 102430.5, 102416.6, 102405.2, 102383.2, 102355.2, 
    102323.7, 102277.4, 102221.3, 102161.5, 102099.3, 102030.7, 101961, 101883,
  102451.1, 102450.4, 102450.2, 102438.4, 102431.2, 102403.8, 102368.2, 
    102323.7, 102272.4, 102212.5, 102149.2, 102086, 102009, 101932.3, 101839.7,
  102482.5, 102481.7, 102478.6, 102455, 102438, 102415.9, 102380.4, 102329.7, 
    102269.2, 102207, 102137.3, 102073.7, 101992.1, 101907.2, 101800,
  102499.9, 102494.6, 102492, 102478.9, 102451.6, 102419.9, 102379.6, 
    102327.8, 102265.3, 102202.4, 102131.7, 102059.2, 101972.7, 101877.9, 
    101759.5,
  102521.9, 102516.8, 102501.2, 102488.6, 102462.3, 102426, 102380.9, 
    102329.3, 102266.7, 102197.3, 102125.3, 102045.7, 101952.1, 101851.4, 
    101720.1,
  102536.9, 102528.7, 102515.7, 102494.8, 102467.1, 102429.5, 102378.8, 
    102325.2, 102268.4, 102195.4, 102115.7, 102029.3, 101928.7, 101818, 
    101679.4,
  102545, 102535.1, 102522.4, 102499.2, 102472.4, 102437, 102383.5, 102325, 
    102262.6, 102190.5, 102105.5, 102008.7, 101902.4, 101782.7, 101635.9,
  102547.6, 102538.1, 102523.9, 102499.8, 102476.2, 102435.8, 102385.4, 
    102327.7, 102261.1, 102181.6, 102090.5, 101985.5, 101873.1, 101742, 101588,
  102555.9, 102536.7, 102524.3, 102505.7, 102479.4, 102436, 102385.7, 
    102325.3, 102255.1, 102168.2, 102070.4, 101959.6, 101839.5, 101697.5, 
    101535,
  101716.4, 101743.3, 101766.2, 101764.4, 101776.8, 101763.3, 101783.6, 
    101808.6, 101823.4, 101839.1, 101858.9, 101882.3, 101906.2, 101940.1, 
    101977.1,
  101771.2, 101801.6, 101796.1, 101788.6, 101777.9, 101757.3, 101768.9, 
    101769.7, 101779, 101792.8, 101808.9, 101823.1, 101842.9, 101867.1, 
    101901.6,
  101757.6, 101794.8, 101782.2, 101782, 101758.1, 101744.1, 101742.4, 101738, 
    101737.2, 101737.5, 101743.1, 101748.7, 101761.5, 101781.1, 101810.8,
  101780.4, 101804.2, 101777.5, 101772, 101733.7, 101726.4, 101711, 101696.2, 
    101684.9, 101677.4, 101672.9, 101670, 101673.4, 101685.9, 101708.3,
  101800.4, 101798.4, 101767.9, 101753.6, 101719.8, 101708.6, 101677.3, 
    101655.3, 101629.5, 101611, 101591.1, 101579.9, 101572.8, 101577.2, 
    101593.6,
  101826.9, 101792.3, 101764.5, 101735.6, 101698.4, 101677, 101634.7, 
    101602.8, 101564.8, 101533.3, 101504, 101482.1, 101462.3, 101460, 101468.1,
  101838.7, 101786.9, 101759.3, 101719.1, 101678.6, 101643.8, 101590.9, 
    101546.7, 101497.8, 101453.4, 101408.5, 101376.4, 101346.7, 101333.3, 
    101326.8,
  101846.9, 101795.1, 101754.4, 101708.2, 101657.2, 101608.9, 101543, 101489, 
    101425.9, 101369.9, 101313.8, 101262.1, 101225, 101193.2, 101175,
  101854.3, 101801.9, 101752.4, 101700.6, 101636.4, 101575.2, 101499.9, 
    101431.8, 101352.9, 101286.7, 101214.3, 101147.2, 101094.8, 101046, 
    101014.3,
  101868.7, 101812.7, 101759.2, 101696.2, 101622, 101546.7, 101461.5, 
    101376.1, 101281.7, 101199, 101112, 101030.3, 100958.7, 100893.6, 100845.1,
  102508.4, 102580.7, 102648.3, 102723.7, 102783.5, 102846.3, 102900.6, 
    102958.6, 103008.5, 103055.1, 103089.3, 103120.8, 103143, 103162.1, 103166,
  102549.2, 102609.7, 102677.2, 102741.4, 102791.9, 102854.1, 102909.6, 
    102962.2, 102998.8, 103037.9, 103068.5, 103092.8, 103110.1, 103118.6, 
    103119.1,
  102554.4, 102619.7, 102684.1, 102744.8, 102801.3, 102852.6, 102897.2, 
    102940, 102975.4, 103007.9, 103033, 103050.9, 103061, 103062.5, 103055,
  102559, 102616.5, 102682.5, 102736.2, 102787.7, 102833.2, 102876.9, 
    102911.6, 102941.1, 102964.7, 102982.7, 102993.3, 102995.2, 102986.9, 
    102970.7,
  102541.5, 102596.5, 102659.1, 102712.3, 102761.7, 102802.8, 102838.1, 
    102867.6, 102892.6, 102911.4, 102923.4, 102925.2, 102915.2, 102898.5, 
    102871.5,
  102519.9, 102568.7, 102628.7, 102679.9, 102721.5, 102760.1, 102789.9, 
    102814, 102830, 102842.6, 102846.2, 102837.9, 102818.8, 102791, 102752.7,
  102486.7, 102532.1, 102587.9, 102634.6, 102671.5, 102705.4, 102728.2, 
    102747.2, 102758.3, 102762.1, 102755.1, 102735, 102706.1, 102665.2, 
    102618.7,
  102445.9, 102488.5, 102538.4, 102579.6, 102613.5, 102639.1, 102656.4, 
    102666.5, 102667.1, 102661.3, 102642.3, 102612.1, 102570.5, 102522, 
    102462.5,
  102393.3, 102432.2, 102475.7, 102512.5, 102540.3, 102560.3, 102570.4, 
    102571.8, 102563, 102545.6, 102514.1, 102469.9, 102418.1, 102356.8, 
    102285.8,
  102331.3, 102365.5, 102402.3, 102432.8, 102455.4, 102467, 102468.7, 102459, 
    102439.5, 102409.4, 102363.8, 102309.1, 102244.5, 102170, 102089.3,
  102917.7, 102952.5, 103010.7, 103052.9, 103094.8, 103145.4, 103175, 
    103208.7, 103229.6, 103244, 103245.8, 103247.4, 103248.6, 103247.7, 
    103232.5,
  102973.5, 103006.4, 103056, 103101.8, 103136.4, 103168.3, 103195, 103213, 
    103216.4, 103220.3, 103219.6, 103214.3, 103206.3, 103195.9, 103184.6,
  103006.8, 103058, 103089.2, 103123.2, 103152.2, 103175.3, 103188, 103193.3, 
    103194.6, 103191, 103184.4, 103178.7, 103168, 103158.9, 103144.4,
  103044.1, 103077.4, 103103.5, 103131.6, 103151.8, 103159.2, 103162, 
    103160.3, 103155.9, 103143.8, 103134, 103124.6, 103113.4, 103100.2, 
    103086.9,
  103068.1, 103075.6, 103105.7, 103113.9, 103126.4, 103125.7, 103124.8, 
    103112, 103101.1, 103089.1, 103077.6, 103065.7, 103053.7, 103041.5, 103024,
  103065.5, 103060.7, 103087.5, 103083.9, 103087.6, 103075.3, 103065.5, 
    103049.7, 103037.3, 103022.1, 103007.5, 102992.5, 102978.9, 102963.6, 
    102947.4,
  103041.6, 103032.9, 103048.8, 103036.9, 103032.6, 103016.2, 103001.7, 
    102981.7, 102962.9, 102943.2, 102927.1, 102910.5, 102895, 102873.7, 
    102850.1,
  103004.9, 102996.1, 103000.9, 102979.1, 102965.2, 102941.4, 102920, 
    102894.2, 102873.4, 102851.3, 102832, 102811.5, 102791.1, 102768.2, 
    102740.8,
  102960, 102940.4, 102932.8, 102903.6, 102883.9, 102855.8, 102829.3, 
    102798.9, 102773, 102748.4, 102724.1, 102698, 102672.1, 102643.6, 102615,
  102899.8, 102873.6, 102850.5, 102817.9, 102791.7, 102756.9, 102723.8, 
    102687.5, 102655.8, 102625.4, 102596.3, 102565.9, 102534.8, 102503.1, 
    102469.2,
  102598.7, 102628.5, 102648.3, 102705.4, 102770.7, 102829.6, 102848.7, 
    102921.5, 102962.7, 102995.2, 103010.7, 103006.9, 103010.9, 103011.4, 
    103020.9,
  102718.3, 102750.3, 102797.6, 102872.7, 102895.2, 102901.3, 102918.6, 
    102971.2, 102977.9, 102997.1, 103007.5, 103012.6, 103009.2, 103006.5, 
    102999.3,
  102837.2, 102866.8, 102897.6, 102933.7, 102936.4, 102939.5, 102953.3, 
    102988.3, 103002.4, 103019.3, 103023.5, 103019.2, 103013.4, 103000.5, 
    102985.6,
  102950.9, 102966.7, 102988.6, 102997.5, 102986.8, 102985.8, 102996.3, 
    103019.9, 103027.3, 103030.8, 103029.6, 103023.3, 103015.3, 102990.6, 
    102970.2,
  103020.4, 103035.3, 103045.9, 103036.1, 103021.2, 103025, 103027.2, 103033, 
    103038, 103038.3, 103034.2, 103021.8, 103007.9, 102976.6, 102951.2,
  103072.7, 103079.6, 103072, 103059.2, 103048.7, 103044, 103042.2, 103039.8, 
    103048, 103043.6, 103036.1, 103015, 102992, 102955.4, 102923.8,
  103099.9, 103083.1, 103074.7, 103068.1, 103064.9, 103053.5, 103049, 
    103045.4, 103040.5, 103030.1, 103016.9, 102994.1, 102962, 102924.4, 
    102882.2,
  103093.5, 103084.5, 103079.6, 103073.7, 103070, 103052.9, 103043.9, 
    103035.5, 103025.2, 103011.1, 102990.6, 102964.6, 102925.3, 102881.5, 
    102832.4,
  103076.2, 103083.4, 103071.8, 103068.7, 103057.8, 103046.3, 103035.6, 
    103018.8, 102999.1, 102980.4, 102954.1, 102915.9, 102872.4, 102824.8, 
    102768.3,
  103064.7, 103067.2, 103060.4, 103052.3, 103039.4, 103027.5, 103009.9, 
    102991.1, 102964.6, 102937.7, 102903, 102859.7, 102810.4, 102756.4, 
    102693.5,
  102246.5, 102268.8, 102306.3, 102416, 102509.5, 102594.2, 102689.7, 
    102749.7, 102803.1, 102849.8, 102899.8, 102922.5, 102944.8, 102969, 
    102979.3,
  102202.5, 102221.6, 102252.3, 102403.9, 102536.4, 102616.2, 102697.4, 
    102747.4, 102793.2, 102826.8, 102864.8, 102894.7, 102918.4, 102934.7, 
    102939.9,
  102171.5, 102192.9, 102201.2, 102415.3, 102500.2, 102590.1, 102680.5, 
    102736, 102788.8, 102821.8, 102856.4, 102871.3, 102888.1, 102897.6, 
    102895.3,
  102135.7, 102177.8, 102192.2, 102431.7, 102500, 102598.7, 102673.4, 
    102724.6, 102769.5, 102796.6, 102820.9, 102840.6, 102850.8, 102852.5, 
    102848.4,
  102123.8, 102184.8, 102227.6, 102437.6, 102488.7, 102589.3, 102649.3, 
    102709.2, 102749.1, 102775.5, 102794.3, 102805.5, 102803.7, 102799.7, 
    102793.1,
  102133.1, 102201.6, 102299.1, 102468, 102494.2, 102588.2, 102633, 102684.4, 
    102719.3, 102741.5, 102752, 102751.8, 102748.3, 102742.9, 102732.5,
  102175, 102232.3, 102368.9, 102467.5, 102495, 102575.7, 102614.1, 102657.8, 
    102683.6, 102699, 102702.2, 102695.6, 102684.9, 102670.6, 102658,
  102222.9, 102317, 102435, 102468.6, 102511.9, 102565.6, 102592.9, 102622.5, 
    102642, 102649.2, 102646.6, 102631.2, 102612.3, 102593.8, 102569.1,
  102287.4, 102435.1, 102463.1, 102468.3, 102517.8, 102539.9, 102571.9, 
    102590.9, 102598.8, 102593.9, 102579.2, 102556.3, 102528.3, 102501.8, 
    102472.5,
  102405.9, 102495.1, 102478.7, 102479.9, 102512, 102519.7, 102538.4, 
    102542.1, 102539.5, 102526, 102502.4, 102470, 102435.5, 102403, 102363.4,
  102689.5, 102735.4, 102782.8, 102827, 102865.4, 102901.3, 102944.8, 
    102963.3, 102990.7, 103014.4, 103026.8, 103030.2, 103023.8, 103028.7, 
    103034.8,
  102713.1, 102752.7, 102803.5, 102839.2, 102874.3, 102907.3, 102943.6, 
    102969.5, 102990.8, 103008, 103024, 103040.1, 103038.3, 103044, 103037.8,
  102695.2, 102743.7, 102794.1, 102832, 102873.6, 102907.7, 102936.8, 
    102959.3, 102977.8, 102994.1, 103007.8, 103021.4, 103023.8, 103045.4, 
    103050.3,
  102689.9, 102738, 102784.2, 102821.9, 102857.4, 102890.4, 102920.1, 
    102943.3, 102961.6, 102984.6, 103006.9, 103025.6, 103043, 103059.4, 
    103050.7,
  102659.1, 102708.4, 102757, 102798.6, 102837.3, 102869, 102895.1, 102916, 
    102936.5, 102963.6, 102986.1, 103006.1, 103017.8, 103034.5, 103036.9,
  102619, 102673.1, 102722.3, 102764.6, 102801, 102833.9, 102862.2, 102886.9, 
    102910.1, 102938, 102959.8, 102977.3, 102990.3, 102994.9, 102995.9,
  102566.1, 102626.7, 102677, 102723.5, 102762.7, 102798.8, 102823, 102848.8, 
    102871.4, 102892.5, 102911.6, 102929.2, 102943, 102953.1, 102954.4,
  102511.5, 102578.2, 102628.7, 102678.6, 102718.1, 102755.2, 102782.2, 
    102805.6, 102825.6, 102846.7, 102864.4, 102883, 102893.4, 102894.1, 102889,
  102452.9, 102524.4, 102578.5, 102628.3, 102667.9, 102705.2, 102732.5, 
    102754.2, 102773.4, 102789.9, 102807.9, 102821, 102830.1, 102831.6, 
    102826.8,
  102394.4, 102468.1, 102529.3, 102574.7, 102611.8, 102646.1, 102672.4, 
    102695.2, 102713.2, 102730.5, 102745, 102758.6, 102762.5, 102758.4, 
    102749.5,
  102782.9, 102804.8, 102821.6, 102825.3, 102823.1, 102820, 102819.8, 
    102819.1, 102811.2, 102796.4, 102778.1, 102760.3, 102735.9, 102709.9, 
    102676.6,
  102835.6, 102853.9, 102865.7, 102868.2, 102872.2, 102875.2, 102875.5, 
    102873.8, 102864.9, 102856, 102839.2, 102818.2, 102788.8, 102756.4, 
    102719.2,
  102862, 102878.3, 102897.9, 102908.4, 102916.9, 102912.7, 102912.7, 
    102914.7, 102904.6, 102890.8, 102878, 102867.9, 102836.9, 102806.3, 
    102757.9,
  102881.4, 102905.1, 102923.7, 102936.1, 102951.4, 102952.3, 102957.1, 
    102950.5, 102968.1, 102961.6, 102956.5, 102932, 102896.4, 102859.1, 
    102806.8,
  102906.1, 102924.9, 102951.6, 102969.7, 102985.9, 102988.6, 102985.8, 
    103001.4, 103008.8, 103000.4, 102989.6, 102974.1, 102941, 102901.9, 
    102840.5,
  102920.5, 102940.9, 102967.6, 102989, 103006.1, 103019.8, 103022, 103027.9, 
    103023.9, 103015.3, 103001.9, 102980.5, 102950.5, 102912.9, 102863.2,
  102927.3, 102955, 102976.9, 102999.4, 103016.6, 103026.1, 103026.7, 
    103025.7, 103018.3, 103008.4, 102995.2, 102977.4, 102948.1, 102909.5, 
    102863,
  102923.7, 102947.2, 102972.6, 102991.1, 103006.1, 103015.7, 103020.4, 
    103016.7, 103007.4, 103000.3, 102985.9, 102959.8, 102930.4, 102888, 
    102841.6,
  102921.4, 102946.3, 102965.9, 102981.6, 102994.6, 103003.9, 102999, 
    102994.2, 102985.3, 102974.6, 102949.6, 102923.1, 102894.9, 102858.7, 
    102808.8,
  102909.1, 102935.8, 102953.9, 102963.6, 102975.1, 102978.5, 102974.1, 
    102966, 102954, 102937, 102911.8, 102886.2, 102854.7, 102818.1, 102767.5,
  102543.6, 102521.5, 102475.1, 102428.1, 102377, 102320.5, 102255.1, 102177, 
    102084.2, 101983.1, 101895.3, 101846, 101819.7, 101792.1, 101746.6,
  102655.6, 102622.9, 102576.4, 102529.7, 102485.4, 102439.2, 102386.7, 
    102322.6, 102246.6, 102165.6, 102082.9, 102024.5, 101974.1, 101936.9, 
    101884.2,
  102736.8, 102698.9, 102672.7, 102631.9, 102587.9, 102539, 102489, 102433.3, 
    102368.9, 102294.9, 102219.5, 102151.1, 102084.7, 102031, 101968.7,
  102803.6, 102785, 102764.8, 102724.7, 102685.1, 102636.5, 102591.2, 
    102540.7, 102484.4, 102419.8, 102345, 102272.9, 102198.1, 102128.5, 
    102061.6,
  102876.9, 102861.7, 102850.1, 102827.6, 102789.9, 102744.6, 102689.1, 
    102632.8, 102578.5, 102520.3, 102451.5, 102378.5, 102298.6, 102217.1, 
    102136.8,
  102918.2, 102918, 102911, 102898.9, 102868.1, 102831.3, 102785.9, 102736.6, 
    102676.2, 102612.2, 102547.2, 102470.2, 102388.6, 102302.6, 102207.9,
  102964.8, 102969.8, 102957.9, 102943.6, 102919.8, 102890.2, 102850.1, 
    102804.3, 102750.6, 102687.1, 102617.6, 102544.9, 102460.3, 102369.5, 
    102270.2,
  103009.6, 103012.8, 103001.1, 102986.2, 102964.6, 102933.3, 102899.9, 
    102854.1, 102802.1, 102743.7, 102675, 102598.6, 102512, 102418.8, 102317.1,
  103054.4, 103052.5, 103041.8, 103025.2, 103002.1, 102970.8, 102936.4, 
    102891.5, 102841.1, 102783.7, 102713.8, 102637.2, 102551, 102454.3, 
    102346.2,
  103080.2, 103076.5, 103069.7, 103055.5, 103034.4, 103002.3, 102965.2, 
    102922.3, 102869.1, 102809.5, 102740.7, 102663.6, 102576.5, 102477.3, 
    102363.4,
  101939.3, 101809, 101651.8, 101487.5, 101315.2, 101129.8, 100925.7, 
    100706.3, 100506.6, 100310.4, 100161, 100003, 99996.14, 100060.1, 100265.3,
  102053.6, 101931.4, 101776.6, 101611.8, 101433.2, 101242.6, 101035, 
    100807.7, 100584.1, 100364.9, 100197.3, 100050.8, 100040.4, 100076, 100249,
  102167, 102042.2, 101891.7, 101727.3, 101551.9, 101360.8, 101153.3, 
    100921.9, 100682.6, 100450.5, 100266.5, 100117, 100070.1, 100078.8, 
    100221.1,
  102271.7, 102151.1, 102009.6, 101850.5, 101673.5, 101487.1, 101277.7, 
    101045.8, 100797.3, 100552.3, 100344.6, 100191.9, 100109.4, 100108.4, 
    100213.1,
  102374.9, 102259.4, 102121.6, 101966.1, 101798.2, 101615.6, 101413.8, 
    101185.6, 100935.6, 100686.2, 100463, 100296.6, 100178.3, 100166.3, 
    100216.2,
  102478, 102366.3, 102233.1, 102084.5, 101921.5, 101743.3, 101548.3, 
    101328.6, 101082.2, 100827.5, 100588.4, 100403.2, 100250.7, 100222.8, 
    100245.8,
  102578.4, 102468.8, 102341.7, 102195.8, 102038.4, 101867.5, 101681.3, 
    101472.6, 101235.9, 100984.6, 100736.6, 100535, 100352.7, 100299.2, 
    100297.8,
  102670.1, 102569.9, 102447.2, 102307.5, 102152.6, 101989, 101810.8, 
    101612.4, 101385.2, 101141, 100884.8, 100665.5, 100461.2, 100385.7, 
    100367.3,
  102753.2, 102663.2, 102551.5, 102414.2, 102267.3, 102105.3, 101933.6, 
    101745.9, 101527.6, 101292.2, 101037.9, 100810.1, 100583.3, 100483.4, 
    100445.9,
  102833.9, 102748.9, 102647.7, 102519.5, 102377.3, 102220.6, 102053.2, 
    101870.8, 101661.3, 101434, 101181.1, 100952.6, 100708.5, 100588, 100530.9,
  101662.6, 101559.5, 101590.9, 101596.7, 101637, 101677, 101725.3, 101759.5, 
    101786.4, 101797, 101795.8, 101792.6, 101798.8, 101801.4, 101810,
  101681.9, 101573, 101615.6, 101585.5, 101633.7, 101659.6, 101694, 101715.3, 
    101733, 101746, 101744.7, 101743.5, 101745.4, 101744.5, 101747,
  101719.5, 101600.4, 101626, 101571.4, 101604.7, 101620.6, 101648.8, 
    101668.2, 101684.8, 101690.2, 101690.5, 101690.7, 101686, 101682.9, 
    101682.9,
  101749.9, 101630, 101624.5, 101559, 101580.5, 101582.2, 101603.9, 101611.2, 
    101621.3, 101628.1, 101630.9, 101629, 101621.9, 101614.9, 101613.4,
  101784.8, 101667.7, 101627.4, 101559.6, 101552.9, 101539.6, 101549.9, 
    101552.4, 101559.2, 101565.6, 101567.2, 101564.5, 101554.5, 101544.4, 
    101543.9,
  101825.7, 101708, 101634.9, 101564.7, 101533.7, 101508.5, 101499.8, 
    101489.4, 101484.8, 101486.6, 101489.8, 101486.8, 101477.9, 101468.4, 
    101466.4,
  101881.2, 101752.3, 101648.7, 101571, 101519.1, 101476.7, 101451.1, 
    101429.1, 101411.2, 101403.5, 101402.3, 101403.6, 101395.1, 101388.3, 
    101384.8,
  101946.5, 101800.7, 101676.2, 101579.6, 101510.2, 101452, 101405.8, 
    101368.2, 101333.3, 101311.7, 101303, 101300.1, 101294.1, 101293.3, 
    101290.2,
  102009, 101851, 101706.8, 101593.8, 101509.7, 101430.8, 101364.4, 101307.1, 
    101256.8, 101220, 101197.5, 101189.1, 101188.1, 101189.6, 101196,
  102064.6, 101900, 101744.6, 101612.1, 101507.9, 101414.9, 101329.5, 
    101251.8, 101181.8, 101127.3, 101092.8, 101072.8, 101073.6, 101084, 
    101089.3,
  101572.8, 101668.8, 101777.8, 101850.9, 101961.1, 102048.6, 102120.3, 
    102180.3, 102240.8, 102284.7, 102333, 102393.4, 102451.3, 102508.9, 
    102565.5,
  101612.1, 101687.3, 101772, 101845.3, 101964, 102025.9, 102094.8, 102151.1, 
    102206.5, 102246.3, 102297.3, 102351.9, 102406.1, 102460.2, 102513.1,
  101630.9, 101707.4, 101790, 101849.5, 101959.6, 102010.9, 102080.7, 
    102125.7, 102173.4, 102206.7, 102252.9, 102302.8, 102351.3, 102402.2, 
    102445.2,
  101660.5, 101715.3, 101796, 101847.6, 101952.4, 101990.7, 102055.9, 102091, 
    102130.6, 102161, 102201.5, 102246.4, 102292.6, 102337.4, 102375.8,
  101663.9, 101712.2, 101791.9, 101839.7, 101936.9, 101971.8, 102028.8, 
    102055.1, 102085.5, 102110.9, 102148.1, 102181.7, 102222.8, 102260.8, 
    102291.9,
  101649.2, 101701.9, 101780.8, 101826.5, 101916.6, 101945.6, 101996.6, 
    102013.6, 102035.1, 102051.4, 102083.4, 102115.6, 102147.8, 102178.9, 
    102202.1,
  101624.2, 101677.5, 101751.7, 101801.3, 101882.8, 101912.8, 101957.9, 
    101968, 101982, 101994.1, 102019.4, 102042.4, 102068.7, 102090.6, 102104.4,
  101598.8, 101648.8, 101720.8, 101776.6, 101843.2, 101878.1, 101912.6, 
    101919.5, 101922.7, 101928.7, 101946.5, 101963.3, 101979.3, 101992.2, 
    101996.5,
  101574.2, 101616.9, 101686.1, 101746.1, 101800.8, 101836.9, 101858.7, 
    101859, 101857.4, 101859.4, 101869.9, 101875.3, 101883, 101883.8, 101878.3,
  101561.1, 101583.5, 101648.8, 101711.1, 101762.5, 101792.9, 101803.9, 
    101800.7, 101789.4, 101783.2, 101781.6, 101779.8, 101775.7, 101764.5, 
    101747.3,
  101653.2, 101799.8, 101949.2, 102072.5, 102180.7, 102277.6, 102369.6, 
    102451.1, 102528.2, 102604.5, 102679.2, 102754.2, 102823.7, 102890.4, 
    102952.8,
  101602.7, 101756.9, 101918.4, 102039.2, 102145, 102238.8, 102327.1, 
    102408.7, 102487.2, 102562.3, 102636.2, 102710.5, 102778.9, 102843.6, 
    102904.3,
  101572.1, 101724.9, 101886, 102006.4, 102111.6, 102200.3, 102283.5, 
    102360.5, 102438, 102515.4, 102589.7, 102663.8, 102730.8, 102792, 102852.7,
  101553.2, 101710.2, 101859.9, 101979.2, 102079.5, 102162.2, 102238, 
    102311.8, 102387.3, 102464.4, 102540, 102609, 102672.9, 102731, 102790,
  101546.6, 101707.5, 101839.5, 101956.9, 102048.6, 102125.8, 102192.4, 
    102261.9, 102334.6, 102408.7, 102481.8, 102548.6, 102609.2, 102666, 
    102721.9,
  101560.5, 101720.8, 101824.4, 101935.7, 102016.5, 102084.7, 102145.2, 
    102208.9, 102276, 102348, 102416.1, 102478.8, 102532.1, 102585.3, 102638.2,
  101592.7, 101726.3, 101820.3, 101917.6, 101989, 102045.8, 102097.2, 102153, 
    102213.9, 102280.6, 102343, 102398.6, 102448.1, 102496, 102543,
  101643, 101736.1, 101821.7, 101897.9, 101955.8, 102004.6, 102046.6, 102093, 
    102146.2, 102206.4, 102263.3, 102310.2, 102353.4, 102395.1, 102438,
  101676.4, 101744, 101814.1, 101878.5, 101922, 101960.5, 101993.8, 102030.1, 
    102074.3, 102124, 102170.7, 102212.7, 102249.4, 102284.1, 102320.8,
  101708.2, 101748.8, 101801.1, 101854, 101881.8, 101912.2, 101933.6, 
    101960.9, 101995.6, 102034.2, 102073.1, 102104.6, 102135.1, 102163.5, 
    102194.9,
  101833.7, 101963.5, 102086.1, 102195.6, 102303.9, 102407, 102513.2, 
    102606.3, 102698.4, 102781.9, 102861, 102934.6, 103004.9, 103067.3, 
    103125.2,
  101781, 101914.8, 102041.9, 102154.4, 102266.3, 102369.5, 102476.5, 
    102572.1, 102666, 102750.9, 102832.8, 102907, 102977.3, 103041, 103099.3,
  101717.7, 101854.4, 101992, 102110.6, 102225.3, 102330.5, 102437.6, 
    102535.8, 102630.8, 102719.6, 102801.8, 102876.3, 102945.3, 103013.7, 
    103074,
  101658.8, 101800.5, 101947, 102068.8, 102186.8, 102292.5, 102399.6, 
    102499.2, 102592.7, 102683, 102767.8, 102845.2, 102916.6, 102981, 103043.5,
  101599.9, 101746.8, 101898, 102023.7, 102145.5, 102254.6, 102359.8, 102461, 
    102556.1, 102645.9, 102732.3, 102812.8, 102884.9, 102953.9, 103014.2,
  101543.2, 101700.8, 101853.3, 101981.9, 102106.8, 102216.3, 102323.1, 
    102421.9, 102517.3, 102608, 102694.5, 102775.7, 102849.5, 102921.9, 
    102982.1,
  101492.1, 101662, 101811.9, 101943, 102069.2, 102180.8, 102286, 102383.7, 
    102478.1, 102568.9, 102656.4, 102737.9, 102812.5, 102882.9, 102945.4,
  101465.1, 101635.1, 101778.2, 101911.7, 102033.9, 102147.1, 102251.3, 
    102345.6, 102438.6, 102528.8, 102615.8, 102699.2, 102775.5, 102845.9, 
    102906.6,
  101454.6, 101614, 101753.8, 101883.2, 102000.2, 102112, 102214.7, 102308.4, 
    102400.3, 102486.4, 102572.1, 102655.2, 102732.7, 102802.6, 102862.3,
  101459.4, 101603.9, 101736.4, 101858.5, 101969, 102076.5, 102177, 102269.1, 
    102356.6, 102443.2, 102526.3, 102608.1, 102684.2, 102755.1, 102819.5,
  102051.8, 102165.2, 102273.6, 102373.8, 102459, 102535.9, 102604.6, 102667, 
    102717.8, 102758.6, 102790.7, 102820, 102840.2, 102834, 102829.2,
  102034.4, 102147.1, 102275.9, 102376, 102466, 102543.9, 102615.5, 102677.9, 
    102728.6, 102770.8, 102805.8, 102833.7, 102846.9, 102839.5, 102823.3,
  102011.9, 102131.5, 102264.6, 102370, 102469.9, 102554.6, 102629.1, 
    102693.3, 102746, 102786.1, 102813.5, 102840.6, 102843.9, 102841.9, 
    102822.7,
  101998.8, 102122.1, 102263.7, 102375.1, 102481.4, 102569.5, 102647.8, 
    102714.1, 102768.1, 102804.8, 102829.5, 102849.3, 102857.4, 102858.2, 
    102829,
  101989.7, 102119.4, 102264.6, 102380.8, 102491.5, 102586.7, 102669.3, 
    102736.4, 102787, 102828.6, 102851.8, 102863.4, 102874, 102870.5, 102836.5,
  101981.2, 102123.4, 102270, 102394, 102504.8, 102604.5, 102686.1, 102752.9, 
    102806.7, 102848.1, 102878.4, 102894.7, 102888.6, 102877.1, 102839.2,
  101977.8, 102133, 102274.7, 102405.6, 102520.3, 102618.9, 102704.3, 
    102771.3, 102828.1, 102870.5, 102898.9, 102912.3, 102910.1, 102886.7, 
    102844.2,
  101961.1, 102130.9, 102280.6, 102416.9, 102533.3, 102636.1, 102721.7, 
    102790.8, 102843.7, 102889.8, 102917.4, 102929.6, 102928.2, 102902.5, 
    102854.1,
  101953.8, 102128.5, 102284.4, 102422.9, 102547.9, 102650.6, 102739.5, 
    102808.6, 102867.1, 102909.1, 102934.6, 102942, 102937.8, 102912.3, 
    102856.6,
  101941.8, 102122.2, 102288.9, 102429.9, 102560.9, 102666.7, 102756.4, 
    102830.5, 102887.4, 102921.9, 102947.5, 102953.5, 102938.9, 102913.7, 
    102861.7,
  101923.6, 101969.5, 102011, 102043, 102046.4, 102045.5, 102036.7, 102021.6, 
    101983.4, 101945.2, 101885.7, 101817.1, 101749.1, 101678.5, 101616.3,
  101908.3, 101954.9, 101998.5, 102025.4, 102027.2, 102031.7, 102024.1, 
    102003.6, 101963.2, 101916.8, 101855.2, 101784.7, 101709.2, 101625.5, 
    101562.5,
  101870.6, 101928.4, 101964.6, 102001.3, 102014.4, 102017.1, 102009.4, 
    101983.5, 101950.5, 101891.6, 101824.8, 101753, 101667.2, 101580.3, 
    101515.8,
  101836.6, 101898.6, 101944.8, 101985.3, 102000.4, 102001.4, 101995.3, 
    101982.2, 101930.8, 101870.8, 101796, 101718.3, 101626.9, 101533.7, 
    101466.8,
  101789.5, 101858.6, 101912.7, 101953.6, 101981.7, 101990.7, 101988.5, 
    101972, 101910.9, 101848.5, 101768, 101683.1, 101589.5, 101494.1, 101419.8,
  101735.6, 101815.8, 101876.5, 101926.4, 101962.2, 101979.7, 101981.3, 
    101962.1, 101901, 101831.3, 101748.2, 101650.6, 101548.9, 101447.4, 
    101364.7,
  101670.9, 101766.7, 101834.7, 101894.8, 101937.9, 101964.3, 101975.8, 
    101952.4, 101891.6, 101819.4, 101726.6, 101621.4, 101513.9, 101404.3, 
    101311.6,
  101593.7, 101707.5, 101787.2, 101864.5, 101915.4, 101955.5, 101964.7, 
    101942.9, 101886, 101805.5, 101711.1, 101595.8, 101477, 101359.1, 101256.8,
  101506.4, 101636.9, 101734.6, 101829.3, 101887.5, 101937.9, 101950.6, 
    101933.7, 101875.2, 101794.7, 101694.8, 101573.9, 101445.8, 101315.6, 
    101201.8,
  101403.5, 101554.1, 101669.6, 101788.5, 101858.7, 101915.4, 101933.8, 
    101922.4, 101872.8, 101790.6, 101685.7, 101556.3, 101417.7, 101275.9, 
    101150.5,
  102021.1, 101962.4, 101900, 101838.6, 101771.4, 101712.2, 101664.3, 
    101625.7, 101599.8, 101584.8, 101586.4, 101605.8, 101640, 101684.5, 
    101739.1,
  102020.9, 101950.6, 101882.6, 101811.2, 101733.1, 101671.1, 101618.7, 
    101569.8, 101537.8, 101519.8, 101514.4, 101526, 101554.2, 101603.5, 
    101652.7,
  102008.8, 101938.5, 101860.1, 101781.4, 101698.9, 101628, 101567.2, 
    101509.8, 101468.1, 101440.3, 101427.3, 101435.7, 101464.6, 101506.8, 
    101542.6,
  101992.4, 101920.5, 101838.4, 101751.8, 101660.9, 101582.4, 101512.5, 
    101447.7, 101397.2, 101361.4, 101343, 101348.5, 101371.1, 101408.2, 
    101433.3,
  101977.4, 101900.5, 101820.5, 101725.2, 101627, 101538.5, 101458.6, 101386, 
    101324.4, 101281.4, 101257.6, 101255.3, 101272.7, 101298.5, 101312.8,
  101960.1, 101881, 101796.9, 101694.6, 101591.9, 101493.2, 101405.6, 
    101322.6, 101250.9, 101201.3, 101168.6, 101162.8, 101173, 101188.4, 
    101190.4,
  101940.4, 101860.4, 101773, 101666.1, 101556.2, 101450.5, 101353, 101260.3, 
    101177.5, 101117.1, 101076.5, 101062.8, 101064.9, 101065.8, 101055.9,
  101919.3, 101840.2, 101747.5, 101638.6, 101522, 101408.4, 101302.1, 
    101197.2, 101105.3, 101034.6, 100986.3, 100965.1, 100957.6, 100945.9, 
    100923.8,
  101895, 101818.8, 101724.5, 101614.4, 101494.1, 101371.2, 101254.5, 
    101139.8, 101035.3, 100950.8, 100893.3, 100860.2, 100837.3, 100815.9, 
    100780.5,
  101868.2, 101795.6, 101701.7, 101595.5, 101467.6, 101337.8, 101209.9, 
    101081.4, 100967.4, 100868.5, 100799.3, 100753.4, 100718.8, 100685.5, 
    100638.5,
  102429.2, 102439.5, 102460.4, 102495.2, 102531.8, 102571, 102610.9, 102643, 
    102674.1, 102709.7, 102738.9, 102766.3, 102791.4, 102811.6, 102825.8,
  102434.7, 102436.7, 102461.7, 102488.6, 102528.9, 102562.8, 102594.5, 
    102624.9, 102653.6, 102683.1, 102710.9, 102738.5, 102762.9, 102779.7, 
    102787.8,
  102422.4, 102425.4, 102449.4, 102472.2, 102508.2, 102537.6, 102570.6, 
    102601.3, 102630.5, 102659.3, 102684.7, 102705.7, 102722.3, 102733.8, 
    102743.1,
  102412.6, 102417.2, 102434.9, 102459.1, 102488.9, 102516.4, 102546, 102574, 
    102599.1, 102623.9, 102644.9, 102662.2, 102672.8, 102679.9, 102685.3,
  102398.5, 102401.4, 102412.4, 102433.6, 102463.2, 102488.8, 102516.8, 
    102542.3, 102565.1, 102586.9, 102605.3, 102619.3, 102625.6, 102630.9, 
    102631.5,
  102385.2, 102383.2, 102390.3, 102407.2, 102433.1, 102456, 102480.2, 
    102499.6, 102522.7, 102539.1, 102552.3, 102562.2, 102568.3, 102568.1, 
    102566.5,
  102363.5, 102355.3, 102365.7, 102373.8, 102398, 102416, 102437.6, 102453.3, 
    102471, 102485.2, 102494.7, 102499.6, 102500.7, 102497.2, 102492.3,
  102348.4, 102332.7, 102335, 102338.1, 102358.5, 102373.3, 102387.5, 
    102400.5, 102413.6, 102423.9, 102427.4, 102427.3, 102423, 102418, 102407.2,
  102325, 102303.9, 102301.5, 102297.9, 102312.3, 102321.2, 102330.9, 
    102337.6, 102344.9, 102350, 102349.8, 102345.3, 102336.4, 102324.8, 
    102311.2,
  102305.5, 102277.4, 102263.5, 102253.9, 102259.2, 102265.4, 102268.6, 
    102269.2, 102270.6, 102269.7, 102264.3, 102252, 102238.2, 102220.7, 
    102202.7,
  102954.5, 103036.5, 103093.9, 103154.3, 103221.1, 103276.6, 103315.4, 
    103366, 103400.1, 103429.3, 103446.7, 103461.8, 103481.2, 103497.4, 
    103503.8,
  102988.7, 103060.4, 103129.7, 103198.1, 103259.6, 103297.8, 103341.3, 
    103381, 103409, 103440.5, 103461.2, 103477.4, 103478.3, 103475, 103490.1,
  103018.4, 103092.3, 103159.2, 103219.2, 103286.1, 103322.8, 103362.3, 
    103397.3, 103421.8, 103440, 103447.1, 103453.2, 103463.9, 103482.5, 
    103497.5,
  103044.4, 103118, 103185.2, 103242.2, 103301.4, 103330.8, 103366.7, 
    103390.5, 103416.1, 103434.3, 103442.3, 103445.7, 103451.5, 103464.4, 
    103479.5,
  103065, 103136.6, 103199.4, 103251.7, 103304.6, 103332.5, 103364.7, 
    103385.4, 103404.4, 103417.3, 103424.9, 103430.8, 103439.2, 103448.6, 
    103460.8,
  103078, 103147.1, 103205.8, 103255.6, 103299.2, 103325.1, 103350.7, 
    103363.7, 103379.7, 103390.2, 103399.2, 103405.3, 103412.3, 103421.7, 
    103426.9,
  103080.8, 103147.1, 103200.9, 103247.8, 103283, 103306.4, 103323.9, 
    103334.8, 103346.5, 103352.9, 103359.6, 103363.5, 103369.5, 103376.5, 
    103381.9,
  103081.5, 103141.6, 103187.1, 103230.2, 103256.7, 103276.2, 103289.4, 
    103297.1, 103304.2, 103309.3, 103313, 103315.9, 103317.1, 103317.9, 
    103319.4,
  103073.8, 103128.6, 103167.9, 103201.1, 103224.4, 103238.3, 103247.3, 
    103251.1, 103252.3, 103254.5, 103253.8, 103253, 103251, 103248.4, 103243.6,
  103063.3, 103110.8, 103140.2, 103168.3, 103182.2, 103193.5, 103196.3, 
    103193.9, 103190.8, 103188.1, 103182.5, 103176.4, 103168, 103158.9, 
    103148.8,
  102918.2, 103018.3, 103074, 103162.6, 103213.6, 103273.3, 103319.5, 103368, 
    103404, 103444.1, 103480.8, 103517.3, 103541.6, 103558.4, 103555.7,
  103000.4, 103069.1, 103128.9, 103205.8, 103246.1, 103303.1, 103344.6, 
    103398.6, 103435, 103471.8, 103499.4, 103525, 103546.3, 103562.5, 103570.5,
  103057.2, 103110.8, 103174.1, 103235.4, 103274, 103331.6, 103369.8, 
    103416.1, 103445.8, 103481.9, 103513.4, 103541.3, 103568.8, 103584.9, 
    103589.6,
  103103.4, 103140.1, 103203.1, 103250.7, 103300, 103342.5, 103378.5, 
    103424.2, 103454.5, 103487.4, 103518.2, 103539.8, 103557.5, 103574.1, 
    103563.2,
  103121.1, 103156.1, 103218, 103260.2, 103308, 103346.2, 103381.3, 103415.7, 
    103443, 103475.7, 103504.2, 103524.2, 103538.1, 103543.7, 103542,
  103123.3, 103164.1, 103215.9, 103258.4, 103304.4, 103336.9, 103365.9, 
    103395.2, 103424.9, 103454.2, 103478.7, 103498.6, 103511, 103515.9, 
    103509.4,
  103118.6, 103153.8, 103203.1, 103242.6, 103281.9, 103311.2, 103343.2, 
    103370.1, 103396.2, 103422.6, 103444.1, 103459.8, 103469.2, 103473.7, 
    103470.1,
  103104.9, 103135.8, 103183.4, 103213.2, 103249.2, 103280.2, 103308.2, 
    103333.1, 103359.8, 103381.3, 103401.2, 103415.3, 103424.1, 103426.2, 
    103420.9,
  103077.8, 103105.4, 103149.3, 103175.8, 103209.9, 103234.4, 103263.8, 
    103287.5, 103309.6, 103330.8, 103348.8, 103361.3, 103369.5, 103371.3, 
    103362.6,
  103041.4, 103069.3, 103106.5, 103130.3, 103160.7, 103184.4, 103208.4, 
    103229.2, 103252.4, 103271.1, 103286.3, 103298.3, 103305.8, 103302.1, 
    103292.1,
  102441.7, 102510.8, 102539.9, 102622.1, 102709, 102773.4, 102835.9, 
    102908.1, 102950.7, 102994.2, 103035.6, 103070.4, 103094.4, 103103.5, 
    103094.9,
  102565.8, 102617, 102634.5, 102701.8, 102769.8, 102830.7, 102893, 102944.7, 
    102979.6, 103020, 103060.6, 103085.4, 103102.5, 103098.9, 103083.5,
  102639.5, 102675.6, 102714.5, 102779.3, 102833.8, 102882.8, 102945, 
    102984.6, 103014.3, 103041.9, 103072, 103089.4, 103103.8, 103093.5, 
    103065.9,
  102721.2, 102763.8, 102790.2, 102836.5, 102877, 102928.1, 102974.2, 
    102998.5, 103025.4, 103054.7, 103073.9, 103078.1, 103084.2, 103066.6, 
    103032.8,
  102792.4, 102823.5, 102853.2, 102885.4, 102917.1, 102964.5, 102997.2, 
    103011.5, 103035.6, 103052.8, 103060.2, 103049.9, 103046, 103021.6, 
    102982.5,
  102882.7, 102869.1, 102896.9, 102913.4, 102951.8, 102985.3, 103009.6, 
    103017.8, 103034.5, 103041.7, 103034.7, 103019.2, 103002.9, 102968.7, 
    102925.9,
  102909.3, 102895, 102926.8, 102940.3, 102977.7, 102989.8, 103006.8, 
    103012.4, 103012.2, 103007.5, 102991.5, 102972, 102948.4, 102904, 102854.8,
  102909.7, 102919.1, 102936.9, 102946.1, 102976.9, 102984.2, 102985.2, 
    102984.2, 102977.5, 102961.9, 102944.2, 102918.8, 102882.4, 102831, 
    102773.8,
  102899.2, 102912.3, 102927.4, 102944.9, 102957.7, 102961.8, 102960.8, 
    102944.2, 102930, 102911.6, 102885.7, 102848.6, 102802.8, 102746.9, 
    102682.2,
  102887.9, 102906.6, 102918.6, 102924.1, 102926.4, 102921.9, 102910.3, 
    102894.9, 102872.9, 102849.4, 102814.9, 102772.1, 102718.2, 102655.4, 
    102579.8,
  101375.1, 101473.7, 101623.1, 101831.3, 101947.9, 102094.1, 102192.4, 
    102278.1, 102336.9, 102387.2, 102429.2, 102468.1, 102476.3, 102480.4, 
    102488.1,
  101434.4, 101492, 101606.4, 101832, 101943, 102087.3, 102196.7, 102283.1, 
    102343.6, 102380.8, 102414.9, 102433.3, 102429.5, 102425.8, 102439.7,
  101537.8, 101571.9, 101598, 101848.1, 101959.1, 102080.3, 102208.4, 
    102277.9, 102337.5, 102364.4, 102382, 102386.9, 102385.7, 102376.3, 
    102383.8,
  101673.9, 101696.6, 101678.6, 101854.8, 102014.8, 102087.6, 102219.8, 
    102276.5, 102329.3, 102346.7, 102355.4, 102349.2, 102337.2, 102324.4, 
    102325.6,
  101826, 101808.5, 101790.4, 101890, 102070.7, 102114.3, 102225.6, 102275.5, 
    102315.3, 102323.5, 102319.3, 102304.8, 102285.4, 102265.3, 102267.8,
  101962.7, 101916.2, 101906.9, 101975.8, 102125.3, 102147.9, 102228.3, 
    102269.3, 102287.1, 102296, 102274.8, 102250.6, 102225, 102207.5, 102202.1,
  102075.6, 102028.7, 102026, 102072.2, 102166.9, 102183.6, 102226.2, 
    102262.4, 102256.9, 102256.9, 102224.8, 102196.3, 102165.4, 102140.6, 
    102131.1,
  102187.3, 102138.9, 102137.3, 102164.7, 102207.3, 102207.9, 102224.8, 
    102239.3, 102222, 102204.9, 102169.2, 102131.5, 102096.7, 102066.1, 102055,
  102271.4, 102229.4, 102222, 102227, 102236.1, 102214.8, 102213.6, 102204.9, 
    102180, 102151.9, 102105, 102064.3, 102023.5, 101989.7, 101968.2,
  102338.4, 102296.7, 102276.5, 102262.2, 102244.7, 102212.4, 102196.9, 
    102167.9, 102130.1, 102089.3, 102034.5, 101985.6, 101940.9, 101904.7, 
    101877.9,
  101632.2, 101728.5, 101800.8, 101880.1, 101940.9, 102008.3, 102067.5, 
    102119.6, 102167, 102218.2, 102278.2, 102336.8, 102397.5, 102460.2, 
    102522.1,
  101548.3, 101658.9, 101744.5, 101831.7, 101906.1, 101980.9, 102045, 
    102104.2, 102162.1, 102222.4, 102284.2, 102358.8, 102427.9, 102497, 
    102561.5,
  101453.4, 101575, 101675.9, 101788.5, 101873, 101962.6, 102033.3, 102098.1, 
    102161.4, 102231.4, 102305.1, 102382, 102452.9, 102520.3, 102586.4,
  101364.4, 101492.5, 101602.3, 101738, 101835.3, 101936, 102010.7, 102082.9, 
    102151.8, 102230.4, 102311.1, 102396.4, 102475.7, 102547.8, 102619,
  101277.2, 101416.6, 101529.4, 101681.3, 101799.5, 101909.3, 101996.2, 
    102072.3, 102151.9, 102236.3, 102326.5, 102412.8, 102490.9, 102560.3, 
    102623,
  101204.2, 101349.7, 101461.1, 101629.3, 101760, 101875, 101971.6, 102054, 
    102138, 102227.5, 102321.2, 102411.9, 102492.5, 102562.3, 102628,
  101149, 101288.1, 101405.2, 101575.8, 101722.5, 101840.4, 101946.8, 
    102031.1, 102121.8, 102213.8, 102307.2, 102396.5, 102475.7, 102546.1, 
    102610.9,
  101099.4, 101234.5, 101352.6, 101530.9, 101683, 101800, 101910, 101999.4, 
    102091.6, 102182.5, 102276.9, 102365.4, 102442.2, 102515.2, 102574.6,
  101052.9, 101187.7, 101305.9, 101499.2, 101647.3, 101763.9, 101871.7, 
    101962.2, 102051.4, 102145.2, 102233.3, 102321.1, 102395.3, 102461.4, 
    102514.4,
  101026.5, 101157.7, 101286.9, 101485.5, 101613.8, 101727.8, 101828.8, 
    101919.1, 102003.8, 102094.1, 102181, 102265, 102334.4, 102394.3, 102437.3,
  102059.4, 102114.8, 102172.8, 102224.2, 102274.9, 102329, 102384.7, 
    102428.8, 102472.5, 102518.6, 102566.8, 102614.9, 102656.6, 102698.9, 
    102739.6,
  102064.1, 102119.3, 102184.3, 102231.2, 102279.3, 102330, 102389.7, 102437, 
    102485.3, 102534.7, 102582.6, 102634, 102676.6, 102722, 102763.6,
  102050.2, 102106.4, 102171.7, 102218.1, 102272.1, 102322.9, 102380.7, 
    102423.7, 102476.4, 102532.8, 102584.4, 102630.4, 102676.9, 102725.6, 
    102771.4,
  102031.6, 102086.3, 102146.7, 102198.4, 102247.7, 102302.9, 102352.3, 
    102408.3, 102456.9, 102509.5, 102562.4, 102613.5, 102661.3, 102708, 102756,
  102009.2, 102058.4, 102113.9, 102161.4, 102214.8, 102265.9, 102319.1, 
    102368.2, 102419.3, 102475, 102527.8, 102578.4, 102628.7, 102675.6, 
    102728.1,
  101977.5, 102026, 102075.4, 102120.4, 102169, 102217.4, 102268.3, 102313.4, 
    102362, 102412.7, 102464.5, 102514.8, 102565, 102616.3, 102669.5,
  101936.4, 101983.5, 102027.4, 102066.2, 102114.6, 102158.6, 102199.2, 
    102240.6, 102288.4, 102337.1, 102384.3, 102433.6, 102481.7, 102534, 
    102590.7,
  101888.4, 101935.8, 101972, 102010.1, 102046.8, 102085, 102120.6, 102157.6, 
    102197.9, 102240.7, 102283.5, 102327, 102373.4, 102427.5, 102484.7,
  101840, 101881.5, 101911.7, 101943.2, 101971.3, 102003.8, 102028.1, 
    102057.5, 102089.9, 102126.4, 102166.7, 102211, 102256.2, 102307.2, 
    102362.2,
  101788.3, 101823.4, 101844.7, 101870.9, 101888.2, 101912, 101929.8, 
    101949.9, 101972.9, 102003.2, 102036.5, 102072.4, 102114.8, 102164.5, 
    102220.2,
  102437.5, 102493.7, 102548.5, 102604, 102652.5, 102702.7, 102754.5, 
    102796.7, 102833.9, 102871.2, 102905.4, 102935.1, 102959.1, 102978.6, 
    102995.7,
  102441.2, 102499.9, 102554.2, 102609.2, 102663.4, 102718, 102770.4, 
    102814.5, 102853.8, 102887.8, 102919.2, 102950.9, 102976.2, 103001, 
    103023.6,
  102433.7, 102495.9, 102552.7, 102608.9, 102664.1, 102716.2, 102767.6, 
    102809.6, 102848.1, 102886.4, 102923.1, 102956.6, 102988, 103013.1, 
    103036.5,
  102425.3, 102480.5, 102536, 102592.2, 102646.1, 102696.7, 102746.4, 
    102788.3, 102826, 102861.3, 102898.8, 102932.3, 102965.2, 102995.1, 
    103027.4,
  102404.1, 102459.2, 102516.3, 102566.8, 102618.8, 102663.8, 102710.2, 
    102750.3, 102786.3, 102821.2, 102856, 102890.1, 102925.8, 102952.6, 
    102983.1,
  102372.3, 102423.2, 102478.8, 102526.6, 102575.9, 102617.2, 102658.2, 
    102693, 102726.3, 102755.7, 102787.5, 102819.3, 102850.8, 102881.6, 
    102909.3,
  102332.7, 102381.7, 102432.2, 102476.3, 102521.9, 102558.9, 102593, 
    102620.7, 102650, 102675.2, 102700, 102727.3, 102755.7, 102781, 102806.9,
  102276.9, 102328.1, 102376, 102415.3, 102455, 102487.4, 102515.6, 102535.5, 
    102557.9, 102577.5, 102598.6, 102615.6, 102635.4, 102655.2, 102675.2,
  102213.4, 102262.1, 102305, 102338.8, 102370.8, 102400.2, 102421, 102434, 
    102448.2, 102461.1, 102473.3, 102481.6, 102490.4, 102500.8, 102514.4,
  102141.6, 102188.8, 102226.2, 102257.7, 102281.8, 102299.4, 102311.4, 
    102318.1, 102324, 102325, 102324.6, 102322.1, 102322.7, 102324.6, 102331.2,
  102203.5, 102288.1, 102366.3, 102433.9, 102502.9, 102571.9, 102639.6, 
    102699.9, 102761.6, 102820, 102869.2, 102909.9, 102944.1, 102967.6, 
    102982.3,
  102133.6, 102202.4, 102276.4, 102347.4, 102423.8, 102497.4, 102569.8, 
    102635.4, 102700.4, 102765.1, 102825.5, 102882.5, 102928.6, 102968.3, 
    102998.3,
  102027.9, 102097.4, 102173.8, 102248, 102324.6, 102401.6, 102480.4, 
    102557.9, 102634.6, 102706.2, 102774.2, 102836.5, 102895.5, 102946.2, 
    102991.2,
  101905.2, 101970.3, 102041.7, 102117.3, 102199.5, 102284.4, 102369.2, 
    102452.2, 102534.7, 102618, 102697.9, 102772, 102839.1, 102902.3, 102956.7,
  101762.3, 101828.3, 101897.8, 101972.9, 102054.1, 102140.9, 102232.9, 
    102327, 102421.3, 102517, 102608.1, 102696.7, 102777.4, 102850.8, 102916.2,
  101604.8, 101660.5, 101724.4, 101798.2, 101881.4, 101971.7, 102069, 
    102171.1, 102274.4, 102380.8, 102485.1, 102587.5, 102684, 102771.8, 
    102854.6,
  101433.9, 101484.7, 101537.8, 101609.3, 101688.2, 101779.7, 101881.3, 
    101989.7, 102106.9, 102222, 102342.1, 102456.7, 102570.9, 102677.5, 
    102775.4,
  101254.1, 101292.7, 101334.6, 101397.1, 101473.2, 101566.6, 101670.3, 
    101785, 101908.3, 102037.1, 102167.6, 102297.5, 102426.9, 102549.2, 
    102667.1,
  101074.6, 101093, 101126, 101176.4, 101245.8, 101333.9, 101433.9, 101553.4, 
    101686.8, 101826.6, 101969.6, 102118.4, 102262.3, 102404.3, 102537.8,
  100896.6, 100902.9, 100911.7, 100950.4, 101004.2, 101086.3, 101186.3, 
    101304.9, 101438.8, 101587, 101746.3, 101903.6, 102069.5, 102228.6, 
    102380.1,
  102174.2, 102246.7, 102309.6, 102359.9, 102399.1, 102424.9, 102435.5, 
    102433.8, 102416.5, 102386.7, 102339.7, 102273, 102187.9, 102089.4, 
    101980.2,
  102123.6, 102198.8, 102269.4, 102331, 102385.5, 102427.6, 102456.9, 
    102470.4, 102468.7, 102452.9, 102425.3, 102382.6, 102328.1, 102258.3, 
    102176.4,
  102049.4, 102134.9, 102222.4, 102294, 102356.9, 102410.9, 102454.7, 
    102484.7, 102499.1, 102500.4, 102492.2, 102469.1, 102432.5, 102382.6, 
    102322.9,
  101970.9, 102062.3, 102154.7, 102237.1, 102313.6, 102380.6, 102438, 
    102483.5, 102515.1, 102531.3, 102541.5, 102537.5, 102520.9, 102490.6, 
    102448.7,
  101868.3, 101973.5, 102079, 102169.8, 102256.5, 102335.6, 102405, 102465.8, 
    102513.4, 102551.2, 102577, 102590.8, 102590.8, 102576.9, 102548.4,
  101746.9, 101866.1, 101982, 102084.7, 102181.9, 102273, 102356.2, 102428.6, 
    102490.6, 102542.2, 102582.7, 102611.6, 102627.9, 102629.8, 102619.9,
  101610, 101737.4, 101861.4, 101979.1, 102088.4, 102190.3, 102283.5, 
    102369.2, 102445.9, 102510.7, 102562.8, 102607.3, 102639, 102659, 102668,
  101460.7, 101590.7, 101723.2, 101847, 101968.6, 102082.9, 102190.4, 
    102286.4, 102375.7, 102451, 102519.9, 102576.5, 102625.6, 102661.2, 
    102686.3,
  101293.4, 101428.3, 101567.5, 101695.2, 101826.4, 101949.7, 102066.2, 
    102176.2, 102279.6, 102370.3, 102449.8, 102517.3, 102581.2, 102631.9, 
    102669.7,
  101113.3, 101251.2, 101394.8, 101528.6, 101665.1, 101797.1, 101922.9, 
    102043, 102156.1, 102257.7, 102352.2, 102434.4, 102508.1, 102572.8, 
    102624.3,
  101939.9, 101913, 101863.7, 101794.1, 101708.2, 101609.9, 101502.6, 
    101376.3, 101245.8, 101100.6, 100951.7, 100800.3, 100651.2, 100502.9, 
    100354,
  101976.1, 101956.5, 101936.5, 101887.3, 101822.9, 101740.9, 101647.7, 
    101542.4, 101427.6, 101304.3, 101166.1, 101011.2, 100851.7, 100695.9, 
    100542.4,
  101965.1, 101965.4, 101956.6, 101937.8, 101900.4, 101843.5, 101773.7, 
    101688.1, 101593.7, 101489.7, 101372.1, 101243.4, 101095.3, 100936.9, 
    100778.7,
  101935.2, 101955.3, 101965.2, 101956.2, 101944.7, 101912.4, 101869, 101808, 
    101730.8, 101640.9, 101546.7, 101439.6, 101317, 101184.2, 101039.9,
  101887.6, 101913.3, 101941.2, 101953.9, 101956.7, 101951.1, 101926.5, 
    101893.9, 101842.2, 101775.6, 101693.5, 101605, 101502, 101394, 101277,
  101823, 101863.6, 101898.2, 101926.1, 101944.6, 101955.3, 101953.4, 
    101938.9, 101914.4, 101876.4, 101821.4, 101754.3, 101673.5, 101581.3, 
    101482.2,
  101740.8, 101793.8, 101837.7, 101882, 101916.1, 101942.1, 101957.1, 
    101963.5, 101958.9, 101943.4, 101915.6, 101877.6, 101822.8, 101759.3, 
    101681.5,
  101650.3, 101707.7, 101760.5, 101813.1, 101861.6, 101902.1, 101932.9, 
    101953.4, 101965.2, 101972.8, 101969.7, 101954.5, 101930.2, 101890.4, 
    101837.4,
  101549.2, 101610.2, 101671.4, 101732.2, 101789.6, 101846.1, 101892.7, 
    101928.9, 101956.1, 101978.5, 101989.5, 101995.4, 101995.2, 101977, 
    101953.6,
  101438.4, 101504.6, 101570.7, 101638.2, 101703.1, 101767.2, 101826.6, 
    101878, 101918.9, 101958.1, 101986.6, 102005.1, 102015, 102021.5, 102019.6,
  101284.3, 101200.9, 101101.8, 101017, 100930.7, 100852.7, 100780.6, 
    100713.7, 100653.3, 100590.2, 100519.5, 100440.3, 100344.6, 100241.8, 
    100130.3,
  101415.8, 101317.8, 101214.5, 101123.3, 101027.9, 100934.7, 100849.8, 
    100766.2, 100687.3, 100609.4, 100535.6, 100457.1, 100366.1, 100262.2, 
    100150,
  101584.6, 101472, 101367.6, 101262.6, 101161.6, 101054, 100949.2, 100847.4, 
    100749.9, 100660.4, 100575.9, 100492.2, 100401.5, 100302.6, 100191.8,
  101736.3, 101634.7, 101524, 101409.2, 101312.3, 101206, 101098.8, 100990.8, 
    100882.5, 100775.7, 100675.4, 100583.6, 100487.2, 100378.6, 100264.7,
  101876.5, 101782.7, 101686.5, 101573.4, 101468.6, 101359.6, 101253, 
    101146.6, 101036.8, 100928.6, 100823.8, 100719.1, 100618.3, 100514.4, 
    100397.1,
  101983.3, 101912.4, 101821.6, 101723.6, 101627.5, 101525.4, 101426.4, 
    101329.5, 101224.1, 101113.1, 101002.9, 100897.5, 100795.5, 100690.6, 
    100576.7,
  102073.1, 102017.1, 101945.9, 101867.7, 101781.4, 101687.8, 101597, 
    101504.3, 101407.8, 101304.7, 101197.1, 101090.1, 100988.8, 100890.6, 
    100787.2,
  102143, 102094.2, 102037.3, 101974.1, 101908.2, 101832.6, 101758.9, 
    101677.6, 101593.3, 101497.9, 101398.1, 101298.5, 101198.5, 101103.6, 
    101006.9,
  102199.6, 102160, 102122.5, 102071.5, 102018.2, 101956.4, 101894.7, 
    101827.1, 101756.4, 101679, 101592.8, 101504.8, 101414.4, 101324.5, 
    101233.8,
  102233.8, 102205.6, 102181.7, 102143.5, 102105.6, 102057.2, 102008.6, 
    101956.7, 101899, 101835.2, 101766.9, 101689.9, 101611.7, 101530.9, 
    101447.1,
  101226.5, 101172.9, 101103.3, 101038, 100973.5, 100908.1, 100833.4, 
    100766.8, 100698, 100631.5, 100577.3, 100516.5, 100471.7, 100424, 100390,
  101218.7, 101163.9, 101091.8, 101027.3, 100960.2, 100892.9, 100822.4, 
    100750.4, 100672, 100609.5, 100535.9, 100475.9, 100414.1, 100358.2, 
    100302.9,
  101200.3, 101150.8, 101078.1, 101016, 100950.6, 100881.7, 100819.8, 
    100741.2, 100658.6, 100586.6, 100506.3, 100434.5, 100361.9, 100290.6, 
    100219.1,
  101187.1, 101135.7, 101067.3, 101001.5, 100934.7, 100874.1, 100813.1, 
    100740.1, 100658.8, 100582.4, 100498.5, 100416.6, 100333.6, 100249.2, 
    100160.9,
  101199.8, 101137.9, 101064.8, 100994.5, 100923.5, 100867.7, 100808.2, 
    100743.1, 100666.3, 100584, 100499.3, 100409.3, 100318.8, 100224.1, 
    100120.5,
  101243.8, 101167.2, 101085.4, 101006.6, 100926.9, 100866.4, 100806.7, 
    100751.6, 100680.5, 100602.3, 100516.7, 100422.7, 100328.4, 100223.3, 
    100110.8,
  101314.3, 101228.7, 101139, 101052.4, 100965.1, 100895.2, 100826.7, 
    100772.2, 100702.9, 100629.4, 100545.7, 100452.8, 100352, 100244.8, 
    100128.9,
  101403.3, 101314.6, 101219.2, 101126.4, 101037.8, 100960.6, 100883, 
    100824.4, 100753.8, 100679, 100593.2, 100500.7, 100400.2, 100292.6, 
    100172.4,
  101506.5, 101416.4, 101320, 101225.3, 101136.9, 101051.4, 100969.2, 
    100899.6, 100830, 100759.5, 100677.7, 100579.7, 100476.6, 100368.8, 
    100252.4,
  101612.3, 101521.9, 101426.7, 101334, 101244.6, 101155.7, 101073.3, 
    100996.7, 100926.9, 100859.2, 100785.9, 100695.3, 100590.4, 100481.4, 
    100366.6,
  101251.1, 101236.3, 101213.8, 101204.8, 101191.2, 101184.2, 101178.7, 
    101170.8, 101167.5, 101156.3, 101143.5, 101126.1, 101103.9, 101088.7, 
    101070,
  101217.1, 101191.7, 101172, 101156.2, 101143.8, 101139.2, 101128, 101121.1, 
    101113.1, 101108.3, 101099.1, 101086.4, 101068.7, 101045.9, 101021.2,
  101182.6, 101145.5, 101119.1, 101094.5, 101077.3, 101061.6, 101055.2, 
    101044.1, 101040.9, 101040.6, 101035.3, 101029.1, 101014.5, 100995.6, 
    100969.2,
  101147.9, 101106.5, 101074, 101049.1, 101026.2, 101005.4, 100989.7, 
    100976.1, 100970, 100967.2, 100966.4, 100960.5, 100949.4, 100933.5, 
    100909.9,
  101117.1, 101070.1, 101034.8, 101000.1, 100971.2, 100943, 100918.7, 
    100900.4, 100890.9, 100888.5, 100884.4, 100879, 100869.9, 100857.7, 
    100835.1,
  101091.1, 101041.5, 100997.3, 100958.5, 100920.9, 100891.8, 100861.8, 
    100840.1, 100820.7, 100810.7, 100800.6, 100795.5, 100783.5, 100767.5, 
    100748.2,
  101073.6, 101015, 100963.8, 100923.6, 100875.8, 100848.4, 100812, 100783.3, 
    100755.3, 100738.8, 100722.3, 100709.2, 100691.6, 100672.8, 100652.5,
  101057.1, 100995.3, 100939.9, 100892, 100842.5, 100802.5, 100768.5, 
    100733.6, 100706, 100678, 100653.1, 100629.2, 100605.2, 100578.4, 100549.8,
  101043.7, 100982.7, 100920.6, 100866.8, 100809, 100769.4, 100736.5, 
    100697.5, 100662.7, 100627.5, 100596.1, 100565.8, 100531.1, 100494.6, 
    100459.6,
  101021.3, 100966.5, 100904.7, 100848.2, 100791.4, 100754.8, 100719.9, 
    100672.8, 100626.2, 100590.7, 100551.6, 100513.2, 100466.1, 100415.7, 
    100368.2,
  101610.5, 101581.3, 101538.7, 101489.3, 101430.3, 101374.9, 101314.2, 
    101264.5, 101225.7, 101202.1, 101190.6, 101183.9, 101188.8, 101201.4, 
    101211.9,
  101618.5, 101582.2, 101538.6, 101485.5, 101429.2, 101369.7, 101315, 
    101256.3, 101210.8, 101174.7, 101149.9, 101135.5, 101125.5, 101122, 
    101121.6,
  101614.7, 101580.9, 101544.6, 101494.4, 101440.5, 101381, 101324.9, 
    101258.2, 101204.9, 101158.3, 101119.6, 101087, 101066.6, 101041.8, 
    101023.5,
  101594.4, 101570.3, 101538.3, 101489.9, 101441.7, 101383.3, 101329.7, 
    101267.7, 101205.4, 101155.6, 101106.7, 101065.3, 101029.1, 100994.7, 
    100951.3,
  101567, 101550.4, 101520.7, 101483.9, 101439.4, 101393.3, 101340.6, 
    101283.4, 101223.4, 101161.3, 101107, 101060.6, 101008.9, 100957.8, 
    100898.8,
  101528.3, 101516.7, 101490, 101464.3, 101427.2, 101392.5, 101344.5, 
    101292.9, 101234.6, 101176.5, 101118.8, 101065.4, 101011.2, 100956.4, 
    100883.7,
  101490.1, 101481.4, 101454.7, 101438.9, 101408.7, 101384.2, 101342.8, 
    101299.8, 101250.1, 101199.3, 101142.7, 101091.2, 101031.8, 100968.1, 
    100904.9,
  101445.3, 101435.3, 101413.7, 101402.1, 101381.1, 101361.3, 101329.4, 
    101294.3, 101256.4, 101211.9, 101168.6, 101114.7, 101066.4, 101000.8, 
    100935.1,
  101401.1, 101387.2, 101365.9, 101351.5, 101337.4, 101322.2, 101298.9, 
    101271.6, 101241.3, 101214.4, 101179.8, 101142.9, 101097.6, 101048.8, 
    100988.5,
  101362.3, 101341.5, 101320.6, 101296.5, 101283.1, 101269.8, 101254.5, 
    101235.1, 101209.7, 101188.4, 101163.2, 101135.4, 101109, 101070.2, 
    101019.7,
  101720.7, 101700.4, 101667.3, 101655.6, 101641.5, 101637.5, 101630.6, 
    101612.9, 101583.7, 101555.6, 101536.3, 101520.5, 101522, 101529.9, 
    101553.2,
  101739.1, 101701.3, 101664.4, 101635.7, 101612.5, 101599.1, 101583.5, 
    101559.4, 101524.9, 101498.9, 101468.7, 101438.7, 101424, 101420.6, 
    101436.3,
  101778, 101717.9, 101670, 101628, 101596.8, 101574.5, 101556.9, 101525.6, 
    101485.8, 101439.8, 101390.7, 101342.9, 101307.3, 101285.9, 101285.5,
  101816.2, 101746, 101684.8, 101620, 101581.4, 101544.4, 101518.8, 101486.8, 
    101445.8, 101391.1, 101327.2, 101261.1, 101197.2, 101143, 101115.8,
  101874, 101796.6, 101716.3, 101646.6, 101586.4, 101536.1, 101505.6, 
    101468.1, 101416.9, 101348.7, 101275, 101187.6, 101097, 101013, 100956.7,
  101919, 101860.4, 101770.3, 101676.3, 101595.2, 101540.6, 101480.5, 
    101445.8, 101389.7, 101322.7, 101245, 101145.2, 101035.1, 100933.4, 
    100853.7,
  101970.9, 101921, 101827.1, 101741.5, 101630.8, 101558.3, 101486.5, 
    101440.7, 101380.4, 101307.8, 101228.9, 101131.9, 101016.4, 100907.4, 
    100808.9,
  102022.8, 101976.2, 101891.5, 101803.6, 101689, 101596.2, 101508.2, 101440, 
    101378.5, 101306.9, 101229.2, 101137.3, 101029.2, 100923.6, 100822.5,
  102064.7, 102018.5, 101952.6, 101873.4, 101767.1, 101660.1, 101560.4, 
    101472.2, 101400.1, 101331.4, 101251, 101166, 101075, 100972.4, 100879.6,
  102101.4, 102059.6, 102005, 101934.1, 101840.9, 101738.2, 101625.7, 
    101529.4, 101440.5, 101370.7, 101295.5, 101214.7, 101134.3, 101048.5, 
    100966.8,
  101950.8, 101996.4, 102009.8, 102020.4, 102024.5, 102023.6, 102025.5, 
    102029.7, 102034.5, 102035.2, 102034.1, 102027.8, 102020.9, 102015.3, 
    102007.7,
  101919.4, 101953.2, 101969.6, 101977.4, 101970, 101968.4, 101966.8, 
    101966.5, 101969.4, 101972.5, 101974.4, 101978.6, 101978, 101970.1, 
    101955.9,
  101876.8, 101913.5, 101926.9, 101933.7, 101925.3, 101910.3, 101896, 
    101890.7, 101890.1, 101896, 101902.3, 101911.3, 101920, 101929.8, 101935,
  101865.7, 101881.5, 101891.8, 101888.8, 101873.7, 101852, 101829.7, 101813, 
    101801.7, 101798.2, 101804.5, 101816.9, 101835.9, 101854.3, 101872.8,
  101851.6, 101846.2, 101846, 101847.7, 101826.5, 101798.9, 101763.8, 
    101733.5, 101710, 101699.6, 101694, 101703.9, 101723.2, 101751.9, 101784.4,
  101859.1, 101827.6, 101824.4, 101808.1, 101782.1, 101749.5, 101707.8, 
    101668.4, 101635.4, 101608.2, 101595.1, 101597.7, 101615.7, 101646.6, 
    101684.2,
  101872.6, 101824, 101796.8, 101769.5, 101751, 101708.1, 101666.4, 101614.5, 
    101566.2, 101524.2, 101498.3, 101491, 101508.9, 101544.6, 101594.6,
  101891.1, 101844.7, 101797.2, 101751.5, 101721.8, 101677.3, 101633.6, 
    101573.5, 101515.4, 101459.8, 101419, 101396.9, 101403.2, 101436.5, 
    101500.7,
  101926.6, 101873.5, 101812.6, 101751.8, 101706.6, 101660.2, 101610.8, 
    101549.2, 101486.3, 101421.8, 101372.1, 101329.7, 101324.9, 101351.2, 
    101413.6,
  101969, 101925.6, 101852.1, 101783.2, 101711.3, 101650.9, 101603, 101541, 
    101479.8, 101411.7, 101359.5, 101316.6, 101300.9, 101315, 101366.1,
  102178.3, 102234.5, 102279.1, 102307.7, 102326.6, 102340.7, 102337, 102324, 
    102309.4, 102301.7, 102290.5, 102269.9, 102236.7, 102181.9, 102107.1,
  102161.4, 102202.2, 102238.9, 102272.8, 102296.2, 102308.1, 102316.3, 
    102323.7, 102302.9, 102295.1, 102265.7, 102238.3, 102196.3, 102133.5, 
    102063.8,
  102117.4, 102161.6, 102206, 102243.2, 102268.5, 102282.2, 102288.1, 
    102290.3, 102276.4, 102263.6, 102238.6, 102210.7, 102168.2, 102108.9, 
    102039.5,
  102070.8, 102115, 102155.9, 102189.5, 102216.2, 102238, 102250.2, 102256.8, 
    102253.8, 102246.6, 102223.5, 102191.4, 102142.1, 102081.6, 102006.2,
  102020.7, 102062, 102100.3, 102133.3, 102158.9, 102182.5, 102200.1, 
    102210.2, 102210.3, 102206.1, 102193.7, 102165.8, 102119.2, 102061.8, 
    101982.5,
  101961.1, 101998.5, 102030.8, 102059.7, 102084, 102108.8, 102131.9, 102151, 
    102165, 102173.7, 102165.3, 102140.1, 102097.7, 102035.3, 101955.5,
  101895.8, 101929.8, 101957.7, 101984.1, 102001.1, 102024.7, 102052.3, 
    102073.2, 102092.7, 102107.2, 102108.1, 102089.2, 102054.4, 101999.1, 
    101928,
  101823.6, 101852, 101875.1, 101895.5, 101909.1, 101931.8, 101957.2, 
    101980.7, 102009.8, 102035.3, 102048.3, 102039.7, 102014.6, 101966.4, 
    101900.6,
  101750.1, 101773.1, 101792.4, 101805.3, 101812.1, 101832.9, 101854.6, 
    101877.4, 101906.9, 101936.3, 101960.1, 101966.9, 101956, 101918.9, 
    101858.8,
  101675.9, 101686.6, 101708.3, 101713.2, 101716.5, 101731.7, 101744.2, 
    101766.2, 101792, 101827.8, 101860.1, 101880.2, 101882.1, 101859.2, 
    101814.5,
  102245.5, 102271.2, 102279.4, 102272.9, 102252.7, 102215.1, 102162.8, 
    102090.6, 102012.5, 101918.9, 101821.3, 101728.5, 101642.8, 101581, 
    101529.7,
  102244.3, 102262.8, 102271.1, 102268.2, 102244.1, 102198.5, 102144.4, 
    102067, 101970.9, 101867.2, 101758.3, 101665.1, 101582.4, 101508.4, 
    101457.8,
  102239.4, 102259.2, 102270.2, 102265.2, 102234.6, 102186.3, 102126.2, 
    102044.1, 101937.6, 101827.4, 101709.5, 101613.2, 101528.6, 101458.9, 
    101411.3,
  102230, 102246.5, 102258.9, 102256.5, 102234.5, 102181.5, 102112.3, 
    102024.7, 101911.9, 101792.6, 101666.1, 101560.8, 101479.9, 101405.7, 
    101341.3,
  102221, 102238.2, 102256, 102248.7, 102225.2, 102177.1, 102095.8, 102002.2, 
    101888.4, 101768.1, 101637, 101525.5, 101443.4, 101355.3, 101271.9,
  102197.8, 102223.4, 102237, 102230.7, 102208.7, 102163.9, 102090.8, 
    101993.1, 101868.1, 101746.9, 101604.3, 101493.9, 101404.7, 101300.5, 
    101201.9,
  102169.7, 102196.7, 102213.8, 102215, 102192.1, 102153.6, 102085.7, 
    101982.6, 101858.7, 101733.3, 101586.5, 101470.8, 101367.2, 101248.3, 
    101137.7,
  102130.6, 102159.4, 102175.7, 102181.7, 102163.3, 102133.3, 102068.3, 
    101974.6, 101847, 101722.4, 101573.8, 101446.9, 101330.8, 101201.8, 
    101076.3,
  102091.2, 102117.9, 102132.7, 102144.8, 102131.5, 102104.2, 102048.6, 
    101960.7, 101845.8, 101717.4, 101563.7, 101430.9, 101301.6, 101157.5, 
    101018.6,
  102036.6, 102065.9, 102086.1, 102095.7, 102092.9, 102072.6, 102023.1, 
    101945.4, 101835.3, 101713.6, 101561.4, 101419.7, 101275.6, 101116.9, 
    100960,
  102078.7, 102084.2, 102084.8, 102078, 102080.7, 102094.3, 102114.8, 
    102136.7, 102165, 102190.2, 102218.6, 102233.5, 102240.4, 102235.3, 
    102226.4,
  102073.6, 102056, 102060.5, 102050.2, 102052, 102062.2, 102079.2, 102099.4, 
    102125.9, 102155.8, 102189.4, 102206.6, 102216, 102211.1, 102203.6,
  102065, 102037.4, 102034.2, 102016.4, 102009.4, 102010.5, 102026.2, 
    102044.8, 102072.9, 102107.4, 102142.2, 102163.1, 102178.5, 102181, 
    102174.6,
  102053.4, 102020.6, 102006.5, 101985.8, 101971.4, 101964, 101972.8, 
    101988.8, 102017.5, 102053.9, 102097, 102116.2, 102130.4, 102135.8, 
    102142.4,
  102046.2, 102004.6, 101972.9, 101947.7, 101923.4, 101905.9, 101907.2, 
    101920.4, 101950.8, 101988.8, 102035, 102063.3, 102079.5, 102091.1, 
    102097.8,
  102038.8, 101989, 101945.3, 101907.2, 101876.8, 101847.8, 101840.7, 
    101850.6, 101883.2, 101924.1, 101973.8, 102007.8, 102023.4, 102038.2, 
    102046.5,
  102041.7, 101978.2, 101918.5, 101864.6, 101826.2, 101788.4, 101772.5, 
    101777.9, 101813.7, 101854.8, 101907, 101943.7, 101957.5, 101979.1, 101985,
  102043.7, 101976.5, 101902.6, 101824.2, 101778.4, 101733.6, 101712.9, 
    101714.3, 101746.4, 101787.1, 101840.9, 101876.2, 101890.5, 101905.7, 
    101910.3,
  102056.3, 101990.4, 101904, 101805.2, 101736.9, 101692.7, 101664.8, 
    101660.5, 101682.3, 101718.8, 101768.3, 101797.9, 101810, 101821.3, 101822,
  102067.4, 102004.4, 101920.8, 101814.8, 101722.8, 101667.6, 101636.8, 
    101621.6, 101625.4, 101655, 101695.1, 101719.6, 101724.6, 101728.9, 
    101722.4,
  102425, 102482.7, 102515, 102533.7, 102538.9, 102528.8, 102502.6, 102460.6, 
    102402.2, 102324.3, 102230.6, 102113, 101969.3, 101799.2, 101609.3,
  102423.6, 102488.1, 102520.2, 102547.9, 102556.4, 102550.7, 102527.1, 
    102487.7, 102430.4, 102356.8, 102266.9, 102154.1, 102014.8, 101847.1, 
    101655.7,
  102398.4, 102471.1, 102510.7, 102549.4, 102568.1, 102568.3, 102548.9, 
    102512.1, 102461.4, 102387.7, 102297.1, 102186.1, 102050.2, 101890.5, 
    101700,
  102375.6, 102455.2, 102507.8, 102548.8, 102574, 102577.8, 102562, 102529.4, 
    102479.2, 102413, 102324.7, 102214.5, 102077.2, 101916.2, 101731.2,
  102341.6, 102428.3, 102490.7, 102536.3, 102574.7, 102586.6, 102573.7, 
    102544, 102501, 102434.4, 102341.5, 102235.8, 102103.8, 101945.5, 101765.5,
  102307.8, 102393.4, 102468.6, 102520.7, 102568.1, 102584.1, 102576.2, 
    102548.6, 102505.2, 102438.4, 102354.8, 102253.9, 102121.3, 101966, 
    101792.4,
  102276, 102347.7, 102435.4, 102496.7, 102547.2, 102572.2, 102571.9, 
    102546.6, 102503.9, 102443.2, 102357.2, 102260.4, 102139.7, 101992, 
    101819.8,
  102257.7, 102309.3, 102397, 102467.4, 102525, 102554.1, 102559.9, 102536.3, 
    102499.9, 102447.2, 102367.4, 102267, 102143.5, 102002.4, 101841.5,
  102243.8, 102278.8, 102357.2, 102427.6, 102490.8, 102524.4, 102536.8, 
    102519.2, 102490.1, 102436.6, 102360, 102265.1, 102148.3, 102009.7, 
    101853.5,
  102237, 102262.3, 102320, 102383.1, 102452.6, 102491, 102509.2, 102497.8, 
    102469.6, 102419.8, 102350.6, 102256.2, 102140.9, 102006, 101856.7,
  102403.4, 102369.5, 102331, 102274.8, 102202.5, 102113.5, 102006.3, 
    101878.4, 101735.8, 101573.7, 101403.1, 101241.7, 101061.6, 100908.5, 
    100767.8,
  102426.4, 102394.9, 102356.8, 102300.2, 102229.1, 102137.9, 102031.9, 
    101902.5, 101761.1, 101592.8, 101417.2, 101238.8, 101049.8, 100887.5, 
    100738.5,
  102449.6, 102425.4, 102383.5, 102323.8, 102252.1, 102159.6, 102052.4, 
    101921.3, 101778.6, 101610.8, 101426.2, 101240.6, 101049.1, 100881.6, 
    100726.1,
  102471.7, 102445.1, 102407.2, 102348.8, 102274.8, 102180.1, 102068, 
    101934.3, 101782.9, 101609.8, 101417.6, 101223.1, 101025.7, 100850.5, 
    100687.1,
  102489.9, 102465, 102428.1, 102373.8, 102297.3, 102202.4, 102086.8, 
    101951.6, 101798.1, 101616.7, 101422.6, 101223.3, 101019.6, 100840.8, 
    100666.4,
  102510, 102483, 102445.8, 102391.3, 102316.8, 102220.9, 102100.1, 101962.4, 
    101805.9, 101619.9, 101424.7, 101217.2, 101007.9, 100821.8, 100635.7,
  102527.4, 102502.3, 102463.8, 102407.2, 102333.6, 102238.6, 102115.7, 
    101974.6, 101816, 101625.9, 101429.9, 101214.7, 101004.5, 100809.6, 
    100611.1,
  102544.9, 102517.2, 102477.9, 102421.2, 102346.4, 102251.4, 102129.6, 
    101984.8, 101824.5, 101632.4, 101437.6, 101212.3, 100996.7, 100788.8, 
    100580.2,
  102564.7, 102536.7, 102491.1, 102432.5, 102357.7, 102260.5, 102139.5, 
    101996, 101831.8, 101640.3, 101441.1, 101209.2, 100989.3, 100767.7, 
    100549.8,
  102581.8, 102552, 102505.3, 102443.1, 102364.6, 102266.7, 102145.8, 
    102000.7, 101834, 101643.9, 101439.3, 101200.2, 100976.6, 100739.2, 
    100514.6,
  101870.8, 101789, 101711.9, 101626.6, 101550.1, 101475.6, 101410.1, 
    101365.3, 101331.6, 101318.6, 101311, 101308.8, 101317.1, 101328.6, 
    101341.3,
  101888.5, 101795.3, 101710.5, 101620.3, 101530.6, 101443.8, 101362.5, 
    101306.4, 101259, 101240.9, 101222.1, 101206.7, 101208, 101209.3, 101214.1,
  101900.6, 101802.2, 101711.3, 101611.6, 101515.2, 101422.6, 101335.5, 
    101269.1, 101208.6, 101178.4, 101144.9, 101117.6, 101107.3, 101097, 
    101089.6,
  101910.4, 101810.9, 101704.8, 101590.5, 101483.5, 101379.9, 101284.8, 
    101203, 101136.7, 101088.3, 101044.6, 101005.3, 100986.1, 100963.1, 
    100945.4,
  101928.2, 101824.8, 101712.5, 101587.1, 101471.2, 101355.4, 101253.3, 
    101158.6, 101082.4, 101012.1, 100958.7, 100904.2, 100874.5, 100837.9, 
    100806.1,
  101948.4, 101835.4, 101718.7, 101583.3, 101456.5, 101330.1, 101216.8, 
    101106.6, 101018.3, 100931.8, 100863.3, 100795.6, 100752.3, 100703.4, 
    100658.1,
  101966.7, 101849.3, 101729.8, 101586.1, 101448.6, 101312.4, 101190.1, 
    101063.1, 100958.9, 100858.8, 100773.4, 100693.8, 100634.5, 100572.7, 
    100511.6,
  101985.9, 101866.5, 101739.3, 101592.7, 101443.4, 101298.6, 101162.9, 
    101021.3, 100902.4, 100787.6, 100683.2, 100588.8, 100514.6, 100440.2, 
    100364,
  102002.9, 101884.9, 101752.8, 101601.1, 101446.9, 101290, 101144.1, 
    100986.4, 100853.3, 100720.7, 100601.6, 100488.7, 100399.2, 100308.8, 
    100216.4,
  102020.1, 101901.4, 101768.9, 101612.3, 101452.7, 101281.4, 101129.9, 
    100954.4, 100808.4, 100657.7, 100525.4, 100391.9, 100286.5, 100179, 
    100070.7,
  101982.7, 102037.2, 102076.1, 102111.2, 102138.3, 102161.2, 102177, 
    102189.7, 102200.6, 102211.9, 102223.8, 102237.8, 102253.7, 102270.4, 
    102290.3,
  101905.9, 101942.3, 101972.9, 101998.3, 102022.7, 102041.1, 102049.5, 
    102055.2, 102061.9, 102068.4, 102076.5, 102085.1, 102096.3, 102110.4, 
    102127.6,
  101808.9, 101842.6, 101870.1, 101891.4, 101905.9, 101916.7, 101918.2, 
    101917.2, 101918.3, 101918.9, 101920.7, 101924.1, 101931.9, 101941.3, 
    101955.8,
  101715.1, 101739.7, 101760.2, 101776.7, 101782.4, 101787, 101782, 101775.5, 
    101769.8, 101763.6, 101758.6, 101755, 101756.3, 101760.2, 101769.4,
  101618.5, 101636.1, 101649.1, 101660.5, 101659.3, 101655.4, 101642.4, 
    101627.3, 101614.5, 101599.8, 101588, 101578.6, 101572.5, 101570, 101572.6,
  101523.8, 101534.8, 101536.3, 101541, 101533, 101519.6, 101499.2, 101476.1, 
    101454.7, 101433.3, 101413.6, 101394.8, 101380.1, 101369.3, 101365.4,
  101431.1, 101431.3, 101422.6, 101420.2, 101407.3, 101383.8, 101354.9, 
    101323.4, 101292, 101262.6, 101233.1, 101205.8, 101183.1, 101162.5, 
    101147.8,
  101343.3, 101330.1, 101312.8, 101298, 101281.9, 101246.5, 101213.2, 
    101170.8, 101130.1, 101092.2, 101053.2, 101014.9, 100980.1, 100950.4, 
    100924.5,
  101260.7, 101233.5, 101204.8, 101174.8, 101153.8, 101111, 101069.8, 
    101020.2, 100968.8, 100920.3, 100870.5, 100822.2, 100776.3, 100733.7, 
    100696.3,
  101183.3, 101142.6, 101102.1, 101059.6, 101029.2, 100980.6, 100930.5, 
    100871.1, 100808.9, 100749, 100689.2, 100627.5, 100567.8, 100514.7, 
    100463.7,
  101917.4, 101934.9, 101957.7, 101983.1, 102015.3, 102052.4, 102091, 
    102132.4, 102180.8, 102234.7, 102294.2, 102358.4, 102426.9, 102498.5, 
    102574.4,
  101808, 101815.1, 101834.1, 101853.8, 101882.1, 101913, 101951.2, 101991.2, 
    102038.3, 102087.7, 102144.3, 102205.4, 102273.3, 102344.9, 102420.8,
  101679.8, 101686.2, 101698, 101712.8, 101736.7, 101766.9, 101802.6, 
    101840.8, 101884.3, 101931.9, 101985.8, 102044.3, 102109.6, 102180.5, 
    102256,
  101551, 101552.1, 101555.6, 101565.5, 101582.9, 101607.9, 101639.5, 
    101675.6, 101714.2, 101762.5, 101814.6, 101873.9, 101938.8, 102009.4, 
    102084.8,
  101415.6, 101408.8, 101404.3, 101406.9, 101416, 101435.2, 101460.4, 
    101490.5, 101527.9, 101571.8, 101624.5, 101683.6, 101750.2, 101822.7, 
    101901.1,
  101277.4, 101261.1, 101246.1, 101238.7, 101239.6, 101250, 101267.2, 
    101290.8, 101321.5, 101362, 101411.5, 101471.4, 101540.5, 101616.3, 
    101698.1,
  101135.8, 101109.1, 101083.3, 101066.3, 101055.9, 101057.7, 101063.4, 
    101076.6, 101099.7, 101132.5, 101177.4, 101234.4, 101303.5, 101382.5, 
    101469.5,
  100992, 100955, 100913.7, 100885.6, 100864.8, 100855.1, 100850.4, 100853.5, 
    100868.3, 100891.5, 100929.1, 100980.9, 101046.6, 101126.3, 101216.8,
  100851.9, 100801.6, 100747.6, 100706.9, 100676.5, 100654.1, 100637.8, 
    100629, 100632.6, 100645.1, 100671.5, 100713.1, 100774.1, 100850.2, 
    100941.1,
  100714, 100651.2, 100584.4, 100534.7, 100486.7, 100454.8, 100426.2, 
    100405.9, 100399.5, 100402.3, 100416.3, 100449.6, 100497.9, 100567.5, 
    100654.1,
  101873.2, 101927.6, 101986.6, 102050, 102120.4, 102198.9, 102283.3, 
    102371.7, 102464.5, 102559.4, 102652.8, 102743.4, 102831.5, 102916.1, 
    102999.3,
  101739.5, 101784.8, 101837.1, 101896.5, 101963.6, 102039.9, 102123.4, 
    102212.1, 102306.5, 102404, 102501.3, 102597.2, 102690.1, 102779.8, 
    102866.2,
  101577.9, 101628, 101675.7, 101734.3, 101797.8, 101872.1, 101953.1, 
    102042.7, 102138.3, 102238.6, 102340.3, 102441, 102538.3, 102632.6, 
    102724.7,
  101412.4, 101463.8, 101507, 101564.7, 101622.9, 101695.3, 101773.4, 
    101859.9, 101954.7, 102055, 102156, 102260, 102362.6, 102461.2, 102557.4,
  101230.3, 101284.1, 101323.8, 101380.4, 101436.9, 101507.4, 101582.2, 
    101669.2, 101760.8, 101860.3, 101962.4, 102065.5, 102169.6, 102273.8, 
    102375.7,
  101042.5, 101094.7, 101128.5, 101185.3, 101238.7, 101307, 101381.1, 
    101466.2, 101557.4, 101656.6, 101754.5, 101857.2, 101961.4, 102064.8, 
    102167.4,
  100847.7, 100894.9, 100922.5, 100977.2, 101027, 101095.6, 101167, 101251.9, 
    101343.9, 101443.8, 101542.5, 101643.3, 101744.4, 101848.9, 101950.7,
  100653.5, 100693.1, 100716.7, 100766, 100812.4, 100879.1, 100947.7, 
    101031.5, 101121.2, 101221.4, 101319.1, 101420.2, 101520.6, 101622.7, 
    101723.9,
  100466.9, 100492.8, 100510.4, 100553.3, 100596.5, 100658.3, 100727.6, 
    100805.7, 100891.7, 100990.9, 101090.7, 101191.8, 101291.3, 101392.5, 
    101490.8,
  100291, 100300.4, 100311.8, 100347.7, 100385, 100442.6, 100504.4, 100583.1, 
    100664.4, 100757.8, 100854, 100953.1, 101052.7, 101153, 101250.6,
  102119.6, 102160.3, 102209.3, 102257.9, 102311.9, 102367.1, 102424.3, 
    102481.2, 102543.1, 102609.2, 102678.3, 102748.9, 102822.9, 102899.3, 
    102977.3,
  102011.4, 102042.1, 102088.4, 102133, 102185, 102237.5, 102293.2, 102348.2, 
    102409.2, 102476.4, 102546.1, 102619, 102695.1, 102772.3, 102851.6,
  101892.2, 101919.8, 101961.8, 102001.1, 102047.3, 102096.2, 102149, 
    102204.5, 102265.8, 102331.8, 102401.4, 102473.8, 102550.2, 102628.9, 
    102709.6,
  101773.1, 101796.4, 101830.6, 101866.1, 101908.5, 101952, 102001.4, 
    102053.1, 102111.4, 102175.2, 102244.1, 102315.5, 102391.4, 102470.2, 
    102552,
  101648.6, 101667.8, 101694.7, 101726.1, 101764.6, 101804.4, 101849.6, 
    101899, 101954.5, 102012.5, 102075.7, 102144.3, 102217.6, 102295.3, 
    102375.7,
  101514.6, 101530.6, 101550.8, 101578.8, 101613.1, 101650.5, 101692.9, 
    101739.4, 101791.5, 101848.2, 101908.7, 101972.8, 102041.1, 102112.7, 
    102188.3,
  101368.2, 101377.8, 101393.6, 101417.4, 101447.5, 101484.7, 101525.7, 
    101571.4, 101623, 101676.4, 101733.6, 101793.5, 101861, 101929.3, 102005.6,
  101207.5, 101211, 101219.2, 101236.3, 101262.3, 101296.7, 101336.2, 
    101382.9, 101437.6, 101493.7, 101553, 101612.3, 101678, 101746.6, 101816.4,
  101027.5, 101022.7, 101020.6, 101031.6, 101049.4, 101080.5, 101118.8, 
    101166.7, 101222.2, 101283.1, 101348.2, 101414.9, 101484.4, 101555.4, 
    101628,
  100831.7, 100817, 100801.9, 100803.9, 100812.1, 100836.5, 100869.7, 100916, 
    100975, 101043.1, 101116.2, 101193, 101271.4, 101351.1, 101429,
  102147.1, 102196.8, 102249.8, 102307.4, 102374, 102445.2, 102522.3, 
    102598.3, 102679.8, 102761.2, 102843.9, 102926.2, 103009.8, 103091.3, 
    103170.7,
  102056.7, 102096.2, 102145.6, 102199.5, 102261.5, 102331.2, 102406.4, 
    102483.9, 102566.8, 102651.1, 102736.8, 102821.9, 102907.6, 102992.5, 
    103074.9,
  101950.4, 101985.2, 102031.5, 102080.6, 102141.5, 102209.1, 102284.8, 
    102363.3, 102447.4, 102531.6, 102619.2, 102706.9, 102794.6, 102883, 
    102969.1,
  101844.1, 101873.3, 101912, 101956.4, 102012.6, 102076.3, 102149.5, 
    102227.6, 102312, 102399.4, 102489.3, 102577.7, 102669.3, 102758.2, 
    102848.8,
  101728.4, 101751.3, 101785.3, 101823.4, 101874.1, 101934, 102002.8, 
    102079.6, 102164, 102252.6, 102344.7, 102436.4, 102528.9, 102622.8, 
    102713.3,
  101610.2, 101626.8, 101651.1, 101683.9, 101727.5, 101781.8, 101846.4, 
    101919.8, 102003.4, 102092.3, 102184.5, 102279.5, 102375.4, 102470.4, 
    102566.9,
  101486.5, 101497.5, 101513.7, 101537.7, 101574.7, 101621.3, 101678.3, 
    101747.1, 101829, 101918.2, 102011.3, 102106.7, 102206.5, 102305.6, 
    102405.5,
  101359.6, 101368.5, 101379.6, 101397.2, 101426, 101463.4, 101512.9, 
    101573.5, 101648.4, 101733, 101825, 101921.5, 102021.7, 102125.4, 102226.5,
  101225.7, 101232.5, 101241.7, 101261.3, 101285.2, 101317.4, 101354.6, 
    101404, 101468, 101545, 101631.6, 101724.7, 101824.5, 101927.2, 102031.5,
  101083.7, 101089.4, 101094, 101113.3, 101138.9, 101175.3, 101211, 101252.1, 
    101300.4, 101363.3, 101437.6, 101525.1, 101617.9, 101719.4, 101822.9,
  102812.6, 102881.2, 102948.9, 103014.1, 103081.3, 103145.7, 103208.6, 
    103269.8, 103334, 103392.5, 103448.5, 103502.9, 103559.4, 103601.6, 
    103635.9,
  102748.6, 102813, 102881.1, 102948.9, 103018.5, 103087.3, 103152.2, 
    103216.2, 103282.6, 103344.4, 103401.5, 103454.5, 103513.1, 103562.1, 
    103599.8,
  102672.6, 102737.5, 102806.6, 102877, 102947.2, 103018.2, 103087.4, 
    103154.7, 103223.8, 103289.5, 103351.3, 103406.7, 103462.1, 103516.4, 
    103559.7,
  102590.9, 102651.4, 102720.5, 102792.2, 102865.2, 102936.5, 103009.7, 
    103080.8, 103153.2, 103223.7, 103287.6, 103348.3, 103404.5, 103457.1, 
    103505.8,
  102504.3, 102561.8, 102628.8, 102698.1, 102773.1, 102846.4, 102919.9, 
    102993.9, 103071, 103144.7, 103212.9, 103276, 103337.7, 103392.2, 103438.8,
  102415.9, 102466, 102530, 102597.9, 102672.6, 102746.3, 102821.7, 102895.5, 
    102973.5, 103050.4, 103124.4, 103191.5, 103257.7, 103315.3, 103363.3,
  102329, 102367.1, 102425.8, 102490.6, 102562.3, 102637.3, 102711.9, 
    102787.4, 102865.3, 102943.7, 103023, 103095, 103165, 103226.3, 103278,
  102243.2, 102272.8, 102320.2, 102376.3, 102443.2, 102517, 102591.6, 
    102667.3, 102748, 102826.5, 102906.8, 102982.4, 103055.3, 103119.5, 
    103175.2,
  102146.8, 102176.1, 102215.3, 102260.3, 102318.1, 102384.4, 102458, 
    102534.1, 102613.3, 102695, 102775.4, 102854.2, 102929.1, 102997.6, 
    103058.2,
  102041.6, 102064.2, 102099.5, 102138.7, 102188.5, 102245.6, 102313.1, 
    102387.6, 102466.3, 102548, 102628.4, 102708.7, 102786.2, 102857.6, 102920,
  103180.7, 103246.2, 103309.9, 103373.3, 103435.2, 103501, 103559.2, 103613, 
    103666.5, 103711.5, 103754.1, 103793.4, 103826.1, 103846.3, 103853,
  103155.8, 103222.5, 103288.3, 103352.9, 103418.1, 103485.8, 103549.3, 
    103603.6, 103651.8, 103701.6, 103744.5, 103782.2, 103810.7, 103830.5, 
    103832.5,
  103125, 103193, 103260.8, 103327.4, 103394.9, 103461.4, 103524.3, 103579.6, 
    103633.6, 103681.1, 103723.9, 103763.3, 103790.8, 103805.6, 103806.8,
  103083.2, 103154.1, 103226.2, 103295.3, 103361.2, 103427.3, 103491.1, 
    103550.5, 103603.2, 103649.5, 103689.9, 103726, 103751.6, 103765, 103764.3,
  103033, 103104.4, 103180.6, 103252.3, 103319.9, 103382.3, 103445.6, 
    103505.2, 103557.4, 103605, 103644.7, 103679.1, 103704.7, 103717.5, 
    103711.3,
  102971.2, 103043.5, 103121.6, 103195.7, 103267.3, 103331.7, 103391.5, 
    103449.1, 103503.4, 103549.7, 103590.1, 103624.5, 103645.1, 103654.8, 
    103654.1,
  102902.6, 102974.3, 103051.9, 103126.5, 103201.6, 103266.7, 103327.6, 
    103383.9, 103436.8, 103484.6, 103523.2, 103557.3, 103579.3, 103587.1, 
    103585.3,
  102827.4, 102898.3, 102975.2, 103047.9, 103121, 103188.8, 103250.9, 
    103307.9, 103361.1, 103409.8, 103448.6, 103479.3, 103500.8, 103507.3, 
    103500.4,
  102744, 102814.3, 102891.6, 102962.6, 103032.4, 103097.2, 103163.2, 
    103221.7, 103275.4, 103321.7, 103358.7, 103388.6, 103410, 103413.9, 
    103402.3,
  102654.3, 102723.7, 102797.2, 102868.3, 102936.6, 103001.9, 103064.6, 
    103124.1, 103176.1, 103220.6, 103258.8, 103284.3, 103299.3, 103302.3, 
    103288.3,
  103175.4, 103233.7, 103287.2, 103336.2, 103382.3, 103429.3, 103473.6, 
    103507.2, 103544.3, 103573.2, 103603.1, 103618.5, 103626.6, 103632.2, 
    103627.2,
  103172.9, 103230.5, 103286.9, 103334.3, 103381.6, 103428.4, 103472.1, 
    103506.9, 103541.3, 103570.2, 103599.2, 103617.2, 103628.7, 103627.2, 
    103612.9,
  103160.1, 103215.1, 103270.4, 103321.1, 103371, 103417.4, 103458.5, 
    103495.3, 103528.8, 103558.8, 103580.9, 103598.2, 103606.7, 103609, 
    103592.6,
  103134.3, 103193.3, 103248.3, 103300.7, 103349, 103394.9, 103434.7, 
    103470.2, 103505.4, 103532.3, 103554.7, 103567.8, 103573.1, 103570.1, 
    103558.7,
  103099.8, 103161.4, 103215.3, 103266.8, 103315.8, 103360.8, 103401.1, 
    103436.7, 103468.6, 103497.8, 103518.7, 103533.4, 103539, 103532.6, 
    103513.1,
  103055.5, 103117.1, 103172.1, 103224.4, 103270.9, 103316.3, 103355.5, 
    103390.8, 103421.4, 103445.9, 103469.9, 103491, 103497.5, 103493.1, 
    103479.5,
  103001.5, 103063, 103116.6, 103169.6, 103216, 103259.8, 103297.3, 103330.1, 
    103361, 103383.3, 103402.9, 103419.4, 103431.6, 103429.8, 103422.3,
  102940.9, 102999.2, 103054, 103104.1, 103151, 103192.6, 103228.4, 103260.9, 
    103289.5, 103311.4, 103328, 103339, 103350.3, 103351.8, 103345.9,
  102874.1, 102929.5, 102984.5, 103032.9, 103079.6, 103119.8, 103156.2, 
    103186, 103210.9, 103230.2, 103243.6, 103251.1, 103254.8, 103251.7, 
    103240.6,
  102801.2, 102851.9, 102906.6, 102952.4, 103000.4, 103041, 103076.9, 
    103105.2, 103126.7, 103145.6, 103159.9, 103165.9, 103164.5, 103158.6, 
    103145.2,
  103146.6, 103186, 103224.8, 103257.9, 103285.2, 103308.8, 103331.7, 
    103347.2, 103353.1, 103355.5, 103352.9, 103341.8, 103328.2, 103301.6, 
    103255.4,
  103172.8, 103215.8, 103256.1, 103286.2, 103312.4, 103336, 103359.5, 
    103375.5, 103385.5, 103389.8, 103388.6, 103382.3, 103370, 103338.6, 
    103289.7,
  103194.4, 103235.4, 103273.4, 103304.5, 103332.1, 103359.8, 103385, 
    103398.3, 103412.2, 103416.6, 103412.5, 103403.7, 103386.3, 103361.2, 
    103313.7,
  103207.9, 103248.8, 103285.6, 103317.8, 103347.2, 103376, 103397.6, 
    103412.6, 103430.1, 103436.2, 103437.7, 103426.4, 103402.4, 103372.7, 
    103322.4,
  103221.1, 103258.6, 103295.9, 103330.6, 103358.4, 103384.6, 103402.8, 
    103411.2, 103421.8, 103432.3, 103444.2, 103435.8, 103409.7, 103371.2, 
    103318.7,
  103227.5, 103267, 103303.9, 103339.4, 103363.7, 103383.5, 103405.3, 
    103408.8, 103412.5, 103422.7, 103436.2, 103433.5, 103410.2, 103366.5, 
    103303,
  103232.1, 103276.2, 103315.2, 103349.6, 103368.7, 103385.5, 103400.5, 
    103407.6, 103407.1, 103409.5, 103423.5, 103418.7, 103396.6, 103349.6, 
    103290.5,
  103228.4, 103277.6, 103316.5, 103354.6, 103380.4, 103395.4, 103406.8, 
    103403.4, 103394.9, 103391.4, 103393.5, 103395, 103374.4, 103327.1, 
    103267.1,
  103222.8, 103275.1, 103318.6, 103360.1, 103387.6, 103402.6, 103418.3, 
    103413.5, 103397.8, 103378.9, 103364.2, 103360.5, 103342.8, 103297.5, 
    103234.3,
  103207.9, 103259, 103311.9, 103360.9, 103389.7, 103409, 103425.3, 103430.2, 
    103404, 103380.9, 103358.6, 103336.4, 103305.9, 103259.8, 103189.3,
  103168.2, 103182.9, 103201.2, 103208.9, 103208.4, 103206.1, 103196.2, 
    103180.8, 103162.9, 103134.7, 103104.3, 103062.3, 103016.4, 102959.8, 
    102889.3,
  103268, 103279.6, 103296.3, 103299.7, 103298.8, 103289.5, 103278.6, 
    103261.4, 103237.5, 103210.4, 103176, 103131.5, 103081.8, 103023, 102949.6,
  103351.4, 103364, 103379.7, 103384.4, 103384.3, 103375.6, 103360.9, 
    103339.5, 103310.6, 103278.2, 103240.8, 103195.8, 103140.2, 103080.6, 
    103005,
  103435.5, 103448.5, 103462.3, 103469.5, 103465.2, 103454.1, 103436.8, 
    103412.2, 103380.4, 103341.8, 103301.5, 103253.2, 103195.2, 103130.6, 
    103052.1,
  103508.7, 103523.5, 103547.9, 103553.2, 103550.9, 103536, 103509.1, 
    103477.5, 103440.2, 103398, 103353.8, 103306.3, 103244.2, 103176, 103091.2,
  103579.6, 103604.1, 103624.9, 103625.6, 103620.8, 103600.1, 103572.2, 
    103537.1, 103492.9, 103446.7, 103396.6, 103347, 103281.8, 103214.3, 
    103121.9,
  103637.8, 103665.8, 103689.9, 103690.3, 103683.1, 103655.1, 103621.9, 
    103585.9, 103537.2, 103482.2, 103436.1, 103380.6, 103311.1, 103238.3, 
    103142,
  103683.3, 103714.9, 103732.7, 103739, 103729.4, 103709.2, 103676.6, 103618, 
    103571.5, 103509.3, 103460.2, 103402, 103331.9, 103250.7, 103153.1,
  103721.6, 103745, 103754.3, 103777.2, 103766.1, 103745.1, 103712.4, 
    103667.7, 103598.9, 103530.4, 103476.8, 103412.5, 103341.1, 103251.8, 
    103149.2,
  103742, 103763.3, 103767.5, 103805.3, 103790.6, 103769.8, 103734, 103687.2, 
    103621, 103543.1, 103480.4, 103418.6, 103340.4, 103244.4, 103133.1,
  101815.9, 101834.2, 101904.6, 101999.7, 102087.9, 102184, 102246, 102277.9, 
    102269.9, 102240, 102194.6, 102117.5, 102029.5, 101916.1, 101790.1,
  102035.7, 102058.1, 102102.9, 102159.4, 102226.6, 102303.3, 102354.7, 
    102383, 102376.8, 102347.9, 102297.9, 102222.6, 102128.5, 102020.4, 
    101901.9,
  102245.7, 102253.4, 102279, 102323.2, 102374.7, 102426.4, 102470.3, 
    102495.1, 102488.6, 102455.8, 102400.3, 102326.4, 102232.6, 102123.3, 
    102003.7,
  102463.5, 102458.3, 102472.7, 102501.9, 102532.6, 102561.8, 102588.6, 
    102603.3, 102598.2, 102565.9, 102510.9, 102431.3, 102333.6, 102220.1, 
    102100.4,
  102656.6, 102647.7, 102652.2, 102667.4, 102687.9, 102704.2, 102718.4, 
    102718.2, 102707, 102665.8, 102608, 102531.2, 102433.2, 102319.1, 102191.7,
  102834.3, 102829.6, 102828.9, 102832.4, 102837.7, 102846.1, 102850.7, 
    102842.5, 102818, 102771.9, 102705.8, 102621.7, 102523.5, 102404.9, 
    102279.2,
  102983.6, 102985.6, 102981.7, 102985.3, 102982, 102981, 102969.8, 102951.2, 
    102920.7, 102870.9, 102798.9, 102713.4, 102609, 102490.8, 102357.4,
  103135.7, 103127.6, 103122.4, 103119.6, 103109.3, 103094.9, 103076.1, 
    103051.4, 103012.3, 102961.5, 102880.7, 102791.4, 102684.1, 102562.4, 
    102426.1,
  103265.6, 103253.2, 103245.3, 103236.3, 103221.9, 103201.1, 103175.2, 
    103141.7, 103097.3, 103036.8, 102961.2, 102858.1, 102747.8, 102624.7, 
    102485.5,
  103378.4, 103366.3, 103351.9, 103337.9, 103323.2, 103299.3, 103265.7, 
    103225.6, 103170.9, 103102.8, 103024.5, 102917.5, 102800.2, 102674, 
    102532.1,
  100001.8, 99705.42, 99508.27, 99405.33, 99396.21, 99437.3, 99511.81, 
    99622.7, 99764.55, 99890.83, 99971.27, 100029.3, 100070, 100065, 100040.3,
  100092.6, 99823.34, 99607.77, 99458.37, 99396.31, 99398.83, 99438.94, 
    99525.44, 99633.91, 99796.37, 99937.66, 100029.4, 100089.3, 100122.1, 
    100139.1,
  100240.4, 99989.96, 99743.22, 99533.17, 99414.29, 99359.18, 99379.12, 
    99433.64, 99528.98, 99671.64, 99842.75, 99995.34, 100099.5, 100164.5, 
    100196,
  100398.3, 100160.4, 99899.87, 99672.1, 99512.3, 99397.48, 99371.2, 
    99386.95, 99470.56, 99587.56, 99760.91, 99949.04, 100093, 100185.8, 
    100247.6,
  100559.8, 100342.9, 100085, 99856.97, 99653, 99497.3, 99409.47, 99391.89, 
    99451.93, 99558.66, 99707.61, 99884.42, 100074.9, 100198, 100280.9,
  100744.9, 100534.9, 100285, 100053, 99834.81, 99650.05, 99517.16, 99459.59, 
    99483.53, 99590.09, 99717.95, 99872.78, 100066.8, 100215.1, 100315.6,
  100940.5, 100735.2, 100502.2, 100271, 100046, 99840.94, 99679.13, 99578.34, 
    99557.91, 99644.07, 99765.67, 99895.56, 100066.3, 100239.1, 100342.1,
  101131.4, 100935.8, 100713.7, 100501.1, 100278.4, 100070.4, 99889.37, 
    99750.66, 99685.56, 99719.97, 99831.49, 99960.11, 100099.9, 100277.9, 
    100383.1,
  101312, 101131.6, 100922.8, 100722.6, 100514.5, 100310.2, 100125.4, 
    99962.45, 99860.91, 99842.09, 99923.67, 100042.2, 100159.5, 100327.9, 
    100434.6,
  101495, 101323.3, 101126.6, 100942, 100748.3, 100554.9, 100373.3, 100205.1, 
    100083.2, 100027.2, 100063.8, 100152.6, 100251.2, 100395.8, 100501.8,
  99940.42, 99970.08, 100023.8, 100093, 100185.7, 100290, 100411.1, 100539.2, 
    100676.4, 100815, 100949, 101080.5, 101208.3, 101333.6, 101457.1,
  99865.8, 99900.09, 99956.65, 100013.9, 100087.1, 100182.8, 100293, 
    100420.2, 100562.1, 100711.3, 100852.4, 100989.7, 101122.1, 101252, 
    101379.4,
  99790.1, 99812.27, 99852.35, 99895.35, 99967.59, 100055.6, 100160.6, 
    100284.3, 100432, 100592, 100741, 100885.8, 101022.3, 101156.4, 101288.7,
  99723.04, 99733.37, 99761.22, 99791.64, 99851.45, 99923.81, 100014.5, 
    100127.5, 100278.8, 100447.8, 100616.5, 100766.8, 100908, 101045.4, 
    101182.6,
  99662.08, 99656.23, 99663.83, 99679.91, 99732.51, 99792.55, 99868.8, 
    99970.38, 100121.1, 100287.7, 100467.2, 100628.2, 100780.3, 100919.8, 
    101061.1,
  99614.04, 99590.04, 99582.95, 99581.15, 99626.66, 99672.71, 99737.93, 
    99824.25, 99967.73, 100132.6, 100300.6, 100466.3, 100627.2, 100776, 
    100922.9,
  99575.3, 99530.28, 99510.23, 99493.82, 99529.27, 99563.52, 99615.74, 
    99688.57, 99818.24, 99965.33, 100124.5, 100294.1, 100459.9, 100616, 
    100765.8,
  99545.45, 99492.8, 99449.94, 99422.52, 99440.62, 99467.39, 99500.23, 
    99558.95, 99662.2, 99795.11, 99950.9, 100113.5, 100281, 100442.4, 100595.7,
  99525.7, 99477.73, 99397.09, 99365.2, 99356.41, 99374.1, 99385.04, 
    99416.79, 99487.66, 99609.02, 99759.26, 99930.14, 100089.8, 100259.9, 
    100411,
  99533.43, 99468.81, 99368.25, 99318.43, 99278.81, 99282.9, 99273.52, 
    99276.59, 99306.44, 99393.02, 99542.49, 99731.53, 99888.66, 100064.6, 
    100218.1,
  101800.7, 101867.4, 101921.3, 101973.1, 102021.6, 102064, 102098.6, 
    102129.7, 102156.8, 102179.8, 102200.7, 102221.4, 102242, 102259.3, 102276,
  101726.7, 101782.8, 101834.5, 101883.2, 101929, 101970, 102005.3, 102036, 
    102063.2, 102086, 102106.5, 102125, 102142.5, 102158.2, 102170.4,
  101631.7, 101686.7, 101735.4, 101780.8, 101822.1, 101861.3, 101893.8, 
    101921.7, 101946.6, 101969.1, 101987.1, 102002.8, 102017.9, 102031.7, 
    102044.7,
  101531.4, 101587.3, 101632.1, 101674.6, 101709, 101744.9, 101775.3, 
    101800.9, 101824, 101844.1, 101861.3, 101875.2, 101887, 101896.9, 101907.5,
  101421.4, 101476.1, 101518.9, 101558.2, 101588.6, 101618.2, 101640.3, 
    101663.9, 101682.7, 101698.8, 101711.7, 101722.3, 101731.5, 101739.3, 
    101744.3,
  101303.3, 101357.1, 101398.4, 101434.8, 101461.5, 101485.4, 101501.3, 
    101516.5, 101530.6, 101543.1, 101551.2, 101558.4, 101562.9, 101565.6, 
    101568.1,
  101177.7, 101228.6, 101267.7, 101302.2, 101324.9, 101343.7, 101352.5, 
    101360.3, 101364.9, 101370.2, 101372.9, 101372.8, 101371.5, 101370.2, 
    101367.7,
  101049.1, 101098.6, 101133, 101164.1, 101179.8, 101192.1, 101193.9, 
    101193.2, 101190.9, 101187.5, 101182.7, 101176.2, 101169, 101163, 101157.5,
  100916.6, 100963.5, 100992.6, 101020.3, 101030.9, 101036.2, 101030.3, 
    101020, 101008.5, 100995.1, 100981.8, 100965.7, 100949.1, 100935, 100925.8,
  100782.1, 100824.8, 100848.6, 100870.5, 100876.3, 100874, 100860.4, 
    100840.9, 100818.8, 100795.4, 100770.2, 100747, 100724, 100702.1, 100689,
  102462, 102486.7, 102495.2, 102505.1, 102511.2, 102515.8, 102517.9, 
    102517.2, 102517.5, 102516.2, 102512, 102503.3, 102493.3, 102474.7, 
    102451.8,
  102402.7, 102419.5, 102426.1, 102436.3, 102443.4, 102450.2, 102452.3, 
    102451.5, 102447.2, 102445, 102441, 102434.7, 102424.7, 102412, 102396.5,
  102333.4, 102341.6, 102351, 102360.9, 102364.1, 102369.5, 102370.2, 
    102368.8, 102368.1, 102365.9, 102363, 102354.1, 102345.8, 102334.8, 
    102319.9,
  102249.2, 102257.5, 102267.1, 102271.6, 102278.9, 102282.1, 102283.1, 
    102280.5, 102276.9, 102272.4, 102267.1, 102262.4, 102252.8, 102241.6, 
    102229.5,
  102168.1, 102170, 102178.1, 102182.5, 102187.2, 102186.6, 102185.9, 
    102181.8, 102178, 102173.4, 102166.5, 102156.6, 102145.5, 102133.4, 
    102120.9,
  102076.5, 102076.8, 102081.8, 102081.5, 102083.9, 102083.6, 102081.8, 
    102076.9, 102073.8, 102066.8, 102061.1, 102052.3, 102043.4, 102032.2, 
    102022.5,
  101978, 101978.2, 101978.8, 101979.6, 101981.6, 101981.1, 101977.2, 
    101972.7, 101969.4, 101965, 101960.6, 101953.9, 101946.9, 101938, 101930.3,
  101883.1, 101881, 101878.5, 101877.2, 101876.9, 101877.6, 101876, 101872.7, 
    101870.4, 101867.6, 101863.6, 101857.6, 101853.2, 101846.6, 101838.4,
  101785.3, 101780.1, 101776.6, 101772.3, 101771, 101769.8, 101768.5, 
    101764.8, 101762.6, 101759.2, 101758.7, 101755, 101749.7, 101744, 101735.9,
  101689.6, 101680.5, 101674.1, 101666, 101662.6, 101662.3, 101661.2, 
    101660.9, 101659.7, 101657.7, 101652.6, 101648.5, 101641.3, 101633.1, 
    101621.2,
  102905.5, 102889.6, 102858.8, 102818.9, 102766.6, 102695.6, 102615, 
    102513.1, 102386.9, 102247.9, 102104.8, 101964.8, 101825.4, 101685.3, 
    101543.9,
  102901.6, 102879.8, 102855.2, 102818.9, 102774.8, 102714.2, 102642.9, 
    102560.5, 102450.5, 102326.1, 102189.4, 102048.4, 101913.5, 101775.2, 
    101637.9,
  102902.1, 102877.9, 102853.7, 102819.4, 102783.6, 102730.5, 102667.3, 
    102594.4, 102502.3, 102390.1, 102261.5, 102123.5, 101986.7, 101848.8, 
    101710.2,
  102885.2, 102860.7, 102840.3, 102806.3, 102770.1, 102721.5, 102673.1, 
    102607.1, 102528.5, 102436.8, 102326.3, 102199, 102065.8, 101930.7, 
    101796.1,
  102870.9, 102850.7, 102829.8, 102797.2, 102759.9, 102711.7, 102662.6, 
    102604.4, 102537.5, 102457, 102361.1, 102254.8, 102132, 102003.7, 101873.3,
  102847.4, 102831.6, 102808.1, 102778.1, 102742.7, 102697.5, 102646.5, 
    102590, 102530.1, 102462.7, 102382.3, 102289.1, 102184.1, 102069.8, 
    101946.9,
  102838.9, 102820.7, 102793.7, 102757.6, 102721, 102680.1, 102635.6, 
    102578.7, 102521.9, 102457.4, 102389.8, 102314.8, 102220, 102120.6, 
    102007.4,
  102823.3, 102799.4, 102776, 102743.1, 102708.1, 102667.5, 102626, 102568.2, 
    102511.4, 102452.3, 102388.9, 102321.6, 102237.4, 102148.5, 102046.2,
  102815.8, 102792.5, 102765.3, 102721.3, 102686.8, 102642.8, 102600.6, 
    102548.2, 102496.5, 102442.2, 102380.6, 102319, 102238.8, 102153, 102062.7,
  102790.7, 102771.2, 102742.9, 102709.6, 102669, 102622.6, 102578.2, 
    102532.4, 102474.7, 102420.9, 102363.1, 102296.9, 102222.1, 102143, 
    102053.7,
  102205.7, 102070.5, 101900.8, 101747.7, 101564.3, 101408.5, 101266, 
    101147.4, 101047.8, 100953.3, 100860.9, 100780.5, 100717.8, 100667.8, 
    100640.6,
  102248.6, 102113.5, 101947.9, 101788.8, 101578.4, 101420.5, 101280.2, 
    101147.6, 101027.8, 100923.6, 100823.4, 100736.8, 100669.3, 100619.8, 
    100578.8,
  102294.5, 102154.2, 102007.6, 101837.2, 101637.7, 101474, 101313.7, 
    101167.6, 101027.3, 100899.1, 100784.4, 100691.8, 100618.2, 100557.1, 
    100502.1,
  102350.3, 102214.3, 102074, 101892.9, 101700.2, 101523.9, 101352.3, 
    101200.3, 101046.4, 100896.9, 100762.1, 100650.6, 100565.5, 100492, 
    100435.1,
  102426.4, 102294.1, 102155.5, 101965.2, 101774.8, 101584, 101417.8, 101251, 
    101082.1, 100919.5, 100761.1, 100625.5, 100515.3, 100424.3, 100356.5,
  102510.4, 102393, 102239.3, 102051.1, 101848.2, 101645.5, 101477.2, 
    101305.5, 101129.6, 100953.9, 100778.4, 100620, 100481.8, 100368.1, 
    100283.3,
  102592.6, 102480.3, 102319, 102138.8, 101934.9, 101727.1, 101550.6, 
    101369.1, 101189, 101006, 100815.2, 100634.1, 100469.9, 100329, 100218,
  102654.6, 102544.9, 102395.8, 102222.1, 102024.7, 101814, 101628.8, 101440, 
    101255.8, 101063.4, 100867.2, 100669.8, 100479.9, 100314.5, 100181.4,
  102707, 102602.9, 102473, 102307.1, 102119.1, 101912.2, 101721.1, 101527.4, 
    101335.1, 101136.1, 100931.4, 100723, 100513.6, 100323.3, 100171.8,
  102773.4, 102663.5, 102537.1, 102380, 102208.9, 102014.9, 101820.1, 101624, 
    101424.7, 101219.6, 101009.4, 100794, 100569.1, 100360.7, 100191.3,
  100538, 100506.3, 100490.3, 100523.1, 100594.1, 100734.6, 100855.2, 
    101010.4, 101186.2, 101360.5, 101538.2, 101709, 101861.8, 102000.5, 102129,
  100635.2, 100506.8, 100460.1, 100503, 100554.9, 100685.5, 100807.6, 100955, 
    101117.7, 101281, 101453, 101617.8, 101765, 101898.6, 102026.1,
  100711.4, 100545.8, 100500.6, 100527.4, 100548.1, 100635.3, 100752.5, 
    100889.1, 101037.1, 101194, 101357.5, 101518.2, 101661.6, 101793.5, 
    101920.5,
  100832, 100668.4, 100555.4, 100522.4, 100551.2, 100577.3, 100709.2, 
    100833.4, 100975.6, 101120.8, 101274.8, 101428.8, 101566.7, 101692.2, 
    101813.5,
  100988.3, 100794.5, 100666.9, 100567.3, 100586.5, 100546.1, 100681.9, 
    100776.3, 100913.8, 101040.4, 101186.3, 101331.5, 101465.9, 101585.4, 
    101700.9,
  101127.3, 100912.2, 100781.4, 100612, 100609.9, 100530.6, 100662.6, 100729, 
    100857.6, 100969.9, 101106.7, 101237, 101364.9, 101476.6, 101584.6,
  101240.9, 101018.9, 100877.1, 100664.8, 100631.7, 100515.4, 100634.4, 
    100682.3, 100797.3, 100894, 101017.7, 101131.2, 101251.2, 101355.4, 
    101459.8,
  101351, 101126.9, 100962.2, 100723.9, 100642.7, 100503.4, 100600.8, 
    100643.2, 100739.8, 100821.2, 100930.4, 101021.7, 101133.1, 101225.5, 
    101326,
  101463, 101242.6, 101051.8, 100791.6, 100668.5, 100500.6, 100568.1, 
    100599.5, 100685.3, 100740, 100833.7, 100903.8, 101001.9, 101087.7, 
    101180.3,
  101576.7, 101356.9, 101161.3, 100877.5, 100713.9, 100523.9, 100534.1, 
    100561.3, 100634.2, 100662.4, 100735.6, 100779.7, 100859.9, 100940, 
    101025.9,
  100894, 101188.4, 101401.7, 101633, 101821.9, 101997.9, 102141.8, 102265.5, 
    102374.8, 102468.6, 102547.4, 102613.4, 102665.6, 102701.6, 102720.9,
  100640.8, 100974.2, 101213.2, 101482.2, 101695.6, 101889.5, 102054.5, 
    102194.4, 102312.4, 102414.3, 102502.9, 102572.6, 102627, 102656.5, 102676,
  100346.1, 100741.9, 101021.2, 101324.4, 101566.3, 101778.2, 101960.7, 
    102113.8, 102248.7, 102356.3, 102451.6, 102526, 102588.8, 102626.3, 
    102644.3,
  100083, 100475.5, 100844.9, 101145.4, 101435, 101663.2, 101863.6, 102032.3, 
    102178.3, 102296.8, 102401, 102477.7, 102540.1, 102577.5, 102600.3,
  99905.37, 100258.6, 100694.4, 100970.5, 101299.3, 101559.3, 101765.7, 
    101946.2, 102104.9, 102229.5, 102342.3, 102424.1, 102490.1, 102529.3, 
    102553.3,
  99817.41, 100104.2, 100562.4, 100861.2, 101160, 101447.8, 101679.8, 
    101858.4, 102034.6, 102161.1, 102278.3, 102364.8, 102435, 102473.1, 102494,
  99820.86, 100008.2, 100429.2, 100779, 101069.2, 101322.8, 101606.3, 
    101769.7, 101960.8, 102094.4, 102209.4, 102298.4, 102368.9, 102415.3, 
    102432.4,
  99863.24, 99988.8, 100330.4, 100687.9, 101008.7, 101213.7, 101519.6, 
    101702.6, 101882.9, 102028.9, 102141.1, 102231.2, 102295.2, 102344.8, 
    102364.8,
  99959.05, 100005.4, 100276.8, 100597.5, 100952.8, 101146.6, 101416.6, 
    101642.1, 101805.8, 101963.6, 102068.2, 102158.9, 102221.4, 102266, 
    102281.5,
  100129.5, 100068.6, 100235.1, 100534.2, 100886.4, 101105.2, 101328.2, 
    101578.4, 101737.6, 101896.8, 102001.3, 102083.4, 102141.2, 102178.9, 
    102190.2,
  101815.4, 101961.4, 102074.8, 102186.1, 102274.6, 102354.9, 102414.1, 
    102460.9, 102502.9, 102539.8, 102568.1, 102591.6, 102613.4, 102636.9, 
    102663.2,
  101641.8, 101798.3, 101925.5, 102052.1, 102155.1, 102248.6, 102320.6, 
    102374.5, 102422.3, 102456, 102482.7, 102501.6, 102521, 102541, 102563.9,
  101423.7, 101605.4, 101752.9, 101905.5, 102024.6, 102134.1, 102218.7, 
    102282.4, 102330.7, 102368, 102396.9, 102413.3, 102424.1, 102434.3, 
    102449.2,
  101188.2, 101385.7, 101558.3, 101734.7, 101873.3, 102000, 102097.9, 102177, 
    102233.8, 102275.6, 102300.8, 102316.5, 102325.2, 102331.5, 102338.4,
  100920, 101140.4, 101342.3, 101541.5, 101707.6, 101856, 101971.6, 102064.5, 
    102130, 102178.2, 102207.6, 102221, 102223.9, 102221.2, 102218.6,
  100624.5, 100871, 101097.6, 101324.2, 101521.8, 101693.8, 101828.6, 
    101939.8, 102016.8, 102068.9, 102102, 102114.1, 102114.7, 102105.7, 
    102094.6,
  100308.1, 100573.5, 100830.1, 101087.8, 101315.4, 101517.5, 101679.1, 
    101805.6, 101900, 101959.9, 101994.3, 102005.3, 102000.4, 101982.5, 
    101961.2,
  99979.47, 100253.8, 100531.9, 100820.8, 101088.8, 101324.6, 101519.5, 
    101667.6, 101775.8, 101847.3, 101883.4, 101893.6, 101883, 101859.3, 
    101825.5,
  99655.27, 99904.09, 100223.6, 100519.5, 100839.9, 101116.9, 101349.2, 
    101528.5, 101653.2, 101735.9, 101776.4, 101785, 101765.3, 101729.7, 
    101686.4,
  99394.16, 99555.98, 99878.79, 100190.7, 100559.8, 100891.8, 101168.9, 
    101386.9, 101532.1, 101625.9, 101672.1, 101673.9, 101649.4, 101603.8, 
    101548.9,
  101492.1, 101566.1, 101641, 101715, 101789.8, 101864.1, 101936.8, 102008.6, 
    102081.8, 102152.5, 102222.8, 102291.6, 102357.4, 102422.1, 102483.8,
  101324.1, 101399.8, 101476.5, 101553.4, 101632, 101709.8, 101786.8, 
    101861.5, 101935.2, 102008.8, 102080, 102150.5, 102219.9, 102285.5, 
    102350.1,
  101132.2, 101222.9, 101304.7, 101389.3, 101470.7, 101552.5, 101632.5, 
    101709.4, 101786.1, 101862.1, 101933.7, 102004.2, 102072.6, 102140.4, 
    102206.3,
  100935.4, 101032.2, 101117.7, 101208.6, 101294.7, 101383.9, 101467.8, 
    101551.4, 101631.6, 101709.1, 101784.8, 101855.8, 101925.2, 101990.5, 
    102056.6,
  100719.2, 100829.3, 100919, 101021.3, 101111.2, 101205.2, 101294.1, 
    101383.3, 101469.2, 101551.1, 101628.1, 101702.4, 101772.8, 101840, 
    101903.5,
  100482.2, 100609.1, 100706.1, 100819, 100917, 101018.4, 101109.1, 101204.6, 
    101293.5, 101384, 101465.1, 101543.8, 101616.7, 101684.7, 101751.4,
  100227.3, 100365.6, 100476, 100603.6, 100710.8, 100823.7, 100922.6, 101020, 
    101114.9, 101206.4, 101293.7, 101375.2, 101453.1, 101523.4, 101589.8,
  99966.45, 100110.1, 100231.7, 100374.2, 100493.6, 100617.5, 100721.1, 
    100826.9, 100924.4, 101023.1, 101113.8, 101198.8, 101278.3, 101356.2, 
    101425.2,
  99679.52, 99843.1, 99979.55, 100135.2, 100270.9, 100402.2, 100522.7, 
    100632.4, 100735.5, 100835.5, 100930.1, 101020.7, 101102.9, 101180.1, 
    101251.6,
  99375.62, 99557.61, 99717.7, 99888.7, 100042.5, 100191.2, 100319, 100437, 
    100541.3, 100644.3, 100739.9, 100831.4, 100918.4, 100995.9, 101070.6,
  101626.7, 101656.4, 101687.3, 101712.6, 101739.5, 101765.3, 101793.9, 
    101822.9, 101857, 101894.3, 101933.4, 101974, 102016.1, 102058.9, 102104.5,
  101522.5, 101550.7, 101580, 101604.8, 101631, 101653.6, 101678.1, 101702.9, 
    101733, 101766.8, 101803.6, 101843.1, 101884.4, 101927.6, 101974,
  101402.6, 101433.5, 101463.8, 101491, 101519, 101543, 101563.2, 101586.2, 
    101609.2, 101636.8, 101668.6, 101704.4, 101745.4, 101786.9, 101832.3,
  101286.4, 101312, 101339, 101365.5, 101390.8, 101417.8, 101439.7, 101459.5, 
    101480.9, 101504.6, 101531.1, 101561.9, 101596.9, 101635.9, 101678.6,
  101158.2, 101184.8, 101208.8, 101235.2, 101258.9, 101284, 101304.4, 
    101325.4, 101344, 101366.8, 101388.2, 101414, 101442.8, 101477.5, 101515.7,
  101023.6, 101054.4, 101077, 101101, 101121.7, 101143.3, 101161.9, 101181.1, 
    101199.6, 101218.4, 101235.5, 101254.9, 101277.3, 101305.7, 101338.9,
  100881.4, 100916.7, 100938.7, 100964.3, 100982, 101002.8, 101015.8, 
    101032.6, 101046.5, 101062.4, 101073.6, 101086.7, 101102.4, 101123.5, 
    101150.6,
  100737, 100775.8, 100798.2, 100824.4, 100838.8, 100859.3, 100869.1, 
    100879.7, 100889.7, 100897.7, 100903.9, 100909.3, 100917.2, 100931.9, 
    100952.3,
  100585.8, 100625.4, 100652.2, 100681.7, 100696.9, 100712.7, 100722.2, 
    100727.1, 100728.7, 100729.7, 100727.3, 100724.3, 100723.2, 100729.4, 
    100740.3,
  100424.1, 100473.2, 100504.8, 100533.7, 100551.1, 100564.9, 100570.5, 
    100571.1, 100566.4, 100561.5, 100551.2, 100540.3, 100529.9, 100525.2, 
    100527.7,
  101310.6, 101319.6, 101330.6, 101345.5, 101367, 101397.1, 101430, 101472.7, 
    101518, 101570, 101623.3, 101682.6, 101743.9, 101810.4, 101872.5,
  101225.1, 101223.2, 101230.6, 101245.3, 101270.2, 101299.7, 101336.1, 
    101372.9, 101418.1, 101468.2, 101524.1, 101583.4, 101645.1, 101709.4, 
    101775.8,
  101119.1, 101118.4, 101122.7, 101131.6, 101150, 101171.7, 101200.2, 
    101236.2, 101280.3, 101329.9, 101382.1, 101439.7, 101500, 101565.2, 
    101632.9,
  101020.1, 101014.8, 101012.7, 101017.5, 101032.4, 101050.5, 101076.9, 
    101107.9, 101147.1, 101191.7, 101241.6, 101294.6, 101352.9, 101416.5, 
    101484,
  100920.5, 100906.5, 100901.1, 100899, 100903.7, 100913.4, 100930.6, 
    100955.3, 100988, 101026.8, 101070.8, 101119.9, 101172.6, 101232.9, 
    101299.1,
  100819, 100798.7, 100783.2, 100773.2, 100769.9, 100773.1, 100783.5, 
    100800.4, 100826.4, 100857.9, 100894, 100937.2, 100984.6, 101039.7, 
    101100.9,
  100715.5, 100688.7, 100663.2, 100643.7, 100630.7, 100624.4, 100623.5, 
    100631.9, 100647.4, 100668.8, 100696.4, 100729.7, 100769.8, 100819.2, 
    100871,
  100608.8, 100574.9, 100536.5, 100510.2, 100486.9, 100469.9, 100460.2, 
    100456.8, 100461, 100474.1, 100491.1, 100514.9, 100543.8, 100580.2, 
    100622.9,
  100505.2, 100462.1, 100414.1, 100377.2, 100340.7, 100313.1, 100291.8, 
    100274.4, 100267.5, 100264.3, 100269.9, 100278.6, 100296.9, 100320.5, 
    100353.9,
  100403.1, 100350.2, 100292.9, 100244.3, 100196.9, 100156.3, 100120.5, 
    100089.5, 100066.4, 100050.7, 100043, 100038.4, 100041.5, 100050.4, 100073,
  101677.9, 101679.5, 101677.3, 101681.5, 101685.2, 101691.8, 101702, 
    101717.2, 101741.5, 101770, 101801.9, 101836.9, 101875.3, 101915.6, 
    101959.7,
  101638.3, 101626.8, 101622.6, 101608.9, 101602.7, 101602.3, 101611.6, 
    101623.3, 101643.8, 101668.9, 101699.1, 101731.2, 101767.1, 101804.2, 
    101845.5,
  101571.2, 101544.1, 101533.8, 101515.9, 101510.1, 101505.8, 101509.7, 
    101517.3, 101535, 101555, 101581.4, 101608.6, 101641.8, 101677.1, 101716.4,
  101499.9, 101466.9, 101447.4, 101418.9, 101405.6, 101396.2, 101395.1, 
    101397.5, 101408.2, 101424.1, 101444.5, 101468.8, 101498.5, 101531.1, 
    101567,
  101413.1, 101371.2, 101341, 101310.9, 101292.2, 101276, 101265.8, 101261.2, 
    101265.8, 101274.8, 101289.9, 101308.5, 101335.2, 101365, 101398.5,
  101319.5, 101271.1, 101231.2, 101195, 101164.8, 101140.3, 101120.8, 
    101107.4, 101103.6, 101104.8, 101114.3, 101128.7, 101148.7, 101176, 
    101208.9,
  101216.9, 101159.7, 101112, 101065, 101026.3, 100992.2, 100961.2, 100938.3, 
    100923.5, 100917.9, 100918.1, 100926.1, 100943.1, 100967.5, 100997.6,
  101106.6, 101043.8, 100986.2, 100928.4, 100879.1, 100832.8, 100790.2, 
    100756.2, 100731.8, 100717.7, 100710.4, 100713.9, 100725.2, 100745.4, 
    100772.2,
  100996.2, 100923.7, 100853.7, 100784.2, 100720.3, 100661, 100609.5, 
    100563.9, 100529.7, 100505.3, 100492.1, 100488, 100494.4, 100508.2, 
    100530.7,
  100882.1, 100798.8, 100716.5, 100636.8, 100558.5, 100487.9, 100423.2, 
    100367.2, 100321, 100288.3, 100266.7, 100255.6, 100255.4, 100263.8, 
    100280.8,
  101710.1, 101796.1, 101858.3, 101911.7, 101956, 102003.5, 102051.1, 
    102102.5, 102149.3, 102193.3, 102225.9, 102257.4, 102288.6, 102320.1, 
    102349.5,
  101708.5, 101774.6, 101829, 101880, 101924.3, 101970.8, 102014.7, 102061.8, 
    102105.3, 102147.8, 102179.3, 102210.9, 102236.2, 102264.4, 102290.1,
  101691.7, 101762.7, 101810.7, 101859.9, 101899, 101942.1, 101980, 102021.2, 
    102061.1, 102101.5, 102137.4, 102165, 102189.2, 102216.2, 102246.1,
  101692.8, 101747, 101781.6, 101828.4, 101865.7, 101904.7, 101938.5, 
    101975.4, 102014.3, 102051.3, 102087.5, 102115.4, 102138.7, 102161.4, 
    102192.5,
  101687.9, 101730, 101760.8, 101798.1, 101832, 101864.5, 101892.9, 101926.2, 
    101962.1, 101998.1, 102028.9, 102059.4, 102085.2, 102106.9, 102126.7,
  101685.9, 101710.7, 101734.3, 101761.4, 101789.2, 101815.3, 101838, 
    101869.2, 101902, 101938.5, 101971, 101999.5, 102026.3, 102056.2, 102078.6,
  101674.5, 101689.7, 101703.7, 101723.5, 101741.8, 101757.9, 101777.6, 
    101804.8, 101834.3, 101868.1, 101901.4, 101931.1, 101956.6, 101981, 
    102004.9,
  101658.5, 101665.1, 101665.4, 101675.4, 101684.5, 101693.5, 101707.6, 
    101729.2, 101756.9, 101789.3, 101819, 101847.2, 101874.9, 101902, 101924,
  101637.3, 101633.7, 101624.2, 101620.9, 101620.8, 101623, 101630.4, 
    101643.4, 101664, 101691.9, 101717.7, 101744.3, 101770.6, 101798.2, 
    101825.7,
  101607.8, 101591.2, 101572.6, 101557.8, 101544.1, 101536.8, 101538.5, 
    101545.1, 101559.1, 101579.7, 101603.4, 101627.3, 101651.4, 101676.1, 
    101700.4,
  101685.5, 101790, 101876.2, 101950.8, 102014.9, 102065.9, 102106.5, 
    102139.5, 102174.4, 102208.6, 102238.2, 102270.1, 102306, 102341.9, 
    102378.1,
  101641.1, 101753.5, 101846, 101926.7, 101994.6, 102044.1, 102080.8, 
    102107.9, 102135.7, 102168.2, 102191.8, 102220.1, 102250.6, 102285.6, 
    102319.8,
  101590.7, 101709.5, 101812.6, 101895.3, 101964, 102016, 102055.5, 102085.3, 
    102106, 102121.2, 102143.6, 102165.6, 102188.6, 102214.4, 102245.2,
  101542.2, 101665.6, 101778, 101862.1, 101932.2, 101981, 102018.6, 102043.6, 
    102062.2, 102076.7, 102091.2, 102103.5, 102117.8, 102137.9, 102161.1,
  101492.1, 101621.2, 101741.2, 101822.3, 101896.4, 101941.7, 101976.5, 
    101999.4, 102011, 102017.9, 102023.2, 102029.2, 102035.2, 102048.1, 
    102064.9,
  101442.8, 101582.3, 101707.2, 101792.7, 101861.1, 101906, 101938.3, 
    101952.4, 101956.2, 101955.7, 101954, 101952.4, 101950.2, 101954, 101959.7,
  101405.3, 101547.9, 101675.1, 101766.3, 101835.8, 101877.5, 101901.7, 
    101908, 101905.7, 101894.6, 101882.5, 101870.3, 101858.5, 101850.4, 
    101847.5,
  101369.1, 101510.8, 101647.2, 101740.3, 101808.9, 101846.1, 101866, 
    101866.3, 101852.6, 101831.6, 101807.3, 101780.8, 101756.8, 101737.6, 
    101722.8,
  101339.4, 101483.5, 101623, 101712.4, 101778.7, 101810.7, 101825.6, 
    101822.4, 101799.1, 101766.7, 101728.5, 101689.5, 101650.7, 101617.2, 
    101588.7,
  101310.9, 101465, 101597.6, 101689.4, 101753.7, 101778.3, 101784.5, 
    101773.8, 101740.4, 101696.7, 101644.4, 101589.3, 101535.3, 101485.9, 
    101442.4,
  101798.7, 101831.1, 101859.6, 101889.5, 101923.6, 101958.6, 101995.2, 
    102032.5, 102071.6, 102113.8, 102155.5, 102198.1, 102240.8, 102282.5, 
    102326.1,
  101734.5, 101764.5, 101789.3, 101817.9, 101849.7, 101884.4, 101921.2, 
    101958.3, 101999.7, 102043.2, 102087.1, 102130.8, 102173.7, 102218.4, 
    102263.4,
  101651.1, 101678.9, 101705.3, 101734, 101764.2, 101798.5, 101837, 101875.9, 
    101918.9, 101961.5, 102007, 102051.6, 102099.6, 102145.4, 102191.7,
  101563.4, 101590.3, 101614.5, 101640.4, 101669.1, 101702.7, 101739.6, 
    101780.1, 101825, 101871.6, 101918.4, 101965.4, 102013.6, 102063.9, 
    102112.8,
  101472.3, 101491.2, 101514.7, 101537.3, 101564.6, 101597.6, 101635, 
    101675.1, 101719.8, 101767.2, 101816.7, 101867.3, 101916.9, 101966.7, 
    102016.6,
  101373.7, 101388.3, 101409.2, 101427.9, 101453.6, 101485.1, 101521.1, 
    101562.5, 101607.5, 101655.1, 101705.2, 101756.1, 101807.8, 101859.8, 
    101912.1,
  101265.7, 101277.2, 101295.5, 101311.9, 101336.8, 101368, 101403.8, 
    101441.6, 101487.1, 101534.7, 101584.8, 101634.8, 101686.3, 101739.5, 
    101792.3,
  101150.5, 101161.2, 101177.6, 101191.5, 101212, 101241.1, 101274.5, 
    101312.8, 101356.4, 101402.3, 101451.3, 101501, 101553.2, 101608.4, 
    101664.6,
  101030, 101043.7, 101057, 101067.7, 101083.4, 101105.3, 101135.3, 101170.8, 
    101212.3, 101255.6, 101302, 101350.4, 101402.3, 101456.9, 101513.4,
  100905.6, 100917.8, 100933.1, 100939.3, 100948.7, 100965.2, 100990.8, 
    101020.2, 101057.3, 101097, 101139.6, 101185.8, 101236.9, 101291.5, 101350,
  102488.9, 102505.7, 102508.8, 102520, 102523, 102527.3, 102536.4, 102535.5, 
    102538, 102539, 102543.6, 102550.2, 102559.8, 102563.4, 102571.5,
  102473.8, 102487.9, 102492.4, 102496.3, 102507.5, 102511.2, 102519.8, 
    102522.1, 102523.8, 102522.3, 102527, 102537.5, 102540.5, 102542.3, 102545,
  102465.3, 102477.3, 102488.4, 102493.9, 102495.1, 102509.2, 102513.1, 
    102515.2, 102515.6, 102514.2, 102511.8, 102508.9, 102509.3, 102508.4, 
    102508.7,
  102469.5, 102465.1, 102480.5, 102485.4, 102500.7, 102505.2, 102508, 
    102509.1, 102505.4, 102505.7, 102499.5, 102490.9, 102481.7, 102475.3, 
    102467.1,
  102446.5, 102448.8, 102471.2, 102480, 102486, 102492.4, 102492.9, 102492.9, 
    102489.7, 102482.8, 102474.9, 102462.6, 102446.8, 102430.4, 102414.8,
  102411.2, 102434.9, 102442.5, 102450.5, 102456.4, 102460.7, 102459.9, 
    102458.2, 102454.3, 102449, 102437.8, 102420.8, 102400.2, 102377.7, 
    102353.1,
  102374.9, 102398.8, 102401.8, 102411.4, 102415.8, 102415.8, 102412, 
    102406.8, 102400.3, 102392.2, 102376.4, 102357.5, 102333.4, 102308.8, 
    102278.9,
  102337.8, 102351.2, 102357.9, 102361.8, 102363.1, 102361.2, 102356.7, 
    102347.3, 102336.7, 102323.5, 102305.2, 102280.6, 102251.4, 102219.5, 
    102184.9,
  102288.5, 102296.4, 102301.3, 102300.6, 102300.2, 102295.2, 102287, 
    102275.2, 102260.4, 102242.2, 102218.5, 102187.7, 102155.4, 102116.4, 
    102078.6,
  102225.5, 102233.1, 102236.3, 102233.3, 102227.8, 102218.9, 102208.7, 
    102194.8, 102175.1, 102152.9, 102123.2, 102087.1, 102046.1, 102002.2, 
    101953.8,
  102933.5, 102950, 102927.3, 102916.8, 102895, 102880.9, 102866.5, 102852.3, 
    102835.7, 102828.9, 102816.6, 102806.1, 102800.6, 102781.5, 102776.9,
  102991.9, 102985.3, 102960, 102943.4, 102921.4, 102903.5, 102884.5, 
    102864.3, 102841.1, 102827.9, 102815.2, 102805.2, 102790.4, 102780.3, 
    102776.1,
  103005.3, 102985.9, 102970.2, 102948.9, 102927, 102905.7, 102889, 102860.7, 
    102840, 102822.5, 102807, 102789, 102772.8, 102759.7, 102751.1,
  103038.8, 103004.9, 102982.1, 102950.8, 102929.1, 102903.7, 102879.9, 
    102845.9, 102818.8, 102798.3, 102777.1, 102757.7, 102740.7, 102726.8, 
    102716.8,
  103074.6, 103025.6, 103000.7, 102961.9, 102930.4, 102902.2, 102871.1, 
    102828.1, 102794.3, 102768, 102743, 102721, 102700.9, 102679.3, 102662,
  103094.6, 103049.9, 103017.2, 102969.8, 102931.9, 102896, 102852, 102803.2, 
    102761.8, 102728, 102696.6, 102670.1, 102640.6, 102614.6, 102587.9,
  103102.6, 103073.3, 103020.2, 102972, 102922.1, 102877.6, 102825.5, 
    102769.2, 102721.5, 102680.1, 102640.5, 102604.5, 102567.7, 102533.2, 
    102495.7,
  103103.9, 103075.9, 103012.2, 102961, 102902, 102853.2, 102786.2, 102723.9, 
    102671.1, 102619.1, 102570.4, 102526.6, 102478.8, 102432.6, 102392.9,
  103099.2, 103057.7, 102994.2, 102939.3, 102871.9, 102809.3, 102737.3, 
    102670.4, 102607.6, 102545.5, 102488.4, 102430.9, 102372.6, 102324.1, 
    102281.5,
  103087.2, 103029.8, 102971.7, 102905.1, 102829.6, 102755.6, 102679.5, 
    102604.7, 102532.4, 102458.3, 102389.6, 102321.2, 102258.2, 102202.2, 
    102149.7,
  102733.6, 102708.2, 102670.4, 102633.1, 102598.7, 102564.8, 102531.2, 
    102499.6, 102470.8, 102455, 102450, 102447.6, 102450.7, 102451.1, 102454.8,
  102868.1, 102840.1, 102811.7, 102780.8, 102746.8, 102718.5, 102687.6, 
    102656.6, 102625.5, 102603, 102584.5, 102569.8, 102563, 102557.6, 102553.6,
  102955.1, 102932.5, 102911.2, 102882.3, 102857.5, 102826.9, 102797.9, 
    102767.3, 102741.9, 102715.7, 102694.9, 102675.5, 102660, 102649, 102637.9,
  103027.8, 103005.6, 102993.9, 102970, 102940.3, 102910.7, 102882.2, 
    102852.6, 102826.9, 102800.8, 102776.7, 102757.8, 102741.3, 102725, 
    102710.1,
  103079.7, 103052.5, 103039.2, 103013.4, 102996.2, 102972.3, 102942.4, 
    102913.6, 102886.3, 102862.3, 102838.7, 102821.1, 102796.9, 102775.2, 
    102753.5,
  103119.5, 103092.6, 103074.7, 103049.2, 103029.4, 103002.3, 102979.7, 
    102946.8, 102923.4, 102900.1, 102878.6, 102853, 102828.8, 102799.3, 
    102765.6,
  103161.6, 103120.5, 103097.8, 103066.7, 103057.5, 103029.5, 103001, 
    102972.4, 102945.3, 102920.2, 102894.9, 102866.2, 102832.4, 102798.1, 
    102769.8,
  103195.5, 103147.1, 103115.7, 103083.3, 103069.7, 103040.5, 103012.6, 
    102982.7, 102956.3, 102926.4, 102893.1, 102857.3, 102819.7, 102795.7, 
    102770.5,
  103228.6, 103178.7, 103137.5, 103100.6, 103078.5, 103046.2, 103016.1, 
    102986.1, 102951, 102913.3, 102870.9, 102835.1, 102810.3, 102779.7, 
    102739.1,
  103257.3, 103196.5, 103151.3, 103110.5, 103083, 103043, 103013.9, 102973.7, 
    102930.5, 102884.2, 102843.1, 102814.7, 102778.1, 102731.4, 102682.2,
  101106.3, 101071.6, 101062.6, 101096.1, 101151.7, 101219.8, 101296.7, 
    101370.5, 101440.2, 101516, 101573.9, 101611.3, 101618.6, 101614.1, 
    101588.5,
  101335.6, 101311.9, 101322.4, 101362.6, 101412.9, 101476.9, 101529.6, 
    101574.7, 101610.2, 101653.3, 101689.5, 101717.5, 101725.1, 101720.8, 
    101696.2,
  101605.3, 101573.5, 101573.3, 101591.5, 101630.4, 101678.4, 101714.2, 
    101738.1, 101759.9, 101799.3, 101828.4, 101853.3, 101853.4, 101835.5, 
    101804.6,
  101855.1, 101812.2, 101807.1, 101821, 101859.6, 101891.2, 101907.2, 
    101909.7, 101922.9, 101943.5, 101957.8, 101970.8, 101976.5, 101962.5, 
    101924.7,
  102087.3, 102049.5, 102038.4, 102042.2, 102046.5, 102057.2, 102057.6, 
    102061.2, 102071, 102080.1, 102087.4, 102093.4, 102084.8, 102061.6, 
    102023.8,
  102289.4, 102255, 102236, 102221.2, 102218.4, 102218.5, 102212.6, 102213.4, 
    102211.3, 102209.6, 102210.4, 102209, 102195.9, 102165.5, 102120.2,
  102475.1, 102435.2, 102404.7, 102382, 102361.1, 102349.4, 102338.7, 
    102340.8, 102331.3, 102325, 102316.4, 102307.5, 102288.8, 102257.4, 
    102215.1,
  102626.8, 102576.3, 102542.5, 102512, 102486.2, 102471.5, 102460.6, 102455, 
    102442, 102430.2, 102416.2, 102399, 102374.9, 102336.4, 102288.8,
  102768.1, 102714.7, 102676.8, 102637.4, 102610.5, 102585.5, 102567.1, 
    102553.1, 102536.9, 102522, 102501, 102475.5, 102444.2, 102395.4, 102342.2,
  102899.7, 102836.2, 102800, 102752.4, 102723.9, 102688.7, 102678.1, 
    102659.5, 102636.1, 102609.2, 102578.8, 102543.2, 102502.7, 102452, 102385,
  100132, 100096.2, 100085.6, 100076.5, 100081.5, 100114.1, 100175.7, 
    100295.5, 100433.4, 100561.2, 100663.8, 100730.5, 100747.1, 100732.6, 
    100679.2,
  100159.2, 100138.9, 100123.4, 100100.4, 100112.1, 100141.8, 100202.5, 
    100307.5, 100446.2, 100577.6, 100677.6, 100741, 100758.5, 100738.4, 
    100683.6,
  100216.7, 100193.7, 100187.5, 100183.1, 100202.6, 100219.3, 100258, 
    100330.1, 100439.9, 100565.9, 100669.5, 100742.8, 100770.3, 100753.9, 
    100696,
  100317.8, 100296, 100280.8, 100281.2, 100291.9, 100312.5, 100346.2, 
    100394.2, 100480.9, 100596.6, 100695.9, 100767.2, 100793.7, 100777.8, 
    100716.3,
  100434, 100440.8, 100418.2, 100415.6, 100418.8, 100439.2, 100453.8, 
    100479.8, 100544.5, 100632.2, 100718.4, 100786.2, 100818.5, 100805.3, 
    100742.4,
  100560.2, 100590.8, 100582.7, 100585.4, 100583.4, 100593.2, 100588.8, 
    100606.2, 100647.6, 100696.8, 100766.4, 100822.8, 100857, 100837.6, 
    100777.8,
  100709.1, 100748.8, 100753.2, 100765.2, 100765.3, 100767.8, 100753.5, 
    100759.2, 100774.5, 100786, 100827, 100866.3, 100896.7, 100878.4, 100817.1,
  100880.2, 100915.7, 100927.3, 100945, 100946.6, 100938.9, 100932.1, 
    100927.3, 100931.3, 100912.6, 100919.4, 100929.4, 100947.9, 100926.2, 
    100863.2,
  101074.1, 101102.5, 101115.1, 101127.3, 101124.7, 101119.3, 101112.6, 
    101102.8, 101092.9, 101059.9, 101039.8, 101016, 101009.7, 100980.4, 100911,
  101266.3, 101297.3, 101304.6, 101313, 101311.3, 101307.1, 101298.2, 
    101278.4, 101257.3, 101216.3, 101179.2, 101128.9, 101097.3, 101046.6, 
    100967.6,
  100592.2, 100591.3, 100583.5, 100556.5, 100526.2, 100478.3, 100404, 
    100316.1, 100217.5, 100095.8, 99962.78, 99808.34, 99636.59, 99468.3, 
    99291.76,
  100558.8, 100552.9, 100542.2, 100522.5, 100496.6, 100457.7, 100400.1, 
    100323.4, 100234.6, 100125, 99995.85, 99846.24, 99673.19, 99510.16, 
    99339.88,
  100507.7, 100499, 100486.5, 100475.4, 100452, 100421, 100383, 100321.3, 
    100243.2, 100142.3, 100020.7, 99872.86, 99707.47, 99549.3, 99382.26,
  100463.6, 100453.8, 100440.1, 100429.8, 100411.2, 100383.8, 100352.1, 
    100302.9, 100238.5, 100142.1, 100030.5, 99884.19, 99722.75, 99566.41, 
    99407.8,
  100415.8, 100400.7, 100385.3, 100371.8, 100356.9, 100336, 100308.1, 
    100268.7, 100215.1, 100130.2, 100026.3, 99884.98, 99731.58, 99587.13, 
    99447.04,
  100376.1, 100353.4, 100331.6, 100317.2, 100307.5, 100289.6, 100262.7, 
    100224.7, 100178, 100102.6, 100008.8, 99875.59, 99735.81, 99608.1, 
    99478.55,
  100341.3, 100308.1, 100279.1, 100260.2, 100246, 100230.8, 100208.2, 
    100172.8, 100124.5, 100058.2, 99975.54, 99861.86, 99744.39, 99627.52, 
    99516.31,
  100297.8, 100257.9, 100228.6, 100206, 100191.3, 100178.7, 100160.1, 
    100126.5, 100079.4, 100012.7, 99938.09, 99845.39, 99746.28, 99649.18, 
    99546.15,
  100248.7, 100201.3, 100168.6, 100147.2, 100137.1, 100128.9, 100112.8, 
    100085.4, 100037.3, 99972.95, 99900.17, 99823.53, 99739.39, 99660.62, 
    99570.03,
  100187.7, 100143.6, 100101.5, 100075.5, 100069.5, 100071.6, 100068.6, 
    100048.9, 100003.8, 99942.14, 99866.73, 99793.89, 99723.86, 99659.87, 
    99585.99,
  100950.9, 100823, 100656.4, 100458.5, 100277.5, 100078.2, 99905.04, 
    99725.46, 99521.93, 99314.84, 99118.82, 98916.83, 98718.38, 98514.14, 
    98315.45,
  100987.9, 100857.5, 100679.9, 100479.4, 100287.9, 100089.2, 99890.71, 
    99680.53, 99470.78, 99260.32, 99052.27, 98845.99, 98638.11, 98430.52, 
    98225.54,
  101005.5, 100878.9, 100716.4, 100529.8, 100332.6, 100132.9, 99930.12, 
    99716.42, 99498.92, 99276.7, 99054.23, 98829.77, 98605.59, 98382.62, 
    98161.98,
  101022.3, 100894.9, 100733.6, 100552.3, 100352.6, 100151.5, 99945.67, 
    99717.75, 99479.85, 99234.87, 98995.81, 98762.55, 98531.67, 98300.69, 
    98073.73,
  101041, 100911.3, 100752.6, 100578.2, 100382.8, 100179.1, 99969.95, 
    99739.28, 99498.05, 99238.31, 98985.23, 98733.87, 98494.88, 98256.11, 
    98019.25,
  101055.7, 100925.3, 100764.4, 100592, 100396.1, 100190.5, 99980.66, 
    99744.78, 99495.2, 99225.8, 98959.38, 98698.61, 98453.73, 98208.95, 
    97959.61,
  101066.8, 100938.1, 100778.4, 100608.9, 100412.6, 100206.7, 99995.45, 
    99756.86, 99504.85, 99233.8, 98960.3, 98689.7, 98432.09, 98174.56, 97912.7,
  101076.7, 100948.3, 100793.3, 100624.7, 100429.6, 100224, 100005.8, 
    99764.74, 99507.55, 99230.09, 98955.06, 98679.41, 98410.38, 98142.69, 
    97870.67,
  101090.9, 100960.1, 100808.6, 100644.1, 100453, 100247, 100024.9, 99780.98, 
    99521.01, 99243.35, 98966.77, 98685.13, 98405.59, 98123.98, 97842.11,
  101104.1, 100971.4, 100823.8, 100659.4, 100475.7, 100270.9, 100048.7, 
    99804.3, 99544.79, 99266.99, 98989.28, 98703.8, 98412.12, 98121.62, 
    97825.68,
  101403.8, 101306.8, 101211.8, 101122.4, 101044.3, 100986, 100932, 100877, 
    100810.2, 100759.9, 100712.2, 100673.4, 100635.4, 100599.6, 100566.5,
  101413.3, 101312.5, 101216.2, 101117.2, 101040.5, 100962.7, 100888.4, 
    100817.3, 100741.4, 100682, 100624.7, 100579.8, 100533.4, 100493.4, 
    100455.5,
  101404.4, 101313.4, 101215.7, 101102.9, 101010.8, 100910.7, 100827.1, 
    100753.4, 100675.5, 100613.8, 100547.2, 100497.8, 100440.4, 100392.1, 
    100345.6,
  101374.5, 101280.5, 101174.6, 101047.7, 100952.3, 100851.9, 100767.8, 
    100683.8, 100595.6, 100521.1, 100451.7, 100392.4, 100330.5, 100277.3, 
    100223.9,
  101352.4, 101256.2, 101140.2, 101011.5, 100906.1, 100805.2, 100707.4, 
    100615.7, 100522.8, 100439.2, 100365.4, 100296.6, 100226.8, 100162.9, 
    100101.7,
  101330.3, 101228.1, 101110.4, 100966.8, 100852.8, 100742.3, 100636.1, 
    100539.4, 100440.1, 100348.8, 100269.5, 100190.6, 100116.4, 100044.9, 
    99977.52,
  101305.5, 101200.4, 101074.6, 100930, 100804.9, 100688, 100571.8, 100468.7, 
    100361.8, 100262.9, 100173.2, 100086.5, 100003, 99923.92, 99849.5,
  101278.4, 101170, 101037.4, 100889.7, 100753.6, 100626.8, 100501.8, 100390, 
    100275.8, 100168.9, 100070.8, 99975.88, 99884.57, 99801.73, 99726.48,
  101249.4, 101138, 101003.5, 100849.2, 100704.9, 100571.3, 100436.4, 
    100312.3, 100191.9, 100076.6, 99969.73, 99866.46, 99768.78, 99678.38, 
    99599.98,
  101220.1, 101100.7, 100962.9, 100806.8, 100656.8, 100515.8, 100372, 
    100235.6, 100106.1, 99980.77, 99865.57, 99753.07, 99646.78, 99550.71, 
    99473.12,
  102028.9, 102041.1, 102021.1, 102010.7, 101980.7, 101934.6, 101884.2, 
    101818.8, 101733.8, 101634.3, 101515.6, 101380.1, 101225.5, 101061.8, 
    100890.6,
  102034.2, 102042.7, 102021.5, 102010.2, 101973.8, 101934, 101884.2, 
    101819.4, 101733.9, 101633.4, 101513.5, 101376.1, 101221, 101052.3, 
    100871.6,
  102027.6, 102032.1, 102019, 102006.6, 101973.3, 101935.1, 101879.9, 
    101814.5, 101735.8, 101638.1, 101522.6, 101384.5, 101228.8, 101053.1, 
    100869.7,
  102019.3, 102025.6, 102014.5, 101999.7, 101969.6, 101932.1, 101879.3, 
    101814.8, 101736.6, 101640.3, 101527.9, 101390.8, 101233.9, 101053.4, 
    100862.4,
  102004, 102017.6, 102005.8, 101992.9, 101963, 101926.8, 101876.8, 101814.1, 
    101738.8, 101645.8, 101538.8, 101405.2, 101249.6, 101068.7, 100870.1,
  101994.1, 102007.4, 101993.4, 101985, 101955.9, 101922.2, 101877.1, 
    101815.1, 101738, 101650.1, 101546.9, 101416.2, 101262.6, 101083, 100881.1,
  101986.2, 101995.9, 101982.3, 101974.3, 101945.1, 101912.9, 101869, 101811, 
    101736.7, 101653.3, 101551.8, 101426.9, 101277.4, 101100.8, 100901.1,
  101979.9, 101986.3, 101971.6, 101960.7, 101932.7, 101901.6, 101856.3, 
    101806.6, 101734.8, 101653.1, 101554.9, 101436.1, 101288.6, 101115.7, 
    100917.8,
  101967.6, 101974, 101958.2, 101948.3, 101919.2, 101891.3, 101844.9, 
    101798.7, 101730.7, 101653.7, 101556, 101440.6, 101296.9, 101129.7, 
    100934.1,
  101954.5, 101957.1, 101938.7, 101930.6, 101902.2, 101874.2, 101830.4, 
    101786.9, 101721.1, 101647.3, 101550.8, 101439.1, 101300.1, 101138.3, 
    100946.6,
  101490.4, 101397.2, 101292, 101197.5, 101094.2, 100987.4, 100880.7, 
    100770.8, 100662.7, 100562.1, 100475.1, 100404.3, 100343.2, 100294.6, 
    100243.3,
  101480.9, 101370.2, 101256.5, 101153.1, 101042.4, 100927.3, 100807.7, 
    100686.6, 100565.8, 100450.4, 100350.2, 100262.5, 100188.6, 100117.9, 
    100052.4,
  101473.9, 101370.5, 101249.1, 101136.8, 101019.5, 100893.8, 100761.9, 
    100628.2, 100493.2, 100359.3, 100240.4, 100137.4, 100044.1, 99957.58, 
    99872.75,
  101465.9, 101351.2, 101224.2, 101099.5, 100976.9, 100843.4, 100703.4, 
    100563, 100416.2, 100274.3, 100139.3, 100016, 99904.02, 99802.73, 99703.93,
  101468.9, 101354.5, 101216.7, 101089.3, 100954.4, 100815.7, 100672.4, 
    100519.9, 100362.7, 100207.7, 100058, 99917.78, 99784.8, 99665.08, 
    99549.02,
  101477.9, 101356.6, 101213.5, 101080.4, 100940.4, 100795.5, 100645.4, 
    100485.3, 100321.3, 100157, 99993.02, 99837.25, 99685.22, 99546.43, 
    99411.42,
  101495, 101364.6, 101227.3, 101083.3, 100937, 100786.2, 100632.1, 100463.4, 
    100296.1, 100119.6, 99948.63, 99775.79, 99606.55, 99446.58, 99292.38,
  101519.3, 101380.5, 101244.2, 101095.8, 100946, 100787.5, 100628.1, 100455, 
    100279.8, 100095.8, 99918.33, 99732.3, 99552.05, 99370.05, 99200.46,
  101551.1, 101408.6, 101272.3, 101117.6, 100962.4, 100798.4, 100637.3, 
    100458.3, 100280.2, 100087.7, 99903.16, 99708.16, 99516.29, 99317.98, 
    99129.93,
  101582, 101446.6, 101303.3, 101156.9, 100994.1, 100823.6, 100655.2, 
    100473.2, 100293.9, 100095.6, 99900.35, 99701.35, 99496.7, 99290.28, 
    99082.87,
  101502.5, 101455.4, 101405.5, 101364, 101324.8, 101296.9, 101276.3, 101266, 
    101270.7, 101288.9, 101319.6, 101359, 101404.8, 101457.8, 101515.6,
  101416.9, 101350.2, 101288.9, 101232.9, 101180.6, 101137.7, 101103.9, 
    101081.2, 101076.1, 101087, 101112.1, 101148, 101192.6, 101244.1, 101304.5,
  101311.4, 101239.3, 101164.8, 101091.3, 101025.9, 100969.5, 100921.3, 
    100885.8, 100868.3, 100867.1, 100882.7, 100910.2, 100947.8, 100997.6, 
    101059.1,
  101213.9, 101132.4, 101044.2, 100956.1, 100873.9, 100802, 100736.5, 
    100686.5, 100652.9, 100639.2, 100642.7, 100660.6, 100689.4, 100733.7, 
    100791.8,
  101117.2, 101027.9, 100923.1, 100821.3, 100720.8, 100631.8, 100551.9, 
    100483.6, 100434, 100402.1, 100389.9, 100395.1, 100413.8, 100447.6, 
    100501.3,
  101028, 100929, 100808.3, 100695.9, 100576.3, 100472.1, 100369.9, 100282.8, 
    100215, 100162.4, 100133.8, 100121.6, 100128.8, 100154.6, 100200.6,
  100940.8, 100833.9, 100701, 100573.6, 100438.5, 100315.7, 100196.7, 
    100090.8, 99999.88, 99930.05, 99880.02, 99851.49, 99843.31, 99855.88, 
    99890.2,
  100865.4, 100749.1, 100601.6, 100463.3, 100312.7, 100172.6, 100033.9, 
    99911.77, 99799.62, 99709.62, 99638.41, 99592.84, 99568.45, 99568.34, 
    99592.16,
  100800, 100671.5, 100513.3, 100359.6, 100197, 100040.4, 99887.44, 99744.06, 
    99614.51, 99509.52, 99419.91, 99356.73, 99314.4, 99299.32, 99309.82,
  100747.1, 100606.6, 100439.5, 100271.9, 100100, 99922.28, 99758.75, 
    99598.98, 99453.8, 99328.98, 99226.69, 99145.62, 99084.04, 99053.84, 
    99049.22,
  102401.9, 102422.2, 102445.7, 102469.6, 102496.7, 102523.1, 102550.7, 
    102576.3, 102603.2, 102626.2, 102646.7, 102662.5, 102669.2, 102664.2, 
    102650.4,
  102302.2, 102311.8, 102332.7, 102351.4, 102376.8, 102401.4, 102429.1, 
    102456.2, 102484.7, 102513.7, 102539.3, 102559.5, 102574.1, 102578.1, 
    102573,
  102177, 102185.7, 102202.1, 102217.3, 102240.4, 102264.2, 102291.5, 102321, 
    102351.8, 102383.6, 102414, 102440.6, 102463.1, 102476.6, 102481.5,
  102052.1, 102056.8, 102065.5, 102075.7, 102093.7, 102115.4, 102142.2, 
    102171.6, 102206.1, 102242.7, 102278.7, 102311, 102338.9, 102361.5, 
    102374.6,
  101916.1, 101914.1, 101914.8, 101920.5, 101933.5, 101950.4, 101974, 
    102004.4, 102040.9, 102080.3, 102121.6, 102162.2, 102198.5, 102230.2, 
    102252.4,
  101776.3, 101769.5, 101760.3, 101758.5, 101764, 101776.8, 101796.3, 
    101825.2, 101862, 101906.5, 101953.5, 102000.9, 102044.3, 102083.6, 
    102114.9,
  101631.4, 101615.9, 101595, 101586.2, 101584.1, 101592.6, 101608.1, 
    101634.8, 101671.3, 101717.8, 101769.2, 101823.3, 101874.8, 101922.7, 
    101961.8,
  101488.4, 101462.3, 101430, 101412.7, 101400.7, 101405.6, 101413.6, 
    101436.1, 101470.9, 101518.3, 101572.8, 101631.6, 101689.7, 101746.7, 
    101795.2,
  101346, 101307.3, 101262.3, 101237.5, 101215.1, 101212, 101216.4, 101235.2, 
    101266.6, 101311.1, 101367.4, 101427.9, 101492.8, 101556.1, 101613.7,
  101202.4, 101152.8, 101096.2, 101060.6, 101030.6, 101020.8, 101022.2, 
    101037.6, 101062.6, 101105.1, 101157.5, 101221.6, 101288.6, 101357.3, 
    101422,
  103220.8, 103235.4, 103235.6, 103225.1, 103201.3, 103171.2, 103130.4, 
    103075.9, 103003.3, 102910.6, 102796.5, 102659, 102505.7, 102338.3, 
    102161.4,
  103184.5, 103198.2, 103203.2, 103197.8, 103179.1, 103147.9, 103107.9, 
    103052.4, 102977.1, 102885.9, 102775, 102640.8, 102483.7, 102309.7, 102128,
  103135.3, 103152.5, 103163.9, 103162.2, 103148.5, 103120.5, 103081.1, 
    103026, 102953.2, 102862.2, 102752.1, 102622.6, 102469.1, 102296, 102110.6,
  103076.8, 103099.6, 103115.7, 103119.2, 103111.6, 103087.1, 103050.6, 
    102999.9, 102930.5, 102839.3, 102728.5, 102600.3, 102447.5, 102274.4, 
    102084.9,
  103010.6, 103039, 103058.4, 103066.5, 103063.1, 103045.1, 103013.2, 
    102966.6, 102901.2, 102813.3, 102703.4, 102579.3, 102428, 102259.9, 
    102073.2,
  102930.3, 102967.9, 102992.4, 103006, 103007.5, 102997.3, 102969.6, 
    102925.9, 102863, 102777.8, 102671.9, 102550.2, 102402.7, 102236.1, 
    102052.8,
  102839.4, 102877.6, 102908.7, 102930.2, 102939.3, 102935.7, 102911.1, 
    102870.7, 102813.6, 102734.6, 102636.4, 102518.1, 102375.5, 102212.2, 
    102033.2,
  102739.4, 102780.2, 102814.3, 102839.3, 102854.2, 102857.8, 102842.3, 
    102809.9, 102757.5, 102685.5, 102593, 102477.8, 102339, 102181.9, 102007.7,
  102625.9, 102670, 102708.1, 102736.5, 102756.1, 102764.6, 102757.1, 
    102732.8, 102689.4, 102625.2, 102540.3, 102431, 102299.9, 102146.7, 
    101976.3,
  102502.6, 102550.6, 102592, 102624.5, 102648.9, 102663.7, 102664.5, 
    102648.4, 102613.2, 102557.1, 102480.8, 102377.4, 102254, 102107.8, 
    101942.1,
  103018, 102960, 102883.6, 102803.8, 102711.3, 102610.3, 102495.2, 102369, 
    102235.5, 102100.3, 101981.2, 101871.2, 101788.3, 101713, 101644.6,
  103012.6, 102940.8, 102857.2, 102769.4, 102668, 102557.6, 102431.9, 102295, 
    102146.5, 101997.2, 101866.6, 101758.8, 101667.1, 101577.5, 101498.2,
  102990.2, 102915.6, 102828.8, 102735.2, 102624.8, 102504.8, 102369.7, 
    102219.1, 102055.1, 101901.1, 101770.2, 101653.4, 101540.2, 101439.5, 
    101346.1,
  102964.5, 102889.6, 102799.2, 102699.6, 102580.7, 102451.5, 102304.8, 
    102142.4, 101970.3, 101807.1, 101670.5, 101529.4, 101402.2, 101287.1, 
    101179.2,
  102939.6, 102859.6, 102765.4, 102659.9, 102533.4, 102394.9, 102235.8, 
    102063.1, 101884, 101718.8, 101568.2, 101412.4, 101268.8, 101133.3, 
    101012.8,
  102914.6, 102831.1, 102731.8, 102618.9, 102488.2, 102341.5, 102172.8, 
    101991.4, 101802.6, 101632.4, 101461.8, 101288.3, 101128.6, 100977.8, 
    100841,
  102883.8, 102801.8, 102696.7, 102578.1, 102440.6, 102284.3, 102110.8, 
    101920, 101722.2, 101543.8, 101355.6, 101171.1, 100995.3, 100827.8, 100674,
  102853.2, 102767, 102661.2, 102537.3, 102392.2, 102229.4, 102047.6, 
    101851.1, 101650.7, 101459.9, 101260.3, 101064.4, 100869.4, 100687.7, 
    100514.2,
  102816.1, 102729.1, 102621.6, 102494.3, 102344.6, 102176.7, 101989.3, 
    101788.3, 101584, 101384.4, 101173, 100966.8, 100757.6, 100557.1, 100365.2,
  102775.6, 102689, 102578.7, 102449.6, 102297.5, 102126.6, 101934.7, 
    101729.1, 101522.7, 101312.6, 101095.9, 100879.4, 100658.2, 100439.4, 
    100230.6,
  102094, 102090.2, 102082, 102076.7, 102079.3, 102085, 102093.7, 102109.4, 
    102131.1, 102157, 102180.3, 102198.2, 102208.7, 102212.3, 102209.2,
  102016.3, 101998.3, 101980.1, 101969.8, 101966.8, 101970.6, 101982.5, 
    102000.6, 102027.7, 102061, 102091, 102120.6, 102144.2, 102160.2, 102167.2,
  101904.8, 101879.8, 101856.6, 101842.1, 101835.5, 101839, 101851, 101874, 
    101907.9, 101946.9, 101984.6, 102019.8, 102048.3, 102072.8, 102092.7,
  101798.2, 101761.7, 101733.7, 101707, 101693.6, 101688.2, 101696.2, 
    101719.5, 101754.4, 101798.5, 101840, 101881.2, 101920.6, 101955.9, 
    101986.2,
  101676.2, 101631.4, 101590.3, 101556.9, 101535.3, 101525.9, 101530.7, 
    101551.9, 101584.6, 101630, 101673, 101720.8, 101766.2, 101807.5, 101847.5,
  101555.6, 101498.9, 101446.7, 101401, 101367.6, 101346.5, 101339.3, 
    101352.3, 101381.2, 101428.7, 101470.5, 101525.1, 101576.2, 101627.6, 
    101678.1,
  101434.1, 101363.5, 101291.6, 101231.2, 101182.7, 101151.4, 101131.9, 
    101134, 101159.2, 101204.8, 101245, 101298.6, 101356.2, 101411.1, 101468.8,
  101319.8, 101229.9, 101143.6, 101064.4, 100994.6, 100947.7, 100914, 
    100900.3, 100917.1, 100953.4, 100991.9, 101044.7, 101105.7, 101168.4, 
    101232.7,
  101210.6, 101103, 100995.2, 100895.3, 100805.7, 100739, 100690.3, 100656.9, 
    100666.2, 100691.1, 100720.7, 100772.5, 100832.3, 100899.1, 100968.7,
  101106.1, 100981.6, 100853.4, 100734, 100619.6, 100530.2, 100457.7, 
    100410.7, 100404.5, 100415.3, 100434.6, 100478.3, 100535.1, 100606, 
    100678.9,
  102288.7, 102263.2, 102233, 102192.5, 102144, 102089.1, 102025.2, 101957.8, 
    101883.4, 101804, 101714.3, 101609.6, 101494.7, 101372.1, 101242.8,
  102239.8, 102217.4, 102194.7, 102155.4, 102113.1, 102063.9, 102008.8, 
    101945.7, 101873.8, 101795.3, 101704.2, 101602.7, 101485.6, 101358.4, 
    101221.4,
  102178.4, 102169.5, 102150.6, 102118, 102078.1, 102034.8, 101978.1, 
    101918.7, 101850.2, 101777.4, 101689.8, 101589.9, 101473.5, 101345.5, 
    101204.8,
  102099.9, 102105.5, 102098.7, 102076.3, 102042.6, 102000.5, 101948.4, 
    101894.7, 101827.9, 101752.1, 101663.7, 101562.2, 101447.1, 101319.6, 
    101180.3,
  102006.5, 102022.6, 102028.1, 102019, 101999.3, 101965.5, 101915.1, 
    101863.6, 101801.1, 101729.6, 101643, 101542.1, 101427.1, 101300.7, 101164,
  101893.7, 101920.2, 101935.4, 101941.5, 101935.4, 101913.4, 101877.2, 
    101829.4, 101770.1, 101701.2, 101621.9, 101525.3, 101415.9, 101292.1, 
    101155.4,
  101769.4, 101798.3, 101821.6, 101836.7, 101842.8, 101833, 101810.4, 
    101773.1, 101725.2, 101667.2, 101594.9, 101506.7, 101401.8, 101282.9, 
    101149.3,
  101624.4, 101657.8, 101690, 101710.9, 101730.3, 101734.4, 101727.1, 
    101701.7, 101663.8, 101611.9, 101546, 101464.6, 101367.3, 101255.3, 
    101127.2,
  101470.8, 101507.5, 101542.1, 101568.5, 101594, 101609.6, 101614.4, 
    101606.8, 101583, 101544.7, 101489.3, 101417.1, 101328.8, 101222.7, 
    101101.5,
  101303.1, 101342.1, 101380.6, 101413.6, 101445.8, 101470.2, 101488.1, 
    101491.2, 101481.6, 101457, 101416.5, 101357.5, 101279.6, 101185, 101072.5,
  101617.7, 101562.4, 101497.1, 101427.2, 101355, 101277.8, 101203.1, 
    101117.7, 101036.2, 100955.4, 100879.1, 100800.5, 100730.1, 100661.4, 
    100595.3,
  101545.8, 101480.9, 101414.8, 101345.5, 101279.4, 101211.1, 101136.7, 
    101052.6, 100972.9, 100890, 100808.1, 100729.2, 100658, 100590.6, 100528,
  101462.2, 101392.9, 101326.7, 101261.5, 101196.7, 101124.1, 101048.4, 
    100968.6, 100890.8, 100808.3, 100730.3, 100654.8, 100584.7, 100517.4, 
    100454.6,
  101382.2, 101306, 101232.3, 101159.7, 101092.8, 101023.9, 100951.7, 
    100872.2, 100790.7, 100707, 100630.4, 100558.1, 100490.6, 100424.9, 
    100357.9,
  101304.8, 101220.2, 101144.4, 101063.8, 100992.4, 100921.8, 100849, 
    100772.5, 100694.4, 100613.8, 100540.4, 100470.9, 100403.4, 100337.4, 
    100265.6,
  101223.1, 101135.2, 101056.3, 100967.1, 100886.4, 100807.8, 100732.6, 
    100657.4, 100579.6, 100503.6, 100431.9, 100364.6, 100297.9, 100228.7, 
    100159.6,
  101134, 101047.4, 100963.4, 100871.2, 100783.2, 100697.9, 100617, 100540.7, 
    100465.1, 100394.8, 100323.7, 100254.4, 100182.6, 100114, 100043.4,
  101039.9, 100955.5, 100866.6, 100774.1, 100683, 100591.1, 100502.4, 
    100417.5, 100342.8, 100272.8, 100201.7, 100126.5, 100050.2, 99975.41, 
    99909.73,
  100947.9, 100864, 100769.9, 100678.3, 100581.7, 100486.4, 100391.6, 100301, 
    100220, 100141.2, 100063.2, 99982.7, 99905.76, 99834.57, 99768.41,
  100855.7, 100772.4, 100677.2, 100582.3, 100483.5, 100383.4, 100283.7, 
    100187.8, 100096.8, 100006.4, 99922.81, 99841.59, 99768.93, 99699.79, 
    99634.98,
  101303.2, 101300.6, 101284.7, 101274.4, 101261.2, 101244.1, 101218.7, 
    101188.2, 101148.7, 101096.8, 101041.5, 100981.3, 100919.1, 100845.6, 
    100765.1,
  101263.5, 101260.3, 101242.4, 101239.4, 101228.6, 101207.1, 101178.1, 
    101138.4, 101090.7, 101042.9, 100989.1, 100926.4, 100861, 100786.7, 
    100711.9,
  101204.3, 101206.4, 101197.1, 101190.1, 101168.2, 101145.2, 101120.6, 
    101087.8, 101047.6, 101000.9, 100947.3, 100887.6, 100820.9, 100747.4, 
    100671.3,
  101160.7, 101160.4, 101148.8, 101134, 101119.3, 101100.9, 101073.8, 
    101036.6, 100995.4, 100950.3, 100898.3, 100839, 100771.8, 100701.4, 100626,
  101109.6, 101099.7, 101092.7, 101082.2, 101073, 101049.9, 101025.8, 
    100993.2, 100957.1, 100913.9, 100864.1, 100805.7, 100738.6, 100664.4, 
    100589,
  101041.8, 101034.9, 101033.3, 101024.1, 101015.5, 100996.3, 100974.1, 
    100943.5, 100911.3, 100869.6, 100818.8, 100763.7, 100693.5, 100621.3, 
    100547.1,
  100970.4, 100970.1, 100971.4, 100967.6, 100963, 100950.2, 100931.9, 
    100901.7, 100869.6, 100831.3, 100786.1, 100734, 100663.2, 100592.7, 
    100514.6,
  100886, 100887.8, 100891.2, 100892.6, 100894.5, 100891.1, 100879.5, 
    100857.3, 100829.5, 100793.6, 100751.5, 100696, 100630, 100556.1, 100478.9,
  100791.7, 100803.3, 100808.4, 100816.6, 100823.4, 100826.2, 100825.5, 
    100806.8, 100779.5, 100750.1, 100712.3, 100660.7, 100604.8, 100532.8, 
    100458.2,
  100685.5, 100700.1, 100714.4, 100729.1, 100744.5, 100756.1, 100763.2, 
    100763.1, 100753.5, 100732.5, 100697.8, 100653.7, 100605.4, 100549.2, 
    100491.8,
  101508.6, 101499.9, 101470.4, 101444.4, 101407.7, 101373.1, 101334.4, 
    101302.8, 101270.9, 101242.8, 101216.5, 101190.8, 101168.5, 101154, 
    101140.2,
  101455, 101438, 101403.1, 101367.6, 101325.4, 101289.4, 101241.6, 101200.1, 
    101164.5, 101135.4, 101107.9, 101082.1, 101057.5, 101034.5, 101018.8,
  101394.7, 101373.1, 101334.9, 101297.9, 101254.8, 101209.6, 101156.5, 
    101110.1, 101066.9, 101028.4, 100993.6, 100956.7, 100927.9, 100905, 
    100884.2,
  101339.6, 101315.2, 101276.8, 101235.9, 101187.8, 101137.3, 101081.4, 
    101025.3, 100981.3, 100938, 100897.6, 100861.2, 100828.1, 100796.8, 
    100772.9,
  101291.6, 101265.2, 101225.8, 101183.7, 101136.5, 101081.2, 101020.6, 
    100962.7, 100909.9, 100860.5, 100814.9, 100773.5, 100737.2, 100700.1, 
    100671.6,
  101243, 101213.4, 101169.9, 101131.7, 101084.1, 101032.4, 100973.8, 
    100911.7, 100851.6, 100794.4, 100743.7, 100702.2, 100664.7, 100633.8, 
    100608,
  101208.8, 101173.4, 101131, 101092.9, 101047.8, 100993.8, 100938.1, 
    100868.5, 100816.4, 100750.6, 100701.6, 100649.9, 100611.8, 100578.3, 
    100550.4,
  101181.3, 101147.2, 101105.2, 101061.8, 101015.8, 100968.6, 100912.6, 
    100851.8, 100788.7, 100727.6, 100668.9, 100614.6, 100581.3, 100545.9, 
    100523.3,
  101186.7, 101143.6, 101106, 101065.7, 101006.3, 100953.1, 100899.8, 
    100832.6, 100778.7, 100718.6, 100659.5, 100615.7, 100569.5, 100526.7, 
    100488.3,
  101205.8, 101179.1, 101140.7, 101086, 101033.8, 100960.7, 100906.4, 
    100832.5, 100779.2, 100716.9, 100658.7, 100606.1, 100553.2, 100509.8, 
    100457,
  101914.1, 101966.1, 102000.4, 102041, 102076.2, 102108.9, 102136.8, 
    102160.3, 102182.7, 102200.9, 102215.2, 102224, 102225.6, 102217.8, 
    102207.5,
  101822.6, 101871.5, 101903.1, 101946.6, 101982.3, 102016.2, 102046.9, 
    102075.2, 102102.6, 102125.2, 102143.6, 102154.5, 102160.7, 102164.9, 
    102166.6,
  101711.8, 101757.3, 101788.2, 101835.1, 101872.6, 101910.1, 101941.4, 
    101972.6, 102000.8, 102027.5, 102052.3, 102074.2, 102090.7, 102101.5, 
    102104.9,
  101598.7, 101643.9, 101679.3, 101725.8, 101761, 101800.1, 101833.2, 
    101863.5, 101895.4, 101925.9, 101954.5, 101978.5, 101999.2, 102014.4, 
    102027.4,
  101484.6, 101528.7, 101561.2, 101605.4, 101646, 101685.2, 101717.9, 
    101751.3, 101781.2, 101813.5, 101844.6, 101874.9, 101899.7, 101920.8, 
    101938.1,
  101380.3, 101418, 101447.1, 101490.2, 101528.9, 101568.9, 101600.1, 
    101632.7, 101666.3, 101701.7, 101734, 101763.5, 101788.4, 101811.4, 
    101832.8,
  101279.2, 101317.2, 101348.5, 101384.3, 101411.3, 101449.3, 101479.6, 
    101509.8, 101544.3, 101582.2, 101619.7, 101653.8, 101678.7, 101702.9, 
    101721.8,
  101202.6, 101236.7, 101256.8, 101294, 101317.8, 101349.9, 101378.3, 
    101404.8, 101429.6, 101466.4, 101501.7, 101533.4, 101559.4, 101585.5, 
    101605.8,
  101106.4, 101162.5, 101187.7, 101216.3, 101235.8, 101268.6, 101286.1, 
    101311.4, 101328.6, 101355.1, 101385.4, 101417.5, 101442.9, 101463.9, 
    101480.8,
  101054, 101111.3, 101138.2, 101150, 101151.1, 101186, 101211.2, 101233.1, 
    101245.4, 101262.1, 101279, 101299, 101313.8, 101335.7, 101345.2,
  102470, 102520, 102551.8, 102573.2, 102587.6, 102586.7, 102574.7, 102542.7, 
    102492.5, 102419.5, 102324, 102203.3, 102068.6, 101924.7, 101768.5,
  102436.1, 102482.6, 102527.2, 102558.1, 102590.5, 102608.3, 102617.3, 
    102608.1, 102584.4, 102547.4, 102495.5, 102420, 102318.7, 102201.1, 
    102068.4,
  102375.3, 102435.9, 102488.4, 102535, 102582, 102613.7, 102642.8, 102656.4, 
    102656.5, 102637, 102602.1, 102548.2, 102479, 102386.8, 102276.3,
  102305, 102372.1, 102433.4, 102491.5, 102548.8, 102595.9, 102639, 102669.6, 
    102692.7, 102703.3, 102692.8, 102664.7, 102617.5, 102555.6, 102475.7,
  102214.9, 102293.3, 102364.1, 102432.7, 102499.1, 102560.6, 102616.4, 
    102661.9, 102703.5, 102728.9, 102742, 102736.6, 102714.9, 102672.3, 
    102612.6,
  102108, 102194, 102270.2, 102350.1, 102425.9, 102501.3, 102570, 102631.7, 
    102686, 102733.3, 102768.2, 102783.9, 102782.5, 102763.8, 102728.8,
  101993.3, 102082, 102165.8, 102255.9, 102339.2, 102423, 102502.9, 102579.1, 
    102648.7, 102711.4, 102762, 102797, 102816.5, 102817.5, 102804.4,
  101858.8, 101956.4, 102040.9, 102139.1, 102230.6, 102326.7, 102416.8, 
    102507.2, 102591.6, 102668.4, 102733.9, 102784.9, 102824.8, 102847.4, 
    102856.9,
  101716.3, 101818, 101906.8, 102010.3, 102106.8, 102212.8, 102313.9, 102414, 
    102510.4, 102599.3, 102677.8, 102745.5, 102800.5, 102844.9, 102874.7,
  101572, 101665.9, 101757.4, 101866.3, 101971.3, 102085.1, 102195.9, 
    102307.9, 102415.6, 102517.1, 102609.3, 102689.9, 102761.3, 102821.3, 
    102869.3,
  102187.9, 102081.3, 101930.4, 101748.5, 101523.1, 101282.9, 101038.6, 
    100913.6, 100724.3, 100549.1, 100352.2, 100221.4, 100119.1, 99991.49, 
    99846.05,
  102285.5, 102204.5, 102087, 101935.3, 101743.8, 101529.8, 101290.4, 101152, 
    100941.3, 100748.8, 100538.2, 100356.3, 100200.2, 100055.2, 99893.03,
  102363.6, 102313.6, 102235.5, 102119.1, 101957, 101765.5, 101529, 101368.3, 
    101156.4, 100926.2, 100720.1, 100532.3, 100344.5, 100172.4, 99980.52,
  102399, 102377.6, 102333, 102253.6, 102140.2, 101989.8, 101788.7, 101599.4, 
    101422.9, 101188.2, 100944.4, 100731.1, 100530, 100337.2, 100131.8,
  102406.2, 102413.1, 102386.8, 102339.3, 102257.4, 102150.8, 101999.1, 
    101833, 101660.5, 101453.7, 101212.7, 100978.3, 100763.9, 100561.4, 
    100346.5,
  102392.1, 102424.4, 102430.4, 102412.2, 102360.7, 102281.7, 102166.6, 
    102024.2, 101867.1, 101685, 101475.2, 101250.6, 101027.4, 100816.6, 
    100595.9,
  102350.6, 102401.6, 102435.3, 102444.2, 102429, 102381.1, 102305.9, 
    102200.4, 102064.8, 101901.6, 101716.8, 101519.5, 101310.5, 101099.3, 
    100880.7,
  102280.2, 102352.7, 102415.3, 102453.7, 102467.5, 102452.1, 102404.3, 
    102334.2, 102234, 102103.3, 101945.7, 101768, 101581.3, 101386.6, 101176.3,
  102175.3, 102280.4, 102358.2, 102427.5, 102471.2, 102488.8, 102476.8, 
    102438.1, 102365.9, 102268.5, 102145.5, 102000.6, 101835.3, 101657.3, 
    101468.8,
  102037.5, 102168.5, 102274.9, 102373.9, 102442.4, 102491.2, 102509.7, 
    102503.7, 102467.7, 102400.6, 102309.1, 102194.5, 102060.2, 101909.6, 
    101740.9,
  101057.8, 100970.8, 100869.2, 100767, 100643, 100532, 100439.7, 100375.7, 
    100302.9, 100226.9, 100153.6, 100085.3, 100028.4, 99987.72, 99969.81,
  101078.9, 100965.7, 100837.3, 100718.9, 100575, 100437.8, 100312.6, 
    100216.1, 100134.1, 100042.3, 99951.71, 99866.59, 99787.23, 99723.58, 
    99676.47,
  101099.5, 100976.2, 100829.5, 100690.7, 100526.9, 100364.3, 100200.9, 
    100068.9, 99968.08, 99865.57, 99743.86, 99632.05, 99522.59, 99423.52, 
    99344.65,
  101141.7, 101006.1, 100840.4, 100679.8, 100499.4, 100314.1, 100119.4, 
    99958.78, 99828.67, 99703.36, 99572.75, 99427.01, 99288.84, 99163.22, 
    99052.06,
  101206.8, 101065.2, 100885.1, 100711.8, 100515.6, 100313, 100098.1, 
    99888.95, 99725.66, 99568.14, 99414.46, 99252.91, 99087.47, 98931.9, 
    98793.27,
  101284.9, 101142.9, 100955.3, 100768.8, 100561.9, 100347.4, 100116, 
    99883.45, 99677.37, 99495.55, 99309.96, 99126.13, 98938.94, 98760.21, 
    98600.18,
  101369.9, 101233.2, 101045.8, 100854.9, 100641.5, 100419.2, 100180.9, 
    99930.96, 99687.07, 99472.94, 99268.83, 99058.63, 98847.45, 98647.54, 
    98468.21,
  101451.2, 101321.3, 101144.1, 100955.5, 100744.3, 100520.2, 100278.8, 
    100029.1, 99768.77, 99520.22, 99294.22, 99072.75, 98831.68, 98598.05, 
    98402.91,
  101529.8, 101404.8, 101247.3, 101067.8, 100861.4, 100642.2, 100404.9, 
    100154.8, 99896.09, 99630.2, 99379.25, 99140.48, 98902.8, 98656.88, 
    98445.48,
  101618.2, 101488.3, 101338.7, 101178.6, 100988.2, 100779.1, 100551.6, 
    100307.5, 100050.9, 99786.02, 99522.76, 99274.45, 99042.74, 98818.77, 
    98613.76,
  101649.1, 101602.2, 101542.6, 101483.8, 101424.8, 101368.7, 101315.1, 
    101264, 101216.2, 101171.9, 101127.7, 101080.5, 101032.7, 100980.6, 
    100923.7,
  101600.1, 101534.9, 101468.2, 101399.6, 101332, 101267.8, 101204.2, 
    101146.7, 101095.1, 101048.6, 101002.4, 100959.1, 100915.7, 100869.7, 
    100824.6,
  101535.5, 101461.9, 101387.8, 101307.9, 101231.9, 101154.9, 101083.5, 
    101018.4, 100962.6, 100912.4, 100866.7, 100827.5, 100788.8, 100753.3, 
    100719,
  101476.9, 101391.4, 101305.5, 101213.4, 101123.9, 101035.7, 100951, 100877, 
    100811.9, 100754.9, 100705.3, 100661.8, 100624.5, 100594.6, 100569.9,
  101420, 101321.6, 101222.9, 101119.2, 101013.9, 100911.8, 100816.5, 
    100727.8, 100647.4, 100577.6, 100515.5, 100465.2, 100426.6, 100401.2, 
    100386.3,
  101364.6, 101254.8, 101143.4, 101021.6, 100902.5, 100786.3, 100669.1, 
    100558.4, 100459.3, 100369, 100291.3, 100232.3, 100188.5, 100164.7, 
    100154.5,
  101316.1, 101192.8, 101065.2, 100931, 100796.8, 100659.2, 100518.8, 
    100388.1, 100262.7, 100149.6, 100056.8, 99985.03, 99936.96, 99910.21, 
    99901.35,
  101268.8, 101135.4, 100995.4, 100849.4, 100694, 100534, 100369.6, 100213.5, 
    100066.1, 99933.41, 99817.75, 99729.09, 99669.9, 99640.38, 99642.68,
  101225.1, 101089.8, 100936.9, 100774.1, 100600.9, 100421.6, 100235.3, 
    100055.9, 99879.51, 99722.75, 99589.8, 99488.52, 99423.59, 99403.95, 
    99417.13,
  101188.5, 101048.1, 100884.5, 100711.3, 100522.8, 100324.6, 100119.2, 
    99917.52, 99720.98, 99540.78, 99389.17, 99262.44, 99186.81, 99166.19, 
    99184.54,
  101841, 101756.9, 101649.6, 101531.8, 101398.5, 101248, 101085.6, 100915.6, 
    100743.9, 100579.5, 100458.8, 100400.9, 100382.5, 100360.9, 100333.9,
  101842, 101754.2, 101648, 101531, 101396.6, 101250.3, 101093.3, 100928.3, 
    100758, 100599.6, 100471.6, 100429, 100385.1, 100337.7, 100313.6,
  101832.9, 101747.1, 101644.3, 101530.6, 101403.1, 101262.3, 101108.3, 
    100947.8, 100779.8, 100621.7, 100480.8, 100417.4, 100350.4, 100318.1, 
    100282.6,
  101822.1, 101735.5, 101633.2, 101522.4, 101398.2, 101259.9, 101110.6, 
    100952.7, 100786.9, 100630.6, 100487.5, 100409.5, 100339.9, 100309.1, 
    100256.8,
  101807.8, 101719.5, 101619.2, 101509.4, 101388.2, 101254.7, 101109, 
    100959.7, 100794, 100641.7, 100494.4, 100396.4, 100330.8, 100300, 100241,
  101789.3, 101699.6, 101597, 101488.7, 101370.7, 101241.1, 101097.9, 
    100954.6, 100793.3, 100637.9, 100498.8, 100393.7, 100337.6, 100308.2, 
    100244.3,
  101767.9, 101674.2, 101571.8, 101462.9, 101348.2, 101224.4, 101083.2, 
    100945.4, 100787.9, 100636.9, 100505.3, 100398.7, 100350.3, 100306.6, 
    100244.3,
  101740.9, 101645.7, 101541.3, 101431.5, 101315.2, 101192.8, 101058.7, 
    100923.6, 100774.3, 100628.5, 100503.9, 100410.8, 100360.1, 100302.4, 
    100244.7,
  101711.4, 101614.8, 101507.4, 101394.5, 101273.9, 101153.6, 101019.8, 
    100889, 100746.7, 100615.5, 100502.7, 100420.1, 100361.2, 100301.2, 
    100246.5,
  101680.2, 101580.3, 101469.6, 101352, 101228.6, 101101.1, 100969.7, 
    100839.3, 100705.5, 100592.6, 100493, 100412.7, 100350.2, 100290.7, 
    100241.6,
  101322, 101247.5, 101159.5, 101078.5, 100992.6, 100921.9, 100861.8, 
    100815.7, 100791.9, 100785.1, 100782.1, 100767.7, 100739.8, 100708.4, 
    100665.3,
  101305.4, 101221.6, 101125, 101027.7, 100929.2, 100845.7, 100770, 100714.4, 
    100680, 100670.7, 100683.6, 100679.4, 100658.2, 100624.3, 100581.9,
  101295.8, 101204.9, 101097.7, 100989.6, 100874.9, 100771.4, 100680.4, 
    100611.8, 100567.7, 100564.6, 100587.9, 100588.6, 100570.6, 100543.2, 
    100501.1,
  101288.4, 101186.8, 101071.6, 100948.5, 100823, 100703.4, 100599.8, 
    100518.5, 100466.4, 100462.1, 100486, 100500.9, 100486.5, 100462.8, 
    100422.7,
  101290.6, 101181.1, 101055.7, 100920.1, 100784.6, 100651.9, 100532.7, 
    100437.9, 100379.6, 100375.3, 100399.3, 100415.1, 100405.4, 100385.2, 
    100345.1,
  101298.8, 101181.4, 101043.1, 100894.1, 100748.5, 100602.6, 100469.9, 
    100368.1, 100301, 100299, 100307.5, 100321.4, 100327.4, 100304.6, 100267.2,
  101313.7, 101187.4, 101035.4, 100876.2, 100717.6, 100558.9, 100414.3, 
    100303.1, 100217.9, 100211.5, 100204.4, 100218.1, 100244.6, 100226.2, 
    100193,
  101337.6, 101200.2, 101036.1, 100866, 100692.9, 100522.9, 100361.9, 
    100239.7, 100137.4, 100121.2, 100103.1, 100110.5, 100163.3, 100148.9, 
    100120.8,
  101369.6, 101218, 101045.1, 100860.4, 100675.8, 100491.3, 100316.4, 
    100180.2, 100059, 100026.7, 99998.45, 100009.8, 100078.9, 100074.8, 
    100059.1,
  101409.4, 101244.3, 101062, 100866.8, 100668.2, 100471.8, 100286, 100139.5, 
    100002.2, 99947.83, 99909.41, 99928.11, 100001.2, 100005.9, 100004.2,
  101825.6, 101815.9, 101795.2, 101774.3, 101748.6, 101725.2, 101695.7, 
    101659.2, 101618.4, 101572.4, 101523.4, 101471.7, 101414.6, 101356.3, 
    101292,
  101796.6, 101779.6, 101758.9, 101729.5, 101698.6, 101668, 101635.8, 
    101600.7, 101560.6, 101513.7, 101461.5, 101407.5, 101350.4, 101289.5, 
    101223.6,
  101756.4, 101736.8, 101711.4, 101678.3, 101646.8, 101611.9, 101577, 
    101539.4, 101497.6, 101450.9, 101400.2, 101343, 101281.2, 101218.4, 101149,
  101722.2, 101699.6, 101669.7, 101634.9, 101597, 101557.9, 101518.1, 
    101478.9, 101435.9, 101389.9, 101335.3, 101275.5, 101211.5, 101147.1, 
    101080.4,
  101687.2, 101660, 101626.3, 101589.1, 101548.2, 101505.5, 101459.4, 
    101414.9, 101368.8, 101319.8, 101267.1, 101208.9, 101144.3, 101076.3, 
    101004.6,
  101659.4, 101627.5, 101591.2, 101550.6, 101502.1, 101451.7, 101400.4, 
    101354.3, 101308.7, 101255.4, 101198.4, 101135, 101070.6, 101001.9, 100933,
  101628.3, 101593.6, 101553.1, 101506.5, 101457, 101402.6, 101344.8, 
    101290.8, 101236.4, 101180.9, 101119.4, 101065.7, 101002.4, 100937.6, 
    100862.7,
  101594.7, 101556.7, 101516.8, 101471, 101412.1, 101349.7, 101289.7, 
    101229.2, 101170.5, 101113.2, 101050.3, 100991.3, 100924.8, 100859, 
    100779.7,
  101561.8, 101527.4, 101480, 101424.9, 101364.9, 101297.2, 101230.5, 
    101167.1, 101102, 101041.4, 100980.9, 100917.1, 100846.1, 100778.5, 
    100706.3,
  101521.7, 101493.4, 101440, 101386.3, 101313.4, 101243.6, 101172, 101104, 
    101035.1, 100970.3, 100903.1, 100837, 100771.6, 100701.1, 100631.5,
  102381, 102379, 102365.9, 102348.4, 102329.7, 102304.6, 102273.5, 102235.9, 
    102190.6, 102137.2, 102079.9, 102015.9, 101950.9, 101877.6, 101799.2,
  102375.3, 102351.2, 102339.2, 102320.1, 102301.4, 102275.2, 102243.1, 
    102204.5, 102157.4, 102106.1, 102045.7, 101982.9, 101914.9, 101841.8, 
    101762.7,
  102335.3, 102325.5, 102310, 102292.7, 102272.7, 102243.7, 102209.8, 
    102170.1, 102121.7, 102068, 102011.8, 101945.8, 101874.4, 101801.1, 
    101721.4,
  102310.8, 102298.5, 102281.6, 102263.5, 102238.5, 102209.6, 102173.9, 
    102130.2, 102081.1, 102028, 101967.8, 101900.8, 101828.9, 101752.2, 
    101669.2,
  102284.6, 102271.4, 102253.4, 102229.8, 102205, 102173.4, 102133.9, 
    102089.5, 102040.3, 101984.9, 101924.6, 101854.6, 101779.5, 101698.7, 
    101614.3,
  102256.8, 102238.9, 102219.6, 102194.5, 102166.9, 102132.8, 102092, 
    102044.5, 101994.2, 101936, 101872.9, 101802.5, 101724.9, 101641.8, 
    101557.5,
  102223.9, 102205.2, 102185.3, 102156.5, 102127.2, 102090.9, 102048.3, 
    101999.5, 101944.9, 101885.3, 101818.9, 101745.3, 101668.2, 101581.5, 
    101494.3,
  102188.3, 102169.5, 102147.4, 102117.1, 102083.1, 102044.4, 102002.5, 
    101948.5, 101892.4, 101829.6, 101759.8, 101685.4, 101606.3, 101519.7, 
    101426.8,
  102152.7, 102133.6, 102111.2, 102077.2, 102040.5, 102001.7, 101951.2, 
    101897.2, 101837, 101772.4, 101701.9, 101626.5, 101543.7, 101451.6, 
    101355.3,
  102114.3, 102096, 102070.7, 102035, 101993.1, 101944.9, 101894.7, 101840.4, 
    101779.5, 101712.3, 101640.9, 101561.6, 101476.7, 101383.5, 101280.3,
  102899.6, 102882.6, 102868.6, 102834.8, 102801.1, 102748.9, 102685.3, 
    102603.8, 102511.1, 102410, 102306.1, 102184.3, 102049.8, 101899, 101733.2,
  102908.1, 102894.2, 102886.4, 102854.5, 102821.1, 102772.6, 102709.8, 
    102634.3, 102548.7, 102455.4, 102352.1, 102241, 102110.4, 101966.2, 
    101807.3,
  102911.8, 102898.8, 102882.4, 102854.3, 102827, 102783.7, 102730.9, 
    102659.4, 102577.8, 102487.3, 102395.8, 102291.8, 102165.9, 102024.1, 
    101867.4,
  102904.3, 102889.2, 102868.5, 102844.9, 102818.2, 102783, 102732.6, 
    102676.2, 102603.6, 102520.1, 102428.8, 102328.4, 102210.9, 102072.9, 
    101918.1,
  102889.9, 102870.5, 102851.8, 102828.7, 102803.7, 102774.8, 102736.3, 
    102682.7, 102615.6, 102540.2, 102452.6, 102354.6, 102244, 102110.6, 
    101961.8,
  102858.8, 102841.4, 102827.9, 102808, 102789.3, 102761.8, 102727.2, 
    102674.8, 102615.9, 102543.2, 102464.2, 102371.5, 102264.4, 102136.2, 
    101993.1,
  102826.2, 102809.7, 102801.8, 102785.6, 102766.4, 102739.4, 102704.6, 
    102656.2, 102602, 102536, 102458.9, 102374.7, 102274.8, 102153.7, 102018.3,
  102793.3, 102777.7, 102766.8, 102746.1, 102726.5, 102702.6, 102667.5, 
    102625.8, 102572.2, 102510.2, 102441.4, 102365.1, 102272.8, 102162.4, 
    102034,
  102747.4, 102732.1, 102717.5, 102696.1, 102674.7, 102650.3, 102619.2, 
    102576.5, 102532.1, 102479, 102417.9, 102346.5, 102260.2, 102159.7, 
    102042.1,
  102696.7, 102681.4, 102663.7, 102643.3, 102620.1, 102594.5, 102563, 
    102526.9, 102485.2, 102443.2, 102385.9, 102319.5, 102238.3, 102144, 
    102036.6 ;

 sftlf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 time_bnds =
  0, 1,
  1, 2,
  2, 3,
  3, 4,
  4, 5,
  5, 6,
  6, 7,
  7, 8,
  8, 9,
  9, 10,
  10, 11,
  11, 12,
  12, 13,
  13, 14,
  14, 15,
  15, 16,
  16, 17,
  17, 18,
  18, 19,
  19, 20,
  20, 21,
  21, 22,
  22, 23,
  23, 24,
  24, 25,
  25, 26,
  26, 27,
  27, 28,
  28, 29,
  29, 30,
  30, 31,
  31, 32,
  32, 33,
  33, 34,
  34, 35,
  35, 36,
  36, 37,
  37, 38,
  38, 39,
  39, 40,
  40, 41,
  41, 42,
  42, 43,
  43, 44,
  44, 45,
  45, 46,
  46, 47,
  47, 48,
  48, 49,
  49, 50,
  50, 51,
  51, 52,
  52, 53,
  53, 54,
  54, 55,
  55, 56,
  56, 57,
  57, 58,
  58, 59,
  59, 60,
  60, 61,
  61, 62,
  62, 63,
  63, 64,
  64, 65,
  65, 66,
  66, 67,
  67, 68,
  68, 69,
  69, 70,
  70, 71,
  71, 72,
  72, 73,
  73, 74,
  74, 75,
  75, 76,
  76, 77,
  77, 78,
  78, 79,
  79, 80,
  80, 81,
  81, 82,
  82, 83,
  83, 84,
  84, 85,
  85, 86,
  86, 87,
  87, 88,
  88, 89,
  89, 90,
  90, 91,
  91, 92,
  92, 93,
  93, 94,
  94, 95,
  95, 96,
  96, 97,
  97, 98,
  98, 99,
  99, 100,
  100, 101,
  101, 102,
  102, 103,
  103, 104,
  104, 105,
  105, 106,
  106, 107,
  107, 108,
  108, 109,
  109, 110,
  110, 111,
  111, 112,
  112, 113,
  113, 114,
  114, 115,
  115, 116,
  116, 117,
  117, 118,
  118, 119,
  119, 120,
  120, 121,
  121, 122,
  122, 123,
  123, 124,
  124, 125,
  125, 126,
  126, 127,
  127, 128,
  128, 129,
  129, 130,
  130, 131,
  131, 132,
  132, 133,
  133, 134,
  134, 135,
  135, 136,
  136, 137,
  137, 138,
  138, 139,
  139, 140,
  140, 141,
  141, 142,
  142, 143,
  143, 144,
  144, 145,
  145, 146,
  146, 147,
  147, 148,
  148, 149,
  149, 150,
  150, 151,
  151, 152,
  152, 153,
  153, 154,
  154, 155,
  155, 156,
  156, 157,
  157, 158,
  158, 159,
  159, 160,
  160, 161,
  161, 162,
  162, 163,
  163, 164,
  164, 165,
  165, 166,
  166, 167,
  167, 168,
  168, 169,
  169, 170,
  170, 171,
  171, 172,
  172, 173,
  173, 174,
  174, 175,
  175, 176,
  176, 177,
  177, 178,
  178, 179,
  179, 180,
  180, 181,
  181, 182 ;

 zsurf =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 grid_xt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15 ;

 grid_yt = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10 ;

 nv = 1, 2 ;

 pfull = 0.0252729048206747, 0.0885404738757409, 0.213072411383256, 
    0.41190537807884, 0.671080828691593, 0.987471468515016, 1.36790961365676, 
    1.82562112064242, 2.38097588033244, 3.06218961364243, 3.90121721567151, 
    4.9296281825995, 6.18008131929323, 7.68875807563375, 9.49537809361575, 
    11.643153995098, 14.1786857151188, 17.1517875598959, 20.6152476986609, 
    24.6245259348741, 29.237386591333, 34.5134757786445, 40.5138467378254, 
    47.3004421634272, 54.9355325495126, 63.4811392623337, 72.9984371159701, 
    83.5471442618119, 95.1849171805989, 107.966767294215, 121.944503506415, 
    137.166169497631, 153.675572970355, 171.511834307961, 190.708985325578, 
    211.295632932361, 233.294677858721, 256.723099608772, 281.591803639405, 
    307.905555737256, 335.66293113824, 364.856338389786, 395.47216160598, 
    427.490864234311, 460.887168786725, 495.630391513078, 531.761718445649, 
    569.289185351388, 607.768705103107, 646.445374671436, 684.792067788697, 
    722.468679913451, 759.124006783627, 794.401045766566, 827.769968639223, 
    858.597822486016, 886.389109609622, 910.841030891388, 931.860653469283, 
    949.549679924174, 964.159924710431, 976.012345333387, 985.470174132691, 
    992.77226220014, 997.948601287575 ;

 phalf = 0.01, 0.0513470268, 0.1404240036, 0.3072783852, 0.5379505539, 
    0.8245489502, 1.170559845, 1.5862843323, 2.0879000854, 2.700272522, 
    3.4550848389, 4.3841940308, 5.5185266113, 6.8925054932, 8.5440936279, 
    10.5147802734, 12.8495031738, 15.5965148926, 18.8071691895, 
    22.5356542969, 26.8386547852, 31.7749560547, 37.4049951172, 
    43.7903613281, 50.9932617188, 59.0759326172, 68.100078125, 78.1262353516, 
    89.2131933594, 101.4173632812, 114.7922466406, 129.3878501562, 
    145.2501478125, 162.4206823438, 180.9360560938, 200.8276451562, 
    222.1212074219, 244.8367185938, 268.9881007812, 294.5831945312, 
    321.6236510156, 350.1049399219, 380.0163883594, 411.3414303125, 
    444.0575547656, 478.1367280469, 513.5456339062, 550.403556875, 
    588.6019571094, 627.3470909766, 665.9273852344, 704.0097012891, 
    741.2475327734, 777.2856108203, 811.7659041211, 843.9830114648, 
    873.3803854492, 899.5263707422, 922.2501762402, 941.5376650684, 
    957.6070185254, 970.7426572876, 981.30107, 989.65107, 995.9000099865, 1000 ;

 scalar_axis = 0 ;

 time = 0.5, 1.5, 2.5, 3.5, 4.5, 5.5, 6.5, 7.5, 8.5, 9.5, 10.5, 11.5, 12.5, 
    13.5, 14.5, 15.5, 16.5, 17.5, 18.5, 19.5, 20.5, 21.5, 22.5, 23.5, 24.5, 
    25.5, 26.5, 27.5, 28.5, 29.5, 30.5, 31.5, 32.5, 33.5, 34.5, 35.5, 36.5, 
    37.5, 38.5, 39.5, 40.5, 41.5, 42.5, 43.5, 44.5, 45.5, 46.5, 47.5, 48.5, 
    49.5, 50.5, 51.5, 52.5, 53.5, 54.5, 55.5, 56.5, 57.5, 58.5, 59.5, 60.5, 
    61.5, 62.5, 63.5, 64.5, 65.5, 66.5, 67.5, 68.5, 69.5, 70.5, 71.5, 72.5, 
    73.5, 74.5, 75.5, 76.5, 77.5, 78.5, 79.5, 80.5, 81.5, 82.5, 83.5, 84.5, 
    85.5, 86.5, 87.5, 88.5, 89.5, 90.5, 91.5, 92.5, 93.5, 94.5, 95.5, 96.5, 
    97.5, 98.5, 99.5, 100.5, 101.5, 102.5, 103.5, 104.5, 105.5, 106.5, 107.5, 
    108.5, 109.5, 110.5, 111.5, 112.5, 113.5, 114.5, 115.5, 116.5, 117.5, 
    118.5, 119.5, 120.5, 121.5, 122.5, 123.5, 124.5, 125.5, 126.5, 127.5, 
    128.5, 129.5, 130.5, 131.5, 132.5, 133.5, 134.5, 135.5, 136.5, 137.5, 
    138.5, 139.5, 140.5, 141.5, 142.5, 143.5, 144.5, 145.5, 146.5, 147.5, 
    148.5, 149.5, 150.5, 151.5, 152.5, 153.5, 154.5, 155.5, 156.5, 157.5, 
    158.5, 159.5, 160.5, 161.5, 162.5, 163.5, 164.5, 165.5, 166.5, 167.5, 
    168.5, 169.5, 170.5, 171.5, 172.5, 173.5, 174.5, 175.5, 176.5, 177.5, 
    178.5, 179.5, 180.5, 181.5 ;
}
