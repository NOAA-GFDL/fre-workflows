netcdf \00010101.ocean_annual.so {
dimensions:
	time = UNLIMITED ; // (1 currently)
	zl = 75 ;
	yh = 10 ;
	xh = 15 ;
	nv = 2 ;
	xq = 1441 ;
	yq = 1162 ;
	zi = 76 ;
variables:
	double average_DT(time) ;
		average_DT:_FillValue = 1.e+20 ;
		average_DT:missing_value = 1.e+20 ;
		average_DT:units = "days" ;
		average_DT:long_name = "Length of average period" ;
	double average_T1(time) ;
		average_T1:_FillValue = 1.e+20 ;
		average_T1:missing_value = 1.e+20 ;
		average_T1:units = "days since 0001-01-01 00:00:00" ;
		average_T1:long_name = "Start time for average period" ;
	double average_T2(time) ;
		average_T2:_FillValue = 1.e+20 ;
		average_T2:missing_value = 1.e+20 ;
		average_T2:units = "days since 0001-01-01 00:00:00" ;
		average_T2:long_name = "End time for average period" ;
	float so(time, zl, yh, xh) ;
		so:_FillValue = 1.e+20f ;
		so:missing_value = 1.e+20f ;
		so:units = "psu" ;
		so:long_name = "Sea Water Salinity" ;
		so:cell_methods = "area:mean zl:mean yh:mean xh:mean time: mean" ;
		so:cell_measures = "volume: volcello area: areacello" ;
		so:time_avg_info = "average_T1,average_T2,average_DT" ;
		so:standard_name = "sea_water_salinity" ;
	double time_bnds(time, nv) ;
		time_bnds:long_name = "time axis boundaries" ;
	double nv(nv) ;
		nv:long_name = "vertex number" ;
	double time(time) ;
		time:units = "days since 0001-01-01 00:00:00" ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:calendar_type = "NOLEAP" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;
	double xh(xh) ;
		xh:units = "degrees_east" ;
		xh:long_name = "h point nominal longitude" ;
		xh:axis = "X" ;
	double xq(xq) ;
		xq:units = "degrees_east" ;
		xq:long_name = "q point nominal longitude" ;
		xq:axis = "X" ;
	double yh(yh) ;
		yh:units = "degrees_north" ;
		yh:long_name = "h point nominal latitude" ;
		yh:axis = "Y" ;
	double yq(yq) ;
		yq:units = "degrees_north" ;
		yq:long_name = "q point nominal latitude" ;
		yq:axis = "Y" ;
	double zi(zi) ;
		zi:units = "meter" ;
		zi:long_name = "Interface z-rho" ;
		zi:axis = "Z" ;
		zi:positive = "down" ;
	double zl(zl) ;
		zl:units = "meter" ;
		zl:long_name = "Layer z-rho" ;
		zl:axis = "Z" ;
		zl:positive = "down" ;

// global attributes:
		:title = "cm5_c96_am5f7c1r0_b06_piC_galb_noiceinit_alb" ;
		:associated_files = "areacello: 00010101.ocean_static.nc" ;
		:grid_type = "regular" ;
		:grid_tile = "N/A" ;
		:history = "Fri Aug 29 13:42:28 2025: ncks -d xh,532,546 -d yh,526,535 /work/cew/scratch//00010101.ocean_annual.nc -O /work/cew/scratch/workflow-test/ocean_annual//ncks_out//00010101.ocean_annual.nc" ;
		:NCO = "netCDF Operators version 5.1.9 (Homepage = http://nco.sf.net, Code = http://github.com/nco/nco, Citation = 10.1016/j.envsoft.2008.03.004)" ;
data:

 average_DT = 365 ;

 average_T1 = 0 ;

 average_T2 = 365 ;

 so =
  35.38194, 35.38821, 35.39954, 35.41414, 35.42913, 35.44204, 35.45264, 
    35.46775, 35.49113, 35.51057, 35.52499, 35.53934, 35.55696, 35.57177, 
    35.58615,
  35.38625, 35.40103, 35.4178, 35.43279, 35.44572, 35.46037, 35.47413, 
    35.48968, 35.50805, 35.52221, 35.53437, 35.54751, 35.56369, 35.57827, 
    35.59275,
  35.3838, 35.40005, 35.42051, 35.43718, 35.45137, 35.47016, 35.49076, 
    35.50874, 35.52416, 35.5348, 35.54519, 35.55713, 35.57343, 35.58828, 
    35.60341,
  35.37607, 35.39221, 35.41131, 35.43444, 35.45382, 35.48092, 35.50257, 
    35.51928, 35.53342, 35.54388, 35.5533, 35.56441, 35.58146, 35.59866, 
    35.61461,
  35.37418, 35.39106, 35.40664, 35.42981, 35.45753, 35.48639, 35.50614, 
    35.52135, 35.53499, 35.54509, 35.55459, 35.56549, 35.58228, 35.59885, 
    35.61545,
  35.37721, 35.4015, 35.41866, 35.44059, 35.46667, 35.48727, 35.50368, 
    35.51868, 35.53247, 35.54332, 35.55313, 35.56251, 35.57658, 35.59302, 
    35.6111,
  35.38316, 35.40884, 35.42866, 35.44965, 35.47217, 35.48794, 35.50311, 
    35.51721, 35.52999, 35.53999, 35.5494, 35.55816, 35.57151, 35.58783, 
    35.60601,
  35.39457, 35.41843, 35.437, 35.45594, 35.47628, 35.49221, 35.50801, 
    35.52194, 35.53466, 35.54383, 35.55301, 35.56104, 35.57311, 35.58829, 
    35.60509,
  35.40924, 35.4287, 35.44646, 35.46474, 35.48413, 35.49978, 35.5155, 
    35.52979, 35.54054, 35.54808, 35.55649, 35.56492, 35.57736, 35.59256, 
    35.60772,
  35.42995, 35.44503, 35.46258, 35.48032, 35.49793, 35.51563, 35.53004, 
    35.54128, 35.54697, 35.55147, 35.55875, 35.5676, 35.57998, 35.59457, 
    35.61117,
  35.38515, 35.39331, 35.4041, 35.41836, 35.43325, 35.44681, 35.45716, 
    35.4716, 35.49395, 35.51293, 35.52738, 35.54174, 35.55928, 35.57396, 
    35.58816,
  35.38979, 35.40578, 35.42229, 35.43704, 35.44986, 35.46405, 35.4773, 
    35.49271, 35.51057, 35.52448, 35.53669, 35.54977, 35.56575, 35.58005, 
    35.59443,
  35.38698, 35.40525, 35.42514, 35.44158, 35.4551, 35.47254, 35.49311, 
    35.51123, 35.52684, 35.5377, 35.54781, 35.55943, 35.57509, 35.58972, 
    35.60467,
  35.37942, 35.39743, 35.41582, 35.43849, 35.45691, 35.48314, 35.50468, 
    35.52154, 35.53577, 35.54652, 35.5559, 35.56697, 35.58323, 35.60015, 
    35.61584,
  35.37748, 35.39586, 35.4108, 35.43351, 35.46047, 35.4885, 35.50816, 
    35.52341, 35.5372, 35.5477, 35.55688, 35.56778, 35.58395, 35.60012, 
    35.61654,
  35.38161, 35.40561, 35.42241, 35.44406, 35.46995, 35.49122, 35.50698, 
    35.52107, 35.53478, 35.54577, 35.55535, 35.56457, 35.57816, 35.59423, 
    35.61211,
  35.38746, 35.41281, 35.43246, 35.45338, 35.47598, 35.49348, 35.50812, 
    35.52145, 35.53433, 35.54527, 35.55459, 35.56268, 35.5747, 35.59037, 
    35.60786,
  35.39887, 35.42252, 35.4407, 35.45959, 35.47999, 35.49775, 35.51317, 
    35.52628, 35.53896, 35.54946, 35.55837, 35.56607, 35.57674, 35.59154, 
    35.60795,
  35.41398, 35.43335, 35.45085, 35.46898, 35.48827, 35.50565, 35.52086, 
    35.53485, 35.5457, 35.55447, 35.56245, 35.57046, 35.58164, 35.59639, 
    35.61097,
  35.43533, 35.4514, 35.4687, 35.48628, 35.50359, 35.52119, 35.53553, 
    35.54677, 35.55321, 35.55897, 35.56569, 35.57408, 35.58544, 35.59848, 
    35.61447,
  35.38759, 35.39647, 35.40701, 35.42113, 35.4362, 35.44971, 35.45957, 
    35.47409, 35.49628, 35.51489, 35.52929, 35.54372, 35.56107, 35.57567, 
    35.58994,
  35.39242, 35.40969, 35.42556, 35.43981, 35.45267, 35.46642, 35.47935, 
    35.49462, 35.51249, 35.52628, 35.53833, 35.55144, 35.5673, 35.58159, 
    35.59591,
  35.38934, 35.40922, 35.4283, 35.44445, 35.45859, 35.47433, 35.49478, 
    35.51292, 35.5287, 35.5397, 35.54966, 35.56112, 35.57637, 35.59091, 
    35.60585,
  35.38187, 35.40073, 35.41881, 35.44174, 35.4594, 35.48474, 35.50629, 
    35.52319, 35.53765, 35.54839, 35.5576, 35.56869, 35.58455, 35.60133, 
    35.61695,
  35.37993, 35.39923, 35.41389, 35.43633, 35.46284, 35.49025, 35.50989, 
    35.52507, 35.53883, 35.54947, 35.5586, 35.56939, 35.58517, 35.60125, 
    35.61755,
  35.38394, 35.40785, 35.42452, 35.44617, 35.472, 35.49337, 35.50922, 
    35.52296, 35.53647, 35.54775, 35.55714, 35.56628, 35.57942, 35.59536, 
    35.61312,
  35.38981, 35.41516, 35.4346, 35.45557, 35.47816, 35.49652, 35.51133, 
    35.52434, 35.5374, 35.54901, 35.55788, 35.56575, 35.57675, 35.59178, 
    35.60912,
  35.40145, 35.4249, 35.4431, 35.46185, 35.48241, 35.50124, 35.51651, 
    35.52953, 35.54233, 35.55322, 35.56188, 35.56924, 35.57892, 35.59325, 
    35.60945,
  35.41686, 35.4363, 35.4537, 35.47172, 35.49105, 35.50947, 35.52461, 
    35.53833, 35.54909, 35.55825, 35.56608, 35.57374, 35.5842, 35.59825, 
    35.61262,
  35.43799, 35.45456, 35.47185, 35.48933, 35.50647, 35.52436, 35.53834, 
    35.54925, 35.55607, 35.56235, 35.56894, 35.57715, 35.58799, 35.60083, 
    35.61628,
  35.39022, 35.39939, 35.40999, 35.42385, 35.43894, 35.45296, 35.46236, 
    35.4767, 35.49872, 35.51712, 35.53144, 35.546, 35.56322, 35.57791, 
    35.59226,
  35.39487, 35.41328, 35.42914, 35.44313, 35.45627, 35.4695, 35.4814, 
    35.49657, 35.51424, 35.52798, 35.54004, 35.55335, 35.56907, 35.5834, 
    35.59774,
  35.39198, 35.41296, 35.4323, 35.44832, 35.4635, 35.47623, 35.49639, 
    35.51448, 35.53022, 35.54136, 35.55115, 35.56262, 35.5776, 35.59215, 
    35.60712,
  35.38443, 35.40448, 35.42234, 35.4463, 35.46192, 35.48634, 35.5078, 
    35.52464, 35.53909, 35.54985, 35.55898, 35.57006, 35.58556, 35.6022, 
    35.6179,
  35.38251, 35.40257, 35.41682, 35.439, 35.46504, 35.49168, 35.51128, 
    35.52651, 35.54025, 35.55093, 35.56001, 35.57076, 35.58625, 35.6022, 
    35.61861,
  35.38623, 35.41003, 35.42627, 35.44793, 35.47373, 35.49487, 35.51075, 
    35.52463, 35.53786, 35.54925, 35.55862, 35.5677, 35.58055, 35.59639, 
    35.61416,
  35.39183, 35.41718, 35.43639, 35.4573, 35.47985, 35.49874, 35.51383, 
    35.52681, 35.54004, 35.55221, 35.56124, 35.5685, 35.57862, 35.59303, 
    35.61028,
  35.40367, 35.42701, 35.44506, 35.46374, 35.48434, 35.50396, 35.51941, 
    35.532, 35.54488, 35.55626, 35.56517, 35.57224, 35.58108, 35.59471, 
    35.61072,
  35.41907, 35.43877, 35.45606, 35.47398, 35.49312, 35.51196, 35.52718, 
    35.54054, 35.55153, 35.56076, 35.56879, 35.5765, 35.58645, 35.59967, 
    35.61388,
  35.44025, 35.45715, 35.4742, 35.49174, 35.50872, 35.5264, 35.54067, 
    35.55132, 35.55817, 35.56467, 35.57134, 35.57949, 35.58998, 35.60239, 
    35.61771,
  35.39338, 35.40301, 35.41418, 35.42779, 35.44289, 35.45768, 35.46548, 
    35.47967, 35.50157, 35.51947, 35.53351, 35.54811, 35.56537, 35.58018, 
    35.59461,
  35.39782, 35.41719, 35.43385, 35.44789, 35.46135, 35.47403, 35.48367, 
    35.49896, 35.51661, 35.53027, 35.54222, 35.55568, 35.57131, 35.5858, 
    35.6002,
  35.39471, 35.41727, 35.43816, 35.45432, 35.46898, 35.47877, 35.49829, 
    35.51624, 35.53178, 35.54309, 35.5529, 35.56445, 35.57919, 35.59385, 
    35.60887,
  35.38764, 35.40955, 35.42739, 35.45205, 35.46508, 35.48827, 35.50935, 
    35.52617, 35.54051, 35.55124, 35.56038, 35.57152, 35.58678, 35.60332, 
    35.61906,
  35.38667, 35.40683, 35.42012, 35.4421, 35.46761, 35.49334, 35.51279, 
    35.52801, 35.54162, 35.55235, 35.56152, 35.57234, 35.5875, 35.60332, 
    35.61974,
  35.39, 35.41349, 35.42841, 35.44989, 35.47547, 35.49641, 35.51234, 
    35.52629, 35.53953, 35.55128, 35.56058, 35.56943, 35.58201, 35.59778, 
    35.61551,
  35.39456, 35.41962, 35.43848, 35.45926, 35.48185, 35.50085, 35.51611, 
    35.5294, 35.54262, 35.55544, 35.56471, 35.57177, 35.58102, 35.59494, 
    35.61198,
  35.4062, 35.42967, 35.44743, 35.46596, 35.48641, 35.50637, 35.52216, 
    35.53467, 35.54729, 35.55929, 35.56849, 35.57555, 35.58379, 35.59672, 
    35.61258,
  35.42136, 35.44138, 35.4586, 35.47637, 35.49535, 35.51436, 35.52981, 
    35.54316, 35.55395, 35.56364, 35.57177, 35.57925, 35.58916, 35.60183, 
    35.61577,
  35.44261, 35.45968, 35.4767, 35.49423, 35.51123, 35.5288, 35.54304, 
    35.55363, 35.56043, 35.56707, 35.57375, 35.5819, 35.59242, 35.60452, 
    35.61955,
  35.39748, 35.40808, 35.41943, 35.43211, 35.44796, 35.46293, 35.4688, 
    35.4828, 35.50446, 35.5218, 35.53569, 35.5504, 35.56744, 35.58234, 
    35.59693,
  35.40298, 35.42355, 35.44011, 35.45369, 35.46664, 35.47842, 35.48639, 
    35.5015, 35.51915, 35.53266, 35.54471, 35.55813, 35.5736, 35.58823, 
    35.60276,
  35.3993, 35.42487, 35.44577, 35.46075, 35.47342, 35.48173, 35.50065, 
    35.5184, 35.53364, 35.54493, 35.55491, 35.56662, 35.58128, 35.59574, 
    35.61068,
  35.39365, 35.41742, 35.43492, 35.45781, 35.46891, 35.491, 35.5115, 
    35.52815, 35.54218, 35.55286, 35.56203, 35.57332, 35.58838, 35.60465, 
    35.62033,
  35.39393, 35.41348, 35.42454, 35.4459, 35.47084, 35.49566, 35.51484, 
    35.53004, 35.54337, 35.55408, 35.56321, 35.57412, 35.58909, 35.60462, 
    35.62098,
  35.39642, 35.41848, 35.43121, 35.45254, 35.4777, 35.49837, 35.51411, 
    35.52811, 35.54174, 35.55377, 35.563, 35.57197, 35.58405, 35.59942, 
    35.61691,
  35.399, 35.42308, 35.44109, 35.46165, 35.48402, 35.5032, 35.51847, 35.5318, 
    35.54519, 35.55878, 35.5684, 35.57567, 35.58434, 35.59764, 35.61423,
  35.40951, 35.43277, 35.44997, 35.46843, 35.48869, 35.50874, 35.5248, 
    35.53748, 35.55007, 35.56285, 35.57232, 35.57944, 35.58751, 35.59985, 
    35.61543,
  35.42385, 35.44407, 35.46128, 35.47905, 35.49789, 35.51712, 35.53263, 
    35.54597, 35.55672, 35.56731, 35.57567, 35.58295, 35.59279, 35.6048, 
    35.61863,
  35.44493, 35.46237, 35.47932, 35.49692, 35.51403, 35.53148, 35.54579, 
    35.55642, 35.5631, 35.57004, 35.57699, 35.58535, 35.59598, 35.60759, 
    35.6225,
  35.40371, 35.41476, 35.42598, 35.43792, 35.454, 35.46828, 35.47289, 
    35.48745, 35.50883, 35.52496, 35.53866, 35.55363, 35.57043, 35.58474, 
    35.59925,
  35.41017, 35.4311, 35.44705, 35.46022, 35.47197, 35.48264, 35.48979, 
    35.50479, 35.52203, 35.53536, 35.54763, 35.5613, 35.5761, 35.59038, 
    35.60502,
  35.40627, 35.43262, 35.45218, 35.46656, 35.47798, 35.48511, 35.50334, 
    35.52085, 35.53597, 35.5472, 35.55747, 35.56944, 35.58398, 35.59818, 
    35.61309,
  35.4015, 35.42493, 35.44188, 35.46292, 35.47326, 35.49436, 35.51408, 
    35.53056, 35.5443, 35.55466, 35.56387, 35.57536, 35.59046, 35.60637, 
    35.62201,
  35.40141, 35.42012, 35.43002, 35.45048, 35.47498, 35.49847, 35.5172, 
    35.53244, 35.54548, 35.55603, 35.56538, 35.57644, 35.59131, 35.60656, 
    35.62284,
  35.40412, 35.42381, 35.43562, 35.45634, 35.48064, 35.50068, 35.51624, 
    35.5303, 35.54424, 35.5571, 35.5666, 35.57536, 35.58688, 35.60189, 
    35.61908,
  35.40458, 35.42718, 35.44452, 35.46462, 35.48649, 35.50572, 35.52105, 
    35.53449, 35.54823, 35.56287, 35.57292, 35.58049, 35.58854, 35.60102, 
    35.61729,
  35.41342, 35.43602, 35.45293, 35.47121, 35.49116, 35.51138, 35.52765, 
    35.54041, 35.5536, 35.56741, 35.57776, 35.58521, 35.5927, 35.60395, 
    35.61901,
  35.42694, 35.4472, 35.46439, 35.48205, 35.50066, 35.52023, 35.53579, 
    35.54894, 35.55991, 35.57192, 35.5814, 35.58916, 35.5986, 35.60949, 
    35.62266,
  35.44735, 35.46529, 35.48211, 35.49969, 35.51683, 35.53434, 35.54893, 
    35.5596, 35.56642, 35.57407, 35.58213, 35.59129, 35.60222, 35.61272, 
    35.62709,
  35.41132, 35.42319, 35.43436, 35.44541, 35.46131, 35.47488, 35.47903, 
    35.4944, 35.51513, 35.52913, 35.54248, 35.55779, 35.57424, 35.58796, 
    35.60238,
  35.41821, 35.43888, 35.4544, 35.46683, 35.47787, 35.488, 35.49442, 
    35.50908, 35.52568, 35.53857, 35.55107, 35.56443, 35.57904, 35.59302, 
    35.60761,
  35.41416, 35.43983, 35.45826, 35.4721, 35.48269, 35.48898, 35.50692, 
    35.52414, 35.53907, 35.55001, 35.56062, 35.57258, 35.58707, 35.60109, 
    35.61605,
  35.40874, 35.43158, 35.44838, 35.46796, 35.47793, 35.49799, 35.51742, 
    35.53382, 35.54735, 35.55741, 35.56678, 35.57856, 35.59356, 35.60915, 
    35.6246,
  35.40783, 35.4264, 35.43619, 35.45574, 35.47931, 35.502, 35.52054, 
    35.53593, 35.54893, 35.55909, 35.56868, 35.58037, 35.59535, 35.61, 
    35.62591,
  35.4113, 35.42902, 35.44099, 35.46158, 35.48473, 35.50434, 35.52004, 
    35.53421, 35.54872, 35.56136, 35.57145, 35.58076, 35.59187, 35.606, 
    35.62242,
  35.41088, 35.43225, 35.44919, 35.46906, 35.49037, 35.50962, 35.52494, 
    35.53836, 35.55246, 35.56789, 35.57841, 35.58656, 35.59497, 35.60615, 
    35.62152,
  35.4185, 35.44075, 35.45695, 35.47528, 35.4953, 35.51554, 35.5317, 
    35.54421, 35.55851, 35.57329, 35.58406, 35.59173, 35.59995, 35.61002, 
    35.62377,
  35.43111, 35.45103, 35.46848, 35.48608, 35.50466, 35.52424, 35.53986, 
    35.55307, 35.56464, 35.57757, 35.58784, 35.5961, 35.6062, 35.61674, 
    35.62868,
  35.4506, 35.46871, 35.48538, 35.50272, 35.51989, 35.53763, 35.55254, 
    35.56341, 35.57045, 35.57915, 35.5882, 35.59803, 35.60956, 35.62032, 
    35.63381,
  35.4214, 35.43402, 35.44509, 35.45608, 35.47091, 35.48351, 35.48805, 
    35.50413, 35.52351, 35.53478, 35.54755, 35.56267, 35.57875, 35.59224, 
    35.60659,
  35.42753, 35.44772, 35.46276, 35.47486, 35.48583, 35.49529, 35.5009, 
    35.51492, 35.53045, 35.54303, 35.55532, 35.56858, 35.58269, 35.5964, 
    35.61095,
  35.42237, 35.44725, 35.46466, 35.47804, 35.48811, 35.49408, 35.51131, 
    35.52819, 35.54306, 35.55421, 35.5648, 35.57671, 35.59112, 35.60485, 
    35.61963,
  35.41616, 35.43847, 35.45497, 35.47345, 35.48329, 35.50291, 35.52174, 
    35.53793, 35.55146, 35.56171, 35.57112, 35.58307, 35.598, 35.61313, 
    35.62814,
  35.41428, 35.43286, 35.44263, 35.4615, 35.48462, 35.5064, 35.5247, 
    35.54025, 35.55383, 35.56406, 35.57401, 35.58577, 35.60026, 35.61433, 
    35.62964,
  35.41756, 35.43445, 35.44652, 35.46734, 35.48969, 35.50891, 35.52509, 
    35.53964, 35.55425, 35.56722, 35.57751, 35.58712, 35.59813, 35.61139, 
    35.62684,
  35.41626, 35.4378, 35.45436, 35.47467, 35.49524, 35.51416, 35.52989, 
    35.54362, 35.5574, 35.57332, 35.58397, 35.59225, 35.60128, 35.61226, 
    35.62683,
  35.42386, 35.44624, 35.46199, 35.48037, 35.50018, 35.5206, 35.53743, 35.55, 
    35.56437, 35.57869, 35.58914, 35.59694, 35.60578, 35.6165, 35.62974,
  35.43582, 35.4554, 35.4729, 35.49073, 35.50951, 35.52932, 35.54512, 
    35.55878, 35.57041, 35.5828, 35.59295, 35.60131, 35.61162, 35.62344, 
    35.63551,
  35.4543, 35.47256, 35.48932, 35.50637, 35.52346, 35.54147, 35.55681, 
    35.5677, 35.57465, 35.58402, 35.59344, 35.60346, 35.6151, 35.62714, 
    35.64123,
  35.43404, 35.44695, 35.45841, 35.4704, 35.48396, 35.49578, 35.50115, 
    35.517, 35.53466, 35.54288, 35.5542, 35.56892, 35.58493, 35.59787, 
    35.61174,
  35.43664, 35.45628, 35.47151, 35.48476, 35.49633, 35.50665, 35.51189, 
    35.52461, 35.53816, 35.54919, 35.56069, 35.5739, 35.58807, 35.60135, 
    35.61563,
  35.43, 35.45441, 35.47169, 35.4856, 35.49551, 35.50125, 35.51786, 35.5342, 
    35.54846, 35.55902, 35.56923, 35.58136, 35.59584, 35.60954, 35.62378,
  35.42323, 35.44531, 35.46241, 35.48072, 35.49038, 35.50944, 35.52764, 
    35.54381, 35.55697, 35.5667, 35.57595, 35.58776, 35.60247, 35.61756, 
    35.63175,
  35.42041, 35.43966, 35.44967, 35.46805, 35.49132, 35.51238, 35.53076, 
    35.54641, 35.56008, 35.56984, 35.57955, 35.59106, 35.60507, 35.61872, 
    35.63314,
  35.42367, 35.44001, 35.45217, 35.47351, 35.49572, 35.51443, 35.53144, 
    35.54628, 35.56041, 35.57281, 35.58309, 35.59278, 35.60363, 35.61634, 
    35.63113,
  35.42196, 35.44363, 35.46043, 35.48107, 35.50089, 35.51906, 35.53546, 
    35.54958, 35.5631, 35.57758, 35.58802, 35.59684, 35.60613, 35.61753, 
    35.6316,
  35.42967, 35.45213, 35.46773, 35.48634, 35.5055, 35.52557, 35.54339, 
    35.55652, 35.57038, 35.58306, 35.59304, 35.60112, 35.61046, 35.62202, 
    35.63549,
  35.44097, 35.46001, 35.47729, 35.49581, 35.51454, 35.53447, 35.55122, 
    35.56537, 35.57605, 35.58716, 35.59681, 35.6053, 35.61605, 35.62891, 
    35.64224,
  35.45854, 35.47688, 35.49408, 35.51107, 35.52793, 35.54575, 35.56142, 
    35.57247, 35.57911, 35.58813, 35.59776, 35.60812, 35.61985, 35.63283, 
    35.64795,
  35.46367, 35.47913, 35.49454, 35.51041, 35.52511, 35.53779, 35.54404, 
    35.55817, 35.57444, 35.58356, 35.59171, 35.60253, 35.6149, 35.625, 
    35.63302,
  35.46526, 35.48658, 35.50508, 35.52135, 35.5351, 35.54605, 35.55135, 
    35.56496, 35.57801, 35.58714, 35.59546, 35.6058, 35.61772, 35.62798, 
    35.63661,
  35.46383, 35.48794, 35.50554, 35.52269, 35.53536, 35.54178, 35.55716, 
    35.57193, 35.58513, 35.59415, 35.60211, 35.61179, 35.62382, 35.63439, 
    35.64422,
  35.4623, 35.48477, 35.50164, 35.51923, 35.52897, 35.54757, 35.56455, 
    35.57892, 35.59099, 35.59953, 35.60698, 35.61678, 35.62902, 35.64104, 
    35.65157,
  35.4649, 35.48375, 35.49405, 35.50994, 35.53181, 35.55028, 35.56694, 
    35.58159, 35.59473, 35.60525, 35.61419, 35.62429, 35.63596, 35.64648, 
    35.65704,
  35.47129, 35.4877, 35.49852, 35.51867, 35.53897, 35.55632, 35.57219, 
    35.58722, 35.60175, 35.61351, 35.62304, 35.63188, 35.64124, 35.65104, 
    35.66209,
  35.47478, 35.49442, 35.50984, 35.52837, 35.54671, 35.56364, 35.57985, 
    35.59502, 35.60872, 35.62126, 35.63101, 35.63919, 35.6487, 35.65894, 
    35.66998,
  35.48294, 35.50336, 35.51824, 35.53573, 35.55445, 35.57288, 35.58878, 
    35.60322, 35.61639, 35.62752, 35.6363, 35.64435, 35.65532, 35.66787, 
    35.67995,
  35.49294, 35.51126, 35.52752, 35.54615, 35.56522, 35.58351, 35.5987, 
    35.61309, 35.62428, 35.63486, 35.64303, 35.65252, 35.66538, 35.67977, 
    35.69238,
  35.50781, 35.5262, 35.54406, 35.56216, 35.57942, 35.59765, 35.61362, 
    35.62522, 35.63479, 35.64477, 35.65263, 35.66215, 35.67567, 35.68943, 
    35.70259,
  35.61591, 35.62823, 35.63593, 35.64046, 35.64555, 35.6553, 35.66605, 
    35.68121, 35.69635, 35.70611, 35.71249, 35.71703, 35.72203, 35.72918, 
    35.74265,
  35.60758, 35.61864, 35.6242, 35.62963, 35.63731, 35.64869, 35.65959, 
    35.67375, 35.68835, 35.70103, 35.71082, 35.71749, 35.72482, 35.73354, 
    35.74843,
  35.5928, 35.60505, 35.61435, 35.62479, 35.63669, 35.64672, 35.66137, 
    35.67566, 35.69138, 35.70538, 35.71632, 35.72566, 35.73658, 35.74806, 
    35.76314,
  35.59107, 35.60541, 35.61771, 35.63318, 35.64513, 35.65993, 35.67307, 
    35.68597, 35.70054, 35.71351, 35.7253, 35.73772, 35.75473, 35.771, 
    35.78662,
  35.60744, 35.62018, 35.63205, 35.64725, 35.66281, 35.67516, 35.68544, 
    35.69675, 35.71151, 35.72484, 35.73765, 35.75182, 35.7704, 35.78775, 
    35.80278,
  35.63252, 35.64525, 35.65531, 35.6689, 35.68135, 35.69183, 35.7007, 
    35.70928, 35.72142, 35.73416, 35.74863, 35.76547, 35.78383, 35.7989, 
    35.81183,
  35.65594, 35.6687, 35.67881, 35.69003, 35.70057, 35.71005, 35.71645, 
    35.72281, 35.73306, 35.7466, 35.76342, 35.78146, 35.79855, 35.81266, 
    35.82308,
  35.67915, 35.68884, 35.69681, 35.70649, 35.716, 35.72437, 35.72794, 
    35.73292, 35.74356, 35.75917, 35.77784, 35.79696, 35.81298, 35.82481, 
    35.83245,
  35.70298, 35.70962, 35.71702, 35.72618, 35.7348, 35.73997, 35.74075, 
    35.74635, 35.7584, 35.77603, 35.79522, 35.81397, 35.82784, 35.83566, 
    35.83949,
  35.72671, 35.73546, 35.74551, 35.75286, 35.75587, 35.75701, 35.75868, 
    35.76543, 35.77987, 35.79815, 35.81772, 35.8329, 35.84159, 35.84379, 
    35.84662,
  35.87261, 35.88245, 35.89123, 35.89799, 35.90428, 35.90997, 35.91418, 
    35.91978, 35.92666, 35.9332, 35.93613, 35.93682, 35.93798, 35.93755, 
    35.9336,
  35.87671, 35.88725, 35.89692, 35.90517, 35.9119, 35.91579, 35.91845, 
    35.92332, 35.93021, 35.93565, 35.93863, 35.94177, 35.94553, 35.94726, 
    35.94553,
  35.87537, 35.88596, 35.8961, 35.90672, 35.91527, 35.91993, 35.9237, 
    35.92741, 35.93311, 35.93828, 35.94358, 35.94973, 35.95598, 35.95996, 
    35.9599,
  35.87941, 35.88991, 35.89951, 35.90886, 35.91691, 35.92424, 35.929, 
    35.93354, 35.9385, 35.94421, 35.95116, 35.95942, 35.96664, 35.97158, 
    35.9729,
  35.88681, 35.89621, 35.90453, 35.9136, 35.92279, 35.93, 35.93439, 35.93827, 
    35.94281, 35.9486, 35.95637, 35.96579, 35.97359, 35.97867, 35.98034,
  35.89351, 35.90137, 35.90934, 35.91836, 35.92752, 35.9341, 35.93829, 
    35.94221, 35.94809, 35.95567, 35.96362, 35.97069, 35.9774, 35.98215, 
    35.98368,
  35.89652, 35.90358, 35.91104, 35.91903, 35.92752, 35.9337, 35.9386, 
    35.94377, 35.9517, 35.96061, 35.96827, 35.97434, 35.97924, 35.98267, 
    35.98404,
  35.90192, 35.90737, 35.91356, 35.92049, 35.92871, 35.93541, 35.94161, 
    35.94823, 35.95751, 35.96676, 35.97349, 35.97838, 35.98217, 35.98439, 
    35.9856,
  35.9049, 35.91131, 35.91867, 35.92707, 35.93651, 35.94493, 35.95135, 
    35.9585, 35.96803, 35.97548, 35.97986, 35.98295, 35.98581, 35.98762, 
    35.98897,
  35.9132, 35.92097, 35.93108, 35.94237, 35.95231, 35.95974, 35.96569, 
    35.9725, 35.9793, 35.98374, 35.98617, 35.98861, 35.99117, 35.9923, 
    35.99397,
  36.08649, 36.08541, 36.08355, 36.08089, 36.07905, 36.07779, 36.07631, 
    36.07544, 36.07571, 36.07628, 36.07699, 36.07733, 36.07734, 36.07651, 
    36.07449,
  36.08912, 36.08736, 36.08541, 36.08337, 36.08196, 36.08118, 36.08081, 
    36.08079, 36.08138, 36.08233, 36.08376, 36.08507, 36.08558, 36.0849, 
    36.08409,
  36.09042, 36.08922, 36.08792, 36.08643, 36.08562, 36.08601, 36.08627, 
    36.08658, 36.08708, 36.0882, 36.08979, 36.09104, 36.09166, 36.09196, 
    36.09288,
  36.09302, 36.09176, 36.0911, 36.09106, 36.09169, 36.09216, 36.09217, 
    36.09205, 36.09258, 36.09366, 36.09511, 36.0966, 36.09805, 36.09941, 
    36.10178,
  36.09854, 36.09698, 36.09615, 36.09592, 36.09602, 36.0965, 36.09705, 
    36.09766, 36.09899, 36.10091, 36.10296, 36.10491, 36.1069, 36.10922, 
    36.11218,
  36.10544, 36.10288, 36.10104, 36.10044, 36.10104, 36.10237, 36.10392, 
    36.10568, 36.10828, 36.11136, 36.11426, 36.11689, 36.11925, 36.12167, 
    36.12432,
  36.10839, 36.10747, 36.10637, 36.10623, 36.1077, 36.11036, 36.11358, 
    36.11731, 36.12169, 36.12606, 36.1295, 36.132, 36.134, 36.13544, 36.13628,
  36.1057, 36.10702, 36.10855, 36.11051, 36.11327, 36.117, 36.12123, 
    36.12653, 36.13217, 36.1371, 36.14038, 36.14245, 36.14377, 36.14467, 
    36.14518,
  36.10406, 36.1064, 36.10913, 36.11306, 36.11761, 36.12269, 36.12796, 
    36.13361, 36.13902, 36.14315, 36.14594, 36.14761, 36.14907, 36.15066, 
    36.15179,
  36.10365, 36.10722, 36.11144, 36.11653, 36.12208, 36.12749, 36.13289, 
    36.1376, 36.14206, 36.14595, 36.14874, 36.15118, 36.15359, 36.15616, 
    36.15803,
  36.24342, 36.24233, 36.23996, 36.23811, 36.23769, 36.23864, 36.23965, 
    36.24114, 36.2419, 36.24332, 36.24358, 36.24232, 36.23986, 36.23903, 
    36.23878,
  36.24905, 36.24865, 36.24831, 36.24835, 36.24966, 36.25127, 36.25268, 
    36.25323, 36.25302, 36.25283, 36.25172, 36.2515, 36.25144, 36.25085, 
    36.24983,
  36.25885, 36.25887, 36.25937, 36.26018, 36.26091, 36.26094, 36.26084, 
    36.25976, 36.2596, 36.25964, 36.26055, 36.26112, 36.26112, 36.26045, 
    36.25999,
  36.26834, 36.26795, 36.26782, 36.26765, 36.26717, 36.26713, 36.26698, 
    36.26711, 36.26752, 36.26838, 36.26923, 36.26926, 36.2694, 36.26921, 
    36.26859,
  36.27652, 36.27528, 36.2745, 36.27457, 36.27493, 36.2756, 36.27612, 
    36.27667, 36.27715, 36.27776, 36.27822, 36.27824, 36.27797, 36.27737, 
    36.27627,
  36.28183, 36.2821, 36.28276, 36.2837, 36.28444, 36.28548, 36.28643, 
    36.28731, 36.2881, 36.28875, 36.28885, 36.28831, 36.28736, 36.28617, 
    36.2849,
  36.28657, 36.28785, 36.28925, 36.29074, 36.2922, 36.29385, 36.29565, 
    36.29718, 36.29812, 36.29821, 36.29762, 36.29656, 36.29507, 36.29375, 
    36.29245,
  36.29065, 36.29196, 36.29353, 36.29548, 36.29772, 36.30013, 36.30235, 
    36.30381, 36.30435, 36.30417, 36.30327, 36.30197, 36.30065, 36.29939, 
    36.29853,
  36.2937, 36.29537, 36.29729, 36.29934, 36.30163, 36.30381, 36.30558, 
    36.30658, 36.30683, 36.30632, 36.30514, 36.30398, 36.30278, 36.30164, 
    36.30173,
  36.29692, 36.2983, 36.29993, 36.30168, 36.30327, 36.30453, 36.30547, 
    36.30627, 36.30679, 36.3066, 36.30581, 36.30482, 36.30415, 36.30472, 
    36.30479,
  36.32001, 36.3204, 36.32088, 36.3215, 36.3223, 36.32296, 36.3232, 36.32299, 
    36.32263, 36.32195, 36.32091, 36.31959, 36.31826, 36.31739, 36.31757,
  36.3333, 36.33434, 36.33526, 36.33599, 36.3364, 36.33624, 36.33559, 
    36.33473, 36.33386, 36.33305, 36.33215, 36.33116, 36.33015, 36.32979, 
    36.33075,
  36.34534, 36.34621, 36.34671, 36.34675, 36.34648, 36.34592, 36.34514, 
    36.34446, 36.34399, 36.34384, 36.34368, 36.34329, 36.34296, 36.34317, 
    36.34414,
  36.35593, 36.35616, 36.35616, 36.35592, 36.35552, 36.35503, 36.35458, 
    36.35431, 36.35434, 36.35459, 36.35476, 36.35476, 36.35462, 36.35459, 
    36.35498,
  36.36464, 36.36485, 36.36494, 36.3649, 36.36478, 36.36465, 36.36464, 
    36.36484, 36.36519, 36.36551, 36.36563, 36.36547, 36.36523, 36.36516, 
    36.36552,
  36.37172, 36.37238, 36.37295, 36.37347, 36.37394, 36.37439, 36.37486, 
    36.37539, 36.37584, 36.37605, 36.37601, 36.37581, 36.37577, 36.37606, 
    36.3768,
  36.37794, 36.37912, 36.3802, 36.38117, 36.38207, 36.38293, 36.38373, 
    36.3844, 36.38485, 36.38506, 36.38511, 36.38519, 36.38552, 36.38625, 
    36.38741,
  36.3834, 36.38468, 36.38596, 36.38722, 36.3884, 36.38953, 36.39051, 
    36.39127, 36.39178, 36.39216, 36.39256, 36.39315, 36.39398, 36.39508, 
    36.39642,
  36.38774, 36.38903, 36.3904, 36.39179, 36.39315, 36.39445, 36.39561, 
    36.39657, 36.39736, 36.39814, 36.39901, 36.40003, 36.40108, 36.4022, 
    36.40326,
  36.39085, 36.39209, 36.39338, 36.39471, 36.39606, 36.39743, 36.39878, 
    36.40007, 36.40133, 36.40253, 36.40369, 36.40487, 36.406, 36.4069, 
    36.40771,
  36.33389, 36.334, 36.33434, 36.33488, 36.33546, 36.33578, 36.33566, 
    36.33523, 36.33455, 36.3337, 36.33262, 36.33146, 36.3305, 36.33047, 
    36.33141,
  36.34822, 36.34874, 36.34911, 36.34922, 36.34895, 36.34832, 36.34742, 
    36.34641, 36.34532, 36.34431, 36.34338, 36.34251, 36.34203, 36.34261, 
    36.34424,
  36.35993, 36.36012, 36.35999, 36.35955, 36.35886, 36.35806, 36.35722, 
    36.35652, 36.356, 36.35563, 36.35515, 36.35468, 36.35473, 36.35557, 
    36.3569,
  36.36987, 36.36978, 36.36943, 36.36896, 36.36843, 36.36798, 36.36767, 
    36.36754, 36.36752, 36.36743, 36.36727, 36.36709, 36.36707, 36.36734, 
    36.36786,
  36.3788, 36.37879, 36.37865, 36.37848, 36.37836, 36.37835, 36.37849, 
    36.3787, 36.37886, 36.37887, 36.37872, 36.37848, 36.37832, 36.37837, 
    36.37858,
  36.387, 36.38716, 36.38727, 36.38742, 36.38765, 36.38799, 36.38839, 
    36.38874, 36.38894, 36.38891, 36.38865, 36.38838, 36.38826, 36.38842, 
    36.38906,
  36.39417, 36.39456, 36.39488, 36.39519, 36.39554, 36.39591, 36.39624, 
    36.39643, 36.39646, 36.39635, 36.39623, 36.39627, 36.39666, 36.39745, 
    36.39875,
  36.3995, 36.40005, 36.40057, 36.40107, 36.40155, 36.40201, 36.40238, 
    36.40263, 36.40281, 36.40302, 36.4034, 36.40408, 36.40509, 36.40639, 
    36.40794,
  36.40327, 36.40393, 36.40471, 36.40558, 36.40649, 36.40736, 36.40814, 
    36.40881, 36.40945, 36.41022, 36.41118, 36.41234, 36.4136, 36.41493, 
    36.41632,
  36.40588, 36.4067, 36.40775, 36.40899, 36.41034, 36.4117, 36.41299, 
    36.41419, 36.41537, 36.4166, 36.4179, 36.41921, 36.42048, 36.42168, 
    36.42284,
  36.27679, 36.27632, 36.27592, 36.2755, 36.27495, 36.27422, 36.27346, 
    36.27268, 36.27192, 36.2712, 36.27046, 36.26988, 36.26962, 36.26994, 
    36.27069,
  36.2877, 36.28706, 36.2863, 36.28542, 36.28443, 36.28346, 36.28248, 
    36.28166, 36.28099, 36.28043, 36.27993, 36.27957, 36.27971, 36.28054, 
    36.28163,
  36.29667, 36.29606, 36.2953, 36.29439, 36.29342, 36.29253, 36.29187, 
    36.29135, 36.29093, 36.29056, 36.29027, 36.2902, 36.29059, 36.29126, 
    36.29163,
  36.30551, 36.30498, 36.30433, 36.30367, 36.30305, 36.30255, 36.30219, 
    36.30191, 36.30164, 36.30142, 36.30133, 36.30129, 36.3012, 36.30099, 
    36.30062,
  36.3141, 36.31367, 36.31321, 36.31284, 36.31258, 36.31247, 36.31242, 
    36.31232, 36.31219, 36.31205, 36.31186, 36.31149, 36.31099, 36.31041, 
    36.30977,
  36.32233, 36.32183, 36.32139, 36.32103, 36.32074, 36.3205, 36.32026, 
    36.31998, 36.31969, 36.31925, 36.31871, 36.31829, 36.31778, 36.31739, 
    36.31732,
  36.32932, 36.32853, 36.32784, 36.32721, 36.32661, 36.32601, 36.32537, 
    36.32468, 36.32397, 36.3233, 36.32277, 36.32255, 36.32257, 36.32294, 
    36.32365,
  36.33437, 36.33346, 36.33258, 36.33174, 36.33096, 36.33016, 36.32937, 
    36.32863, 36.328, 36.32755, 36.3274, 36.32758, 36.32813, 36.32902, 
    36.33016,
  36.33766, 36.33694, 36.33624, 36.3356, 36.33504, 36.33451, 36.33404, 
    36.33369, 36.33354, 36.3336, 36.33391, 36.33449, 36.33531, 36.33628, 
    36.33736,
  36.34029, 36.33979, 36.33944, 36.33929, 36.33933, 36.33946, 36.33961, 
    36.33979, 36.34006, 36.34045, 36.34099, 36.34166, 36.34244, 36.34328, 
    36.3441,
  36.09129, 36.09025, 36.08921, 36.08807, 36.08679, 36.08544, 36.08415, 
    36.08301, 36.08207, 36.08132, 36.0808, 36.08047, 36.08046, 36.08087, 
    36.08149,
  36.0994, 36.09812, 36.09681, 36.09539, 36.09387, 36.09245, 36.09117, 
    36.09016, 36.08941, 36.08881, 36.08843, 36.0882, 36.08822, 36.08855, 
    36.08905,
  36.10646, 36.10527, 36.10397, 36.10262, 36.10131, 36.10011, 36.09904, 
    36.09821, 36.09752, 36.09691, 36.09634, 36.09597, 36.09594, 36.09612, 
    36.09618,
  36.11314, 36.11198, 36.11072, 36.10948, 36.10832, 36.10734, 36.10653, 
    36.10578, 36.10508, 36.10443, 36.104, 36.10375, 36.10355, 36.10329, 
    36.10272,
  36.11908, 36.11782, 36.11657, 36.1154, 36.11431, 36.11335, 36.11251, 
    36.1118, 36.11122, 36.11074, 36.11032, 36.10993, 36.10945, 36.10865, 
    36.10765,
  36.12434, 36.12278, 36.1213, 36.11992, 36.11866, 36.1175, 36.11634, 
    36.11525, 36.11434, 36.11347, 36.11258, 36.11168, 36.11082, 36.11001, 
    36.10918,
  36.12823, 36.12624, 36.12438, 36.12262, 36.12094, 36.11929, 36.11765, 
    36.11602, 36.11449, 36.11316, 36.11201, 36.11104, 36.11023, 36.10966, 
    36.10929,
  36.13068, 36.12828, 36.12599, 36.1238, 36.12166, 36.11958, 36.11759, 
    36.11572, 36.11404, 36.11261, 36.11141, 36.11049, 36.10983, 36.10946, 
    36.10939,
  36.13213, 36.1296, 36.12719, 36.12485, 36.12255, 36.12035, 36.1183, 
    36.11645, 36.11483, 36.11347, 36.11243, 36.11173, 36.11142, 36.11138, 
    36.11154,
  36.13384, 36.1313, 36.1289, 36.12659, 36.12447, 36.12254, 36.12081, 
    36.11928, 36.11797, 36.11689, 36.11612, 36.11565, 36.11543, 36.11544, 
    36.11559,
  35.84835, 35.84627, 35.84442, 35.84262, 35.84058, 35.83823, 35.8357, 
    35.8332, 35.8308, 35.82863, 35.82678, 35.82533, 35.8245, 35.82428, 
    35.82453,
  35.85585, 35.85389, 35.85178, 35.84945, 35.84692, 35.84431, 35.84173, 
    35.83928, 35.837, 35.83497, 35.83329, 35.83195, 35.83107, 35.83069, 
    35.83067,
  35.86289, 35.86059, 35.85814, 35.85558, 35.85296, 35.85037, 35.84782, 
    35.84542, 35.84332, 35.84137, 35.83971, 35.83834, 35.83731, 35.83665, 
    35.8363,
  35.86813, 35.86557, 35.86289, 35.86016, 35.85747, 35.85488, 35.85247, 
    35.85025, 35.84822, 35.8463, 35.84457, 35.84315, 35.84205, 35.84138, 
    35.84066,
  35.87239, 35.86959, 35.86679, 35.86404, 35.86135, 35.85872, 35.8562, 
    35.85382, 35.85154, 35.84944, 35.84764, 35.84618, 35.84499, 35.8438, 
    35.8425,
  35.87637, 35.87308, 35.86992, 35.86689, 35.86401, 35.86121, 35.85849, 
    35.8558, 35.85317, 35.85068, 35.84842, 35.84638, 35.84454, 35.84282, 
    35.84115,
  35.87927, 35.87548, 35.87186, 35.86839, 35.86501, 35.86168, 35.85839, 
    35.85518, 35.8521, 35.84921, 35.84657, 35.84418, 35.84204, 35.84011, 
    35.83838,
  35.88031, 35.87614, 35.87222, 35.86835, 35.86453, 35.86078, 35.85707, 
    35.85349, 35.85013, 35.84701, 35.84415, 35.84159, 35.83932, 35.83733, 
    35.8356,
  35.88014, 35.87588, 35.87178, 35.86775, 35.86375, 35.8598, 35.85594, 
    35.85225, 35.8488, 35.84561, 35.8427, 35.84009, 35.83781, 35.8359, 
    35.83432,
  35.8801, 35.87579, 35.87164, 35.86758, 35.86357, 35.85966, 35.85593, 
    35.85242, 35.84915, 35.8461, 35.84332, 35.84091, 35.83887, 35.8372, 
    35.83581,
  35.60096, 35.5981, 35.59537, 35.5928, 35.59027, 35.58757, 35.58463, 
    35.58142, 35.57809, 35.57474, 35.57158, 35.56875, 35.56641, 35.56466, 
    35.56369,
  35.60706, 35.60444, 35.60178, 35.599, 35.59605, 35.59284, 35.58948, 
    35.58604, 35.58266, 35.57937, 35.57631, 35.5736, 35.5714, 35.56974, 
    35.5687,
  35.61383, 35.61084, 35.60768, 35.60437, 35.60099, 35.59759, 35.59419, 
    35.59083, 35.58754, 35.58437, 35.58144, 35.57888, 35.57671, 35.57492, 
    35.57363,
  35.61986, 35.61636, 35.61272, 35.60907, 35.60543, 35.60183, 35.59829, 
    35.59485, 35.59153, 35.58838, 35.58547, 35.58286, 35.58054, 35.57857, 
    35.57695,
  35.62538, 35.6213, 35.61718, 35.61314, 35.60924, 35.60548, 35.60183, 
    35.59825, 35.59474, 35.59137, 35.58823, 35.58536, 35.58276, 35.58042, 
    35.57835,
  35.63127, 35.62654, 35.62185, 35.61731, 35.61298, 35.60886, 35.60482, 
    35.60082, 35.59692, 35.59319, 35.58969, 35.58644, 35.58347, 35.58072, 
    35.57824,
  35.63669, 35.63144, 35.6263, 35.62135, 35.61662, 35.612, 35.6074, 35.6029, 
    35.59853, 35.59431, 35.59027, 35.58649, 35.58303, 35.57991, 35.57711,
  35.64036, 35.63477, 35.62939, 35.62423, 35.61915, 35.61407, 35.60905, 
    35.60416, 35.59943, 35.59486, 35.59051, 35.58643, 35.58267, 35.57924, 
    35.57615,
  35.64198, 35.63636, 35.63092, 35.62559, 35.62024, 35.61497, 35.60977, 
    35.60472, 35.59986, 35.5952, 35.59076, 35.5866, 35.58273, 35.57919, 
    35.57602,
  35.64274, 35.6372, 35.63179, 35.62644, 35.62111, 35.6158, 35.61059, 
    35.60556, 35.60072, 35.59609, 35.59169, 35.5876, 35.58389, 35.58055, 
    35.57762,
  35.4043, 35.40101, 35.39772, 35.39449, 35.39143, 35.38848, 35.38556, 
    35.38259, 35.37946, 35.37623, 35.37303, 35.36997, 35.36719, 35.36478, 
    35.36279,
  35.40738, 35.40409, 35.40082, 35.39758, 35.39438, 35.39119, 35.38797, 
    35.38469, 35.38135, 35.37802, 35.37479, 35.37173, 35.36898, 35.36663, 
    35.36473,
  35.41187, 35.40844, 35.40495, 35.40141, 35.39786, 35.3943, 35.39075, 
    35.38725, 35.38379, 35.38044, 35.37724, 35.37425, 35.37159, 35.36937, 
    35.36761,
  35.4174, 35.41359, 35.40964, 35.40563, 35.40167, 35.39779, 35.39397, 
    35.39029, 35.38674, 35.38337, 35.38019, 35.37724, 35.37458, 35.37231, 
    35.37044,
  35.42424, 35.41993, 35.41544, 35.41091, 35.40643, 35.40208, 35.39791, 
    35.39394, 35.39019, 35.38662, 35.3832, 35.38003, 35.37716, 35.3746, 
    35.37233,
  35.43226, 35.42747, 35.42246, 35.41738, 35.41236, 35.4075, 35.40285, 
    35.39843, 35.39421, 35.39014, 35.38631, 35.38272, 35.37942, 35.37639, 
    35.37366,
  35.44016, 35.43493, 35.42948, 35.42396, 35.41851, 35.41322, 35.4081, 
    35.40314, 35.39839, 35.39384, 35.38952, 35.38546, 35.38168, 35.3782, 
    35.37509,
  35.4465, 35.44093, 35.4352, 35.42944, 35.42374, 35.41811, 35.41258, 
    35.40721, 35.40205, 35.39709, 35.39238, 35.38796, 35.3839, 35.38021, 
    35.37691,
  35.45059, 35.44487, 35.43905, 35.43323, 35.42736, 35.42148, 35.41568, 
    35.41004, 35.40461, 35.39943, 35.39454, 35.39002, 35.38587, 35.38208, 
    35.37864,
  35.45336, 35.44761, 35.44179, 35.43594, 35.43003, 35.42406, 35.41813, 
    35.41236, 35.40685, 35.40163, 35.39674, 35.39217, 35.38795, 35.3841, 
    35.38065,
  35.26357, 35.26066, 35.25769, 35.25474, 35.25188, 35.24913, 35.24646, 
    35.24381, 35.24107, 35.23821, 35.23534, 35.23258, 35.23, 35.22763, 
    35.22549,
  35.26489, 35.26182, 35.25878, 35.25581, 35.25293, 35.25011, 35.24732, 
    35.2445, 35.24162, 35.2387, 35.23581, 35.23302, 35.2304, 35.228, 35.22586,
  35.26701, 35.26387, 35.26076, 35.2577, 35.25469, 35.2517, 35.24871, 
    35.24571, 35.24271, 35.23974, 35.23685, 35.23407, 35.23146, 35.22905, 
    35.22692,
  35.27023, 35.26691, 35.2636, 35.26031, 35.25706, 35.25385, 35.25067, 
    35.24752, 35.24443, 35.24141, 35.23851, 35.23576, 35.23315, 35.23075, 
    35.22864,
  35.27512, 35.27151, 35.26785, 35.2642, 35.26058, 35.25703, 35.25357, 
    35.25021, 35.24696, 35.24382, 35.24081, 35.23796, 35.23532, 35.23287, 
    35.23064,
  35.28146, 35.2775, 35.27343, 35.26931, 35.26523, 35.26123, 35.25736, 
    35.25365, 35.25012, 35.24675, 35.24357, 35.24057, 35.23774, 35.2351, 
    35.23264,
  35.28828, 35.28398, 35.27952, 35.27498, 35.27045, 35.26598, 35.26164, 
    35.25753, 35.25364, 35.24996, 35.2465, 35.24326, 35.24021, 35.23736, 
    35.23473,
  35.2945, 35.28992, 35.28518, 35.28033, 35.27543, 35.27057, 35.26585, 
    35.26134, 35.25708, 35.25305, 35.24926, 35.24574, 35.2425, 35.23954, 
    35.23685,
  35.29957, 35.29477, 35.28982, 35.28478, 35.27967, 35.27454, 35.26952, 
    35.26472, 35.26018, 35.25586, 35.25182, 35.24813, 35.24477, 35.24173, 
    35.23898,
  35.30379, 35.29886, 35.29376, 35.2886, 35.28335, 35.27806, 35.27285, 
    35.26785, 35.2631, 35.25863, 35.25449, 35.25071, 35.24725, 35.24409, 
    35.24122,
  35.15041, 35.148, 35.14554, 35.14307, 35.14067, 35.13835, 35.13613, 
    35.13394, 35.13169, 35.12929, 35.12679, 35.12434, 35.12205, 35.11995, 
    35.118,
  35.1521, 35.14947, 35.14686, 35.14433, 35.14189, 35.13955, 35.13727, 
    35.13494, 35.1325, 35.12999, 35.12746, 35.12499, 35.12265, 35.12047, 
    35.11847,
  35.15429, 35.15156, 35.14889, 35.14632, 35.14385, 35.14144, 35.13904, 
    35.1366, 35.13409, 35.13155, 35.12905, 35.1266, 35.12424, 35.12199, 
    35.1199,
  35.15734, 35.15449, 35.1517, 35.149, 35.14639, 35.14386, 35.14137, 35.1389, 
    35.13642, 35.13394, 35.13147, 35.12904, 35.12662, 35.12429, 35.12213,
  35.16171, 35.15868, 35.15568, 35.15273, 35.14988, 35.14711, 35.14444, 
    35.14182, 35.13926, 35.13671, 35.1342, 35.13173, 35.12933, 35.12701, 
    35.12482,
  35.16723, 35.16402, 35.16076, 35.15751, 35.15432, 35.15119, 35.14817, 
    35.14526, 35.14246, 35.13972, 35.13707, 35.13449, 35.13204, 35.12971, 
    35.12753,
  35.17321, 35.16982, 35.16632, 35.16279, 35.15926, 35.15575, 35.15232, 
    35.14905, 35.1459, 35.14288, 35.13999, 35.13726, 35.1347, 35.13231, 
    35.13004,
  35.17874, 35.17519, 35.17152, 35.1678, 35.16402, 35.16022, 35.15648, 
    35.15287, 35.1494, 35.14606, 35.1429, 35.13994, 35.1372, 35.13467, 
    35.13234,
  35.18356, 35.17986, 35.17604, 35.17218, 35.16825, 35.16426, 35.16029, 
    35.15644, 35.15275, 35.1492, 35.14585, 35.14274, 35.13987, 35.13726, 
    35.1349,
  35.18786, 35.18403, 35.1801, 35.17613, 35.17208, 35.16795, 35.16383, 
    35.15985, 35.15605, 35.15243, 35.14901, 35.14585, 35.14295, 35.14029, 
    35.13783,
  35.05313, 35.05111, 35.04909, 35.0471, 35.04518, 35.04334, 35.0416, 
    35.03996, 35.03837, 35.03674, 35.035, 35.0331, 35.03117, 35.02934, 
    35.02765,
  35.05491, 35.05264, 35.0504, 35.04825, 35.04623, 35.04434, 35.04261, 
    35.04096, 35.03928, 35.03752, 35.03563, 35.03367, 35.03174, 35.02992, 
    35.02824,
  35.05722, 35.05478, 35.05241, 35.05016, 35.04807, 35.04615, 35.04434, 
    35.04259, 35.04084, 35.03905, 35.03722, 35.03538, 35.03357, 35.03175, 
    35.03,
  35.06039, 35.05782, 35.05531, 35.05294, 35.05072, 35.04866, 35.04673, 
    35.04489, 35.04313, 35.04142, 35.03974, 35.03808, 35.03639, 35.03464, 
    35.03285,
  35.06486, 35.06215, 35.05949, 35.05693, 35.05449, 35.05218, 35.05001, 
    35.048, 35.04614, 35.0444, 35.04275, 35.04113, 35.0395, 35.03782, 35.03613,
  35.07059, 35.06779, 35.06498, 35.0622, 35.05948, 35.05685, 35.05437, 
    35.05207, 35.04994, 35.04797, 35.04612, 35.04431, 35.04254, 35.04084, 
    35.03925,
  35.07682, 35.07398, 35.07106, 35.06813, 35.06522, 35.06234, 35.05955, 
    35.05693, 35.05446, 35.05213, 35.04991, 35.04779, 35.04579, 35.04397, 
    35.0423,
  35.08284, 35.07997, 35.07699, 35.07398, 35.07094, 35.06788, 35.06488, 
    35.06199, 35.05923, 35.05655, 35.05396, 35.0515, 35.04922, 35.04715, 
    35.04525,
  35.08847, 35.08555, 35.08251, 35.07943, 35.07631, 35.07314, 35.06997, 
    35.06688, 35.06389, 35.06095, 35.05811, 35.05542, 35.05293, 35.05066, 
    35.04862,
  35.09382, 35.09085, 35.08775, 35.0846, 35.08141, 35.07813, 35.07481, 
    35.07155, 35.06839, 35.06531, 35.06236, 35.05959, 35.05705, 35.05476, 
    35.0527,
  34.97135, 34.96986, 34.96836, 34.96688, 34.96545, 34.96408, 34.96278, 
    34.96153, 34.96037, 34.95928, 34.95816, 34.95691, 34.9555, 34.95393, 
    34.95234,
  34.97268, 34.97094, 34.96924, 34.96761, 34.96606, 34.96462, 34.96329, 
    34.96208, 34.96097, 34.95989, 34.95877, 34.95754, 34.95616, 34.95465, 
    34.95312,
  34.97462, 34.97268, 34.97079, 34.969, 34.96733, 34.96581, 34.96444, 
    34.9632, 34.96205, 34.96097, 34.95992, 34.95884, 34.95768, 34.95638, 
    34.955,
  34.97731, 34.97517, 34.97312, 34.97118, 34.96939, 34.96775, 34.96626, 
    34.96489, 34.96365, 34.96257, 34.96163, 34.96078, 34.95988, 34.95889, 
    34.9577,
  34.98126, 34.97898, 34.97677, 34.97467, 34.97269, 34.97084, 34.96914, 
    34.96756, 34.96619, 34.96504, 34.9641, 34.96331, 34.96251, 34.96163, 
    34.96059,
  34.98651, 34.98415, 34.98183, 34.97958, 34.97742, 34.97535, 34.97339, 
    34.97158, 34.96997, 34.96862, 34.96749, 34.9665, 34.96552, 34.96454, 
    34.9636,
  34.99223, 34.98985, 34.98746, 34.98512, 34.98283, 34.98061, 34.97846, 
    34.97647, 34.97466, 34.97306, 34.97163, 34.97029, 34.96901, 34.9678, 
    34.96672,
  34.99798, 34.99559, 34.99316, 34.99076, 34.98839, 34.98606, 34.9838, 
    34.9817, 34.97976, 34.97794, 34.97622, 34.97455, 34.97294, 34.97146, 
    34.97015,
  35.00368, 35.00129, 34.99883, 34.99637, 34.99395, 34.99154, 34.98919, 
    34.98698, 34.9849, 34.98289, 34.98092, 34.97899, 34.97715, 34.97546, 
    34.97396,
  35.00943, 35.00706, 35.00461, 35.00214, 34.99968, 34.99719, 34.99472, 
    34.99236, 34.9901, 34.98788, 34.98571, 34.98363, 34.9817, 34.97998, 
    34.97852,
  34.90573, 34.90471, 34.90364, 34.90255, 34.90145, 34.90036, 34.89927, 
    34.89816, 34.89704, 34.896, 34.89505, 34.89414, 34.89315, 34.892, 34.89065,
  34.90704, 34.90582, 34.90457, 34.90333, 34.90212, 34.90094, 34.89978, 
    34.89865, 34.89758, 34.89661, 34.89573, 34.89486, 34.89394, 34.89288, 
    34.89163,
  34.90863, 34.90724, 34.90585, 34.90448, 34.90316, 34.9019, 34.90071, 
    34.89961, 34.89857, 34.89764, 34.89679, 34.89599, 34.89522, 34.89436, 
    34.89336,
  34.91069, 34.90915, 34.90763, 34.90616, 34.90478, 34.90348, 34.90226, 
    34.90111, 34.90004, 34.89907, 34.89825, 34.89757, 34.89699, 34.89639, 
    34.89565,
  34.91372, 34.91211, 34.91051, 34.90897, 34.90749, 34.9061, 34.90476, 
    34.90349, 34.90231, 34.90128, 34.90047, 34.89985, 34.89932, 34.8988, 
    34.89819,
  34.91777, 34.91612, 34.91449, 34.91291, 34.91139, 34.90992, 34.90849, 
    34.9071, 34.9058, 34.90469, 34.9038, 34.90308, 34.90245, 34.9018, 34.90111,
  34.92236, 34.92069, 34.91903, 34.91742, 34.91588, 34.91436, 34.91288, 
    34.91144, 34.91011, 34.90895, 34.90797, 34.90709, 34.9062, 34.90531, 
    34.90443,
  34.9272, 34.92548, 34.92378, 34.92213, 34.92054, 34.91899, 34.91747, 
    34.91604, 34.91474, 34.91357, 34.91251, 34.91147, 34.91039, 34.90928, 
    34.90824,
  34.93225, 34.93048, 34.92874, 34.92703, 34.92539, 34.92379, 34.92223, 
    34.92079, 34.91948, 34.91829, 34.91714, 34.91596, 34.91473, 34.9135, 
    34.91237,
  34.93747, 34.9357, 34.93395, 34.93224, 34.93059, 34.92895, 34.92736, 
    34.92588, 34.92451, 34.92323, 34.92196, 34.92065, 34.91932, 34.91805, 
    34.91695,
  34.84925, 34.84875, 34.84822, 34.84767, 34.84711, 34.84656, 34.84601, 
    34.84544, 34.84483, 34.84421, 34.84363, 34.84312, 34.84267, 34.84219, 
    34.84155,
  34.85178, 34.85111, 34.85038, 34.84963, 34.84889, 34.84816, 34.84744, 
    34.84673, 34.84601, 34.84531, 34.84468, 34.84414, 34.84364, 34.84315, 
    34.84255,
  34.85448, 34.85366, 34.85278, 34.85186, 34.85096, 34.85009, 34.84924, 
    34.84842, 34.84762, 34.84687, 34.84618, 34.84557, 34.84504, 34.84457, 
    34.84406,
  34.85732, 34.85641, 34.85541, 34.85437, 34.85336, 34.85239, 34.85145, 
    34.85054, 34.84966, 34.84883, 34.84807, 34.84742, 34.84689, 34.84644, 
    34.84599,
  34.86052, 34.85957, 34.85852, 34.85743, 34.85636, 34.85533, 34.85433, 
    34.85335, 34.85238, 34.85146, 34.85063, 34.84993, 34.84936, 34.84888, 
    34.84841,
  34.86415, 34.86319, 34.86213, 34.86104, 34.85998, 34.85895, 34.85794, 
    34.85693, 34.85592, 34.85495, 34.85407, 34.85332, 34.85267, 34.85208, 
    34.85145,
  34.86801, 34.86702, 34.86597, 34.8649, 34.86387, 34.86287, 34.86188, 
    34.8609, 34.85993, 34.859, 34.85816, 34.85739, 34.85663, 34.85583, 34.855,
  34.87198, 34.87096, 34.8699, 34.86884, 34.86782, 34.86683, 34.86587, 
    34.86493, 34.86404, 34.86321, 34.86245, 34.86168, 34.86086, 34.85995, 
    34.85899,
  34.87611, 34.87506, 34.87399, 34.87294, 34.87192, 34.87093, 34.86997, 
    34.86906, 34.86823, 34.86747, 34.86676, 34.86601, 34.86515, 34.8642, 
    34.86322,
  34.88044, 34.87938, 34.87832, 34.8773, 34.87632, 34.87537, 34.87443, 
    34.87355, 34.87275, 34.87202, 34.87132, 34.87055, 34.86968, 34.86871, 
    34.86775,
  34.79794, 34.79773, 34.79755, 34.79738, 34.79722, 34.79708, 34.79701, 
    34.79696, 34.79688, 34.79678, 34.79669, 34.79662, 34.79663, 34.79679, 
    34.7971,
  34.80126, 34.801, 34.80076, 34.80051, 34.80026, 34.80003, 34.79985, 
    34.79969, 34.79951, 34.79935, 34.79924, 34.79918, 34.79917, 34.79927, 
    34.79949,
  34.80472, 34.80445, 34.80417, 34.80385, 34.80352, 34.80321, 34.80294, 
    34.80269, 34.80244, 34.80222, 34.80207, 34.80199, 34.80196, 34.802, 
    34.80214,
  34.8083, 34.80802, 34.8077, 34.80733, 34.80694, 34.80657, 34.80624, 
    34.80593, 34.80562, 34.80535, 34.80515, 34.80502, 34.80495, 34.80494, 
    34.80499,
  34.8121, 34.81183, 34.8115, 34.81109, 34.81067, 34.81027, 34.80992, 
    34.80958, 34.80924, 34.80893, 34.80867, 34.80849, 34.80836, 34.80827, 
    34.8082,
  34.81616, 34.8159, 34.81557, 34.81516, 34.81473, 34.81434, 34.814, 
    34.81368, 34.81335, 34.81303, 34.81276, 34.81255, 34.81236, 34.81216, 
    34.8119,
  34.82037, 34.82011, 34.81977, 34.81936, 34.81893, 34.81854, 34.81821, 
    34.81792, 34.81763, 34.81736, 34.81713, 34.81694, 34.81672, 34.8164, 
    34.81597,
  34.82462, 34.82433, 34.82399, 34.82357, 34.82315, 34.82275, 34.8224, 
    34.82211, 34.82186, 34.82165, 34.82148, 34.82132, 34.82106, 34.82067, 
    34.82015,
  34.82886, 34.82855, 34.8282, 34.82779, 34.82738, 34.82698, 34.82662, 
    34.82631, 34.82605, 34.82587, 34.82573, 34.82556, 34.82529, 34.82487, 
    34.82433,
  34.83308, 34.83276, 34.83242, 34.83204, 34.83167, 34.83131, 34.83096, 
    34.83064, 34.83039, 34.8302, 34.83005, 34.82987, 34.82958, 34.82915, 
    34.82863,
  34.74962, 34.74927, 34.74894, 34.74861, 34.74826, 34.74793, 34.74768, 
    34.7475, 34.74732, 34.74717, 34.74709, 34.74706, 34.74709, 34.74728, 
    34.74789,
  34.75447, 34.75415, 34.75385, 34.75352, 34.75317, 34.75282, 34.75254, 
    34.7523, 34.75205, 34.75183, 34.75169, 34.75162, 34.75161, 34.75171, 
    34.75214,
  34.7591, 34.75886, 34.75864, 34.7584, 34.75809, 34.75778, 34.75751, 
    34.75728, 34.75702, 34.75679, 34.75664, 34.75655, 34.75651, 34.75653, 
    34.75681,
  34.7635, 34.76335, 34.76326, 34.76311, 34.76289, 34.76264, 34.76244, 
    34.76226, 34.76208, 34.76191, 34.76178, 34.76171, 34.76166, 34.76163, 
    34.76177,
  34.76779, 34.76775, 34.76777, 34.76773, 34.76761, 34.76745, 34.76736, 
    34.76729, 34.76722, 34.76716, 34.76712, 34.76712, 34.76711, 34.76708, 
    34.76709,
  34.7721, 34.77215, 34.77223, 34.77229, 34.77229, 34.77225, 34.77227, 
    34.77233, 34.7724, 34.77249, 34.77261, 34.77275, 34.77285, 34.77287, 
    34.77279,
  34.77643, 34.77652, 34.77665, 34.77676, 34.77686, 34.77694, 34.77706, 
    34.77723, 34.77743, 34.77766, 34.77796, 34.7783, 34.77856, 34.77866, 
    34.77859,
  34.78075, 34.78087, 34.78103, 34.78119, 34.78134, 34.78149, 34.78169, 
    34.78193, 34.78222, 34.78257, 34.783, 34.78349, 34.78388, 34.78408, 
    34.78407,
  34.7851, 34.78523, 34.78542, 34.78563, 34.78583, 34.78603, 34.78627, 
    34.78655, 34.78688, 34.78729, 34.7878, 34.78834, 34.78879, 34.78907, 
    34.78915,
  34.78952, 34.78965, 34.78986, 34.79012, 34.79038, 34.79064, 34.79092, 
    34.79122, 34.79157, 34.79201, 34.79254, 34.79309, 34.79358, 34.7939, 
    34.79407,
  34.70416, 34.70354, 34.703, 34.70254, 34.7021, 34.70167, 34.70133, 34.7011, 
    34.7009, 34.70073, 34.70066, 34.70071, 34.70087, 34.70113, 34.70169,
  34.70859, 34.70803, 34.70757, 34.70718, 34.7068, 34.70641, 34.7061, 
    34.70588, 34.70567, 34.70549, 34.70539, 34.70542, 34.70555, 34.70576, 
    34.70621,
  34.71302, 34.71257, 34.71224, 34.71201, 34.71174, 34.71144, 34.71119, 
    34.71101, 34.71085, 34.7107, 34.71063, 34.71067, 34.71078, 34.71094, 
    34.71128,
  34.71751, 34.71722, 34.71705, 34.71698, 34.71685, 34.71666, 34.7165, 
    34.71641, 34.71634, 34.71629, 34.71629, 34.71638, 34.7165, 34.71662, 
    34.71684,
  34.72217, 34.72202, 34.72202, 34.72208, 34.72211, 34.72204, 34.72202, 
    34.72204, 34.72211, 34.72219, 34.72232, 34.72252, 34.72269, 34.72282, 
    34.72295,
  34.72703, 34.72699, 34.72711, 34.7273, 34.72744, 34.72755, 34.72766, 
    34.72783, 34.72803, 34.72826, 34.72857, 34.72892, 34.72924, 34.72945, 
    34.72955,
  34.73206, 34.73211, 34.7323, 34.73257, 34.73283, 34.73306, 34.73331, 
    34.7336, 34.73392, 34.73429, 34.73475, 34.73528, 34.73578, 34.73612, 
    34.73628,
  34.73717, 34.73729, 34.73755, 34.73788, 34.73823, 34.73857, 34.73891, 
    34.73929, 34.7397, 34.74017, 34.74075, 34.74141, 34.74203, 34.74249, 
    34.74275,
  34.74232, 34.74248, 34.74279, 34.74319, 34.74362, 34.74406, 34.74448, 
    34.74493, 34.74539, 34.74592, 34.74656, 34.74729, 34.74797, 34.7485, 
    34.74887,
  34.7475, 34.74768, 34.74803, 34.74849, 34.74899, 34.74951, 34.75002, 
    34.75051, 34.75103, 34.75161, 34.75228, 34.75303, 34.75375, 34.75436, 
    34.75481,
  34.67008, 34.66946, 34.66888, 34.66833, 34.66774, 34.66708, 34.66645, 
    34.66589, 34.66536, 34.66485, 34.6644, 34.66408, 34.6639, 34.66388, 
    34.66407,
  34.67577, 34.67516, 34.67461, 34.67409, 34.67354, 34.67293, 34.67233, 
    34.67177, 34.67125, 34.67073, 34.67027, 34.66991, 34.66968, 34.66957, 
    34.66965,
  34.68106, 34.6805, 34.68002, 34.67959, 34.67915, 34.67865, 34.67813, 
    34.67764, 34.67716, 34.6767, 34.67628, 34.67596, 34.67572, 34.67556, 
    34.67553,
  34.68602, 34.68554, 34.68516, 34.68484, 34.68454, 34.68416, 34.68374, 
    34.68335, 34.68296, 34.6826, 34.68229, 34.68206, 34.68187, 34.6817, 
    34.68158,
  34.69071, 34.69033, 34.69003, 34.68983, 34.68963, 34.68938, 34.68909, 
    34.68881, 34.68856, 34.68834, 34.68818, 34.68809, 34.68801, 34.68792, 
    34.68781,
  34.69527, 34.69493, 34.69468, 34.69456, 34.69445, 34.69432, 34.69415, 
    34.69402, 34.6939, 34.69384, 34.69385, 34.69394, 34.69405, 34.69411, 
    34.6941,
  34.69973, 34.69938, 34.69917, 34.69908, 34.69905, 34.69901, 34.69897, 
    34.69897, 34.69899, 34.69907, 34.69923, 34.6995, 34.69982, 34.70007, 
    34.7002,
  34.70409, 34.70374, 34.70353, 34.70348, 34.70351, 34.70355, 34.70363, 
    34.70375, 34.7039, 34.70409, 34.70438, 34.70479, 34.70525, 34.70565, 
    34.70593,
  34.70836, 34.70801, 34.70782, 34.7078, 34.70789, 34.70803, 34.70821, 
    34.70844, 34.70869, 34.70898, 34.70937, 34.70987, 34.71043, 34.71092, 
    34.7113,
  34.71257, 34.71224, 34.71209, 34.71211, 34.71227, 34.71251, 34.7128, 
    34.71312, 34.71347, 34.71385, 34.71431, 34.71488, 34.71549, 34.71607, 
    34.71656,
  34.63477, 34.63394, 34.63317, 34.63245, 34.63173, 34.63092, 34.6301, 
    34.62941, 34.62883, 34.6283, 34.62786, 34.62754, 34.62737, 34.62737, 
    34.62753,
  34.64103, 34.64021, 34.63944, 34.63873, 34.638, 34.63721, 34.63642, 
    34.63571, 34.63509, 34.63452, 34.63403, 34.63367, 34.63342, 34.63331, 
    34.63335,
  34.64706, 34.64625, 34.64552, 34.64486, 34.64422, 34.64351, 34.64278, 
    34.64211, 34.64151, 34.64095, 34.64047, 34.64011, 34.63984, 34.63967, 
    34.63959,
  34.65287, 34.65212, 34.65147, 34.65093, 34.6504, 34.6498, 34.64917, 
    34.64855, 34.64799, 34.64747, 34.64703, 34.64671, 34.64648, 34.64629, 
    34.64614,
  34.65851, 34.65786, 34.65733, 34.6569, 34.65647, 34.65597, 34.65543, 
    34.65488, 34.65437, 34.65392, 34.65356, 34.65332, 34.65316, 34.65302, 
    34.65287,
  34.66402, 34.66348, 34.66304, 34.66267, 34.66232, 34.66192, 34.66146, 
    34.66099, 34.66055, 34.66016, 34.65989, 34.65975, 34.65971, 34.65969, 
    34.65963,
  34.66946, 34.66896, 34.66856, 34.66823, 34.66793, 34.66761, 34.66724, 
    34.66686, 34.66649, 34.66617, 34.66597, 34.66593, 34.66602, 34.66614, 
    34.66621,
  34.67474, 34.67425, 34.67385, 34.67353, 34.67327, 34.67302, 34.67275, 
    34.67245, 34.67218, 34.67193, 34.6718, 34.67184, 34.67202, 34.67224, 
    34.6724,
  34.67969, 34.67921, 34.6788, 34.6785, 34.67828, 34.67809, 34.67791, 
    34.67773, 34.67754, 34.67739, 34.67733, 34.67744, 34.67767, 34.67794, 
    34.67815,
  34.68427, 34.6838, 34.68341, 34.68314, 34.68296, 34.68284, 34.68275, 
    34.68266, 34.68259, 34.68254, 34.68257, 34.68274, 34.68301, 34.68331, 
    34.68358,
  34.61554, 34.61493, 34.61435, 34.61383, 34.61336, 34.61288, 34.61242, 
    34.61205, 34.61178, 34.61156, 34.61139, 34.61132, 34.61137, 34.61155, 
    34.61189,
  34.6208, 34.62019, 34.61961, 34.6191, 34.61863, 34.61814, 34.61769, 
    34.61731, 34.61703, 34.6168, 34.61663, 34.61657, 34.6166, 34.61674, 34.617,
  34.62593, 34.62529, 34.62472, 34.62423, 34.6238, 34.62337, 34.62297, 
    34.62264, 34.62237, 34.62216, 34.62203, 34.62199, 34.62204, 34.62215, 
    34.62234,
  34.63095, 34.63029, 34.62974, 34.62932, 34.62896, 34.6286, 34.62827, 
    34.62797, 34.62774, 34.62756, 34.62747, 34.62748, 34.62755, 34.62767, 
    34.62782,
  34.63592, 34.63525, 34.63474, 34.63438, 34.63406, 34.63376, 34.63346, 
    34.6332, 34.63299, 34.63284, 34.63279, 34.63285, 34.63298, 34.63313, 
    34.6333,
  34.64088, 34.64022, 34.63973, 34.63937, 34.63907, 34.63878, 34.6385, 
    34.63826, 34.63806, 34.63792, 34.63791, 34.63801, 34.6382, 34.63842, 
    34.63866,
  34.64583, 34.6452, 34.6447, 34.64429, 34.64397, 34.64367, 34.64339, 
    34.64315, 34.64296, 34.64284, 34.64284, 34.64298, 34.64322, 34.64352, 
    34.64383,
  34.65068, 34.65006, 34.64954, 34.64911, 34.64875, 34.64843, 34.64815, 
    34.6479, 34.64773, 34.64763, 34.64766, 34.64783, 34.64812, 34.64846, 
    34.64881,
  34.6553, 34.65467, 34.65414, 34.6537, 34.65334, 34.65303, 34.65274, 
    34.65252, 34.65237, 34.65231, 34.65237, 34.65257, 34.65289, 34.65325, 
    34.65361,
  34.65963, 34.659, 34.65847, 34.65804, 34.6577, 34.65741, 34.65716, 
    34.65697, 34.65688, 34.65687, 34.65698, 34.65722, 34.65755, 34.65792, 
    34.65829,
  34.61257, 34.61216, 34.61177, 34.61144, 34.61115, 34.61088, 34.61063, 
    34.61045, 34.61032, 34.61025, 34.61023, 34.61029, 34.61043, 34.61066, 
    34.61102,
  34.61723, 34.61683, 34.61646, 34.61613, 34.61584, 34.61558, 34.61534, 
    34.61516, 34.61504, 34.61498, 34.61499, 34.61506, 34.61519, 34.6154, 
    34.61572,
  34.62178, 34.62136, 34.621, 34.62069, 34.62043, 34.62022, 34.62003, 
    34.61989, 34.61981, 34.61979, 34.61983, 34.61993, 34.62009, 34.6203, 
    34.62056,
  34.62624, 34.6258, 34.62545, 34.62518, 34.62498, 34.62482, 34.6247, 
    34.62461, 34.62457, 34.62458, 34.62466, 34.62481, 34.625, 34.62521, 
    34.62545,
  34.63063, 34.63018, 34.62984, 34.62962, 34.62947, 34.62936, 34.62926, 
    34.62921, 34.62919, 34.62923, 34.62933, 34.62951, 34.62973, 34.62997, 
    34.63023,
  34.63501, 34.63455, 34.63422, 34.63402, 34.63388, 34.63377, 34.63368, 
    34.63362, 34.63361, 34.63364, 34.63375, 34.63395, 34.63421, 34.63449, 
    34.63481,
  34.63943, 34.63896, 34.63863, 34.6384, 34.63824, 34.6381, 34.63798, 
    34.6379, 34.63786, 34.6379, 34.63801, 34.63821, 34.6385, 34.63884, 
    34.63921,
  34.64384, 34.64337, 34.643, 34.64273, 34.64252, 34.64235, 34.64219, 
    34.64208, 34.64203, 34.64206, 34.64218, 34.6424, 34.64272, 34.64309, 
    34.64349,
  34.64801, 34.64756, 34.64719, 34.6469, 34.64667, 34.64647, 34.64629, 
    34.64617, 34.64612, 34.64616, 34.64631, 34.64655, 34.64688, 34.64727, 
    34.64768,
  34.65185, 34.65145, 34.65111, 34.65083, 34.65061, 34.65041, 34.65025, 
    34.65015, 34.65014, 34.65022, 34.6504, 34.65068, 34.65103, 34.65142, 
    34.65183,
  34.61934, 34.619, 34.61871, 34.61845, 34.61824, 34.61805, 34.6179, 
    34.61778, 34.61773, 34.61774, 34.61782, 34.61795, 34.61814, 34.6184, 
    34.61874,
  34.62331, 34.62298, 34.6227, 34.62247, 34.62227, 34.62209, 34.62196, 
    34.62187, 34.62185, 34.62188, 34.62197, 34.62212, 34.62231, 34.62254, 
    34.62284,
  34.6272, 34.62687, 34.62659, 34.62637, 34.62619, 34.62605, 34.62595, 
    34.62592, 34.62595, 34.62604, 34.62618, 34.62636, 34.62658, 34.62681, 
    34.62708,
  34.631, 34.63065, 34.63037, 34.63016, 34.63002, 34.62993, 34.6299, 
    34.62993, 34.63002, 34.63016, 34.63034, 34.63056, 34.6308, 34.63105, 
    34.6313,
  34.63468, 34.63433, 34.63407, 34.6339, 34.6338, 34.63376, 34.63377, 
    34.63385, 34.63397, 34.63414, 34.63434, 34.63459, 34.63485, 34.63512, 
    34.63538,
  34.63828, 34.63795, 34.63771, 34.63758, 34.63751, 34.6375, 34.63754, 
    34.63762, 34.63775, 34.63792, 34.63814, 34.63839, 34.63868, 34.63897, 
    34.63927,
  34.64181, 34.64152, 34.64132, 34.64121, 34.64116, 34.64116, 34.64119, 
    34.64127, 34.64139, 34.64156, 34.64177, 34.64203, 34.64232, 34.64265, 
    34.64299,
  34.64528, 34.64502, 34.64486, 34.64476, 34.64472, 34.64472, 34.64475, 
    34.64481, 34.64492, 34.64509, 34.6453, 34.64556, 34.64586, 34.64621, 
    34.64658,
  34.64865, 34.6484, 34.64825, 34.64817, 34.64814, 34.64815, 34.64817, 
    34.64823, 34.64834, 34.64851, 34.64873, 34.64899, 34.64931, 34.64966, 
    34.65003,
  34.65191, 34.65167, 34.6515, 34.65142, 34.6514, 34.65141, 34.65143, 
    34.65151, 34.65165, 34.65184, 34.65207, 34.65235, 34.65267, 34.65302, 
    34.65339,
  34.63158, 34.63139, 34.63122, 34.63109, 34.631, 34.63093, 34.63089, 
    34.63089, 34.63093, 34.631, 34.63111, 34.63126, 34.63147, 34.63173, 
    34.63206,
  34.63458, 34.63442, 34.6343, 34.63422, 34.63417, 34.63414, 34.63414, 
    34.63417, 34.63425, 34.63436, 34.6345, 34.63469, 34.63492, 34.63519, 
    34.63552,
  34.63754, 34.63741, 34.63731, 34.63726, 34.63725, 34.63726, 34.63732, 
    34.63742, 34.63755, 34.63771, 34.6379, 34.63815, 34.63842, 34.63872, 
    34.63905,
  34.64045, 34.64032, 34.64025, 34.64023, 34.64025, 34.64032, 34.64043, 
    34.64059, 34.64077, 34.641, 34.64124, 34.64153, 34.64185, 34.64218, 
    34.64251,
  34.64328, 34.64317, 34.64311, 34.64312, 34.64317, 34.64328, 34.64343, 
    34.64363, 34.64387, 34.64413, 34.64441, 34.64474, 34.64508, 34.64544, 
    34.64579,
  34.64603, 34.64594, 34.6459, 34.64592, 34.64601, 34.64614, 34.64632, 
    34.64655, 34.64681, 34.64709, 34.64739, 34.64772, 34.64808, 34.64845, 
    34.64883,
  34.64873, 34.64865, 34.64864, 34.64868, 34.64878, 34.64892, 34.64912, 
    34.64936, 34.64963, 34.64992, 34.65023, 34.65056, 34.65092, 34.6513, 
    34.6517,
  34.65134, 34.6513, 34.65131, 34.65137, 34.65149, 34.65165, 34.65185, 
    34.6521, 34.65238, 34.65267, 34.65298, 34.65332, 34.65367, 34.65405, 
    34.65444,
  34.65382, 34.65382, 34.65387, 34.65397, 34.65411, 34.65428, 34.6545, 
    34.65476, 34.65504, 34.65534, 34.65565, 34.65598, 34.65632, 34.65668, 
    34.65706,
  34.65616, 34.65622, 34.65631, 34.65645, 34.65661, 34.65681, 34.65704, 
    34.6573, 34.65759, 34.65789, 34.65819, 34.6585, 34.65882, 34.65916, 
    34.65952,
  34.65057, 34.65036, 34.65019, 34.65007, 34.64999, 34.64995, 34.64993, 
    34.64996, 34.65002, 34.65013, 34.65027, 34.65044, 34.65064, 34.65087, 
    34.65114,
  34.65264, 34.65246, 34.65232, 34.65224, 34.65221, 34.6522, 34.65222, 
    34.65229, 34.6524, 34.65255, 34.65273, 34.65294, 34.65317, 34.65342, 
    34.6537,
  34.65465, 34.65449, 34.65437, 34.65432, 34.65431, 34.65434, 34.65441, 
    34.65453, 34.6547, 34.6549, 34.65512, 34.65538, 34.65565, 34.65594, 
    34.65623,
  34.65662, 34.65647, 34.65636, 34.65632, 34.65634, 34.65641, 34.65654, 
    34.65671, 34.65693, 34.65717, 34.65744, 34.65773, 34.65804, 34.65836, 
    34.65867,
  34.65855, 34.6584, 34.65831, 34.65828, 34.65833, 34.65843, 34.6586, 
    34.65882, 34.65907, 34.65934, 34.65963, 34.65994, 34.66027, 34.66059, 
    34.66091,
  34.66043, 34.66029, 34.66021, 34.66021, 34.66027, 34.6604, 34.6606, 
    34.66085, 34.66112, 34.6614, 34.66169, 34.662, 34.66232, 34.66265, 
    34.66298,
  34.66227, 34.66216, 34.6621, 34.66212, 34.66221, 34.66236, 34.66257, 
    34.66283, 34.6631, 34.66338, 34.66367, 34.66396, 34.66426, 34.66458, 
    34.66489,
  34.66409, 34.66401, 34.66399, 34.66403, 34.66415, 34.66431, 34.66454, 
    34.66479, 34.66506, 34.66533, 34.6656, 34.66589, 34.66617, 34.66647, 
    34.66676,
  34.66589, 34.66584, 34.66586, 34.66594, 34.66607, 34.66626, 34.66648, 
    34.66673, 34.667, 34.66725, 34.66751, 34.66777, 34.66804, 34.66831, 
    34.66859,
  34.66768, 34.66768, 34.66772, 34.66783, 34.66797, 34.66815, 34.66837, 
    34.66862, 34.66888, 34.66913, 34.66938, 34.66962, 34.66987, 34.67012, 
    34.67038,
  34.6684, 34.6682, 34.66801, 34.66784, 34.66772, 34.66762, 34.66756, 
    34.66754, 34.66757, 34.66763, 34.66772, 34.66781, 34.66793, 34.66806, 
    34.66821,
  34.67007, 34.6699, 34.66974, 34.66962, 34.66955, 34.6695, 34.66948, 
    34.66951, 34.66958, 34.66967, 34.66978, 34.66991, 34.67005, 34.67021, 
    34.67037,
  34.67172, 34.67156, 34.67143, 34.67134, 34.67131, 34.6713, 34.67133, 
    34.67141, 34.67152, 34.67164, 34.67178, 34.67194, 34.67211, 34.6723, 
    34.67249,
  34.67336, 34.67321, 34.6731, 34.67303, 34.67302, 34.67306, 34.67313, 
    34.67325, 34.67338, 34.67353, 34.67368, 34.67385, 34.67405, 34.67426, 
    34.67445,
  34.67498, 34.67484, 34.67474, 34.67469, 34.67471, 34.67477, 34.67487, 
    34.67501, 34.67517, 34.67532, 34.67547, 34.67564, 34.67583, 34.67604, 
    34.67625,
  34.67657, 34.67645, 34.67636, 34.67633, 34.67637, 34.67645, 34.67657, 
    34.67672, 34.67687, 34.67702, 34.67715, 34.6773, 34.67747, 34.67765, 
    34.67784,
  34.67813, 34.67803, 34.67797, 34.67796, 34.67801, 34.6781, 34.67823, 
    34.67838, 34.67852, 34.67864, 34.67876, 34.67888, 34.67902, 34.67918, 
    34.67935,
  34.67966, 34.6796, 34.67957, 34.67959, 34.67965, 34.67974, 34.67986, 34.68, 
    34.68012, 34.68022, 34.68031, 34.6804, 34.68052, 34.68065, 34.6808,
  34.68118, 34.68115, 34.68115, 34.68118, 34.68125, 34.68134, 34.68146, 
    34.68158, 34.68167, 34.68176, 34.68182, 34.6819, 34.68199, 34.6821, 
    34.68223,
  34.68267, 34.68267, 34.6827, 34.68274, 34.6828, 34.68288, 34.68299, 
    34.68309, 34.68317, 34.68324, 34.68329, 34.68335, 34.68342, 34.68352, 
    34.68364,
  34.68723, 34.68703, 34.68685, 34.68667, 34.68652, 34.68638, 34.68628, 
    34.68622, 34.6862, 34.68618, 34.68618, 34.68618, 34.6862, 34.68621, 
    34.68624,
  34.68832, 34.68814, 34.68798, 34.68784, 34.68772, 34.68762, 34.68756, 
    34.68754, 34.68755, 34.68756, 34.68758, 34.68762, 34.68768, 34.68774, 
    34.6878,
  34.68941, 34.68924, 34.68909, 34.68897, 34.68888, 34.68882, 34.68879, 
    34.68881, 34.68884, 34.68888, 34.68894, 34.68901, 34.68912, 34.68921, 
    34.68932,
  34.69052, 34.69036, 34.69021, 34.69011, 34.69004, 34.69, 34.69001, 
    34.69004, 34.6901, 34.69016, 34.69024, 34.69035, 34.69048, 34.69061, 
    34.69075,
  34.69165, 34.69149, 34.69135, 34.69125, 34.6912, 34.69118, 34.69121, 
    34.69126, 34.69133, 34.6914, 34.69148, 34.69159, 34.69172, 34.69186, 
    34.69201,
  34.69279, 34.69264, 34.69251, 34.69242, 34.69237, 34.69237, 34.6924, 
    34.69246, 34.69252, 34.69259, 34.69267, 34.69276, 34.69289, 34.69302, 
    34.69318,
  34.69392, 34.69379, 34.69368, 34.6936, 34.69356, 34.69357, 34.6936, 
    34.69365, 34.6937, 34.69375, 34.69381, 34.6939, 34.694, 34.69411, 34.69424,
  34.69505, 34.69494, 34.69485, 34.69478, 34.69475, 34.69476, 34.69478, 
    34.69482, 34.69486, 34.69489, 34.69494, 34.69501, 34.6951, 34.6952, 
    34.69534,
  34.69616, 34.69607, 34.696, 34.69595, 34.69593, 34.69593, 34.69595, 
    34.69598, 34.69601, 34.69603, 34.69607, 34.69613, 34.6962, 34.6963, 
    34.69642,
  34.69726, 34.69719, 34.69714, 34.6971, 34.69708, 34.69708, 34.6971, 
    34.69712, 34.69715, 34.69717, 34.6972, 34.69725, 34.69731, 34.6974, 
    34.69752,
  34.70597, 34.70581, 34.70566, 34.70552, 34.7054, 34.70531, 34.70523, 
    34.70517, 34.70512, 34.70509, 34.70507, 34.70506, 34.70505, 34.70503, 
    34.70501,
  34.70692, 34.7068, 34.70668, 34.70658, 34.7065, 34.70644, 34.70639, 
    34.70637, 34.70636, 34.70636, 34.70638, 34.70642, 34.70646, 34.7065, 
    34.70653,
  34.7079, 34.7078, 34.7077, 34.70762, 34.70757, 34.70753, 34.70752, 
    34.70753, 34.70756, 34.7076, 34.70766, 34.70774, 34.70782, 34.70792, 
    34.708,
  34.70889, 34.70881, 34.70872, 34.70866, 34.70861, 34.7086, 34.70862, 
    34.70866, 34.70872, 34.70879, 34.70888, 34.70897, 34.70908, 34.70921, 
    34.70931,
  34.70988, 34.70981, 34.70974, 34.70967, 34.70964, 34.70965, 34.70969, 
    34.70975, 34.70983, 34.70992, 34.71001, 34.7101, 34.71021, 34.71034, 
    34.71048,
  34.71083, 34.71078, 34.71072, 34.71067, 34.71065, 34.71067, 34.71073, 
    34.7108, 34.71088, 34.71097, 34.71106, 34.71114, 34.71124, 34.71134, 
    34.71144,
  34.71177, 34.71173, 34.71169, 34.71165, 34.71165, 34.71169, 34.71175, 
    34.71182, 34.7119, 34.71198, 34.71206, 34.71214, 34.71222, 34.71231, 
    34.71242,
  34.71267, 34.71266, 34.71264, 34.71263, 34.71265, 34.7127, 34.71276, 
    34.71284, 34.71291, 34.71299, 34.71305, 34.71313, 34.71319, 34.71326, 
    34.71335,
  34.71356, 34.71357, 34.71358, 34.71359, 34.71363, 34.71368, 34.71375, 
    34.71383, 34.7139, 34.71397, 34.71403, 34.71409, 34.71415, 34.71421, 
    34.71429,
  34.71443, 34.71446, 34.71449, 34.71453, 34.71458, 34.71464, 34.71471, 
    34.71479, 34.71486, 34.71493, 34.71498, 34.71503, 34.71508, 34.71515, 
    34.71523,
  34.72516, 34.72504, 34.72491, 34.7248, 34.7247, 34.72462, 34.72457, 
    34.72453, 34.72449, 34.72447, 34.72445, 34.72443, 34.7244, 34.72435, 
    34.72429,
  34.72576, 34.72566, 34.72556, 34.72548, 34.72541, 34.72537, 34.72535, 
    34.72534, 34.72533, 34.72534, 34.72535, 34.72536, 34.72538, 34.72539, 
    34.72538,
  34.72639, 34.72631, 34.72623, 34.72616, 34.72612, 34.7261, 34.7261, 
    34.72612, 34.72615, 34.72618, 34.72623, 34.72628, 34.72634, 34.72639, 
    34.72645,
  34.72705, 34.72698, 34.72691, 34.72685, 34.72681, 34.72681, 34.72683, 
    34.72688, 34.72693, 34.72699, 34.72706, 34.72712, 34.7272, 34.72729, 
    34.7274,
  34.72775, 34.72768, 34.72761, 34.72755, 34.72752, 34.72752, 34.72756, 
    34.72762, 34.72768, 34.72776, 34.72783, 34.7279, 34.72797, 34.72804, 
    34.72812,
  34.72845, 34.7284, 34.72833, 34.72828, 34.72824, 34.72825, 34.72829, 
    34.72835, 34.72842, 34.72849, 34.72857, 34.72863, 34.72869, 34.72875, 
    34.72884,
  34.72915, 34.72911, 34.72906, 34.72902, 34.72899, 34.729, 34.72904, 
    34.7291, 34.72916, 34.72922, 34.72928, 34.72934, 34.72938, 34.72942, 
    34.72945,
  34.72982, 34.72981, 34.72978, 34.72975, 34.72974, 34.72976, 34.7298, 
    34.72985, 34.7299, 34.72995, 34.73, 34.73003, 34.73006, 34.73009, 34.73013,
  34.7305, 34.7305, 34.73048, 34.73047, 34.73048, 34.7305, 34.73055, 
    34.73059, 34.73064, 34.73068, 34.73071, 34.73074, 34.73076, 34.73078, 
    34.73082,
  34.73117, 34.73118, 34.73119, 34.73119, 34.73121, 34.73124, 34.73128, 
    34.73133, 34.73137, 34.7314, 34.73143, 34.73145, 34.73146, 34.73148, 
    34.73152,
  34.74409, 34.74399, 34.7439, 34.74381, 34.74374, 34.74368, 34.74364, 
    34.7436, 34.74358, 34.74355, 34.74353, 34.7435, 34.74347, 34.74342, 
    34.74337,
  34.74441, 34.74432, 34.74424, 34.74417, 34.74412, 34.74408, 34.74405, 
    34.74403, 34.74402, 34.74402, 34.74403, 34.74404, 34.74405, 34.74406, 
    34.74405,
  34.74477, 34.74469, 34.74461, 34.74455, 34.74451, 34.74448, 34.74446, 
    34.74446, 34.74446, 34.74448, 34.74451, 34.74454, 34.74458, 34.74463, 
    34.74466,
  34.74517, 34.74509, 34.74502, 34.74495, 34.74491, 34.74489, 34.74488, 
    34.74489, 34.74492, 34.74495, 34.74498, 34.74503, 34.74506, 34.74511, 
    34.74514,
  34.74563, 34.74555, 34.74547, 34.7454, 34.74535, 34.74532, 34.74532, 
    34.74533, 34.74537, 34.74541, 34.74545, 34.7455, 34.74553, 34.74559, 
    34.74568,
  34.74611, 34.74604, 34.74596, 34.74589, 34.74583, 34.7458, 34.7458, 
    34.74582, 34.74585, 34.74588, 34.74593, 34.74597, 34.74599, 34.74601, 
    34.74599,
  34.7466, 34.74654, 34.74647, 34.7464, 34.74635, 34.74632, 34.74632, 
    34.74633, 34.74636, 34.74639, 34.74643, 34.74646, 34.74648, 34.74649, 
    34.74651,
  34.74707, 34.74703, 34.74698, 34.74692, 34.74687, 34.74685, 34.74685, 
    34.74687, 34.74689, 34.74691, 34.74694, 34.74696, 34.74697, 34.74697, 
    34.74699,
  34.74755, 34.74752, 34.74748, 34.74744, 34.7474, 34.74738, 34.74739, 
    34.74741, 34.74743, 34.74744, 34.74745, 34.74746, 34.74746, 34.74746, 
    34.74747,
  34.74804, 34.74802, 34.74799, 34.74796, 34.74794, 34.74792, 34.74793, 
    34.74795, 34.74797, 34.74798, 34.74798, 34.74798, 34.74798, 34.74798, 
    34.748,
  34.76316, 34.76305, 34.76296, 34.76288, 34.76281, 34.76276, 34.76271, 
    34.76269, 34.76267, 34.76266, 34.76266, 34.76267, 34.76266, 34.76266, 
    34.76265,
  34.76334, 34.76324, 34.76315, 34.76308, 34.76302, 34.76298, 34.76295, 
    34.76294, 34.76293, 34.76293, 34.76295, 34.76297, 34.76298, 34.763, 34.763,
  34.76357, 34.76347, 34.76338, 34.76331, 34.76325, 34.76322, 34.7632, 
    34.76319, 34.7632, 34.76321, 34.76324, 34.76328, 34.76333, 34.76339, 
    34.76346,
  34.76385, 34.76374, 34.76365, 34.76357, 34.76351, 34.76347, 34.76344, 
    34.76343, 34.76343, 34.76344, 34.76346, 34.76349, 34.76355, 34.76361, 
    34.76369,
  34.7642, 34.76409, 34.76398, 34.76389, 34.76381, 34.76376, 34.76372, 
    34.7637, 34.76369, 34.76369, 34.7637, 34.76372, 34.76375, 34.76373, 
    34.76364,
  34.76461, 34.7645, 34.76439, 34.76428, 34.76418, 34.76411, 34.76407, 
    34.76405, 34.76404, 34.76405, 34.76407, 34.76411, 34.76415, 34.76415, 
    34.76418,
  34.76502, 34.76492, 34.76482, 34.76471, 34.76461, 34.76453, 34.76448, 
    34.76447, 34.76447, 34.76449, 34.76452, 34.76455, 34.76458, 34.7646, 
    34.7646,
  34.76543, 34.76534, 34.76524, 34.76514, 34.76504, 34.76496, 34.76492, 
    34.7649, 34.76491, 34.76492, 34.76493, 34.76494, 34.76495, 34.76495, 
    34.76496,
  34.76584, 34.76576, 34.76567, 34.76557, 34.76548, 34.7654, 34.76536, 
    34.76535, 34.76535, 34.76535, 34.76535, 34.76535, 34.76535, 34.76535, 
    34.76538,
  34.76625, 34.76618, 34.76609, 34.76601, 34.76593, 34.76587, 34.76583, 
    34.76582, 34.76581, 34.76581, 34.76581, 34.7658, 34.7658, 34.76581, 
    34.76584,
  34.78043, 34.78032, 34.78021, 34.78011, 34.78002, 34.77994, 34.77988, 
    34.77983, 34.77979, 34.77977, 34.77977, 34.77975, 34.77974, 34.77973, 
    34.77972,
  34.78053, 34.78041, 34.78031, 34.78022, 34.78013, 34.78006, 34.78001, 
    34.77998, 34.77994, 34.77991, 34.7799, 34.77989, 34.77988, 34.77987, 
    34.77986,
  34.78067, 34.78056, 34.78046, 34.78037, 34.7803, 34.78027, 34.78025, 
    34.78025, 34.78024, 34.78022, 34.7802, 34.78019, 34.78017, 34.78016, 
    34.78017,
  34.78088, 34.78077, 34.78066, 34.78057, 34.78051, 34.78049, 34.78052, 
    34.78056, 34.78062, 34.78067, 34.7807, 34.78074, 34.78082, 34.78098, 
    34.78112,
  34.78116, 34.78105, 34.78094, 34.78083, 34.78076, 34.78072, 34.78074, 
    34.78078, 34.78086, 34.78094, 34.781, 34.78106, 34.78117, 34.78145, 
    34.78187,
  34.7815, 34.7814, 34.78129, 34.78118, 34.78108, 34.78101, 34.78098, 34.781, 
    34.78104, 34.78109, 34.78113, 34.78116, 34.7812, 34.78131, 34.78136,
  34.78185, 34.78176, 34.78167, 34.78156, 34.78146, 34.78136, 34.7813, 
    34.78128, 34.78128, 34.7813, 34.78131, 34.7813, 34.78128, 34.78127, 
    34.78123,
  34.78219, 34.78211, 34.78203, 34.78194, 34.78183, 34.78174, 34.78166, 
    34.78162, 34.7816, 34.78159, 34.78157, 34.78154, 34.7815, 34.78146, 
    34.78144,
  34.78254, 34.78246, 34.78238, 34.7823, 34.7822, 34.78211, 34.78204, 
    34.78199, 34.78197, 34.78194, 34.78191, 34.78188, 34.78184, 34.7818, 
    34.78179,
  34.78289, 34.78281, 34.78274, 34.78265, 34.78257, 34.78249, 34.78242, 
    34.78239, 34.78237, 34.78234, 34.78232, 34.7823, 34.78228, 34.78227, 
    34.78228,
  34.79328, 34.7932, 34.79311, 34.79304, 34.79297, 34.7929, 34.79285, 
    34.7928, 34.79277, 34.79276, 34.79274, 34.79273, 34.79271, 34.79269, 
    34.79267,
  34.79337, 34.79329, 34.7932, 34.79312, 34.79305, 34.79298, 34.79292, 
    34.79287, 34.79284, 34.79281, 34.7928, 34.79279, 34.79277, 34.79277, 
    34.79277,
  34.7935, 34.79341, 34.79332, 34.79324, 34.79316, 34.79309, 34.79303, 
    34.79297, 34.79291, 34.79286, 34.79282, 34.79279, 34.79276, 34.79274, 
    34.79273,
  34.79368, 34.79359, 34.7935, 34.7934, 34.79332, 34.79324, 34.79318, 
    34.79313, 34.79307, 34.79301, 34.79294, 34.79287, 34.79278, 34.79261, 
    34.79247,
  34.79393, 34.79384, 34.79375, 34.79364, 34.79355, 34.79346, 34.7934, 
    34.79337, 34.79335, 34.79333, 34.7933, 34.79325, 34.79318, 34.79302, 
    34.79274,
  34.7942, 34.79413, 34.79405, 34.79396, 34.79386, 34.79377, 34.7937, 
    34.79366, 34.79367, 34.7937, 34.79373, 34.79374, 34.79375, 34.79377, 
    34.79389,
  34.7945, 34.79443, 34.79437, 34.79429, 34.7942, 34.79411, 34.79403, 
    34.79398, 34.79399, 34.79401, 34.79404, 34.79403, 34.79402, 34.79404, 
    34.79407,
  34.7948, 34.79473, 34.79467, 34.79461, 34.79453, 34.79444, 34.79436, 
    34.7943, 34.79428, 34.79427, 34.79425, 34.79421, 34.79415, 34.79409, 
    34.79403,
  34.79508, 34.79502, 34.79497, 34.7949, 34.79483, 34.79475, 34.79467, 
    34.7946, 34.79456, 34.79452, 34.79448, 34.79443, 34.79437, 34.79432, 
    34.7943,
  34.79536, 34.7953, 34.79525, 34.79518, 34.7951, 34.79503, 34.79496, 
    34.7949, 34.79486, 34.79482, 34.79479, 34.79476, 34.79474, 34.79474, 
    34.79476,
  34.80344, 34.8034, 34.80336, 34.80332, 34.80329, 34.80326, 34.80325, 
    34.80324, 34.80324, 34.80325, 34.80326, 34.80327, 34.80328, 34.80328, 
    34.80328,
  34.80351, 34.80347, 34.80343, 34.80339, 34.80336, 34.80333, 34.80331, 
    34.8033, 34.80331, 34.80332, 34.80333, 34.80335, 34.80336, 34.80336, 
    34.80336,
  34.80359, 34.80355, 34.80351, 34.80347, 34.80344, 34.80341, 34.80338, 
    34.80336, 34.80335, 34.80334, 34.80334, 34.80334, 34.80333, 34.80332, 
    34.80333,
  34.8037, 34.80365, 34.80361, 34.80357, 34.80353, 34.80349, 34.80346, 
    34.80344, 34.80342, 34.80339, 34.80337, 34.80335, 34.80333, 34.80333, 
    34.80336,
  34.80383, 34.80379, 34.80375, 34.80371, 34.80366, 34.80362, 34.80358, 
    34.80355, 34.80352, 34.80349, 34.80346, 34.80341, 34.80335, 34.8033, 
    34.8034,
  34.80399, 34.80395, 34.80392, 34.80388, 34.80384, 34.8038, 34.80376, 
    34.80372, 34.80369, 34.80366, 34.80362, 34.80357, 34.80348, 34.80331, 
    34.80307,
  34.80415, 34.80412, 34.80409, 34.80406, 34.80403, 34.80399, 34.80396, 
    34.80392, 34.8039, 34.80389, 34.80387, 34.80383, 34.80375, 34.80363, 
    34.80356,
  34.80433, 34.80429, 34.80427, 34.80424, 34.80421, 34.80418, 34.80414, 
    34.80411, 34.80408, 34.80408, 34.80408, 34.80405, 34.80402, 34.80401, 
    34.80405,
  34.8045, 34.80447, 34.80444, 34.80441, 34.80437, 34.80434, 34.8043, 
    34.80426, 34.80424, 34.80423, 34.80422, 34.80421, 34.8042, 34.80418, 
    34.8042,
  34.80466, 34.80463, 34.8046, 34.80456, 34.80453, 34.80449, 34.80445, 
    34.80442, 34.80438, 34.80436, 34.80436, 34.80436, 34.80437, 34.80438, 
    34.80441,
  34.81174, 34.81173, 34.81173, 34.81173, 34.81175, 34.81177, 34.81179, 
    34.81182, 34.81186, 34.81189, 34.81193, 34.81196, 34.81199, 34.81202, 
    34.81205,
  34.81184, 34.81183, 34.81183, 34.81184, 34.81184, 34.81186, 34.81188, 
    34.8119, 34.81194, 34.81197, 34.812, 34.81203, 34.81205, 34.81207, 
    34.81209,
  34.81195, 34.81193, 34.81192, 34.81192, 34.81192, 34.81193, 34.81194, 
    34.81196, 34.81198, 34.812, 34.81202, 34.81203, 34.81203, 34.81203, 
    34.81205,
  34.81205, 34.81204, 34.81202, 34.81201, 34.812, 34.812, 34.812, 34.812, 
    34.812, 34.812, 34.812, 34.812, 34.81197, 34.81197, 34.81193,
  34.81218, 34.81216, 34.81213, 34.81212, 34.8121, 34.81209, 34.81207, 
    34.81206, 34.81205, 34.81203, 34.81201, 34.81199, 34.81195, 34.81199, 
    34.81185,
  34.81233, 34.81229, 34.81227, 34.81225, 34.81224, 34.81222, 34.81221, 
    34.81219, 34.81216, 34.81213, 34.81209, 34.81205, 34.81202, 34.8121, 
    34.81229,
  34.8125, 34.81246, 34.81243, 34.8124, 34.81239, 34.81238, 34.81237, 
    34.81235, 34.81233, 34.81229, 34.81226, 34.81222, 34.81218, 34.81219, 
    34.81224,
  34.81268, 34.81263, 34.8126, 34.81257, 34.81255, 34.81254, 34.81253, 
    34.81251, 34.81249, 34.81246, 34.81244, 34.81242, 34.81239, 34.81239, 
    34.81241,
  34.81284, 34.81281, 34.81277, 34.81274, 34.81272, 34.81269, 34.81268, 
    34.81265, 34.81262, 34.8126, 34.81259, 34.81258, 34.81257, 34.81258, 
    34.81261,
  34.813, 34.81296, 34.81292, 34.81289, 34.81286, 34.81284, 34.81281, 
    34.81277, 34.81274, 34.81273, 34.81272, 34.81273, 34.81274, 34.81276, 
    34.81281,
  34.81851, 34.81852, 34.81853, 34.81856, 34.8186, 34.81865, 34.8187, 
    34.81874, 34.8188, 34.81885, 34.8189, 34.81894, 34.81898, 34.81901, 
    34.81904,
  34.81863, 34.81864, 34.81866, 34.8187, 34.81874, 34.81878, 34.81884, 
    34.81889, 34.81895, 34.819, 34.81906, 34.8191, 34.81914, 34.81916, 
    34.81919,
  34.81875, 34.81876, 34.81877, 34.8188, 34.81884, 34.81889, 34.81894, 
    34.819, 34.81905, 34.81909, 34.81913, 34.81917, 34.8192, 34.81923, 
    34.81926,
  34.81886, 34.81886, 34.81887, 34.81889, 34.81892, 34.81896, 34.819, 
    34.81905, 34.81911, 34.81916, 34.81919, 34.81922, 34.81924, 34.81925, 
    34.81934,
  34.81897, 34.81897, 34.81897, 34.81899, 34.819, 34.81903, 34.81906, 
    34.81909, 34.81913, 34.81917, 34.81921, 34.81921, 34.81919, 34.81918, 
    34.8194,
  34.8191, 34.81909, 34.81909, 34.8191, 34.81911, 34.81913, 34.81916, 
    34.81918, 34.8192, 34.81921, 34.81922, 34.8192, 34.81918, 34.81917, 
    34.81928,
  34.81925, 34.81924, 34.81923, 34.81923, 34.81924, 34.81926, 34.81929, 
    34.81932, 34.81932, 34.81932, 34.81931, 34.81928, 34.81927, 34.81928, 
    34.81933,
  34.81942, 34.8194, 34.81939, 34.81938, 34.81939, 34.81941, 34.81945, 
    34.81947, 34.81948, 34.81947, 34.81945, 34.81944, 34.81943, 34.81939, 
    34.81933,
  34.81958, 34.81957, 34.81956, 34.81955, 34.81956, 34.81958, 34.8196, 
    34.81963, 34.81963, 34.81963, 34.81963, 34.81964, 34.81963, 34.8196, 
    34.81956,
  34.81975, 34.81974, 34.81973, 34.81973, 34.81973, 34.81974, 34.81976, 
    34.81977, 34.81978, 34.81979, 34.8198, 34.81983, 34.81985, 34.81989, 
    34.81994,
  34.82449, 34.82448, 34.82449, 34.8245, 34.82454, 34.82457, 34.8246, 
    34.82464, 34.82468, 34.82472, 34.82475, 34.82478, 34.82479, 34.82481, 
    34.82483,
  34.8246, 34.8246, 34.82461, 34.82463, 34.82467, 34.8247, 34.82474, 
    34.82478, 34.82483, 34.82487, 34.82491, 34.82495, 34.82498, 34.825, 
    34.82502,
  34.82472, 34.82472, 34.82473, 34.82475, 34.82478, 34.82481, 34.82485, 
    34.82489, 34.82493, 34.82497, 34.825, 34.82504, 34.82507, 34.8251, 
    34.82514,
  34.82483, 34.82482, 34.82483, 34.82484, 34.82487, 34.8249, 34.82494, 
    34.82497, 34.82501, 34.82504, 34.82507, 34.82508, 34.8251, 34.82508, 
    34.82504,
  34.82494, 34.82492, 34.82492, 34.82493, 34.82494, 34.82497, 34.825, 
    34.82503, 34.82507, 34.82511, 34.82514, 34.82515, 34.82513, 34.82505, 
    34.82483,
  34.82505, 34.82504, 34.82502, 34.82502, 34.82503, 34.82504, 34.82507, 
    34.8251, 34.82514, 34.82517, 34.8252, 34.8252, 34.82517, 34.82509, 
    34.82494,
  34.82517, 34.82516, 34.82515, 34.82514, 34.82514, 34.82515, 34.82517, 
    34.8252, 34.82523, 34.82524, 34.82525, 34.82524, 34.8252, 34.82512, 
    34.82502,
  34.8253, 34.82529, 34.82529, 34.82528, 34.82527, 34.82528, 34.8253, 
    34.82533, 34.82534, 34.82534, 34.82532, 34.82529, 34.82527, 34.82522, 
    34.8252,
  34.82543, 34.82542, 34.82542, 34.82542, 34.82541, 34.82542, 34.82544, 
    34.82545, 34.82546, 34.82545, 34.82543, 34.82541, 34.82542, 34.82542, 
    34.82544,
  34.82555, 34.82555, 34.82555, 34.82554, 34.82554, 34.82555, 34.82556, 
    34.82557, 34.82558, 34.82557, 34.82556, 34.82557, 34.8256, 34.82563, 
    34.82567,
  34.82911, 34.82911, 34.82912, 34.82915, 34.8292, 34.82925, 34.8293, 
    34.82935, 34.8294, 34.82944, 34.82948, 34.8295, 34.82952, 34.82955, 
    34.82961,
  34.82924, 34.82925, 34.82928, 34.82932, 34.82937, 34.82942, 34.82947, 
    34.82952, 34.82959, 34.82966, 34.82972, 34.82977, 34.8298, 34.82983, 
    34.82986,
  34.82937, 34.82938, 34.82941, 34.82946, 34.82952, 34.82957, 34.82962, 
    34.82968, 34.82975, 34.82982, 34.82989, 34.82996, 34.83001, 34.83006, 
    34.8301,
  34.8295, 34.82951, 34.82953, 34.82957, 34.82962, 34.82968, 34.82973, 
    34.8298, 34.82987, 34.82994, 34.83001, 34.83009, 34.83016, 34.83021, 
    34.83023,
  34.82961, 34.82962, 34.82964, 34.82967, 34.82971, 34.82976, 34.82982, 
    34.82988, 34.82996, 34.83004, 34.83012, 34.83018, 34.83025, 34.83026, 
    34.83027,
  34.82974, 34.82974, 34.82975, 34.82976, 34.82978, 34.82983, 34.82989, 
    34.82996, 34.83005, 34.83014, 34.83023, 34.83028, 34.83032, 34.83032, 
    34.83031,
  34.82988, 34.82988, 34.82988, 34.82988, 34.82989, 34.82992, 34.82998, 
    34.83006, 34.83016, 34.83027, 34.83035, 34.83039, 34.83041, 34.83049, 
    34.83062,
  34.83002, 34.83002, 34.83003, 34.83002, 34.83003, 34.83005, 34.8301, 
    34.83019, 34.8303, 34.8304, 34.83047, 34.83052, 34.83057, 34.83075, 34.831,
  34.83016, 34.83017, 34.83017, 34.83017, 34.83017, 34.83019, 34.83024, 
    34.83033, 34.83044, 34.83053, 34.8306, 34.83068, 34.83078, 34.83097, 
    34.83117,
  34.83029, 34.8303, 34.8303, 34.8303, 34.8303, 34.83032, 34.83038, 34.83047, 
    34.83057, 34.83066, 34.83075, 34.83083, 34.83093, 34.83107, 34.83119,
  34.83331, 34.83333, 34.83337, 34.83342, 34.83348, 34.83354, 34.8336, 
    34.83364, 34.83369, 34.83373, 34.83376, 34.83376, 34.83377, 34.83378, 
    34.83382,
  34.83344, 34.83347, 34.83352, 34.83359, 34.83366, 34.83371, 34.83376, 
    34.83381, 34.83385, 34.8339, 34.83394, 34.83397, 34.83398, 34.83399, 
    34.83399,
  34.83356, 34.8336, 34.83366, 34.83374, 34.83381, 34.83387, 34.83392, 
    34.83397, 34.83403, 34.83408, 34.83413, 34.83418, 34.83422, 34.83425, 
    34.83426,
  34.83366, 34.8337, 34.83376, 34.83384, 34.83392, 34.83399, 34.83406, 
    34.83413, 34.83419, 34.83427, 34.83435, 34.83444, 34.83453, 34.83463, 
    34.83471,
  34.83375, 34.83379, 34.83385, 34.83391, 34.83398, 34.83405, 34.83414, 
    34.83422, 34.83432, 34.83442, 34.83453, 34.83463, 34.83472, 34.83485, 
    34.83508,
  34.83384, 34.83388, 34.83393, 34.83398, 34.83403, 34.8341, 34.83417, 
    34.83427, 34.8344, 34.83455, 34.83469, 34.83479, 34.83484, 34.83494, 
    34.83518,
  34.83393, 34.83397, 34.83401, 34.83406, 34.8341, 34.83416, 34.83422, 
    34.83432, 34.83447, 34.83466, 34.83485, 34.83496, 34.83503, 34.83514, 
    34.83537,
  34.83403, 34.83406, 34.8341, 34.83415, 34.83419, 34.83424, 34.83432, 
    34.83442, 34.83458, 34.83479, 34.83499, 34.83512, 34.83525, 34.83545, 
    34.83566,
  34.83413, 34.83416, 34.8342, 34.83424, 34.83429, 34.83434, 34.83442, 
    34.83454, 34.83471, 34.83492, 34.83511, 34.83528, 34.83547, 34.83569, 
    34.83582,
  34.83424, 34.83426, 34.8343, 34.83434, 34.83438, 34.83443, 34.83452, 
    34.83465, 34.83482, 34.83501, 34.83522, 34.83541, 34.83558, 34.8357, 
    34.83576,
  34.83692, 34.83691, 34.83691, 34.83694, 34.83698, 34.83706, 34.83717, 
    34.83728, 34.83737, 34.83743, 34.83747, 34.83751, 34.83755, 34.83763, 
    34.83772,
  34.83698, 34.83698, 34.837, 34.83704, 34.8371, 34.8372, 34.83733, 34.83745, 
    34.83756, 34.83766, 34.83775, 34.83781, 34.83787, 34.83792, 34.83797,
  34.83705, 34.83706, 34.83709, 34.83714, 34.8372, 34.8373, 34.83742, 
    34.83755, 34.8377, 34.83785, 34.83801, 34.83813, 34.83823, 34.83834, 
    34.83844,
  34.83711, 34.83713, 34.83716, 34.83721, 34.83726, 34.83733, 34.83743, 
    34.83757, 34.83773, 34.83793, 34.83818, 34.8384, 34.83857, 34.83875, 
    34.8389,
  34.83717, 34.83718, 34.83722, 34.83726, 34.8373, 34.83735, 34.83741, 
    34.8375, 34.83763, 34.83784, 34.83813, 34.83843, 34.83864, 34.83877, 
    34.83894,
  34.83722, 34.83723, 34.83727, 34.8373, 34.83734, 34.83738, 34.83743, 
    34.83747, 34.83755, 34.83771, 34.83801, 34.83835, 34.83859, 34.8387, 
    34.839,
  34.83727, 34.83728, 34.83731, 34.83735, 34.83738, 34.83741, 34.83746, 
    34.8375, 34.83756, 34.83771, 34.83798, 34.83833, 34.8386, 34.83882, 
    34.8392,
  34.83732, 34.83734, 34.83736, 34.83739, 34.83743, 34.83746, 34.83751, 
    34.83756, 34.83765, 34.83781, 34.83808, 34.83842, 34.83871, 34.83891, 
    34.83889,
  34.83737, 34.83739, 34.83742, 34.83745, 34.83749, 34.83752, 34.83756, 
    34.83763, 34.83774, 34.83792, 34.8382, 34.83852, 34.83876, 34.8389, 
    34.83902,
  34.83743, 34.83745, 34.83748, 34.83752, 34.83755, 34.83758, 34.83762, 
    34.83772, 34.83784, 34.83804, 34.83829, 34.83856, 34.83873, 34.83877, 
    34.83863,
  34.84045, 34.8405, 34.84058, 34.84068, 34.84081, 34.84095, 34.84112, 
    34.8413, 34.84145, 34.84157, 34.84165, 34.84172, 34.84177, 34.84184, 
    34.84192,
  34.84053, 34.84059, 34.84068, 34.8408, 34.84093, 34.84109, 34.84127, 
    34.84146, 34.84163, 34.84177, 34.8419, 34.84201, 34.84209, 34.84216, 
    34.8422,
  34.84059, 34.84066, 34.84075, 34.84087, 34.841, 34.84115, 34.84133, 
    34.84152, 34.8417, 34.84189, 34.84209, 34.84228, 34.84243, 34.84255, 
    34.84259,
  34.84062, 34.84069, 34.84078, 34.8409, 34.84101, 34.84114, 34.84128, 
    34.84145, 34.84163, 34.84185, 34.84212, 34.8424, 34.8426, 34.84272, 
    34.84274,
  34.84064, 34.84071, 34.84079, 34.84089, 34.84099, 34.8411, 34.8412, 
    34.8413, 34.84141, 34.84161, 34.84192, 34.84232, 34.84262, 34.8428, 
    34.84262,
  34.84064, 34.8407, 34.84077, 34.84086, 34.84095, 34.84104, 34.84112, 
    34.84118, 34.84124, 34.84135, 34.84163, 34.84214, 34.84258, 34.8428, 
    34.84242,
  34.84064, 34.84069, 34.84075, 34.84083, 34.84091, 34.84099, 34.84106, 
    34.84111, 34.84116, 34.84126, 34.84154, 34.84209, 34.84258, 34.84278, 
    34.84243,
  34.84064, 34.84067, 34.84072, 34.84079, 34.84086, 34.84093, 34.841, 
    34.84107, 34.84113, 34.84126, 34.84157, 34.84213, 34.84261, 34.84277, 
    34.84189,
  34.84064, 34.84066, 34.8407, 34.84076, 34.84083, 34.84091, 34.84098, 
    34.84104, 34.84111, 34.84129, 34.84166, 34.8422, 34.84259, 34.8427, 
    34.84231,
  34.84065, 34.84067, 34.84072, 34.84078, 34.84085, 34.84092, 34.84096, 
    34.84102, 34.84113, 34.84133, 34.84169, 34.84215, 34.84245, 34.84242, 
    34.84211,
  34.84324, 34.84328, 34.84334, 34.8434, 34.84347, 34.84355, 34.84363, 
    34.8437, 34.84376, 34.84378, 34.84378, 34.84378, 34.84382, 34.84391, 
    34.84399,
  34.84331, 34.84336, 34.84342, 34.84349, 34.84357, 34.84366, 34.84375, 
    34.84384, 34.84391, 34.84396, 34.844, 34.84402, 34.84408, 34.84414, 
    34.84417,
  34.84336, 34.84341, 34.84348, 34.84355, 34.84364, 34.84373, 34.84383, 
    34.84392, 34.84401, 34.8441, 34.84419, 34.84428, 34.84434, 34.84437, 
    34.84436,
  34.8434, 34.84345, 34.84351, 34.84359, 34.84367, 34.84376, 34.84385, 
    34.84393, 34.84402, 34.84414, 34.84429, 34.84447, 34.84457, 34.84457, 
    34.84452,
  34.84342, 34.84347, 34.84354, 34.84361, 34.84369, 34.84378, 34.84385, 
    34.84391, 34.84396, 34.84404, 34.84423, 34.84456, 34.8448, 34.84479, 
    34.84454,
  34.84344, 34.84349, 34.84356, 34.84363, 34.8437, 34.84378, 34.84385, 
    34.84389, 34.84392, 34.84396, 34.84412, 34.84451, 34.84492, 34.84496, 
    34.84428,
  34.84346, 34.8435, 34.84356, 34.84362, 34.84369, 34.84377, 34.84383, 
    34.84387, 34.84389, 34.84394, 34.8441, 34.84451, 34.84498, 34.84502, 
    34.8437,
  34.84347, 34.8435, 34.84354, 34.8436, 34.84367, 34.84373, 34.84379, 
    34.84384, 34.84388, 34.84395, 34.84414, 34.84458, 34.84504, 34.84518, 
    34.84221,
  34.84348, 34.84349, 34.84353, 34.84359, 34.84364, 34.8437, 34.84375, 
    34.84381, 34.84388, 34.84398, 34.84422, 34.84467, 34.84507, 34.84526, 
    34.84521,
  34.84349, 34.84351, 34.84356, 34.84361, 34.84366, 34.84373, 34.8438, 
    34.84384, 34.84391, 34.84405, 34.84433, 34.8447, 34.84498, 34.8451, 
    34.84487,
  34.84626, 34.84621, 34.84616, 34.8461, 34.84604, 34.84597, 34.8459, 
    34.84583, 34.84575, 34.84566, 34.84557, 34.84547, 34.84536, 34.8453, 
    34.84531,
  34.84623, 34.84619, 34.84615, 34.84609, 34.84603, 34.84595, 34.84586, 
    34.84579, 34.84571, 34.84563, 34.84552, 34.84541, 34.84532, 34.84526, 
    34.84527,
  34.84622, 34.84618, 34.84615, 34.84611, 34.84605, 34.84597, 34.8459, 
    34.84584, 34.8458, 34.84575, 34.84568, 34.8456, 34.84548, 34.84536, 
    34.84527,
  34.84623, 34.8462, 34.84617, 34.84614, 34.8461, 34.84605, 34.84599, 
    34.84595, 34.84592, 34.84592, 34.84593, 34.84595, 34.84591, 34.8457, 
    34.84541,
  34.84624, 34.84621, 34.8462, 34.84619, 34.84617, 34.84614, 34.8461, 
    34.84605, 34.84603, 34.84603, 34.84609, 34.8462, 34.8463, 34.84599, 
    34.84536,
  34.84624, 34.84623, 34.84623, 34.84623, 34.84623, 34.84622, 34.84619, 
    34.84615, 34.84612, 34.84613, 34.84619, 34.84635, 34.84655, 34.84623, 
    34.84463,
  34.84623, 34.84622, 34.84623, 34.84624, 34.84626, 34.84627, 34.84626, 
    34.84624, 34.84623, 34.84624, 34.84631, 34.84649, 34.84673, 34.8465, 
    34.84397,
  34.84621, 34.8462, 34.84621, 34.84623, 34.84626, 34.84629, 34.8463, 
    34.8463, 34.84631, 34.84634, 34.84642, 34.84663, 34.84687, 34.84682, 
    34.84222,
  34.84622, 34.8462, 34.8462, 34.84622, 34.84626, 34.84628, 34.8463, 
    34.84633, 34.84637, 34.84643, 34.84654, 34.84679, 34.847, 34.84708, 
    34.84597,
  34.84623, 34.84621, 34.84622, 34.84626, 34.84629, 34.84631, 34.84636, 
    34.84641, 34.84645, 34.84652, 34.84665, 34.84689, 34.84705, 34.84719, 
    34.84748,
  34.84874, 34.84859, 34.84842, 34.84824, 34.84806, 34.84789, 34.84774, 
    34.84762, 34.8475, 34.8474, 34.84728, 34.84717, 34.84702, 34.84684, 
    34.84672,
  34.84861, 34.84846, 34.8483, 34.84813, 34.84794, 34.84775, 34.84755, 
    34.84739, 34.84723, 34.84707, 34.84691, 34.84679, 34.84673, 34.84666, 
    34.8466,
  34.84855, 34.8484, 34.84825, 34.8481, 34.84793, 34.84773, 34.84752, 
    34.84731, 34.84711, 34.84694, 34.84679, 34.8467, 34.84672, 34.84665, 
    34.84655,
  34.84855, 34.84841, 34.84827, 34.84813, 34.84798, 34.84782, 34.84761, 
    34.84739, 34.8472, 34.84707, 34.847, 34.84706, 34.84721, 34.84713, 
    34.84693,
  34.84859, 34.84845, 34.84833, 34.84821, 34.84809, 34.84796, 34.84779, 
    34.84757, 34.84737, 34.84725, 34.84723, 34.84738, 34.84757, 34.84755, 
    34.84644,
  34.84861, 34.8485, 34.8484, 34.84831, 34.84821, 34.8481, 34.84795, 
    34.84775, 34.84754, 34.84743, 34.84745, 34.84762, 34.84782, 34.84784, 
    34.84463,
  34.84862, 34.84853, 34.84845, 34.84837, 34.84829, 34.84819, 34.84807, 
    34.84792, 34.84774, 34.84768, 34.84772, 34.84791, 34.84807, 34.84811, 
    34.84397,
  34.84863, 34.84855, 34.84848, 34.84843, 34.84836, 34.84827, 34.84817, 
    34.84807, 34.84798, 34.84797, 34.84803, 34.84819, 34.84828, 34.84833, 
    34.84222,
  34.84866, 34.84859, 34.84853, 34.84848, 34.84845, 34.8484, 34.84835, 
    34.8483, 34.84828, 34.8483, 34.84836, 34.84843, 34.84849, 34.8486, 
    34.84598,
  34.84869, 34.84864, 34.84858, 34.84858, 34.8486, 34.84861, 34.84856, 
    34.84849, 34.8485, 34.84854, 34.84865, 34.84874, 34.84877, 34.84887, 
    34.84837,
  34.85201, 34.85188, 34.85169, 34.85146, 34.8512, 34.85095, 34.85073, 
    34.85055, 34.85038, 34.85018, 34.84994, 34.84971, 34.84951, 34.84926, 
    34.84899,
  34.85184, 34.85167, 34.85149, 34.85128, 34.85103, 34.85076, 34.8505, 
    34.85027, 34.85006, 34.84983, 34.84957, 34.84935, 34.84925, 34.84917, 
    34.84902,
  34.85175, 34.85156, 34.85138, 34.85119, 34.85099, 34.85075, 34.85048, 
    34.8502, 34.84992, 34.84964, 34.84937, 34.84919, 34.84921, 34.84911, 
    34.84896,
  34.85173, 34.85153, 34.85135, 34.85118, 34.85102, 34.85084, 34.85062, 
    34.85034, 34.85004, 34.84974, 34.84951, 34.84945, 34.84963, 34.84955, 
    34.8494,
  34.85174, 34.85156, 34.85139, 34.85125, 34.8511, 34.85096, 34.8508, 
    34.85057, 34.85027, 34.84991, 34.8497, 34.84978, 34.84998, 34.84981, 
    34.84662,
  34.85172, 34.85156, 34.85141, 34.85128, 34.85117, 34.85104, 34.8509, 
    34.85071, 34.85044, 34.85009, 34.84993, 34.85004, 34.85029, 34.85011, 
    34.84463,
  34.85168, 34.85154, 34.85141, 34.85128, 34.85116, 34.85103, 34.85089, 
    34.85072, 34.8505, 34.85024, 34.85019, 34.85035, 34.85057, 34.85046, 
    34.84397,
  34.85166, 34.85151, 34.85139, 34.85127, 34.85117, 34.85103, 34.85089, 
    34.85074, 34.8506, 34.8505, 34.85052, 34.85062, 34.85078, 34.85071, 
    34.84222,
  34.85165, 34.85152, 34.8514, 34.8513, 34.85125, 34.85114, 34.85102, 
    34.85089, 34.85082, 34.85085, 34.85092, 34.85096, 34.85098, 34.85087, 
    34.84598,
  34.85163, 34.85151, 34.85142, 34.85134, 34.85134, 34.8513, 34.85123, 
    34.85116, 34.85117, 34.85126, 34.85129, 34.85125, 34.85095, 34.85129, 
    34.84838,
  34.85669, 34.85645, 34.85617, 34.85576, 34.85525, 34.85471, 34.85418, 
    34.85371, 34.85331, 34.85289, 34.85245, 34.85204, 34.85169, 34.85136, 
    34.85107,
  34.85637, 34.85605, 34.85573, 34.85536, 34.85491, 34.85437, 34.85382, 
    34.85331, 34.85292, 34.85255, 34.85213, 34.85175, 34.85154, 34.85135, 
    34.85114,
  34.8562, 34.85582, 34.85549, 34.85516, 34.85481, 34.85438, 34.8539, 
    34.85338, 34.8529, 34.85245, 34.85202, 34.85178, 34.85171, 34.85149, 
    34.85126,
  34.85612, 34.85574, 34.85541, 34.85511, 34.85482, 34.85453, 34.8542, 
    34.85378, 34.85324, 34.85271, 34.85226, 34.85212, 34.85213, 34.85167, 
    34.85138,
  34.85605, 34.85571, 34.85539, 34.85509, 34.85484, 34.85462, 34.85438, 
    34.85409, 34.85363, 34.85304, 34.85249, 34.85243, 34.85241, 34.85144, 
    34.84662,
  34.85591, 34.85563, 34.85532, 34.85502, 34.85476, 34.85452, 34.8543, 
    34.85408, 34.85374, 34.85322, 34.85267, 34.8527, 34.85272, 34.85168, 
    34.84463,
  34.85571, 34.8554, 34.85507, 34.8548, 34.85456, 34.8543, 34.85405, 
    34.85384, 34.8536, 34.85321, 34.85286, 34.85299, 34.85298, 34.85156, 
    34.84397,
  34.85554, 34.85519, 34.85488, 34.85468, 34.85446, 34.85418, 34.85385, 
    34.85359, 34.8534, 34.85318, 34.8531, 34.85327, 34.85321, 34.8519, 
    34.84222,
  34.85548, 34.85514, 34.8549, 34.85475, 34.8546, 34.85437, 34.85401, 
    34.85375, 34.85365, 34.85362, 34.85361, 34.85365, 34.85353, 34.85271, 
    34.84598,
  34.85542, 34.85517, 34.85497, 34.85485, 34.85468, 34.85454, 34.85429, 
    34.85418, 34.85406, 34.85394, 34.85392, 34.85382, 34.8534, 34.85247, 
    34.84838,
  34.86066, 34.86025, 34.85991, 34.85939, 34.85865, 34.85782, 34.85702, 
    34.85635, 34.85583, 34.85537, 34.8549, 34.85448, 34.85418, 34.85403, 
    34.85393,
  34.8602, 34.8597, 34.85926, 34.85877, 34.85815, 34.85744, 34.85671, 
    34.85602, 34.85548, 34.85505, 34.85457, 34.85409, 34.85377, 34.85361, 
    34.85359,
  34.86, 34.85944, 34.85897, 34.85854, 34.85807, 34.85754, 34.85695, 
    34.85631, 34.85563, 34.85501, 34.85446, 34.85397, 34.85364, 34.8533, 
    34.85307,
  34.85996, 34.85938, 34.85889, 34.85849, 34.85812, 34.85779, 34.85744, 
    34.85699, 34.85627, 34.85538, 34.85465, 34.85427, 34.85403, 34.8534, 
    34.8527,
  34.85984, 34.85931, 34.85884, 34.85843, 34.85809, 34.8578, 34.85754, 
    34.85726, 34.85677, 34.85591, 34.85511, 34.85468, 34.85441, 34.85328, 
    34.84662,
  34.85954, 34.85911, 34.85867, 34.85824, 34.85786, 34.85751, 34.85722, 
    34.85703, 34.85677, 34.85622, 34.85543, 34.85498, 34.85466, 34.8536, 
    34.84463,
  34.85919, 34.85886, 34.85846, 34.858, 34.85756, 34.85707, 34.85668, 
    34.85651, 34.8564, 34.85601, 34.85538, 34.85524, 34.85487, 34.8516, 
    34.84397,
  34.85897, 34.85852, 34.85807, 34.85772, 34.85739, 34.85675, 34.85631, 
    34.85611, 34.85599, 34.85576, 34.85552, 34.85559, 34.85513, 34.85194, 
    34.84222,
  34.85886, 34.85843, 34.8578, 34.85777, 34.8575, 34.85689, 34.85643, 
    34.85632, 34.85623, 34.85611, 34.856, 34.85585, 34.85522, 34.85315, 
    34.84598,
  34.85856, 34.85832, 34.858, 34.85777, 34.85754, 34.85719, 34.85686, 
    34.85669, 34.85649, 34.85633, 34.85614, 34.85514, 34.8535, 34.85247, 
    34.84838,
  34.86469, 34.86411, 34.86384, 34.86338, 34.86257, 34.86163, 34.86075, 
    34.85994, 34.85931, 34.85888, 34.85848, 34.8581, 34.85793, 34.85804, 
    34.85832,
  34.86416, 34.86351, 34.86306, 34.86257, 34.86191, 34.86117, 34.86044, 
    34.85967, 34.859, 34.85857, 34.8581, 34.85749, 34.85711, 34.85723, 
    34.85775,
  34.864, 34.86325, 34.8627, 34.86224, 34.86177, 34.86125, 34.86074, 
    34.86015, 34.85934, 34.85856, 34.85783, 34.85695, 34.85635, 34.85612, 
    34.85626,
  34.86393, 34.86317, 34.86256, 34.86211, 34.86174, 34.86139, 34.86102, 
    34.86065, 34.86004, 34.85901, 34.85791, 34.85678, 34.85606, 34.85555, 
    34.85464,
  34.86373, 34.86303, 34.86239, 34.86187, 34.86146, 34.86109, 34.8607, 
    34.86047, 34.8602, 34.85952, 34.85841, 34.85717, 34.85649, 34.85577, 
    34.84662,
  34.86327, 34.86273, 34.86217, 34.86157, 34.86094, 34.86034, 34.8599, 
    34.85979, 34.85989, 34.85964, 34.85887, 34.85754, 34.85675, 34.85607, 
    34.84463,
  34.86285, 34.86255, 34.86222, 34.86154, 34.86056, 34.8597, 34.85929, 
    34.8592, 34.85938, 34.85928, 34.85859, 34.85743, 34.85683, 34.8516, 
    34.84397,
  34.86249, 34.86239, 34.86229, 34.86153, 34.86017, 34.85935, 34.85906, 
    34.85892, 34.85887, 34.85867, 34.85817, 34.85752, 34.85717, 34.85194, 
    34.84222,
  34.86206, 34.86201, 34.86198, 34.86115, 34.85987, 34.85932, 34.859, 
    34.85883, 34.85858, 34.85822, 34.85788, 34.8576, 34.85719, 34.85316, 
    34.84598,
  34.86172, 34.86149, 34.86125, 34.86058, 34.85991, 34.85952, 34.85919, 
    34.85892, 34.85863, 34.85829, 34.85781, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.86683, 34.86624, 34.86604, 34.86571, 34.86496, 34.86404, 34.8633, 
    34.86261, 34.86188, 34.86135, 34.86101, 34.86074, 34.86049, 34.86057, 
    34.86104,
  34.86637, 34.86563, 34.8652, 34.86481, 34.86417, 34.86351, 34.86295, 
    34.86236, 34.86169, 34.86119, 34.86087, 34.86049, 34.86039, 34.86074, 
    34.86116,
  34.86633, 34.86537, 34.8648, 34.86439, 34.86395, 34.86351, 34.86306, 
    34.86261, 34.86202, 34.86141, 34.86088, 34.86032, 34.86048, 34.86088, 
    34.86102,
  34.86628, 34.86529, 34.86463, 34.8642, 34.86386, 34.8635, 34.86313, 
    34.8628, 34.8625, 34.86189, 34.86089, 34.86013, 34.86024, 34.86006, 
    34.8601,
  34.86586, 34.86504, 34.86436, 34.86383, 34.8634, 34.86291, 34.86248, 
    34.8622, 34.86227, 34.86212, 34.86108, 34.86035, 34.8605, 34.85934, 
    34.84662,
  34.86534, 34.86478, 34.86412, 34.86343, 34.86263, 34.86192, 34.86156, 
    34.86145, 34.86172, 34.86191, 34.86093, 34.86009, 34.8602, 34.85988, 
    34.84463,
  34.8649, 34.86457, 34.86412, 34.86338, 34.86206, 34.86129, 34.86108, 
    34.86102, 34.86124, 34.86152, 34.86085, 34.85997, 34.85961, 34.8516, 
    34.84397,
  34.86436, 34.86406, 34.86399, 34.86343, 34.8616, 34.86093, 34.86079, 
    34.86084, 34.86093, 34.86088, 34.86031, 34.85978, 34.85934, 34.85194, 
    34.84222,
  34.8637, 34.8634, 34.86356, 34.86292, 34.86126, 34.86087, 34.86069, 
    34.86058, 34.86038, 34.86003, 34.85973, 34.85949, 34.85799, 34.85316, 
    34.84598,
  34.86344, 34.86292, 34.86264, 34.86194, 34.86125, 34.86082, 34.86054, 
    34.86035, 34.86012, 34.85984, 34.85965, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.86985, 34.86932, 34.86918, 34.86894, 34.86834, 34.86757, 34.86705, 
    34.8667, 34.86623, 34.86555, 34.86501, 34.86462, 34.86413, 34.86361, 
    34.86357,
  34.86979, 34.86888, 34.86848, 34.86822, 34.86767, 34.86711, 34.86675, 
    34.86636, 34.86599, 34.86553, 34.86507, 34.86446, 34.86378, 34.86345, 
    34.86333,
  34.87011, 34.86881, 34.86818, 34.86785, 34.86745, 34.86707, 34.86672, 
    34.86635, 34.866, 34.86564, 34.86518, 34.86435, 34.86404, 34.8642, 
    34.86418,
  34.86988, 34.86869, 34.86802, 34.86766, 34.86738, 34.86703, 34.86656, 
    34.86605, 34.86573, 34.86555, 34.86506, 34.86404, 34.86386, 34.86415, 
    34.86431,
  34.86917, 34.86838, 34.86779, 34.86732, 34.86685, 34.86624, 34.8656, 
    34.86513, 34.86504, 34.86533, 34.86499, 34.86339, 34.8627, 34.86378, 
    34.84662,
  34.86862, 34.86814, 34.86752, 34.86668, 34.86573, 34.86504, 34.86465, 
    34.86449, 34.86462, 34.86509, 34.86483, 34.86304, 34.86223, 34.86126, 
    34.84463,
  34.86822, 34.86789, 34.86734, 34.86611, 34.86496, 34.86448, 34.86438, 
    34.86444, 34.86461, 34.86486, 34.86438, 34.8629, 34.86232, 34.8516, 
    34.84397,
  34.86752, 34.86695, 34.86646, 34.86546, 34.86464, 34.86435, 34.8643, 
    34.86438, 34.8644, 34.8642, 34.86338, 34.8627, 34.86226, 34.85194, 
    34.84222,
  34.867, 34.86623, 34.86366, 34.86509, 34.86454, 34.86418, 34.86393, 
    34.86376, 34.86355, 34.86326, 34.86306, 34.86304, 34.85808, 34.85316, 
    34.84598,
  34.8667, 34.86604, 34.86551, 34.86492, 34.86444, 34.86399, 34.86374, 
    34.86362, 34.86337, 34.86303, 34.86014, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87115, 34.87074, 34.87058, 34.87036, 34.8698, 34.86912, 34.86862, 
    34.86834, 34.8681, 34.86781, 34.86741, 34.86705, 34.86656, 34.86609, 
    34.86554,
  34.87162, 34.87057, 34.87012, 34.8699, 34.86939, 34.86885, 34.86849, 
    34.86823, 34.86792, 34.86768, 34.86729, 34.86672, 34.86597, 34.86533, 
    34.86498,
  34.87187, 34.87063, 34.86993, 34.86966, 34.86929, 34.86893, 34.8686, 
    34.86827, 34.8679, 34.86754, 34.86711, 34.86644, 34.86567, 34.86546, 
    34.86577,
  34.87148, 34.87034, 34.86976, 34.8695, 34.86923, 34.86893, 34.86854, 
    34.86811, 34.86763, 34.86723, 34.86681, 34.8661, 34.86593, 34.86612, 
    34.8662,
  34.87075, 34.86998, 34.86952, 34.86914, 34.86865, 34.86823, 34.86777, 
    34.86728, 34.86691, 34.86684, 34.86686, 34.86617, 34.86277, 34.8643, 
    34.84662,
  34.8703, 34.8698, 34.86926, 34.86848, 34.86778, 34.86745, 34.86711, 
    34.86675, 34.86654, 34.8667, 34.86687, 34.86631, 34.86582, 34.86133, 
    34.84463,
  34.86998, 34.86962, 34.86899, 34.86798, 34.8674, 34.86723, 34.86701, 
    34.86669, 34.86648, 34.86663, 34.86668, 34.86622, 34.86547, 34.8516, 
    34.84397,
  34.86972, 34.8693, 34.86872, 34.86794, 34.86737, 34.86717, 34.86697, 
    34.86671, 34.86654, 34.8665, 34.86642, 34.86598, 34.86443, 34.85194, 
    34.84222,
  34.8698, 34.86954, 34.86366, 34.86809, 34.86748, 34.8672, 34.86699, 
    34.8668, 34.8667, 34.86672, 34.86656, 34.86642, 34.85808, 34.85316, 
    34.84598,
  34.86974, 34.86927, 34.86889, 34.86816, 34.86773, 34.86758, 34.86755, 
    34.86742, 34.86732, 34.86771, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87171, 34.87134, 34.87115, 34.87094, 34.87048, 34.86996, 34.86958, 
    34.86943, 34.86951, 34.86957, 34.86933, 34.86872, 34.86831, 34.86816, 
    34.86793,
  34.87211, 34.87134, 34.87088, 34.87062, 34.87016, 34.86972, 34.86945, 
    34.86923, 34.8692, 34.86906, 34.86884, 34.8683, 34.86736, 34.86693, 
    34.86747,
  34.87216, 34.8713, 34.87074, 34.87048, 34.8701, 34.86979, 34.86956, 
    34.86932, 34.86918, 34.86886, 34.86838, 34.86763, 34.86703, 34.86718, 
    34.86806,
  34.87183, 34.87088, 34.87046, 34.87028, 34.87004, 34.86979, 34.86956, 
    34.86928, 34.86905, 34.86873, 34.86835, 34.86781, 34.86771, 34.86724, 
    34.86717,
  34.87131, 34.87057, 34.8702, 34.86997, 34.8697, 34.86941, 34.86916, 
    34.86887, 34.86858, 34.86832, 34.86837, 34.86843, 34.86277, 34.86431, 
    34.84662,
  34.87095, 34.87045, 34.87008, 34.86971, 34.86929, 34.86907, 34.86882, 
    34.86836, 34.86819, 34.86821, 34.86847, 34.86892, 34.86874, 34.86133, 
    34.84463,
  34.87077, 34.8705, 34.87023, 34.86973, 34.86916, 34.86898, 34.86878, 
    34.86833, 34.86822, 34.86829, 34.86864, 34.86911, 34.86754, 34.8516, 
    34.84397,
  34.87074, 34.87055, 34.87033, 34.86981, 34.86925, 34.86899, 34.86877, 
    34.86842, 34.86832, 34.8685, 34.86881, 34.86903, 34.86523, 34.85194, 
    34.84222,
  34.87095, 34.87086, 34.86366, 34.86996, 34.86945, 34.86927, 34.86926, 
    34.86919, 34.86921, 34.86934, 34.8693, 34.8679, 34.85808, 34.85316, 
    34.84598,
  34.87119, 34.87085, 34.87044, 34.87008, 34.86977, 34.86986, 34.87002, 
    34.86989, 34.86921, 34.86953, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87204, 34.87187, 34.87168, 34.8716, 34.87147, 34.87137, 34.87129, 
    34.87119, 34.8713, 34.87144, 34.87112, 34.87084, 34.87029, 34.86988, 
    34.86995,
  34.87219, 34.87199, 34.87166, 34.87145, 34.87128, 34.87108, 34.87095, 
    34.87106, 34.87122, 34.87144, 34.87086, 34.8698, 34.86935, 34.86923, 
    34.86964,
  34.87226, 34.87199, 34.87165, 34.87141, 34.87121, 34.87099, 34.87085, 
    34.87079, 34.87082, 34.87098, 34.87042, 34.8698, 34.86938, 34.8695, 
    34.86942,
  34.87214, 34.87173, 34.87152, 34.87134, 34.8711, 34.87086, 34.87072, 
    34.87069, 34.87054, 34.87038, 34.87013, 34.8705, 34.87077, 34.86738, 
    34.86717,
  34.8719, 34.87144, 34.87127, 34.87118, 34.87098, 34.87083, 34.87077, 
    34.87074, 34.87062, 34.87028, 34.87037, 34.87117, 34.86277, 34.86431, 
    34.84662,
  34.87177, 34.87137, 34.87121, 34.87114, 34.87097, 34.87083, 34.8708, 
    34.87082, 34.87073, 34.87053, 34.87077, 34.87138, 34.86932, 34.86133, 
    34.84463,
  34.87173, 34.87151, 34.87139, 34.87128, 34.87099, 34.87091, 34.86894, 
    34.87083, 34.87082, 34.87098, 34.87109, 34.87109, 34.86936, 34.8516, 
    34.84397,
  34.87174, 34.87167, 34.87161, 34.87135, 34.8711, 34.8712, 34.87116, 
    34.87107, 34.87111, 34.87122, 34.87098, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.8718, 34.87154, 34.86366, 34.87135, 34.87135, 34.87163, 34.87168, 
    34.87164, 34.87121, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87203, 34.87179, 34.8716, 34.87152, 34.87169, 34.87204, 34.87249, 
    34.87169, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87234, 34.87227, 34.87215, 34.87214, 34.87222, 34.87227, 34.87231, 
    34.87228, 34.87235, 34.87244, 34.87224, 34.87164, 34.87073, 34.86993, 
    34.87001,
  34.87243, 34.87244, 34.87234, 34.87224, 34.87228, 34.87223, 34.87213, 
    34.87191, 34.87199, 34.87225, 34.87218, 34.87134, 34.87036, 34.86978, 
    34.86967,
  34.87248, 34.87243, 34.87232, 34.87231, 34.87228, 34.8721, 34.87195, 
    34.87186, 34.8718, 34.87199, 34.87208, 34.87154, 34.87165, 34.87137, 
    34.86942,
  34.87241, 34.87231, 34.87228, 34.87232, 34.87221, 34.87197, 34.87186, 
    34.87194, 34.87189, 34.8719, 34.872, 34.87196, 34.87194, 34.86738, 
    34.86717,
  34.87241, 34.87227, 34.87222, 34.87224, 34.87216, 34.87209, 34.87203, 
    34.87197, 34.87193, 34.87197, 34.87211, 34.87172, 34.86277, 34.86431, 
    34.84662,
  34.87242, 34.87235, 34.87227, 34.87221, 34.87221, 34.87234, 34.87228, 
    34.8717, 34.87202, 34.87202, 34.8721, 34.87162, 34.86932, 34.86133, 
    34.84463,
  34.8724, 34.8725, 34.87249, 34.87241, 34.87246, 34.87255, 34.86894, 
    34.87193, 34.87212, 34.87205, 34.87198, 34.87109, 34.86938, 34.8516, 
    34.84397,
  34.87263, 34.87243, 34.87186, 34.87251, 34.87292, 34.87326, 34.87284, 
    34.87238, 34.87195, 34.87188, 34.87099, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.87277, 34.87161, 34.86366, 34.8724, 34.87335, 34.87366, 34.87381, 
    34.87271, 34.87143, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87305, 34.87294, 34.87284, 34.87263, 34.87321, 34.87379, 34.87362, 
    34.87173, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87234, 34.87227, 34.87215, 34.87214, 34.87223, 34.87227, 34.87232, 
    34.87229, 34.87235, 34.87244, 34.87224, 34.87164, 34.87073, 34.86993, 
    34.87001,
  34.87243, 34.87245, 34.87234, 34.87224, 34.87228, 34.87223, 34.87213, 
    34.87191, 34.87199, 34.87226, 34.87218, 34.87134, 34.87038, 34.86978, 
    34.86967,
  34.87248, 34.87243, 34.87232, 34.87231, 34.87228, 34.8721, 34.87195, 
    34.87186, 34.87181, 34.87202, 34.8721, 34.87154, 34.87165, 34.87137, 
    34.86942,
  34.87241, 34.87231, 34.87229, 34.87232, 34.87221, 34.87197, 34.87186, 
    34.87194, 34.87189, 34.8719, 34.872, 34.87197, 34.87194, 34.86738, 
    34.86717,
  34.87241, 34.87227, 34.87222, 34.87224, 34.87216, 34.87209, 34.87203, 
    34.87197, 34.87193, 34.87197, 34.87212, 34.87172, 34.86277, 34.86431, 
    34.84662,
  34.87242, 34.87235, 34.87227, 34.87221, 34.87221, 34.87234, 34.87228, 
    34.87171, 34.87202, 34.87203, 34.8721, 34.87162, 34.86932, 34.86133, 
    34.84463,
  34.8724, 34.8725, 34.87249, 34.87242, 34.87246, 34.87255, 34.86894, 
    34.87193, 34.87213, 34.87205, 34.87198, 34.87109, 34.86938, 34.8516, 
    34.84397,
  34.87263, 34.87243, 34.87186, 34.87252, 34.87299, 34.87476, 34.87285, 
    34.87238, 34.87195, 34.87188, 34.87099, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.87277, 34.87161, 34.86366, 34.87242, 34.87455, 34.87531, 34.87498, 
    34.87273, 34.87143, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87306, 34.87294, 34.87285, 34.87263, 34.87331, 34.8745, 34.87363, 
    34.87173, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87234, 34.87227, 34.87215, 34.87214, 34.87223, 34.87227, 34.87232, 
    34.87229, 34.87235, 34.87244, 34.87224, 34.87164, 34.87073, 34.86993, 
    34.87001,
  34.87243, 34.87245, 34.87234, 34.87224, 34.87228, 34.87223, 34.87213, 
    34.87191, 34.87199, 34.87226, 34.87218, 34.87134, 34.87038, 34.86978, 
    34.86967,
  34.87248, 34.87243, 34.87232, 34.87231, 34.87228, 34.8721, 34.87195, 
    34.87186, 34.87181, 34.87202, 34.8721, 34.87154, 34.87165, 34.87137, 
    34.86942,
  34.87241, 34.87231, 34.87229, 34.87232, 34.87221, 34.87197, 34.87186, 
    34.87194, 34.87189, 34.8719, 34.872, 34.87197, 34.87194, 34.86738, 
    34.86717,
  34.87241, 34.87227, 34.87222, 34.87224, 34.87216, 34.87209, 34.87203, 
    34.87197, 34.87193, 34.87197, 34.87212, 34.87172, 34.86277, 34.86431, 
    34.84662,
  34.87242, 34.87235, 34.87227, 34.87221, 34.87221, 34.87234, 34.87228, 
    34.87171, 34.87202, 34.87203, 34.8721, 34.87162, 34.86932, 34.86133, 
    34.84463,
  34.8724, 34.8725, 34.87249, 34.87242, 34.87246, 34.87255, 34.86894, 
    34.87193, 34.87213, 34.87205, 34.87198, 34.87109, 34.86938, 34.8516, 
    34.84397,
  34.87263, 34.87243, 34.87186, 34.87252, 34.87299, 34.87476, 34.87285, 
    34.87238, 34.87195, 34.87188, 34.87099, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.87277, 34.87161, 34.86366, 34.87242, 34.87455, 34.87531, 34.87498, 
    34.87273, 34.87143, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87306, 34.87294, 34.87285, 34.87263, 34.87331, 34.8745, 34.87363, 
    34.87173, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87234, 34.87227, 34.87215, 34.87214, 34.87223, 34.87227, 34.87232, 
    34.87229, 34.87235, 34.87244, 34.87224, 34.87164, 34.87073, 34.86993, 
    34.87001,
  34.87243, 34.87245, 34.87234, 34.87224, 34.87228, 34.87223, 34.87213, 
    34.87191, 34.87199, 34.87226, 34.87218, 34.87134, 34.87038, 34.86978, 
    34.86967,
  34.87248, 34.87243, 34.87232, 34.87231, 34.87228, 34.8721, 34.87195, 
    34.87186, 34.87181, 34.87202, 34.8721, 34.87154, 34.87165, 34.87137, 
    34.86942,
  34.87241, 34.87231, 34.87229, 34.87232, 34.87221, 34.87197, 34.87186, 
    34.87194, 34.87189, 34.8719, 34.872, 34.87197, 34.87194, 34.86738, 
    34.86717,
  34.87241, 34.87227, 34.87222, 34.87224, 34.87216, 34.87209, 34.87203, 
    34.87197, 34.87193, 34.87197, 34.87212, 34.87172, 34.86277, 34.86431, 
    34.84662,
  34.87242, 34.87235, 34.87227, 34.87221, 34.87221, 34.87234, 34.87228, 
    34.87171, 34.87202, 34.87203, 34.8721, 34.87162, 34.86932, 34.86133, 
    34.84463,
  34.8724, 34.8725, 34.87249, 34.87242, 34.87246, 34.87255, 34.86894, 
    34.87193, 34.87213, 34.87205, 34.87198, 34.87109, 34.86938, 34.8516, 
    34.84397,
  34.87263, 34.87243, 34.87186, 34.87252, 34.87299, 34.87476, 34.87285, 
    34.87238, 34.87195, 34.87188, 34.87099, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.87277, 34.87161, 34.86366, 34.87242, 34.87455, 34.87531, 34.87498, 
    34.87273, 34.87143, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87306, 34.87294, 34.87285, 34.87263, 34.87331, 34.8745, 34.87363, 
    34.87173, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87234, 34.87227, 34.87215, 34.87214, 34.87223, 34.87227, 34.87232, 
    34.87229, 34.87235, 34.87244, 34.87224, 34.87164, 34.87073, 34.86993, 
    34.87001,
  34.87243, 34.87245, 34.87234, 34.87224, 34.87228, 34.87223, 34.87213, 
    34.87191, 34.87199, 34.87226, 34.87218, 34.87134, 34.87038, 34.86978, 
    34.86967,
  34.87248, 34.87243, 34.87232, 34.87231, 34.87228, 34.8721, 34.87195, 
    34.87186, 34.87181, 34.87202, 34.8721, 34.87154, 34.87165, 34.87137, 
    34.86942,
  34.87241, 34.87231, 34.87229, 34.87232, 34.87221, 34.87197, 34.87186, 
    34.87194, 34.87189, 34.8719, 34.872, 34.87197, 34.87194, 34.86738, 
    34.86717,
  34.87241, 34.87227, 34.87222, 34.87224, 34.87216, 34.87209, 34.87203, 
    34.87197, 34.87193, 34.87197, 34.87212, 34.87172, 34.86277, 34.86431, 
    34.84662,
  34.87242, 34.87235, 34.87227, 34.87221, 34.87221, 34.87234, 34.87228, 
    34.87171, 34.87202, 34.87203, 34.8721, 34.87162, 34.86932, 34.86133, 
    34.84463,
  34.8724, 34.8725, 34.87249, 34.87242, 34.87246, 34.87255, 34.86894, 
    34.87193, 34.87213, 34.87205, 34.87198, 34.87109, 34.86938, 34.8516, 
    34.84397,
  34.87263, 34.87243, 34.87186, 34.87252, 34.87299, 34.87476, 34.87285, 
    34.87238, 34.87195, 34.87188, 34.87099, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.87277, 34.87161, 34.86366, 34.87242, 34.87455, 34.87531, 34.87498, 
    34.87273, 34.87143, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87306, 34.87294, 34.87285, 34.87263, 34.87331, 34.8745, 34.87363, 
    34.87173, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87234, 34.87227, 34.87215, 34.87214, 34.87223, 34.87227, 34.87232, 
    34.87229, 34.87235, 34.87244, 34.87224, 34.87164, 34.87073, 34.86993, 
    34.87001,
  34.87243, 34.87245, 34.87234, 34.87224, 34.87228, 34.87223, 34.87213, 
    34.87191, 34.87199, 34.87226, 34.87218, 34.87134, 34.87038, 34.86978, 
    34.86967,
  34.87248, 34.87243, 34.87232, 34.87231, 34.87228, 34.8721, 34.87195, 
    34.87186, 34.87181, 34.87202, 34.8721, 34.87154, 34.87165, 34.87137, 
    34.86942,
  34.87241, 34.87231, 34.87229, 34.87232, 34.87221, 34.87197, 34.87186, 
    34.87194, 34.87189, 34.8719, 34.872, 34.87197, 34.87194, 34.86738, 
    34.86717,
  34.87241, 34.87227, 34.87222, 34.87224, 34.87216, 34.87209, 34.87203, 
    34.87197, 34.87193, 34.87197, 34.87212, 34.87172, 34.86277, 34.86431, 
    34.84662,
  34.87242, 34.87235, 34.87227, 34.87221, 34.87221, 34.87234, 34.87228, 
    34.87171, 34.87202, 34.87203, 34.8721, 34.87162, 34.86932, 34.86133, 
    34.84463,
  34.8724, 34.8725, 34.87249, 34.87242, 34.87246, 34.87255, 34.86894, 
    34.87193, 34.87213, 34.87205, 34.87198, 34.87109, 34.86938, 34.8516, 
    34.84397,
  34.87263, 34.87243, 34.87186, 34.87252, 34.87299, 34.87476, 34.87285, 
    34.87238, 34.87195, 34.87188, 34.87099, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.87277, 34.87161, 34.86366, 34.87242, 34.87455, 34.87531, 34.87498, 
    34.87273, 34.87143, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87306, 34.87294, 34.87285, 34.87263, 34.87331, 34.8745, 34.87363, 
    34.87173, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87234, 34.87227, 34.87215, 34.87214, 34.87223, 34.87227, 34.87232, 
    34.87229, 34.87235, 34.87244, 34.87224, 34.87164, 34.87073, 34.86993, 
    34.87001,
  34.87243, 34.87245, 34.87234, 34.87224, 34.87228, 34.87223, 34.87213, 
    34.87191, 34.87199, 34.87226, 34.87218, 34.87134, 34.87038, 34.86978, 
    34.86967,
  34.87248, 34.87243, 34.87232, 34.87231, 34.87228, 34.8721, 34.87195, 
    34.87186, 34.87181, 34.87202, 34.8721, 34.87154, 34.87165, 34.87137, 
    34.86942,
  34.87241, 34.87231, 34.87229, 34.87232, 34.87221, 34.87197, 34.87186, 
    34.87194, 34.87189, 34.8719, 34.872, 34.87197, 34.87194, 34.86738, 
    34.86717,
  34.87241, 34.87227, 34.87222, 34.87224, 34.87216, 34.87209, 34.87203, 
    34.87197, 34.87193, 34.87197, 34.87212, 34.87172, 34.86277, 34.86431, 
    34.84662,
  34.87242, 34.87235, 34.87227, 34.87221, 34.87221, 34.87234, 34.87228, 
    34.87171, 34.87202, 34.87203, 34.8721, 34.87162, 34.86932, 34.86133, 
    34.84463,
  34.8724, 34.8725, 34.87249, 34.87242, 34.87246, 34.87255, 34.86894, 
    34.87193, 34.87213, 34.87205, 34.87198, 34.87109, 34.86938, 34.8516, 
    34.84397,
  34.87263, 34.87243, 34.87186, 34.87252, 34.87299, 34.87476, 34.87285, 
    34.87238, 34.87195, 34.87188, 34.87099, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.87277, 34.87161, 34.86366, 34.87242, 34.87455, 34.87531, 34.87498, 
    34.87273, 34.87143, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87306, 34.87294, 34.87285, 34.87263, 34.87331, 34.8745, 34.87363, 
    34.87173, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87234, 34.87227, 34.87215, 34.87214, 34.87223, 34.87227, 34.87232, 
    34.87229, 34.87235, 34.87244, 34.87224, 34.87164, 34.87073, 34.86993, 
    34.87001,
  34.87243, 34.87245, 34.87234, 34.87224, 34.87228, 34.87223, 34.87213, 
    34.87191, 34.87199, 34.87226, 34.87218, 34.87134, 34.87038, 34.86978, 
    34.86967,
  34.87248, 34.87243, 34.87232, 34.87231, 34.87228, 34.8721, 34.87195, 
    34.87186, 34.87181, 34.87202, 34.8721, 34.87154, 34.87165, 34.87137, 
    34.86942,
  34.87241, 34.87231, 34.87229, 34.87232, 34.87221, 34.87197, 34.87186, 
    34.87194, 34.87189, 34.8719, 34.872, 34.87197, 34.87194, 34.86738, 
    34.86717,
  34.87241, 34.87227, 34.87222, 34.87224, 34.87216, 34.87209, 34.87203, 
    34.87197, 34.87193, 34.87197, 34.87212, 34.87172, 34.86277, 34.86431, 
    34.84662,
  34.87242, 34.87235, 34.87227, 34.87221, 34.87221, 34.87234, 34.87228, 
    34.87171, 34.87202, 34.87203, 34.8721, 34.87162, 34.86932, 34.86133, 
    34.84463,
  34.8724, 34.8725, 34.87249, 34.87242, 34.87246, 34.87255, 34.86894, 
    34.87193, 34.87213, 34.87205, 34.87198, 34.87109, 34.86938, 34.8516, 
    34.84397,
  34.87263, 34.87243, 34.87186, 34.87252, 34.87299, 34.87476, 34.87285, 
    34.87238, 34.87195, 34.87188, 34.87099, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.87277, 34.87161, 34.86366, 34.87242, 34.87455, 34.87531, 34.87498, 
    34.87273, 34.87143, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87306, 34.87294, 34.87285, 34.87263, 34.87331, 34.8745, 34.87363, 
    34.87173, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838,
  34.87234, 34.87227, 34.87215, 34.87214, 34.87223, 34.87227, 34.87232, 
    34.87229, 34.87235, 34.87244, 34.87224, 34.87164, 34.87073, 34.86993, 
    34.87001,
  34.87243, 34.87245, 34.87234, 34.87224, 34.87228, 34.87223, 34.87213, 
    34.87191, 34.87199, 34.87226, 34.87218, 34.87134, 34.87038, 34.86978, 
    34.86967,
  34.87248, 34.87243, 34.87232, 34.87231, 34.87228, 34.8721, 34.87195, 
    34.87186, 34.87181, 34.87202, 34.8721, 34.87154, 34.87165, 34.87137, 
    34.86942,
  34.87241, 34.87231, 34.87229, 34.87232, 34.87221, 34.87197, 34.87186, 
    34.87194, 34.87189, 34.8719, 34.872, 34.87197, 34.87194, 34.86738, 
    34.86717,
  34.87241, 34.87227, 34.87222, 34.87224, 34.87216, 34.87209, 34.87203, 
    34.87197, 34.87193, 34.87197, 34.87212, 34.87172, 34.86277, 34.86431, 
    34.84662,
  34.87242, 34.87235, 34.87227, 34.87221, 34.87221, 34.87234, 34.87228, 
    34.87171, 34.87202, 34.87203, 34.8721, 34.87162, 34.86932, 34.86133, 
    34.84463,
  34.8724, 34.8725, 34.87249, 34.87242, 34.87246, 34.87255, 34.86894, 
    34.87193, 34.87213, 34.87205, 34.87198, 34.87109, 34.86938, 34.8516, 
    34.84397,
  34.87263, 34.87243, 34.87186, 34.87252, 34.87299, 34.87476, 34.87285, 
    34.87238, 34.87195, 34.87188, 34.87099, 34.86976, 34.86523, 34.85194, 
    34.84222,
  34.87277, 34.87161, 34.86366, 34.87242, 34.87455, 34.87531, 34.87498, 
    34.87273, 34.87143, 34.87102, 34.87074, 34.86804, 34.85808, 34.85316, 
    34.84598,
  34.87306, 34.87294, 34.87285, 34.87263, 34.87331, 34.8745, 34.87363, 
    34.87173, 34.86929, 34.86967, 34.86018, 34.85518, 34.8535, 34.85247, 
    34.84838 ;

 time_bnds =
  0, 365 ;

 nv = 1, 2 ;

 time = 182.5 ;

 xh = -166.875, -166.625, -166.375, -166.125, -165.875, -165.625, -165.375, 
    -165.125, -164.875, -164.625, -164.375, -164.125, -163.875, -163.625, 
    -163.375 ;

 xq = -300, -299.75, -299.5, -299.25, -299, -298.75, -298.5, -298.25, -298, 
    -297.75, -297.5, -297.25, -297, -296.75, -296.5, -296.25, -296, -295.75, 
    -295.5, -295.25, -295, -294.75, -294.5, -294.25, -294, -293.75, -293.5, 
    -293.25, -293, -292.75, -292.5, -292.25, -292, -291.75, -291.5, -291.25, 
    -291, -290.75, -290.5, -290.25, -290, -289.75, -289.5, -289.25, -289, 
    -288.75, -288.5, -288.25, -288, -287.75, -287.5, -287.25, -287, -286.75, 
    -286.5, -286.25, -286, -285.75, -285.5, -285.25, -285, -284.75, -284.5, 
    -284.25, -284, -283.75, -283.5, -283.25, -283, -282.75, -282.5, -282.25, 
    -282, -281.75, -281.5, -281.25, -281, -280.75, -280.5, -280.25, -280, 
    -279.75, -279.5, -279.25, -279, -278.75, -278.5, -278.25, -278, -277.75, 
    -277.5, -277.25, -277, -276.75, -276.5, -276.25, -276, -275.75, -275.5, 
    -275.25, -275, -274.75, -274.5, -274.25, -274, -273.75, -273.5, -273.25, 
    -273, -272.75, -272.5, -272.25, -272, -271.75, -271.5, -271.25, -271, 
    -270.75, -270.5, -270.25, -270, -269.75, -269.5, -269.25, -269, -268.75, 
    -268.5, -268.25, -268, -267.75, -267.5, -267.25, -267, -266.75, -266.5, 
    -266.25, -266, -265.75, -265.5, -265.25, -265, -264.75, -264.5, -264.25, 
    -264, -263.75, -263.5, -263.25, -263, -262.75, -262.5, -262.25, -262, 
    -261.75, -261.5, -261.25, -261, -260.75, -260.5, -260.25, -260, -259.75, 
    -259.5, -259.25, -259, -258.75, -258.5, -258.25, -258, -257.75, -257.5, 
    -257.25, -257, -256.75, -256.5, -256.25, -256, -255.75, -255.5, -255.25, 
    -255, -254.75, -254.5, -254.25, -254, -253.75, -253.5, -253.25, -253, 
    -252.75, -252.5, -252.25, -252, -251.75, -251.5, -251.25, -251, -250.75, 
    -250.5, -250.25, -250, -249.75, -249.5, -249.25, -249, -248.75, -248.5, 
    -248.25, -248, -247.75, -247.5, -247.25, -247, -246.75, -246.5, -246.25, 
    -246, -245.75, -245.5, -245.25, -245, -244.75, -244.5, -244.25, -244, 
    -243.75, -243.5, -243.25, -243, -242.75, -242.5, -242.25, -242, -241.75, 
    -241.5, -241.25, -241, -240.75, -240.5, -240.25, -240, -239.75, -239.5, 
    -239.25, -239, -238.75, -238.5, -238.25, -238, -237.75, -237.5, -237.25, 
    -237, -236.75, -236.5, -236.25, -236, -235.75, -235.5, -235.25, -235, 
    -234.75, -234.5, -234.25, -234, -233.75, -233.5, -233.25, -233, -232.75, 
    -232.5, -232.25, -232, -231.75, -231.5, -231.25, -231, -230.75, -230.5, 
    -230.25, -230, -229.75, -229.5, -229.25, -229, -228.75, -228.5, -228.25, 
    -228, -227.75, -227.5, -227.25, -227, -226.75, -226.5, -226.25, -226, 
    -225.75, -225.5, -225.25, -225, -224.75, -224.5, -224.25, -224, -223.75, 
    -223.5, -223.25, -223, -222.75, -222.5, -222.25, -222, -221.75, -221.5, 
    -221.25, -221, -220.75, -220.5, -220.25, -220, -219.75, -219.5, -219.25, 
    -219, -218.75, -218.5, -218.25, -218, -217.75, -217.5, -217.25, -217, 
    -216.75, -216.5, -216.25, -216, -215.75, -215.5, -215.25, -215, -214.75, 
    -214.5, -214.25, -214, -213.75, -213.5, -213.25, -213, -212.75, -212.5, 
    -212.25, -212, -211.75, -211.5, -211.25, -211, -210.75, -210.5, -210.25, 
    -210, -209.75, -209.5, -209.25, -209, -208.75, -208.5, -208.25, -208, 
    -207.75, -207.5, -207.25, -207, -206.75, -206.5, -206.25, -206, -205.75, 
    -205.5, -205.25, -205, -204.75, -204.5, -204.25, -204, -203.75, -203.5, 
    -203.25, -203, -202.75, -202.5, -202.25, -202, -201.75, -201.5, -201.25, 
    -201, -200.75, -200.5, -200.25, -200, -199.75, -199.5, -199.25, -199, 
    -198.75, -198.5, -198.25, -198, -197.75, -197.5, -197.25, -197, -196.75, 
    -196.5, -196.25, -196, -195.75, -195.5, -195.25, -195, -194.75, -194.5, 
    -194.25, -194, -193.75, -193.5, -193.25, -193, -192.75, -192.5, -192.25, 
    -192, -191.75, -191.5, -191.25, -191, -190.75, -190.5, -190.25, -190, 
    -189.75, -189.5, -189.25, -189, -188.75, -188.5, -188.25, -188, -187.75, 
    -187.5, -187.25, -187, -186.75, -186.5, -186.25, -186, -185.75, -185.5, 
    -185.25, -185, -184.75, -184.5, -184.25, -184, -183.75, -183.5, -183.25, 
    -183, -182.75, -182.5, -182.25, -182, -181.75, -181.5, -181.25, -181, 
    -180.75, -180.5, -180.25, -180, -179.75, -179.5, -179.25, -179, -178.75, 
    -178.5, -178.25, -178, -177.75, -177.5, -177.25, -177, -176.75, -176.5, 
    -176.25, -176, -175.75, -175.5, -175.25, -175, -174.75, -174.5, -174.25, 
    -174, -173.75, -173.5, -173.25, -173, -172.75, -172.5, -172.25, -172, 
    -171.75, -171.5, -171.25, -171, -170.75, -170.5, -170.25, -170, -169.75, 
    -169.5, -169.25, -169, -168.75, -168.5, -168.25, -168, -167.75, -167.5, 
    -167.25, -167, -166.75, -166.5, -166.25, -166, -165.75, -165.5, -165.25, 
    -165, -164.75, -164.5, -164.25, -164, -163.75, -163.5, -163.25, -163, 
    -162.75, -162.5, -162.25, -162, -161.75, -161.5, -161.25, -161, -160.75, 
    -160.5, -160.25, -160, -159.75, -159.5, -159.25, -159, -158.75, -158.5, 
    -158.25, -158, -157.75, -157.5, -157.25, -157, -156.75, -156.5, -156.25, 
    -156, -155.75, -155.5, -155.25, -155, -154.75, -154.5, -154.25, -154, 
    -153.75, -153.5, -153.25, -153, -152.75, -152.5, -152.25, -152, -151.75, 
    -151.5, -151.25, -151, -150.75, -150.5, -150.25, -150, -149.75, -149.5, 
    -149.25, -149, -148.75, -148.5, -148.25, -148, -147.75, -147.5, -147.25, 
    -147, -146.75, -146.5, -146.25, -146, -145.75, -145.5, -145.25, -145, 
    -144.75, -144.5, -144.25, -144, -143.75, -143.5, -143.25, -143, -142.75, 
    -142.5, -142.25, -142, -141.75, -141.5, -141.25, -141, -140.75, -140.5, 
    -140.25, -140, -139.75, -139.5, -139.25, -139, -138.75, -138.5, -138.25, 
    -138, -137.75, -137.5, -137.25, -137, -136.75, -136.5, -136.25, -136, 
    -135.75, -135.5, -135.25, -135, -134.75, -134.5, -134.25, -134, -133.75, 
    -133.5, -133.25, -133, -132.75, -132.5, -132.25, -132, -131.75, -131.5, 
    -131.25, -131, -130.75, -130.5, -130.25, -130, -129.75, -129.5, -129.25, 
    -129, -128.75, -128.5, -128.25, -128, -127.75, -127.5, -127.25, -127, 
    -126.75, -126.5, -126.25, -126, -125.75, -125.5, -125.25, -125, -124.75, 
    -124.5, -124.25, -124, -123.75, -123.5, -123.25, -123, -122.75, -122.5, 
    -122.25, -122, -121.75, -121.5, -121.25, -121, -120.75, -120.5, -120.25, 
    -120, -119.75, -119.5, -119.25, -119, -118.75, -118.5, -118.25, -118, 
    -117.75, -117.5, -117.25, -117, -116.75, -116.5, -116.25, -116, -115.75, 
    -115.5, -115.25, -115, -114.75, -114.5, -114.25, -114, -113.75, -113.5, 
    -113.25, -113, -112.75, -112.5, -112.25, -112, -111.75, -111.5, -111.25, 
    -111, -110.75, -110.5, -110.25, -110, -109.75, -109.5, -109.25, -109, 
    -108.75, -108.5, -108.25, -108, -107.75, -107.5, -107.25, -107, -106.75, 
    -106.5, -106.25, -106, -105.75, -105.5, -105.25, -105, -104.75, -104.5, 
    -104.25, -104, -103.75, -103.5, -103.25, -103, -102.75, -102.5, -102.25, 
    -102, -101.75, -101.5, -101.25, -101, -100.75, -100.5, -100.25, -100, 
    -99.75, -99.5, -99.25, -99, -98.75, -98.5, -98.25, -98, -97.75, -97.5, 
    -97.25, -97, -96.75, -96.5, -96.25, -96, -95.75, -95.5, -95.25, -95, 
    -94.75, -94.5, -94.25, -94, -93.75, -93.5, -93.25, -93, -92.75, -92.5, 
    -92.25, -92, -91.75, -91.5, -91.25, -91, -90.75, -90.5, -90.25, -90, 
    -89.75, -89.5, -89.25, -89, -88.75, -88.5, -88.25, -88, -87.75, -87.5, 
    -87.25, -87, -86.75, -86.5, -86.25, -86, -85.75, -85.5, -85.25, -85, 
    -84.75, -84.5, -84.25, -84, -83.75, -83.5, -83.25, -83, -82.75, -82.5, 
    -82.25, -82, -81.75, -81.5, -81.25, -81, -80.75, -80.5, -80.25, -80, 
    -79.75, -79.5, -79.25, -79, -78.75, -78.5, -78.25, -78, -77.75, -77.5, 
    -77.25, -77, -76.75, -76.5, -76.25, -76, -75.75, -75.5, -75.25, -75, 
    -74.75, -74.5, -74.25, -74, -73.75, -73.5, -73.25, -73, -72.75, -72.5, 
    -72.25, -72, -71.75, -71.5, -71.25, -71, -70.75, -70.5, -70.25, -70, 
    -69.75, -69.5, -69.25, -69, -68.75, -68.5, -68.25, -68, -67.75, -67.5, 
    -67.25, -67, -66.75, -66.5, -66.25, -66, -65.75, -65.5, -65.25, -65, 
    -64.75, -64.5, -64.25, -64, -63.75, -63.5, -63.25, -63, -62.75, -62.5, 
    -62.25, -62, -61.75, -61.5, -61.25, -61, -60.75, -60.5, -60.25, -60, 
    -59.75, -59.5, -59.25, -59, -58.75, -58.5, -58.25, -58, -57.75, -57.5, 
    -57.25, -57, -56.75, -56.5, -56.25, -56, -55.75, -55.5, -55.25, -55, 
    -54.75, -54.5, -54.25, -54, -53.75, -53.5, -53.25, -53, -52.75, -52.5, 
    -52.25, -52, -51.75, -51.5, -51.25, -51, -50.75, -50.5, -50.25, -50, 
    -49.75, -49.5, -49.25, -49, -48.75, -48.5, -48.25, -48, -47.75, -47.5, 
    -47.25, -47, -46.75, -46.5, -46.25, -46, -45.75, -45.5, -45.25, -45, 
    -44.75, -44.5, -44.25, -44, -43.75, -43.5, -43.25, -43, -42.75, -42.5, 
    -42.25, -42, -41.75, -41.5, -41.25, -41, -40.75, -40.5, -40.25, -40, 
    -39.75, -39.5, -39.25, -39, -38.75, -38.5, -38.25, -38, -37.75, -37.5, 
    -37.25, -37, -36.75, -36.5, -36.25, -36, -35.75, -35.5, -35.25, -35, 
    -34.75, -34.5, -34.25, -34, -33.75, -33.5, -33.25, -33, -32.75, -32.5, 
    -32.25, -32, -31.75, -31.5, -31.25, -31, -30.75, -30.5, -30.25, -30, 
    -29.75, -29.5, -29.25, -29, -28.75, -28.5, -28.25, -28, -27.75, -27.5, 
    -27.25, -27, -26.75, -26.5, -26.25, -26, -25.75, -25.5, -25.25, -25, 
    -24.75, -24.5, -24.25, -24, -23.75, -23.5, -23.25, -23, -22.75, -22.5, 
    -22.25, -22, -21.75, -21.5, -21.25, -21, -20.75, -20.5, -20.25, -20, 
    -19.75, -19.5, -19.25, -19, -18.75, -18.5, -18.25, -18, -17.75, -17.5, 
    -17.25, -17, -16.75, -16.5, -16.25, -16, -15.75, -15.5, -15.25, -15, 
    -14.75, -14.5, -14.25, -14, -13.75, -13.5, -13.25, -13, -12.75, -12.5, 
    -12.25, -12, -11.75, -11.5, -11.25, -11, -10.75, -10.5, -10.25, -10, 
    -9.75, -9.5, -9.25, -9, -8.75, -8.5, -8.25, -8, -7.75, -7.5, -7.25, -7, 
    -6.75, -6.5, -6.25, -6, -5.75, -5.5, -5.25, -5, -4.75, -4.5, -4.25, -4, 
    -3.75, -3.5, -3.25, -3, -2.75, -2.5, -2.25, -2, -1.75, -1.5, -1.25, -1, 
    -0.75, -0.5, -0.25, 0, 0.25, 0.5, 0.75, 1, 1.25, 1.5, 1.75, 2, 2.25, 2.5, 
    2.75, 3, 3.25, 3.5, 3.75, 4, 4.25, 4.5, 4.75, 5, 5.25, 5.5, 5.75, 6, 
    6.25, 6.5, 6.75, 7, 7.25, 7.5, 7.75, 8, 8.25, 8.5, 8.75, 9, 9.25, 9.5, 
    9.75, 10, 10.25, 10.5, 10.75, 11, 11.25, 11.5, 11.75, 12, 12.25, 12.5, 
    12.75, 13, 13.25, 13.5, 13.75, 14, 14.25, 14.5, 14.75, 15, 15.25, 15.5, 
    15.75, 16, 16.25, 16.5, 16.75, 17, 17.25, 17.5, 17.75, 18, 18.25, 18.5, 
    18.75, 19, 19.25, 19.5, 19.75, 20, 20.25, 20.5, 20.75, 21, 21.25, 21.5, 
    21.75, 22, 22.25, 22.5, 22.75, 23, 23.25, 23.5, 23.75, 24, 24.25, 24.5, 
    24.75, 25, 25.25, 25.5, 25.75, 26, 26.25, 26.5, 26.75, 27, 27.25, 27.5, 
    27.75, 28, 28.25, 28.5, 28.75, 29, 29.25, 29.5, 29.75, 30, 30.25, 30.5, 
    30.75, 31, 31.25, 31.5, 31.75, 32, 32.25, 32.5, 32.75, 33, 33.25, 33.5, 
    33.75, 34, 34.25, 34.5, 34.75, 35, 35.25, 35.5, 35.75, 36, 36.25, 36.5, 
    36.75, 37, 37.25, 37.5, 37.75, 38, 38.25, 38.5, 38.75, 39, 39.25, 39.5, 
    39.75, 40, 40.25, 40.5, 40.75, 41, 41.25, 41.5, 41.75, 42, 42.25, 42.5, 
    42.75, 43, 43.25, 43.5, 43.75, 44, 44.25, 44.5, 44.75, 45, 45.25, 45.5, 
    45.75, 46, 46.25, 46.5, 46.75, 47, 47.25, 47.5, 47.75, 48, 48.25, 48.5, 
    48.75, 49, 49.25, 49.5, 49.75, 50, 50.25, 50.5, 50.75, 51, 51.25, 51.5, 
    51.75, 52, 52.25, 52.5, 52.75, 53, 53.25, 53.5, 53.75, 54, 54.25, 54.5, 
    54.75, 55, 55.25, 55.5, 55.75, 56, 56.25, 56.5, 56.75, 57, 57.25, 57.5, 
    57.75, 58, 58.25, 58.5, 58.75, 59, 59.25, 59.5, 59.75, 60 ;

 yh = -14.3476556382336, -14.1053228834302, -13.862732304759, 
    -13.6198879813569, -13.3767940148509, -13.1334545290505, 
    -12.889873669635, -12.6460556038367, -12.4020045201193, -12.1577246278516 ;

 yq = -88.57, -88.4717626572265, -88.3735253144531, -88.2752879716797, 
    -88.1770506289062, -88.0788132861328, -87.9805759433593, 
    -87.8823386005859, -87.7841012578124, -87.685863915039, 
    -87.5876265722655, -87.4893892294921, -87.3911518867186, 
    -87.2929145439452, -87.1946772011717, -87.0964398583983, 
    -86.9982025156249, -86.8999651728514, -86.801727830078, 
    -86.7034904873045, -86.6052531445311, -86.5070158017576, 
    -86.4087784589842, -86.3105411162107, -86.2123037734373, 
    -86.1140664306638, -86.0158290878904, -85.917591745117, 
    -85.8193544023435, -85.7211170595701, -85.6228797167966, 
    -85.5246423740232, -85.4264050312497, -85.3281676884763, 
    -85.2299303457028, -85.1316930029294, -85.0334556601559, 
    -84.9352183173825, -84.836980974609, -84.7387436318356, 
    -84.6405062890622, -84.5422689462887, -84.4440316035153, 
    -84.3457942607418, -84.2475569179684, -84.1493195751949, 
    -84.0510822324215, -83.952844889648, -83.8546075468746, 
    -83.7563702041011, -83.6581328613277, -83.5598955185542, 
    -83.4616581757808, -83.3634208330074, -83.2651834902339, 
    -83.1669461474605, -83.068708804687, -82.9704714619136, 
    -82.8722341191401, -82.7739967763667, -82.6757594335932, 
    -82.5775220908198, -82.4792847480463, -82.3810474052729, 
    -82.2828100624995, -82.184572719726, -82.0863353769526, 
    -81.9880980341791, -81.8898606914057, -81.7916233486322, 
    -81.6933860058588, -81.5951486630853, -81.4969113203119, 
    -81.3986739775384, -81.300436634765, -81.2021992919915, 
    -81.1039619492181, -81.0057246064447, -80.9074872636712, 
    -80.8092499208978, -80.7110125781243, -80.6127752353509, 
    -80.5145378925774, -80.416300549804, -80.3180632070305, 
    -80.2198258642571, -80.1215885214836, -80.0233511787102, 
    -79.9251138359367, -79.8268764931633, -79.7286391503899, 
    -79.6304018076164, -79.532164464843, -79.4339271220695, 
    -79.3356897792961, -79.2374524365226, -79.1392150937492, 
    -79.0409777509757, -78.9427404082023, -78.8445030654288, 
    -78.7462657226554, -78.6480283798819, -78.5497910371085, 
    -78.4515536943351, -78.3533163515616, -78.2550790087882, 
    -78.1568416660147, -78.0586043232413, -77.9603669804678, 
    -77.8621296376944, -77.7638922949209, -77.6656549521475, 
    -77.567417609374, -77.4691802666006, -77.3709429238272, 
    -77.2727055810537, -77.1744682382803, -77.0762308955068, 
    -76.9779935527334, -76.8797562099599, -76.7815188671865, 
    -76.683281524413, -76.5850441816396, -76.4868068388661, 
    -76.3885694960927, -76.2903321533192, -76.1920948105458, 
    -76.0938574677724, -75.9956201249989, -75.8973827822255, 
    -75.799145439452, -75.7009080966786, -75.6026707539051, 
    -75.5044334111317, -75.4061960683582, -75.3079587255848, 
    -75.2097213828113, -75.1114840400379, -75.0132466972644, 
    -74.915009354491, -74.8167720117176, -74.7185346689441, 
    -74.6202973261707, -74.5220599833972, -74.4238226406238, 
    -74.3255852978503, -74.2273479550769, -74.1291106123034, -74.03087326953, 
    -73.9326359267565, -73.8343985839831, -73.7361612412097, 
    -73.6379238984362, -73.5396865556628, -73.4414492128893, 
    -73.3432118701159, -73.2449745273424, -73.146737184569, 
    -73.0484998417955, -72.9502624990221, -72.8520251562486, 
    -72.7537878134752, -72.6555504707017, -72.5573131279283, 
    -72.4590757851549, -72.3608384423814, -72.262601099608, 
    -72.1643637568345, -72.0661264140611, -71.9678890712876, 
    -71.8696517285142, -71.7714143857407, -71.6731770429673, 
    -71.5749397001938, -71.4767023574204, -71.3784650146469, 
    -71.2802276718735, -71.1819903291001, -71.0837529863266, 
    -70.9855156435532, -70.8872783007797, -70.7890409580063, 
    -70.6908036152328, -70.5925662724594, -70.4943289296859, 
    -70.3960915869125, -70.297854244139, -70.1996169013656, 
    -70.1013795585922, -70.0031422158187, -69.9049048730453, 
    -69.8066675302718, -69.7084301874984, -69.6101928447249, 
    -69.5119555019515, -69.413718159178, -69.3154808164046, 
    -69.2172434736311, -69.1190061308577, -69.0207687880842, 
    -68.9225314453108, -68.8242941025374, -68.7260567597639, 
    -68.6278194169905, -68.529582074217, -68.4313447314436, 
    -68.3331073886701, -68.2348700458967, -68.1366327031232, 
    -68.0383953603498, -67.9401580175763, -67.8419206748029, 
    -67.7436833320294, -67.645445989256, -67.5472086464826, 
    -67.4489713037091, -67.3507339609357, -67.2524966181622, 
    -67.1542592753888, -67.0560219326153, -66.9577845898419, 
    -66.8595472470684, -66.7611033247456, -66.6622639175771, 
    -66.5630277320751, -66.4633934743105, -66.3633598499694, 
    -66.2629255644095, -66.1620893227181, -66.0608498297698, 
    -65.9592057902861, -65.8571559088953, -65.7546988901932, 
    -65.6518334388049, -65.5485582594471, -65.4448720569916, 
    -65.3407735365292, -65.2362614034349, -65.1313343634339, 
    -65.0259911226682, -64.9202303877641, -64.8140508659012, 
    -64.7074512648812, -64.6004302931986, -64.4929866601119, 
    -64.3851190757157, -64.2768262510133, -64.1681068979915, 
    -64.0589597296948, -63.9493834603014, -63.8393768052001, 
    -63.7289384810678, -63.6180672059484, -63.5067616993321, 
    -63.3950206822365, -63.2828428772874, -63.1702270088021, 
    -63.0571718028725, -62.9436759874495, -62.8297382924289, 
    -62.7153574497375, -62.600532193421, -62.485261259732, -62.3695433872201, 
    -62.2533773168219, -62.1367617919531, -62.0196955586006, 
    -61.9021773654167, -61.7842059638133, -61.6657801080578, 
    -61.5468985553701, -61.4275600660202, -61.3077634034271, 
    -61.1875073342589, -61.0667906285338, -60.9456120597223, 
    -60.8239704048502, -60.701864444603, -60.5792929634313, 
    -60.4562547496572, -60.332748595582, -60.2087732975946, 
    -60.0843276562813, -59.9594104765369, -59.8340205676764, 
    -59.7081567435483, -59.5818178226485, -59.455002628236, 
    -59.3277099884489, -59.1999387364222, -59.0716877104066, 
    -58.9429557538877, -58.8137417157078, -58.6840444501872, 
    -58.5538628172478, -58.4231956825373, -58.2920419175544, 
    -58.160400399776, -58.0282700127841, -57.8956496463955, -57.762538196791, 
    -57.6289345666471, -57.4948376652679, -57.3602464087187, 
    -57.2251597199603, -57.0895765289849, -56.9534957729527, 
    -56.8169163963301, -56.679837351028, -56.5422575965431, 
    -56.4041761000982, -56.265591836785, -56.1265037897078, 
    -55.9869109501277, -55.8468123176089, -55.7062069001651, 
    -55.5650937144078, -55.4234717856951, -55.2813401482819, 
    -55.1386978454716, -54.9955439297677, -54.8518774630279, 
    -54.7076975166181, -54.5630031715685, -54.4177935187296, 
    -54.2720676589303, -54.1258247031364, -53.9790637726108, 
    -53.8317839990738, -53.683984524865, -53.5356645031064, 
    -53.3868230978662, -53.2374594843233, -53.0875728489336, 
    -52.9371623895964, -52.7862273158227, -52.6347668489031, 
    -52.4827802220782, -52.3302666807091, -52.1772254824485, 
    -52.0236558974136, -51.8695572083592, -51.7149287108517, 
    -51.5597697134448, -51.4040795378545, -51.2478575191369, 
    -51.0911030058648, -50.9338153603067, -50.7759939586058, 
    -50.6176381909598, -50.4587474618019, -50.2993211899819, 
    -50.1393588089485, -49.9788597669322, -49.8178235271288, 
    -49.6562495678833, -49.4941373828755, -49.3314864813044, 
    -49.1682963880751, -49.0045666439851, -48.8402968059115, 
    -48.6754864469987, -48.5101351568465, -48.3442425416991, 
    -48.1778082246342, -48.0108318457522, -47.8433130623667, 
    -47.6752515491949, -47.5066469985477, -47.3374991205218, 
    -47.1678076431901, -46.9975723127939, -46.8267928939348, 
    -46.6554691697666, -46.4836009421878, -46.3111880320339, 
    -46.1382302792701, -45.964727543184, -45.790679702578, -45.6160866559627, 
    -45.4409483217492, -45.2652646384418, -45.089035564831, 
    -44.9122610801857, -44.7349411844457, -44.557075898414, 
    -44.3786652639488, -44.1997093441552, -44.0202082235765, 
    -43.8401620083859, -43.6595708265764, -43.4784348281518, 
    -43.2967541853167, -43.1145290926651, -42.9317597673704, 
    -42.7484464493728, -42.5645894015674, -42.3801889099915, 
    -42.1952452840104, -42.0097588565035, -41.8237299840487, 
    -41.6371590471069, -41.4500464502048, -41.262392622117, 
    -41.0741980160475, -40.8854631098099, -40.6961884060064, 
    -40.5063744322059, -40.3160217411211, -40.1251309107839, -39.93370254472, 
    -39.741737272122, -39.5492357480213, -39.3561986534582, 
    -39.1626266956511, -38.9685206081638, -38.7738811510716, 
    -38.578709111125, -38.383005301913, -38.1867705640235, -37.9900057652026, 
    -37.792711800512, -37.5948895924842, -37.3965400912763, 
    -37.1976642748214, -36.998263148978, -36.7983377476777, 
    -36.5978891330702, -36.3969183956667, -36.1954266544803, 
    -35.9934150571649, -35.7908847801515, -35.5878370287813, 
    -35.3842730374377, -35.1801940696746, -34.975601418343, 
    -34.7704964057139, -34.5648803835998, -34.3587547334724, 
    -34.152120866578, -33.94498022405, -33.7373342770182, -33.5291845267155, 
    -33.3205325045815, -33.1113797723624, -32.901727922209, 
    -32.6915785767703, -32.4809333892845, -32.2697940436663, 
    -32.0581622545914, -31.8460397675771, -31.6334283590593, 
    -31.4203298364668, -31.206746038291, -30.9926788341526, 
    -30.7781301248646, -30.5631018424912, -30.3475959504032, 
    -30.1316144433295, -29.9151593474048, -29.6982327202131, 
    -29.4808366508275, -29.2629732598456, -29.0446446994212, 
    -28.825853153292, -28.6066008368019, -28.3868899969211, 
    -28.1667229122599, -27.9461018930793, -27.7250292812972, -27.50350745049, 
    -27.281538805889, -27.0591257843741, -26.8362708544607, 
    -26.6129765162842, -26.3892453015782, -26.1650797736486, 
    -25.9404825273438, -25.7154561890184, -25.4900034164941, 
    -25.2641268990141, -25.0378293571939, -24.8111135429665, 
    -24.5839822395226, -24.3564382612468, -24.1284844536475, 
    -23.9001236932831, -23.671358887682, -23.4421929752584, 
    -23.2126289252224, -22.9826697374859, -22.7523184425622, 
    -22.5215781014612, -22.2904518055793, -22.0589426765843, 
    -21.8270538662944, -21.5947885565529, -21.362149959097, 
    -21.1291413154218, -20.8957658966385, -20.6620270033283, 
    -20.4279279653895, -20.1934721418813, -19.9586629208602, 
    -19.7235037192131, -19.4879979824837, -19.252149184694, -19.015960828161, 
    -18.7794364433077, -18.5425795884684, -18.3053938496899, 
    -18.0678828405262, -17.8300502018287, -17.5918996015312, 
    -17.3534347344289, -17.1146593219533, -16.8755771119409, 
    -16.6361918783977, -16.3965074212573, -16.1565275661354, 
    -15.9162561640777, -15.6756970913041, -15.4348542489463, 
    -15.1937315627822, -14.9523329829638, -14.7106624837407, 
    -14.4687240631789, -14.2265217428746, -13.9840595676627, 
    -13.7413416053212, -13.4983719462701, -13.2551547032665, 
    -13.011694011094, -12.7679940262485, -12.5240589266184, -12.279892911161, 
    -12.0355001995743, -11.7908850319639, -11.5460516685066, 
    -11.3010043891084, -11.0557474930589, -10.810285298682, 
    -10.5646221429814, -10.3187623812829, -10.0727103868724, 
    -9.82647055062974, -9.5800472806593, -9.33344500191614, 
    -9.08666815582889, -8.83972119991878, -8.59260860741517, 
    -8.3453348668676, -8.0979044817544, -7.850321970088, -7.60259186401695, 
    -7.35471870942481, -7.10670706552594, -6.85856150445826, 
    -6.61028661087316, -6.36188698152251, -6.11336722484299, 
    -5.86473196053772, -5.61598581915533, -5.36713344166667, 
    -5.11817947903895, -4.86912859180776, -4.61998544964686, 
    -4.37075473093582, -4.12144112232571, -3.87204931830292, 
    -3.62258402075114, -3.3730499385116, -3.1234517869418, -2.87379428747266, 
    -2.6240821671643, -2.37432015826051, -2.12451299774205, 
    -1.87466542687879, -1.62478219078095, -1.37486803794932, 
    -1.12492771982485, -0.874965990337434, -0.624987605454166, 
    -0.37499732272713, -0.124999900840802, 0.124999900840802, 
    0.37499732272713, 0.624987605454166, 0.874965990337434, 1.12492771982485, 
    1.37486803794932, 1.62478219078095, 1.87466542687879, 2.12451299774205, 
    2.37432015826051, 2.6240821671643, 2.87379428747266, 3.1234517869418, 
    3.3730499385116, 3.62258402075114, 3.87204931830292, 4.12144112232571, 
    4.37075473093582, 4.61998544964686, 4.86912859180776, 5.11817947903895, 
    5.36713344166667, 5.61598581915533, 5.86473196053772, 6.11336722484299, 
    6.36188698152251, 6.61028661087316, 6.85856150445826, 7.10670706552594, 
    7.35471870942481, 7.60259186401695, 7.850321970088, 8.0979044817544, 
    8.3453348668676, 8.59260860741517, 8.83972119991878, 9.08666815582889, 
    9.33344500191614, 9.5800472806593, 9.82647055062974, 10.0727103868724, 
    10.3187623812829, 10.5646221429814, 10.810285298682, 11.0557474930589, 
    11.3010043891084, 11.5460516685066, 11.7908850319639, 12.0355001995743, 
    12.279892911161, 12.5240589266184, 12.7679940262485, 13.011694011094, 
    13.2551547032665, 13.4983719462701, 13.7413416053212, 13.9840595676627, 
    14.2265217428746, 14.4687240631789, 14.7106624837407, 14.9523329829638, 
    15.1937315627822, 15.4348542489463, 15.6756970913041, 15.9162561640777, 
    16.1565275661354, 16.3965074212573, 16.6361918783977, 16.8755771119409, 
    17.1146593219533, 17.3534347344289, 17.5918996015312, 17.8300502018287, 
    18.0678828405262, 18.3053938496899, 18.5425795884684, 18.7794364433077, 
    19.015960828161, 19.252149184694, 19.4879979824837, 19.7235037192131, 
    19.9586629208602, 20.1934721418813, 20.4279279653895, 20.6620270033283, 
    20.8957658966385, 21.1291413154218, 21.362149959097, 21.5947885565529, 
    21.8270538662944, 22.0589426765843, 22.2904518055793, 22.5215781014612, 
    22.7523184425622, 22.9826697374859, 23.2126289252224, 23.4421929752584, 
    23.671358887682, 23.9001236932831, 24.1284844536475, 24.3564382612468, 
    24.5839822395226, 24.8111135429665, 25.0378293571939, 25.2641268990141, 
    25.4900034164941, 25.7154561890184, 25.9404825273438, 26.1650797736486, 
    26.3892453015782, 26.6129765162842, 26.8362708544607, 27.0591257843741, 
    27.281538805889, 27.50350745049, 27.7250292812972, 27.9461018930793, 
    28.1667229122599, 28.3868899969211, 28.6066008368019, 28.825853153292, 
    29.0446446994212, 29.2629732598456, 29.4808366508275, 29.6982327202131, 
    29.9151593474048, 30.1316144433295, 30.3475959504032, 30.5631018424912, 
    30.7781301248646, 30.9926788341526, 31.206746038291, 31.4203298364668, 
    31.6334283590593, 31.8460397675771, 32.0581622545914, 32.2697940436663, 
    32.4809333892845, 32.6915785767703, 32.901727922209, 33.1113797723624, 
    33.3205325045815, 33.5291845267155, 33.7373342770182, 33.94498022405, 
    34.152120866578, 34.3587547334724, 34.5648803835998, 34.7704964057139, 
    34.975601418343, 35.1801940696746, 35.3842730374377, 35.5878370287813, 
    35.7908847801515, 35.9934150571649, 36.1954266544803, 36.3969183956667, 
    36.5978891330702, 36.7983377476777, 36.998263148978, 37.1976642748214, 
    37.3965400912763, 37.5948895924842, 37.792711800512, 37.9900057652026, 
    38.1867705640235, 38.383005301913, 38.578709111125, 38.7738811510716, 
    38.9685206081638, 39.1626266956511, 39.3561986534582, 39.5492357480213, 
    39.741737272122, 39.93370254472, 40.1251309107839, 40.3160217411211, 
    40.5063744322059, 40.6961884060064, 40.8854631098099, 41.0741980160475, 
    41.262392622117, 41.4500464502048, 41.6371590471069, 41.8237299840487, 
    42.0097588565035, 42.1952452840104, 42.3801889099915, 42.5645894015674, 
    42.7484464493728, 42.9317597673704, 43.1145290926651, 43.2967541853167, 
    43.4784348281518, 43.6595708265764, 43.8401620083859, 44.0202082235765, 
    44.1997093441552, 44.3786652639488, 44.557075898414, 44.7349411844457, 
    44.9122610801857, 45.089035564831, 45.2652646384418, 45.4409483217492, 
    45.6160866559627, 45.790679702578, 45.964727543184, 46.1382302792701, 
    46.3111880320339, 46.4836009421878, 46.6554691697666, 46.8267928939348, 
    46.9975723127939, 47.1678076431901, 47.3374991205218, 47.5066469985477, 
    47.6752515491949, 47.8433130623667, 48.0108318457522, 48.1778082246342, 
    48.3442425416991, 48.5101351568465, 48.6754864469987, 48.8402968059115, 
    49.0045666439851, 49.1682963880751, 49.3314864813044, 49.4941373828755, 
    49.6562495678833, 49.8178235271288, 49.9788597669322, 50.1393588089485, 
    50.2993211899819, 50.4587474618019, 50.6176381909598, 50.7759939586058, 
    50.9338153603067, 51.0911030058648, 51.2478575191369, 51.4040795378545, 
    51.5597697134448, 51.7149287108517, 51.8695572083592, 52.0236558974136, 
    52.1772254824485, 52.3302666807091, 52.4827802220782, 52.6347668489031, 
    52.7862273158227, 52.9371623895964, 53.0875728489336, 53.2374594843233, 
    53.3868230978662, 53.5356645031064, 53.683984524865, 53.8317839990738, 
    53.9790637726108, 54.1258247031364, 54.2720676589303, 54.4177935187296, 
    54.5630031715685, 54.7076975166181, 54.8518774630279, 54.9955439297677, 
    55.1386978454716, 55.2813401482819, 55.4234717856951, 55.5650937144078, 
    55.7062069001651, 55.8468123176089, 55.9869109501277, 56.1265037897078, 
    56.265591836785, 56.4041761000982, 56.5422575965431, 56.679837351028, 
    56.8169163963301, 56.9534957729527, 57.0895765289849, 57.2251597199603, 
    57.3602464087187, 57.4948376652679, 57.6289345666471, 57.762538196791, 
    57.8956496463955, 58.0282700127841, 58.160400399776, 58.2920419175544, 
    58.4231956825373, 58.5538628172478, 58.6840444501872, 58.8137417157078, 
    58.9429557538877, 59.0716877104066, 59.1999387364222, 59.3277099884489, 
    59.455002628236, 59.5818178226485, 59.7081567435483, 59.8340205676764, 
    59.9594104765369, 60.0843276562813, 60.2087732975946, 60.332748595582, 
    60.4562547496572, 60.5792929634313, 60.701864444603, 60.8239704048502, 
    60.9456120597223, 61.0667906285338, 61.1875073342589, 61.3077634034271, 
    61.4275600660202, 61.5468985553701, 61.6657801080578, 61.7842059638133, 
    61.9021773654167, 62.0196955586006, 62.1367617919531, 62.2533773168219, 
    62.3695433872201, 62.485261259732, 62.600532193421, 62.7153574497375, 
    62.8297382924289, 62.9436759874495, 63.0571718028725, 63.1702270088021, 
    63.2828428772874, 63.3950206822365, 63.5067616993321, 63.6180672059484, 
    63.7289384810678, 63.8393768052001, 63.9493834603014, 64.0589597296948, 
    64.1670473974877, 64.2751350652807, 64.3832227330736, 64.4913104008666, 
    64.5993980686595, 64.7074857364524, 64.8155734042454, 64.9236610720383, 
    65.0317487398313, 65.1398364076242, 65.2479240754171, 65.3560117432101, 
    65.464099411003, 65.5721870787959, 65.6802747465889, 65.7883624143818, 
    65.8964500821748, 66.0045377499677, 66.1126254177607, 66.2207130855536, 
    66.3288007533465, 66.4368884211394, 66.5449760889324, 66.6530637567253, 
    66.7611514245183, 66.8692390923112, 66.9773267601041, 67.0854144278971, 
    67.19350209569, 67.301589763483, 67.4096774312759, 67.5177650990688, 
    67.6258527668618, 67.7339404346547, 67.8420281024476, 67.9501157702406, 
    68.0582034380335, 68.1662911058265, 68.2743787736194, 68.3824664414123, 
    68.4905541092053, 68.5986417769982, 68.7067294447912, 68.8148171125841, 
    68.922904780377, 69.03099244817, 69.1390801159629, 69.2471677837559, 
    69.3552554515488, 69.4633431193417, 69.5714307871347, 69.6795184549276, 
    69.7876061227205, 69.8956937905135, 70.0037814583064, 70.1118691260994, 
    70.2199567938923, 70.3280444616852, 70.4361321294782, 70.5442197972711, 
    70.652307465064, 70.760395132857, 70.8684828006499, 70.9765704684429, 
    71.0846581362358, 71.1927458040287, 71.3008334718217, 71.4089211396146, 
    71.5170088074075, 71.6250964752005, 71.7331841429934, 71.8412718107864, 
    71.9493594785793, 72.0574471463722, 72.1655348141652, 72.2736224819581, 
    72.3817101497511, 72.489797817544, 72.5978854853369, 72.7059731531299, 
    72.8140608209228, 72.9221484887157, 73.0302361565087, 73.1383238243016, 
    73.2464114920946, 73.3544991598875, 73.4625868276804, 73.5706744954734, 
    73.6787621632663, 73.7868498310593, 73.8949374988522, 74.0030251666451, 
    74.1111128344381, 74.219200502231, 74.3272881700239, 74.4353758378169, 
    74.5434635056098, 74.6515511734028, 74.7596388411957, 74.8677265089886, 
    74.9758141767816, 75.0839018445745, 75.1919895123675, 75.3000771801604, 
    75.4081648479533, 75.5162525157463, 75.6243401835392, 75.7324278513321, 
    75.8405155191251, 75.948603186918, 76.056690854711, 76.1647785225039, 
    76.2728661902968, 76.3809538580898, 76.4890415258827, 76.5971291936756, 
    76.7052168614686, 76.8133045292615, 76.9213921970545, 77.0294798648474, 
    77.1375675326403, 77.2456552004333, 77.3537428682262, 77.4618305360192, 
    77.5699182038121, 77.678005871605, 77.786093539398, 77.8941812071909, 
    78.0022688749839, 78.1103565427768, 78.2184442105697, 78.3265318783627, 
    78.4346195461556, 78.5427072139485, 78.6507948817415, 78.7588825495344, 
    78.8669702173273, 78.9750578851203, 79.0831455529132, 79.1912332207062, 
    79.2993208884991, 79.407408556292, 79.515496224085, 79.6235838918779, 
    79.7316715596709, 79.8397592274638, 79.9478468952567, 80.0559345630497, 
    80.1640222308426, 80.2721098986355, 80.3801975664285, 80.4882852342214, 
    80.5963729020144, 80.7044605698073, 80.8125482376002, 80.9206359053932, 
    81.0287235731861, 81.1368112409791, 81.244898908772, 81.3529865765649, 
    81.4610742443579, 81.5691619121508, 81.6772495799437, 81.7853372477367, 
    81.8934249155296, 82.0015125833226, 82.1096002511155, 82.2176879189084, 
    82.3257755867014, 82.4338632544943, 82.5419509222873, 82.6500385900802, 
    82.7581262578731, 82.8662139256661, 82.974301593459, 83.0823892612519, 
    83.1904769290449, 83.2985645968378, 83.4066522646308, 83.5147399324237, 
    83.6228276002166, 83.7309152680096, 83.8390029358025, 83.9470906035955, 
    84.0551782713884, 84.1632659391813, 84.2713536069743, 84.3794412747672, 
    84.4875289425601, 84.5956166103531, 84.703704278146, 84.811791945939, 
    84.9198796137319, 85.0279672815248, 85.1360549493178, 85.2441426171107, 
    85.3522302849037, 85.4603179526966, 85.5684056204895, 85.6764932882825, 
    85.7845809560754, 85.8926686238683, 86.0007562916613, 86.1088439594542, 
    86.2169316272472, 86.3250192950401, 86.433106962833, 86.541194630626, 
    86.6492822984189, 86.7573699662119, 86.8654576340048, 86.9735453017977, 
    87.0816329695907, 87.1897206373836, 87.2978083051765, 87.4058959729695, 
    87.5139836407624, 87.6220713085554, 87.7301589763483, 87.8382466441412, 
    87.9463343119342, 88.0544219797271, 88.1625096475201, 88.270597315313, 
    88.3786849831059, 88.4867726508989, 88.5948603186918, 88.7029479864847, 
    88.8110356542777, 88.9191233220706, 89.0272109898635, 89.1352986576565, 
    89.2433863254494, 89.3514739932424, 89.4595616610353, 89.5676493288282, 
    89.6757369966212, 89.7838246644141, 89.891912332207, 90 ;

 zi = 0, 2, 4, 6, 8, 10, 12, 14, 16.01, 18.02, 20.04, 22.07, 24.12, 26.2, 
    28.31, 30.46, 32.67, 34.95, 37.32, 39.8, 42.41, 45.18, 48.13, 51.3, 
    54.73, 58.47, 62.56, 67.05, 72, 77.48, 83.55, 90.29, 97.79, 106.13, 
    115.41, 125.74, 137.23, 150, 164.19, 179.93, 197.38, 216.69, 238.04, 
    261.6, 287.57, 316.15, 347.56, 382.03, 419.8, 461.12, 506.26, 555.51, 
    609.16, 667.53, 730.95, 799.76, 874.32, 955, 1042.21, 1136.35, 1237.86, 
    1347.19, 1464.81, 1591.21, 1726.89, 1872.39, 2028.26, 2195.07, 2373.42, 
    2563.93, 2767.24, 2984.02, 3214.95, 3460.75, 3722.17, 6500 ;

 zl = 1, 3, 5, 7, 9, 11, 13, 15.005, 17.015, 19.03, 21.055, 23.095, 25.16, 
    27.255, 29.385, 31.565, 33.81, 36.135, 38.56, 41.105, 43.795, 46.655, 
    49.715, 53.015, 56.6, 60.515, 64.805, 69.525, 74.74, 80.515, 86.92, 
    94.04, 101.96, 110.77, 120.575, 131.485, 143.615, 157.095, 172.06, 
    188.655, 207.035, 227.365, 249.82, 274.585, 301.86, 331.855, 364.795, 
    400.915, 440.46, 483.69, 530.885, 582.335, 638.345, 699.24, 765.355, 
    837.04, 914.66, 998.605, 1089.28, 1187.105, 1292.525, 1406, 1528.01, 
    1659.05, 1799.64, 1950.325, 2111.665, 2284.245, 2468.675, 2665.585, 
    2875.63, 3099.485, 3337.85, 3591.46, 5111.085 ;
}
